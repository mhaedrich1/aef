module dtc_split875_bm61 (
	input  wire [12-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node7;
	wire [11-1:0] node8;
	wire [11-1:0] node9;
	wire [11-1:0] node10;
	wire [11-1:0] node12;
	wire [11-1:0] node15;
	wire [11-1:0] node16;
	wire [11-1:0] node20;
	wire [11-1:0] node21;
	wire [11-1:0] node22;
	wire [11-1:0] node25;
	wire [11-1:0] node28;
	wire [11-1:0] node31;
	wire [11-1:0] node32;
	wire [11-1:0] node33;
	wire [11-1:0] node34;
	wire [11-1:0] node37;
	wire [11-1:0] node40;
	wire [11-1:0] node41;
	wire [11-1:0] node45;
	wire [11-1:0] node46;
	wire [11-1:0] node47;
	wire [11-1:0] node50;
	wire [11-1:0] node53;
	wire [11-1:0] node54;
	wire [11-1:0] node57;
	wire [11-1:0] node60;
	wire [11-1:0] node61;
	wire [11-1:0] node62;
	wire [11-1:0] node63;
	wire [11-1:0] node64;
	wire [11-1:0] node67;
	wire [11-1:0] node70;
	wire [11-1:0] node71;
	wire [11-1:0] node75;
	wire [11-1:0] node76;
	wire [11-1:0] node77;
	wire [11-1:0] node81;
	wire [11-1:0] node82;
	wire [11-1:0] node85;
	wire [11-1:0] node88;
	wire [11-1:0] node89;
	wire [11-1:0] node90;
	wire [11-1:0] node91;
	wire [11-1:0] node94;
	wire [11-1:0] node97;
	wire [11-1:0] node99;
	wire [11-1:0] node102;
	wire [11-1:0] node103;
	wire [11-1:0] node104;
	wire [11-1:0] node108;
	wire [11-1:0] node109;
	wire [11-1:0] node112;
	wire [11-1:0] node115;
	wire [11-1:0] node116;
	wire [11-1:0] node117;
	wire [11-1:0] node118;
	wire [11-1:0] node119;
	wire [11-1:0] node121;
	wire [11-1:0] node124;
	wire [11-1:0] node127;
	wire [11-1:0] node128;
	wire [11-1:0] node129;
	wire [11-1:0] node133;
	wire [11-1:0] node135;
	wire [11-1:0] node138;
	wire [11-1:0] node139;
	wire [11-1:0] node140;
	wire [11-1:0] node141;
	wire [11-1:0] node145;
	wire [11-1:0] node146;
	wire [11-1:0] node150;
	wire [11-1:0] node151;
	wire [11-1:0] node152;
	wire [11-1:0] node155;
	wire [11-1:0] node158;
	wire [11-1:0] node159;
	wire [11-1:0] node162;
	wire [11-1:0] node165;
	wire [11-1:0] node166;
	wire [11-1:0] node167;
	wire [11-1:0] node168;
	wire [11-1:0] node170;
	wire [11-1:0] node173;
	wire [11-1:0] node176;
	wire [11-1:0] node177;
	wire [11-1:0] node178;
	wire [11-1:0] node181;
	wire [11-1:0] node184;
	wire [11-1:0] node187;
	wire [11-1:0] node188;
	wire [11-1:0] node189;
	wire [11-1:0] node190;
	wire [11-1:0] node193;
	wire [11-1:0] node196;
	wire [11-1:0] node197;
	wire [11-1:0] node200;
	wire [11-1:0] node203;
	wire [11-1:0] node204;
	wire [11-1:0] node205;
	wire [11-1:0] node208;
	wire [11-1:0] node211;
	wire [11-1:0] node212;
	wire [11-1:0] node215;
	wire [11-1:0] node218;
	wire [11-1:0] node219;
	wire [11-1:0] node220;
	wire [11-1:0] node221;
	wire [11-1:0] node222;
	wire [11-1:0] node223;
	wire [11-1:0] node224;
	wire [11-1:0] node228;
	wire [11-1:0] node231;
	wire [11-1:0] node232;
	wire [11-1:0] node234;
	wire [11-1:0] node237;
	wire [11-1:0] node238;
	wire [11-1:0] node241;
	wire [11-1:0] node244;
	wire [11-1:0] node245;
	wire [11-1:0] node246;
	wire [11-1:0] node248;
	wire [11-1:0] node251;
	wire [11-1:0] node252;
	wire [11-1:0] node255;
	wire [11-1:0] node258;
	wire [11-1:0] node259;
	wire [11-1:0] node262;
	wire [11-1:0] node263;
	wire [11-1:0] node266;
	wire [11-1:0] node269;
	wire [11-1:0] node270;
	wire [11-1:0] node271;
	wire [11-1:0] node272;
	wire [11-1:0] node273;
	wire [11-1:0] node276;
	wire [11-1:0] node279;
	wire [11-1:0] node280;
	wire [11-1:0] node283;
	wire [11-1:0] node286;
	wire [11-1:0] node287;
	wire [11-1:0] node288;
	wire [11-1:0] node292;
	wire [11-1:0] node293;
	wire [11-1:0] node296;
	wire [11-1:0] node299;
	wire [11-1:0] node300;
	wire [11-1:0] node301;
	wire [11-1:0] node302;
	wire [11-1:0] node305;
	wire [11-1:0] node308;
	wire [11-1:0] node309;
	wire [11-1:0] node312;
	wire [11-1:0] node315;
	wire [11-1:0] node316;
	wire [11-1:0] node317;
	wire [11-1:0] node320;
	wire [11-1:0] node323;
	wire [11-1:0] node325;
	wire [11-1:0] node328;
	wire [11-1:0] node329;
	wire [11-1:0] node330;
	wire [11-1:0] node331;
	wire [11-1:0] node332;
	wire [11-1:0] node333;
	wire [11-1:0] node336;
	wire [11-1:0] node339;
	wire [11-1:0] node340;
	wire [11-1:0] node343;
	wire [11-1:0] node346;
	wire [11-1:0] node347;
	wire [11-1:0] node348;
	wire [11-1:0] node351;
	wire [11-1:0] node354;
	wire [11-1:0] node355;
	wire [11-1:0] node358;
	wire [11-1:0] node361;
	wire [11-1:0] node362;
	wire [11-1:0] node363;
	wire [11-1:0] node364;
	wire [11-1:0] node367;
	wire [11-1:0] node370;
	wire [11-1:0] node373;
	wire [11-1:0] node374;
	wire [11-1:0] node375;
	wire [11-1:0] node378;
	wire [11-1:0] node381;
	wire [11-1:0] node382;
	wire [11-1:0] node385;
	wire [11-1:0] node388;
	wire [11-1:0] node389;
	wire [11-1:0] node390;
	wire [11-1:0] node391;
	wire [11-1:0] node392;
	wire [11-1:0] node395;
	wire [11-1:0] node398;
	wire [11-1:0] node399;
	wire [11-1:0] node402;
	wire [11-1:0] node405;
	wire [11-1:0] node406;
	wire [11-1:0] node407;
	wire [11-1:0] node410;
	wire [11-1:0] node413;
	wire [11-1:0] node414;
	wire [11-1:0] node418;
	wire [11-1:0] node419;
	wire [11-1:0] node420;
	wire [11-1:0] node422;
	wire [11-1:0] node425;
	wire [11-1:0] node427;
	wire [11-1:0] node430;
	wire [11-1:0] node431;
	wire [11-1:0] node432;
	wire [11-1:0] node436;
	wire [11-1:0] node439;
	wire [11-1:0] node440;
	wire [11-1:0] node441;
	wire [11-1:0] node442;
	wire [11-1:0] node443;
	wire [11-1:0] node444;
	wire [11-1:0] node445;
	wire [11-1:0] node446;
	wire [11-1:0] node449;
	wire [11-1:0] node452;
	wire [11-1:0] node453;
	wire [11-1:0] node456;
	wire [11-1:0] node459;
	wire [11-1:0] node460;
	wire [11-1:0] node461;
	wire [11-1:0] node464;
	wire [11-1:0] node467;
	wire [11-1:0] node468;
	wire [11-1:0] node471;
	wire [11-1:0] node474;
	wire [11-1:0] node475;
	wire [11-1:0] node476;
	wire [11-1:0] node477;
	wire [11-1:0] node480;
	wire [11-1:0] node483;
	wire [11-1:0] node484;
	wire [11-1:0] node487;
	wire [11-1:0] node490;
	wire [11-1:0] node491;
	wire [11-1:0] node492;
	wire [11-1:0] node496;
	wire [11-1:0] node498;
	wire [11-1:0] node501;
	wire [11-1:0] node502;
	wire [11-1:0] node503;
	wire [11-1:0] node504;
	wire [11-1:0] node506;
	wire [11-1:0] node509;
	wire [11-1:0] node510;
	wire [11-1:0] node513;
	wire [11-1:0] node516;
	wire [11-1:0] node517;
	wire [11-1:0] node518;
	wire [11-1:0] node521;
	wire [11-1:0] node524;
	wire [11-1:0] node525;
	wire [11-1:0] node528;
	wire [11-1:0] node531;
	wire [11-1:0] node532;
	wire [11-1:0] node533;
	wire [11-1:0] node534;
	wire [11-1:0] node537;
	wire [11-1:0] node540;
	wire [11-1:0] node541;
	wire [11-1:0] node544;
	wire [11-1:0] node547;
	wire [11-1:0] node548;
	wire [11-1:0] node551;
	wire [11-1:0] node552;
	wire [11-1:0] node555;
	wire [11-1:0] node558;
	wire [11-1:0] node559;
	wire [11-1:0] node560;
	wire [11-1:0] node561;
	wire [11-1:0] node562;
	wire [11-1:0] node563;
	wire [11-1:0] node566;
	wire [11-1:0] node569;
	wire [11-1:0] node570;
	wire [11-1:0] node573;
	wire [11-1:0] node576;
	wire [11-1:0] node577;
	wire [11-1:0] node578;
	wire [11-1:0] node581;
	wire [11-1:0] node584;
	wire [11-1:0] node585;
	wire [11-1:0] node589;
	wire [11-1:0] node590;
	wire [11-1:0] node591;
	wire [11-1:0] node594;
	wire [11-1:0] node595;
	wire [11-1:0] node598;
	wire [11-1:0] node601;
	wire [11-1:0] node602;
	wire [11-1:0] node603;
	wire [11-1:0] node606;
	wire [11-1:0] node609;
	wire [11-1:0] node610;
	wire [11-1:0] node613;
	wire [11-1:0] node616;
	wire [11-1:0] node617;
	wire [11-1:0] node618;
	wire [11-1:0] node619;
	wire [11-1:0] node620;
	wire [11-1:0] node623;
	wire [11-1:0] node626;
	wire [11-1:0] node628;
	wire [11-1:0] node631;
	wire [11-1:0] node632;
	wire [11-1:0] node633;
	wire [11-1:0] node636;
	wire [11-1:0] node639;
	wire [11-1:0] node640;
	wire [11-1:0] node644;
	wire [11-1:0] node645;
	wire [11-1:0] node646;
	wire [11-1:0] node647;
	wire [11-1:0] node650;
	wire [11-1:0] node653;
	wire [11-1:0] node654;
	wire [11-1:0] node657;
	wire [11-1:0] node660;
	wire [11-1:0] node661;
	wire [11-1:0] node662;
	wire [11-1:0] node665;
	wire [11-1:0] node668;
	wire [11-1:0] node669;
	wire [11-1:0] node673;
	wire [11-1:0] node674;
	wire [11-1:0] node675;
	wire [11-1:0] node676;
	wire [11-1:0] node677;
	wire [11-1:0] node678;
	wire [11-1:0] node680;
	wire [11-1:0] node683;
	wire [11-1:0] node684;
	wire [11-1:0] node688;
	wire [11-1:0] node689;
	wire [11-1:0] node691;
	wire [11-1:0] node694;
	wire [11-1:0] node697;
	wire [11-1:0] node698;
	wire [11-1:0] node699;
	wire [11-1:0] node700;
	wire [11-1:0] node703;
	wire [11-1:0] node706;
	wire [11-1:0] node707;
	wire [11-1:0] node710;
	wire [11-1:0] node713;
	wire [11-1:0] node714;
	wire [11-1:0] node716;
	wire [11-1:0] node719;
	wire [11-1:0] node720;
	wire [11-1:0] node723;
	wire [11-1:0] node726;
	wire [11-1:0] node727;
	wire [11-1:0] node728;
	wire [11-1:0] node729;
	wire [11-1:0] node730;
	wire [11-1:0] node734;
	wire [11-1:0] node735;
	wire [11-1:0] node738;
	wire [11-1:0] node741;
	wire [11-1:0] node742;
	wire [11-1:0] node743;
	wire [11-1:0] node746;
	wire [11-1:0] node750;
	wire [11-1:0] node751;
	wire [11-1:0] node752;
	wire [11-1:0] node753;
	wire [11-1:0] node757;
	wire [11-1:0] node759;
	wire [11-1:0] node762;
	wire [11-1:0] node763;
	wire [11-1:0] node764;
	wire [11-1:0] node767;
	wire [11-1:0] node770;
	wire [11-1:0] node773;
	wire [11-1:0] node774;
	wire [11-1:0] node775;
	wire [11-1:0] node776;
	wire [11-1:0] node777;
	wire [11-1:0] node779;
	wire [11-1:0] node782;
	wire [11-1:0] node784;
	wire [11-1:0] node787;
	wire [11-1:0] node788;
	wire [11-1:0] node790;
	wire [11-1:0] node793;
	wire [11-1:0] node794;
	wire [11-1:0] node797;
	wire [11-1:0] node800;
	wire [11-1:0] node801;
	wire [11-1:0] node802;
	wire [11-1:0] node803;
	wire [11-1:0] node806;
	wire [11-1:0] node809;
	wire [11-1:0] node810;
	wire [11-1:0] node814;
	wire [11-1:0] node815;
	wire [11-1:0] node816;
	wire [11-1:0] node819;
	wire [11-1:0] node822;
	wire [11-1:0] node823;
	wire [11-1:0] node827;
	wire [11-1:0] node828;
	wire [11-1:0] node829;
	wire [11-1:0] node830;
	wire [11-1:0] node831;
	wire [11-1:0] node835;
	wire [11-1:0] node838;
	wire [11-1:0] node839;
	wire [11-1:0] node841;
	wire [11-1:0] node844;
	wire [11-1:0] node845;
	wire [11-1:0] node848;
	wire [11-1:0] node851;
	wire [11-1:0] node852;
	wire [11-1:0] node853;
	wire [11-1:0] node854;
	wire [11-1:0] node858;
	wire [11-1:0] node860;
	wire [11-1:0] node863;
	wire [11-1:0] node864;
	wire [11-1:0] node867;
	wire [11-1:0] node868;
	wire [11-1:0] node871;
	wire [11-1:0] node874;
	wire [11-1:0] node875;
	wire [11-1:0] node876;
	wire [11-1:0] node877;
	wire [11-1:0] node878;
	wire [11-1:0] node879;
	wire [11-1:0] node880;
	wire [11-1:0] node881;
	wire [11-1:0] node882;
	wire [11-1:0] node885;
	wire [11-1:0] node888;
	wire [11-1:0] node889;
	wire [11-1:0] node892;
	wire [11-1:0] node895;
	wire [11-1:0] node896;
	wire [11-1:0] node899;
	wire [11-1:0] node900;
	wire [11-1:0] node903;
	wire [11-1:0] node906;
	wire [11-1:0] node907;
	wire [11-1:0] node908;
	wire [11-1:0] node911;
	wire [11-1:0] node913;
	wire [11-1:0] node916;
	wire [11-1:0] node917;
	wire [11-1:0] node919;
	wire [11-1:0] node922;
	wire [11-1:0] node923;
	wire [11-1:0] node927;
	wire [11-1:0] node928;
	wire [11-1:0] node929;
	wire [11-1:0] node930;
	wire [11-1:0] node932;
	wire [11-1:0] node935;
	wire [11-1:0] node936;
	wire [11-1:0] node940;
	wire [11-1:0] node941;
	wire [11-1:0] node943;
	wire [11-1:0] node946;
	wire [11-1:0] node949;
	wire [11-1:0] node950;
	wire [11-1:0] node951;
	wire [11-1:0] node954;
	wire [11-1:0] node955;
	wire [11-1:0] node958;
	wire [11-1:0] node961;
	wire [11-1:0] node962;
	wire [11-1:0] node964;
	wire [11-1:0] node967;
	wire [11-1:0] node968;
	wire [11-1:0] node971;
	wire [11-1:0] node974;
	wire [11-1:0] node975;
	wire [11-1:0] node976;
	wire [11-1:0] node977;
	wire [11-1:0] node978;
	wire [11-1:0] node979;
	wire [11-1:0] node983;
	wire [11-1:0] node984;
	wire [11-1:0] node987;
	wire [11-1:0] node990;
	wire [11-1:0] node991;
	wire [11-1:0] node992;
	wire [11-1:0] node995;
	wire [11-1:0] node998;
	wire [11-1:0] node999;
	wire [11-1:0] node1002;
	wire [11-1:0] node1005;
	wire [11-1:0] node1006;
	wire [11-1:0] node1007;
	wire [11-1:0] node1008;
	wire [11-1:0] node1011;
	wire [11-1:0] node1014;
	wire [11-1:0] node1016;
	wire [11-1:0] node1019;
	wire [11-1:0] node1020;
	wire [11-1:0] node1022;
	wire [11-1:0] node1025;
	wire [11-1:0] node1027;
	wire [11-1:0] node1030;
	wire [11-1:0] node1031;
	wire [11-1:0] node1032;
	wire [11-1:0] node1033;
	wire [11-1:0] node1034;
	wire [11-1:0] node1037;
	wire [11-1:0] node1040;
	wire [11-1:0] node1041;
	wire [11-1:0] node1044;
	wire [11-1:0] node1047;
	wire [11-1:0] node1048;
	wire [11-1:0] node1051;
	wire [11-1:0] node1052;
	wire [11-1:0] node1055;
	wire [11-1:0] node1058;
	wire [11-1:0] node1059;
	wire [11-1:0] node1060;
	wire [11-1:0] node1063;
	wire [11-1:0] node1064;
	wire [11-1:0] node1068;
	wire [11-1:0] node1069;
	wire [11-1:0] node1072;
	wire [11-1:0] node1073;
	wire [11-1:0] node1076;
	wire [11-1:0] node1079;
	wire [11-1:0] node1080;
	wire [11-1:0] node1081;
	wire [11-1:0] node1082;
	wire [11-1:0] node1083;
	wire [11-1:0] node1084;
	wire [11-1:0] node1085;
	wire [11-1:0] node1088;
	wire [11-1:0] node1091;
	wire [11-1:0] node1094;
	wire [11-1:0] node1095;
	wire [11-1:0] node1096;
	wire [11-1:0] node1099;
	wire [11-1:0] node1102;
	wire [11-1:0] node1103;
	wire [11-1:0] node1106;
	wire [11-1:0] node1109;
	wire [11-1:0] node1110;
	wire [11-1:0] node1111;
	wire [11-1:0] node1112;
	wire [11-1:0] node1115;
	wire [11-1:0] node1118;
	wire [11-1:0] node1119;
	wire [11-1:0] node1122;
	wire [11-1:0] node1125;
	wire [11-1:0] node1126;
	wire [11-1:0] node1127;
	wire [11-1:0] node1130;
	wire [11-1:0] node1133;
	wire [11-1:0] node1134;
	wire [11-1:0] node1138;
	wire [11-1:0] node1139;
	wire [11-1:0] node1140;
	wire [11-1:0] node1141;
	wire [11-1:0] node1142;
	wire [11-1:0] node1145;
	wire [11-1:0] node1148;
	wire [11-1:0] node1150;
	wire [11-1:0] node1153;
	wire [11-1:0] node1154;
	wire [11-1:0] node1155;
	wire [11-1:0] node1158;
	wire [11-1:0] node1161;
	wire [11-1:0] node1162;
	wire [11-1:0] node1165;
	wire [11-1:0] node1168;
	wire [11-1:0] node1169;
	wire [11-1:0] node1170;
	wire [11-1:0] node1171;
	wire [11-1:0] node1174;
	wire [11-1:0] node1177;
	wire [11-1:0] node1178;
	wire [11-1:0] node1181;
	wire [11-1:0] node1184;
	wire [11-1:0] node1185;
	wire [11-1:0] node1186;
	wire [11-1:0] node1189;
	wire [11-1:0] node1192;
	wire [11-1:0] node1195;
	wire [11-1:0] node1196;
	wire [11-1:0] node1197;
	wire [11-1:0] node1198;
	wire [11-1:0] node1199;
	wire [11-1:0] node1202;
	wire [11-1:0] node1205;
	wire [11-1:0] node1206;
	wire [11-1:0] node1207;
	wire [11-1:0] node1210;
	wire [11-1:0] node1213;
	wire [11-1:0] node1214;
	wire [11-1:0] node1217;
	wire [11-1:0] node1220;
	wire [11-1:0] node1221;
	wire [11-1:0] node1222;
	wire [11-1:0] node1224;
	wire [11-1:0] node1227;
	wire [11-1:0] node1228;
	wire [11-1:0] node1231;
	wire [11-1:0] node1234;
	wire [11-1:0] node1235;
	wire [11-1:0] node1237;
	wire [11-1:0] node1240;
	wire [11-1:0] node1242;
	wire [11-1:0] node1245;
	wire [11-1:0] node1246;
	wire [11-1:0] node1247;
	wire [11-1:0] node1248;
	wire [11-1:0] node1249;
	wire [11-1:0] node1253;
	wire [11-1:0] node1254;
	wire [11-1:0] node1257;
	wire [11-1:0] node1260;
	wire [11-1:0] node1261;
	wire [11-1:0] node1262;
	wire [11-1:0] node1265;
	wire [11-1:0] node1268;
	wire [11-1:0] node1269;
	wire [11-1:0] node1273;
	wire [11-1:0] node1274;
	wire [11-1:0] node1275;
	wire [11-1:0] node1276;
	wire [11-1:0] node1279;
	wire [11-1:0] node1282;
	wire [11-1:0] node1284;
	wire [11-1:0] node1287;
	wire [11-1:0] node1288;
	wire [11-1:0] node1289;
	wire [11-1:0] node1292;
	wire [11-1:0] node1295;
	wire [11-1:0] node1296;
	wire [11-1:0] node1300;
	wire [11-1:0] node1301;
	wire [11-1:0] node1302;
	wire [11-1:0] node1303;
	wire [11-1:0] node1304;
	wire [11-1:0] node1305;
	wire [11-1:0] node1306;
	wire [11-1:0] node1307;
	wire [11-1:0] node1311;
	wire [11-1:0] node1312;
	wire [11-1:0] node1315;
	wire [11-1:0] node1318;
	wire [11-1:0] node1319;
	wire [11-1:0] node1320;
	wire [11-1:0] node1323;
	wire [11-1:0] node1326;
	wire [11-1:0] node1328;
	wire [11-1:0] node1331;
	wire [11-1:0] node1332;
	wire [11-1:0] node1333;
	wire [11-1:0] node1334;
	wire [11-1:0] node1337;
	wire [11-1:0] node1340;
	wire [11-1:0] node1341;
	wire [11-1:0] node1344;
	wire [11-1:0] node1347;
	wire [11-1:0] node1348;
	wire [11-1:0] node1349;
	wire [11-1:0] node1353;
	wire [11-1:0] node1354;
	wire [11-1:0] node1357;
	wire [11-1:0] node1360;
	wire [11-1:0] node1361;
	wire [11-1:0] node1362;
	wire [11-1:0] node1363;
	wire [11-1:0] node1364;
	wire [11-1:0] node1368;
	wire [11-1:0] node1369;
	wire [11-1:0] node1373;
	wire [11-1:0] node1374;
	wire [11-1:0] node1375;
	wire [11-1:0] node1378;
	wire [11-1:0] node1381;
	wire [11-1:0] node1384;
	wire [11-1:0] node1385;
	wire [11-1:0] node1386;
	wire [11-1:0] node1387;
	wire [11-1:0] node1390;
	wire [11-1:0] node1393;
	wire [11-1:0] node1394;
	wire [11-1:0] node1397;
	wire [11-1:0] node1400;
	wire [11-1:0] node1401;
	wire [11-1:0] node1402;
	wire [11-1:0] node1405;
	wire [11-1:0] node1408;
	wire [11-1:0] node1409;
	wire [11-1:0] node1412;
	wire [11-1:0] node1415;
	wire [11-1:0] node1416;
	wire [11-1:0] node1417;
	wire [11-1:0] node1418;
	wire [11-1:0] node1419;
	wire [11-1:0] node1420;
	wire [11-1:0] node1423;
	wire [11-1:0] node1426;
	wire [11-1:0] node1427;
	wire [11-1:0] node1430;
	wire [11-1:0] node1433;
	wire [11-1:0] node1434;
	wire [11-1:0] node1435;
	wire [11-1:0] node1438;
	wire [11-1:0] node1441;
	wire [11-1:0] node1442;
	wire [11-1:0] node1445;
	wire [11-1:0] node1448;
	wire [11-1:0] node1449;
	wire [11-1:0] node1450;
	wire [11-1:0] node1453;
	wire [11-1:0] node1454;
	wire [11-1:0] node1457;
	wire [11-1:0] node1460;
	wire [11-1:0] node1461;
	wire [11-1:0] node1462;
	wire [11-1:0] node1465;
	wire [11-1:0] node1468;
	wire [11-1:0] node1469;
	wire [11-1:0] node1473;
	wire [11-1:0] node1474;
	wire [11-1:0] node1475;
	wire [11-1:0] node1476;
	wire [11-1:0] node1478;
	wire [11-1:0] node1481;
	wire [11-1:0] node1482;
	wire [11-1:0] node1485;
	wire [11-1:0] node1488;
	wire [11-1:0] node1489;
	wire [11-1:0] node1490;
	wire [11-1:0] node1493;
	wire [11-1:0] node1496;
	wire [11-1:0] node1497;
	wire [11-1:0] node1500;
	wire [11-1:0] node1503;
	wire [11-1:0] node1504;
	wire [11-1:0] node1505;
	wire [11-1:0] node1506;
	wire [11-1:0] node1510;
	wire [11-1:0] node1511;
	wire [11-1:0] node1514;
	wire [11-1:0] node1517;
	wire [11-1:0] node1518;
	wire [11-1:0] node1519;
	wire [11-1:0] node1522;
	wire [11-1:0] node1525;
	wire [11-1:0] node1526;
	wire [11-1:0] node1530;
	wire [11-1:0] node1531;
	wire [11-1:0] node1532;
	wire [11-1:0] node1533;
	wire [11-1:0] node1534;
	wire [11-1:0] node1535;
	wire [11-1:0] node1536;
	wire [11-1:0] node1539;
	wire [11-1:0] node1542;
	wire [11-1:0] node1543;
	wire [11-1:0] node1546;
	wire [11-1:0] node1549;
	wire [11-1:0] node1550;
	wire [11-1:0] node1551;
	wire [11-1:0] node1555;
	wire [11-1:0] node1556;
	wire [11-1:0] node1559;
	wire [11-1:0] node1562;
	wire [11-1:0] node1563;
	wire [11-1:0] node1564;
	wire [11-1:0] node1565;
	wire [11-1:0] node1568;
	wire [11-1:0] node1571;
	wire [11-1:0] node1572;
	wire [11-1:0] node1576;
	wire [11-1:0] node1577;
	wire [11-1:0] node1579;
	wire [11-1:0] node1582;
	wire [11-1:0] node1583;
	wire [11-1:0] node1586;
	wire [11-1:0] node1589;
	wire [11-1:0] node1590;
	wire [11-1:0] node1591;
	wire [11-1:0] node1592;
	wire [11-1:0] node1593;
	wire [11-1:0] node1597;
	wire [11-1:0] node1598;
	wire [11-1:0] node1602;
	wire [11-1:0] node1603;
	wire [11-1:0] node1604;
	wire [11-1:0] node1607;
	wire [11-1:0] node1610;
	wire [11-1:0] node1611;
	wire [11-1:0] node1614;
	wire [11-1:0] node1617;
	wire [11-1:0] node1618;
	wire [11-1:0] node1619;
	wire [11-1:0] node1621;
	wire [11-1:0] node1624;
	wire [11-1:0] node1627;
	wire [11-1:0] node1628;
	wire [11-1:0] node1629;
	wire [11-1:0] node1632;
	wire [11-1:0] node1635;
	wire [11-1:0] node1636;
	wire [11-1:0] node1640;
	wire [11-1:0] node1641;
	wire [11-1:0] node1642;
	wire [11-1:0] node1643;
	wire [11-1:0] node1644;
	wire [11-1:0] node1647;
	wire [11-1:0] node1648;
	wire [11-1:0] node1651;
	wire [11-1:0] node1654;
	wire [11-1:0] node1655;
	wire [11-1:0] node1656;
	wire [11-1:0] node1659;
	wire [11-1:0] node1662;
	wire [11-1:0] node1663;
	wire [11-1:0] node1666;
	wire [11-1:0] node1669;
	wire [11-1:0] node1670;
	wire [11-1:0] node1671;
	wire [11-1:0] node1672;
	wire [11-1:0] node1675;
	wire [11-1:0] node1678;
	wire [11-1:0] node1679;
	wire [11-1:0] node1682;
	wire [11-1:0] node1685;
	wire [11-1:0] node1686;
	wire [11-1:0] node1687;
	wire [11-1:0] node1690;
	wire [11-1:0] node1693;
	wire [11-1:0] node1695;
	wire [11-1:0] node1698;
	wire [11-1:0] node1699;
	wire [11-1:0] node1700;
	wire [11-1:0] node1701;
	wire [11-1:0] node1702;
	wire [11-1:0] node1705;
	wire [11-1:0] node1708;
	wire [11-1:0] node1711;
	wire [11-1:0] node1712;
	wire [11-1:0] node1713;
	wire [11-1:0] node1716;
	wire [11-1:0] node1719;
	wire [11-1:0] node1720;
	wire [11-1:0] node1723;
	wire [11-1:0] node1726;
	wire [11-1:0] node1727;
	wire [11-1:0] node1728;
	wire [11-1:0] node1729;
	wire [11-1:0] node1732;
	wire [11-1:0] node1735;
	wire [11-1:0] node1736;
	wire [11-1:0] node1739;
	wire [11-1:0] node1742;
	wire [11-1:0] node1743;
	wire [11-1:0] node1744;
	wire [11-1:0] node1748;
	wire [11-1:0] node1751;
	wire [11-1:0] node1752;
	wire [11-1:0] node1753;
	wire [11-1:0] node1754;
	wire [11-1:0] node1755;
	wire [11-1:0] node1756;
	wire [11-1:0] node1757;
	wire [11-1:0] node1758;
	wire [11-1:0] node1759;
	wire [11-1:0] node1760;
	wire [11-1:0] node1763;
	wire [11-1:0] node1766;
	wire [11-1:0] node1767;
	wire [11-1:0] node1770;
	wire [11-1:0] node1773;
	wire [11-1:0] node1774;
	wire [11-1:0] node1775;
	wire [11-1:0] node1778;
	wire [11-1:0] node1781;
	wire [11-1:0] node1782;
	wire [11-1:0] node1785;
	wire [11-1:0] node1788;
	wire [11-1:0] node1789;
	wire [11-1:0] node1790;
	wire [11-1:0] node1792;
	wire [11-1:0] node1795;
	wire [11-1:0] node1796;
	wire [11-1:0] node1800;
	wire [11-1:0] node1801;
	wire [11-1:0] node1802;
	wire [11-1:0] node1805;
	wire [11-1:0] node1808;
	wire [11-1:0] node1809;
	wire [11-1:0] node1812;
	wire [11-1:0] node1815;
	wire [11-1:0] node1816;
	wire [11-1:0] node1817;
	wire [11-1:0] node1818;
	wire [11-1:0] node1819;
	wire [11-1:0] node1823;
	wire [11-1:0] node1826;
	wire [11-1:0] node1827;
	wire [11-1:0] node1828;
	wire [11-1:0] node1831;
	wire [11-1:0] node1834;
	wire [11-1:0] node1837;
	wire [11-1:0] node1838;
	wire [11-1:0] node1839;
	wire [11-1:0] node1840;
	wire [11-1:0] node1843;
	wire [11-1:0] node1846;
	wire [11-1:0] node1848;
	wire [11-1:0] node1851;
	wire [11-1:0] node1852;
	wire [11-1:0] node1853;
	wire [11-1:0] node1856;
	wire [11-1:0] node1859;
	wire [11-1:0] node1860;
	wire [11-1:0] node1863;
	wire [11-1:0] node1866;
	wire [11-1:0] node1867;
	wire [11-1:0] node1868;
	wire [11-1:0] node1869;
	wire [11-1:0] node1870;
	wire [11-1:0] node1871;
	wire [11-1:0] node1874;
	wire [11-1:0] node1877;
	wire [11-1:0] node1878;
	wire [11-1:0] node1881;
	wire [11-1:0] node1884;
	wire [11-1:0] node1885;
	wire [11-1:0] node1886;
	wire [11-1:0] node1889;
	wire [11-1:0] node1892;
	wire [11-1:0] node1894;
	wire [11-1:0] node1897;
	wire [11-1:0] node1898;
	wire [11-1:0] node1899;
	wire [11-1:0] node1900;
	wire [11-1:0] node1903;
	wire [11-1:0] node1906;
	wire [11-1:0] node1907;
	wire [11-1:0] node1910;
	wire [11-1:0] node1913;
	wire [11-1:0] node1914;
	wire [11-1:0] node1915;
	wire [11-1:0] node1918;
	wire [11-1:0] node1921;
	wire [11-1:0] node1924;
	wire [11-1:0] node1925;
	wire [11-1:0] node1926;
	wire [11-1:0] node1927;
	wire [11-1:0] node1929;
	wire [11-1:0] node1932;
	wire [11-1:0] node1933;
	wire [11-1:0] node1937;
	wire [11-1:0] node1938;
	wire [11-1:0] node1939;
	wire [11-1:0] node1942;
	wire [11-1:0] node1945;
	wire [11-1:0] node1946;
	wire [11-1:0] node1949;
	wire [11-1:0] node1952;
	wire [11-1:0] node1953;
	wire [11-1:0] node1954;
	wire [11-1:0] node1955;
	wire [11-1:0] node1958;
	wire [11-1:0] node1961;
	wire [11-1:0] node1962;
	wire [11-1:0] node1965;
	wire [11-1:0] node1968;
	wire [11-1:0] node1969;
	wire [11-1:0] node1971;
	wire [11-1:0] node1974;
	wire [11-1:0] node1975;
	wire [11-1:0] node1978;
	wire [11-1:0] node1981;
	wire [11-1:0] node1982;
	wire [11-1:0] node1983;
	wire [11-1:0] node1984;
	wire [11-1:0] node1985;
	wire [11-1:0] node1986;
	wire [11-1:0] node1987;
	wire [11-1:0] node1990;
	wire [11-1:0] node1993;
	wire [11-1:0] node1995;
	wire [11-1:0] node1998;
	wire [11-1:0] node1999;
	wire [11-1:0] node2000;
	wire [11-1:0] node2003;
	wire [11-1:0] node2006;
	wire [11-1:0] node2007;
	wire [11-1:0] node2010;
	wire [11-1:0] node2013;
	wire [11-1:0] node2014;
	wire [11-1:0] node2015;
	wire [11-1:0] node2016;
	wire [11-1:0] node2020;
	wire [11-1:0] node2023;
	wire [11-1:0] node2024;
	wire [11-1:0] node2025;
	wire [11-1:0] node2028;
	wire [11-1:0] node2031;
	wire [11-1:0] node2032;
	wire [11-1:0] node2035;
	wire [11-1:0] node2038;
	wire [11-1:0] node2039;
	wire [11-1:0] node2040;
	wire [11-1:0] node2041;
	wire [11-1:0] node2043;
	wire [11-1:0] node2046;
	wire [11-1:0] node2047;
	wire [11-1:0] node2050;
	wire [11-1:0] node2053;
	wire [11-1:0] node2054;
	wire [11-1:0] node2055;
	wire [11-1:0] node2058;
	wire [11-1:0] node2061;
	wire [11-1:0] node2062;
	wire [11-1:0] node2065;
	wire [11-1:0] node2068;
	wire [11-1:0] node2069;
	wire [11-1:0] node2070;
	wire [11-1:0] node2071;
	wire [11-1:0] node2074;
	wire [11-1:0] node2077;
	wire [11-1:0] node2078;
	wire [11-1:0] node2081;
	wire [11-1:0] node2084;
	wire [11-1:0] node2085;
	wire [11-1:0] node2088;
	wire [11-1:0] node2090;
	wire [11-1:0] node2093;
	wire [11-1:0] node2094;
	wire [11-1:0] node2095;
	wire [11-1:0] node2096;
	wire [11-1:0] node2097;
	wire [11-1:0] node2098;
	wire [11-1:0] node2101;
	wire [11-1:0] node2104;
	wire [11-1:0] node2105;
	wire [11-1:0] node2108;
	wire [11-1:0] node2111;
	wire [11-1:0] node2112;
	wire [11-1:0] node2113;
	wire [11-1:0] node2116;
	wire [11-1:0] node2119;
	wire [11-1:0] node2120;
	wire [11-1:0] node2123;
	wire [11-1:0] node2126;
	wire [11-1:0] node2127;
	wire [11-1:0] node2128;
	wire [11-1:0] node2131;
	wire [11-1:0] node2132;
	wire [11-1:0] node2135;
	wire [11-1:0] node2138;
	wire [11-1:0] node2140;
	wire [11-1:0] node2141;
	wire [11-1:0] node2144;
	wire [11-1:0] node2147;
	wire [11-1:0] node2148;
	wire [11-1:0] node2149;
	wire [11-1:0] node2150;
	wire [11-1:0] node2151;
	wire [11-1:0] node2154;
	wire [11-1:0] node2157;
	wire [11-1:0] node2158;
	wire [11-1:0] node2161;
	wire [11-1:0] node2164;
	wire [11-1:0] node2165;
	wire [11-1:0] node2166;
	wire [11-1:0] node2170;
	wire [11-1:0] node2171;
	wire [11-1:0] node2174;
	wire [11-1:0] node2177;
	wire [11-1:0] node2178;
	wire [11-1:0] node2179;
	wire [11-1:0] node2180;
	wire [11-1:0] node2184;
	wire [11-1:0] node2187;
	wire [11-1:0] node2188;
	wire [11-1:0] node2189;
	wire [11-1:0] node2193;
	wire [11-1:0] node2194;
	wire [11-1:0] node2197;
	wire [11-1:0] node2200;
	wire [11-1:0] node2201;
	wire [11-1:0] node2202;
	wire [11-1:0] node2203;
	wire [11-1:0] node2204;
	wire [11-1:0] node2205;
	wire [11-1:0] node2206;
	wire [11-1:0] node2207;
	wire [11-1:0] node2211;
	wire [11-1:0] node2213;
	wire [11-1:0] node2216;
	wire [11-1:0] node2217;
	wire [11-1:0] node2218;
	wire [11-1:0] node2222;
	wire [11-1:0] node2223;
	wire [11-1:0] node2227;
	wire [11-1:0] node2228;
	wire [11-1:0] node2229;
	wire [11-1:0] node2230;
	wire [11-1:0] node2233;
	wire [11-1:0] node2236;
	wire [11-1:0] node2237;
	wire [11-1:0] node2240;
	wire [11-1:0] node2243;
	wire [11-1:0] node2244;
	wire [11-1:0] node2246;
	wire [11-1:0] node2249;
	wire [11-1:0] node2251;
	wire [11-1:0] node2254;
	wire [11-1:0] node2255;
	wire [11-1:0] node2256;
	wire [11-1:0] node2257;
	wire [11-1:0] node2258;
	wire [11-1:0] node2262;
	wire [11-1:0] node2264;
	wire [11-1:0] node2267;
	wire [11-1:0] node2268;
	wire [11-1:0] node2269;
	wire [11-1:0] node2272;
	wire [11-1:0] node2275;
	wire [11-1:0] node2277;
	wire [11-1:0] node2280;
	wire [11-1:0] node2281;
	wire [11-1:0] node2282;
	wire [11-1:0] node2283;
	wire [11-1:0] node2286;
	wire [11-1:0] node2289;
	wire [11-1:0] node2291;
	wire [11-1:0] node2294;
	wire [11-1:0] node2295;
	wire [11-1:0] node2296;
	wire [11-1:0] node2300;
	wire [11-1:0] node2301;
	wire [11-1:0] node2305;
	wire [11-1:0] node2306;
	wire [11-1:0] node2307;
	wire [11-1:0] node2308;
	wire [11-1:0] node2309;
	wire [11-1:0] node2310;
	wire [11-1:0] node2313;
	wire [11-1:0] node2316;
	wire [11-1:0] node2317;
	wire [11-1:0] node2320;
	wire [11-1:0] node2323;
	wire [11-1:0] node2324;
	wire [11-1:0] node2325;
	wire [11-1:0] node2328;
	wire [11-1:0] node2331;
	wire [11-1:0] node2332;
	wire [11-1:0] node2335;
	wire [11-1:0] node2338;
	wire [11-1:0] node2339;
	wire [11-1:0] node2340;
	wire [11-1:0] node2341;
	wire [11-1:0] node2344;
	wire [11-1:0] node2347;
	wire [11-1:0] node2349;
	wire [11-1:0] node2352;
	wire [11-1:0] node2353;
	wire [11-1:0] node2354;
	wire [11-1:0] node2358;
	wire [11-1:0] node2359;
	wire [11-1:0] node2362;
	wire [11-1:0] node2365;
	wire [11-1:0] node2366;
	wire [11-1:0] node2367;
	wire [11-1:0] node2368;
	wire [11-1:0] node2369;
	wire [11-1:0] node2372;
	wire [11-1:0] node2375;
	wire [11-1:0] node2376;
	wire [11-1:0] node2379;
	wire [11-1:0] node2382;
	wire [11-1:0] node2383;
	wire [11-1:0] node2384;
	wire [11-1:0] node2387;
	wire [11-1:0] node2390;
	wire [11-1:0] node2391;
	wire [11-1:0] node2394;
	wire [11-1:0] node2397;
	wire [11-1:0] node2398;
	wire [11-1:0] node2399;
	wire [11-1:0] node2400;
	wire [11-1:0] node2403;
	wire [11-1:0] node2406;
	wire [11-1:0] node2407;
	wire [11-1:0] node2411;
	wire [11-1:0] node2412;
	wire [11-1:0] node2413;
	wire [11-1:0] node2416;
	wire [11-1:0] node2419;
	wire [11-1:0] node2421;
	wire [11-1:0] node2424;
	wire [11-1:0] node2425;
	wire [11-1:0] node2426;
	wire [11-1:0] node2427;
	wire [11-1:0] node2428;
	wire [11-1:0] node2429;
	wire [11-1:0] node2430;
	wire [11-1:0] node2433;
	wire [11-1:0] node2436;
	wire [11-1:0] node2437;
	wire [11-1:0] node2441;
	wire [11-1:0] node2442;
	wire [11-1:0] node2444;
	wire [11-1:0] node2447;
	wire [11-1:0] node2450;
	wire [11-1:0] node2451;
	wire [11-1:0] node2452;
	wire [11-1:0] node2454;
	wire [11-1:0] node2457;
	wire [11-1:0] node2458;
	wire [11-1:0] node2461;
	wire [11-1:0] node2464;
	wire [11-1:0] node2465;
	wire [11-1:0] node2468;
	wire [11-1:0] node2469;
	wire [11-1:0] node2473;
	wire [11-1:0] node2474;
	wire [11-1:0] node2475;
	wire [11-1:0] node2476;
	wire [11-1:0] node2477;
	wire [11-1:0] node2480;
	wire [11-1:0] node2483;
	wire [11-1:0] node2484;
	wire [11-1:0] node2487;
	wire [11-1:0] node2490;
	wire [11-1:0] node2491;
	wire [11-1:0] node2493;
	wire [11-1:0] node2496;
	wire [11-1:0] node2497;
	wire [11-1:0] node2500;
	wire [11-1:0] node2503;
	wire [11-1:0] node2504;
	wire [11-1:0] node2505;
	wire [11-1:0] node2506;
	wire [11-1:0] node2509;
	wire [11-1:0] node2512;
	wire [11-1:0] node2514;
	wire [11-1:0] node2517;
	wire [11-1:0] node2518;
	wire [11-1:0] node2519;
	wire [11-1:0] node2522;
	wire [11-1:0] node2525;
	wire [11-1:0] node2527;
	wire [11-1:0] node2530;
	wire [11-1:0] node2531;
	wire [11-1:0] node2532;
	wire [11-1:0] node2533;
	wire [11-1:0] node2534;
	wire [11-1:0] node2536;
	wire [11-1:0] node2539;
	wire [11-1:0] node2540;
	wire [11-1:0] node2544;
	wire [11-1:0] node2545;
	wire [11-1:0] node2546;
	wire [11-1:0] node2549;
	wire [11-1:0] node2552;
	wire [11-1:0] node2553;
	wire [11-1:0] node2556;
	wire [11-1:0] node2559;
	wire [11-1:0] node2560;
	wire [11-1:0] node2561;
	wire [11-1:0] node2562;
	wire [11-1:0] node2565;
	wire [11-1:0] node2568;
	wire [11-1:0] node2570;
	wire [11-1:0] node2573;
	wire [11-1:0] node2574;
	wire [11-1:0] node2575;
	wire [11-1:0] node2578;
	wire [11-1:0] node2581;
	wire [11-1:0] node2582;
	wire [11-1:0] node2586;
	wire [11-1:0] node2587;
	wire [11-1:0] node2588;
	wire [11-1:0] node2589;
	wire [11-1:0] node2591;
	wire [11-1:0] node2594;
	wire [11-1:0] node2595;
	wire [11-1:0] node2598;
	wire [11-1:0] node2601;
	wire [11-1:0] node2602;
	wire [11-1:0] node2603;
	wire [11-1:0] node2606;
	wire [11-1:0] node2609;
	wire [11-1:0] node2610;
	wire [11-1:0] node2613;
	wire [11-1:0] node2616;
	wire [11-1:0] node2617;
	wire [11-1:0] node2618;
	wire [11-1:0] node2619;
	wire [11-1:0] node2622;
	wire [11-1:0] node2625;
	wire [11-1:0] node2628;
	wire [11-1:0] node2629;
	wire [11-1:0] node2630;
	wire [11-1:0] node2633;
	wire [11-1:0] node2636;
	wire [11-1:0] node2637;
	wire [11-1:0] node2641;
	wire [11-1:0] node2642;
	wire [11-1:0] node2643;
	wire [11-1:0] node2644;
	wire [11-1:0] node2645;
	wire [11-1:0] node2646;
	wire [11-1:0] node2647;
	wire [11-1:0] node2648;
	wire [11-1:0] node2651;
	wire [11-1:0] node2652;
	wire [11-1:0] node2655;
	wire [11-1:0] node2658;
	wire [11-1:0] node2659;
	wire [11-1:0] node2660;
	wire [11-1:0] node2663;
	wire [11-1:0] node2666;
	wire [11-1:0] node2667;
	wire [11-1:0] node2670;
	wire [11-1:0] node2673;
	wire [11-1:0] node2674;
	wire [11-1:0] node2675;
	wire [11-1:0] node2676;
	wire [11-1:0] node2679;
	wire [11-1:0] node2682;
	wire [11-1:0] node2683;
	wire [11-1:0] node2687;
	wire [11-1:0] node2688;
	wire [11-1:0] node2690;
	wire [11-1:0] node2693;
	wire [11-1:0] node2694;
	wire [11-1:0] node2697;
	wire [11-1:0] node2700;
	wire [11-1:0] node2701;
	wire [11-1:0] node2702;
	wire [11-1:0] node2703;
	wire [11-1:0] node2706;
	wire [11-1:0] node2707;
	wire [11-1:0] node2710;
	wire [11-1:0] node2713;
	wire [11-1:0] node2714;
	wire [11-1:0] node2715;
	wire [11-1:0] node2719;
	wire [11-1:0] node2721;
	wire [11-1:0] node2724;
	wire [11-1:0] node2725;
	wire [11-1:0] node2726;
	wire [11-1:0] node2727;
	wire [11-1:0] node2730;
	wire [11-1:0] node2733;
	wire [11-1:0] node2734;
	wire [11-1:0] node2738;
	wire [11-1:0] node2739;
	wire [11-1:0] node2740;
	wire [11-1:0] node2743;
	wire [11-1:0] node2746;
	wire [11-1:0] node2747;
	wire [11-1:0] node2750;
	wire [11-1:0] node2753;
	wire [11-1:0] node2754;
	wire [11-1:0] node2755;
	wire [11-1:0] node2756;
	wire [11-1:0] node2757;
	wire [11-1:0] node2758;
	wire [11-1:0] node2762;
	wire [11-1:0] node2763;
	wire [11-1:0] node2766;
	wire [11-1:0] node2769;
	wire [11-1:0] node2770;
	wire [11-1:0] node2771;
	wire [11-1:0] node2774;
	wire [11-1:0] node2777;
	wire [11-1:0] node2778;
	wire [11-1:0] node2782;
	wire [11-1:0] node2783;
	wire [11-1:0] node2784;
	wire [11-1:0] node2785;
	wire [11-1:0] node2788;
	wire [11-1:0] node2791;
	wire [11-1:0] node2792;
	wire [11-1:0] node2795;
	wire [11-1:0] node2798;
	wire [11-1:0] node2799;
	wire [11-1:0] node2800;
	wire [11-1:0] node2803;
	wire [11-1:0] node2806;
	wire [11-1:0] node2807;
	wire [11-1:0] node2811;
	wire [11-1:0] node2812;
	wire [11-1:0] node2813;
	wire [11-1:0] node2814;
	wire [11-1:0] node2817;
	wire [11-1:0] node2818;
	wire [11-1:0] node2821;
	wire [11-1:0] node2824;
	wire [11-1:0] node2825;
	wire [11-1:0] node2827;
	wire [11-1:0] node2830;
	wire [11-1:0] node2831;
	wire [11-1:0] node2834;
	wire [11-1:0] node2837;
	wire [11-1:0] node2838;
	wire [11-1:0] node2839;
	wire [11-1:0] node2840;
	wire [11-1:0] node2843;
	wire [11-1:0] node2846;
	wire [11-1:0] node2847;
	wire [11-1:0] node2850;
	wire [11-1:0] node2853;
	wire [11-1:0] node2854;
	wire [11-1:0] node2856;
	wire [11-1:0] node2859;
	wire [11-1:0] node2860;
	wire [11-1:0] node2863;
	wire [11-1:0] node2866;
	wire [11-1:0] node2867;
	wire [11-1:0] node2868;
	wire [11-1:0] node2869;
	wire [11-1:0] node2870;
	wire [11-1:0] node2871;
	wire [11-1:0] node2872;
	wire [11-1:0] node2875;
	wire [11-1:0] node2878;
	wire [11-1:0] node2879;
	wire [11-1:0] node2882;
	wire [11-1:0] node2885;
	wire [11-1:0] node2886;
	wire [11-1:0] node2887;
	wire [11-1:0] node2890;
	wire [11-1:0] node2893;
	wire [11-1:0] node2896;
	wire [11-1:0] node2897;
	wire [11-1:0] node2898;
	wire [11-1:0] node2899;
	wire [11-1:0] node2902;
	wire [11-1:0] node2905;
	wire [11-1:0] node2908;
	wire [11-1:0] node2909;
	wire [11-1:0] node2910;
	wire [11-1:0] node2913;
	wire [11-1:0] node2916;
	wire [11-1:0] node2917;
	wire [11-1:0] node2921;
	wire [11-1:0] node2922;
	wire [11-1:0] node2923;
	wire [11-1:0] node2924;
	wire [11-1:0] node2925;
	wire [11-1:0] node2928;
	wire [11-1:0] node2931;
	wire [11-1:0] node2932;
	wire [11-1:0] node2936;
	wire [11-1:0] node2937;
	wire [11-1:0] node2938;
	wire [11-1:0] node2942;
	wire [11-1:0] node2943;
	wire [11-1:0] node2946;
	wire [11-1:0] node2949;
	wire [11-1:0] node2950;
	wire [11-1:0] node2951;
	wire [11-1:0] node2952;
	wire [11-1:0] node2955;
	wire [11-1:0] node2958;
	wire [11-1:0] node2960;
	wire [11-1:0] node2963;
	wire [11-1:0] node2964;
	wire [11-1:0] node2965;
	wire [11-1:0] node2968;
	wire [11-1:0] node2971;
	wire [11-1:0] node2972;
	wire [11-1:0] node2975;
	wire [11-1:0] node2978;
	wire [11-1:0] node2979;
	wire [11-1:0] node2980;
	wire [11-1:0] node2981;
	wire [11-1:0] node2982;
	wire [11-1:0] node2984;
	wire [11-1:0] node2987;
	wire [11-1:0] node2989;
	wire [11-1:0] node2992;
	wire [11-1:0] node2993;
	wire [11-1:0] node2994;
	wire [11-1:0] node2997;
	wire [11-1:0] node3000;
	wire [11-1:0] node3001;
	wire [11-1:0] node3004;
	wire [11-1:0] node3007;
	wire [11-1:0] node3008;
	wire [11-1:0] node3009;
	wire [11-1:0] node3010;
	wire [11-1:0] node3013;
	wire [11-1:0] node3016;
	wire [11-1:0] node3017;
	wire [11-1:0] node3021;
	wire [11-1:0] node3022;
	wire [11-1:0] node3023;
	wire [11-1:0] node3026;
	wire [11-1:0] node3029;
	wire [11-1:0] node3030;
	wire [11-1:0] node3034;
	wire [11-1:0] node3035;
	wire [11-1:0] node3036;
	wire [11-1:0] node3037;
	wire [11-1:0] node3038;
	wire [11-1:0] node3042;
	wire [11-1:0] node3043;
	wire [11-1:0] node3046;
	wire [11-1:0] node3049;
	wire [11-1:0] node3050;
	wire [11-1:0] node3052;
	wire [11-1:0] node3055;
	wire [11-1:0] node3056;
	wire [11-1:0] node3059;
	wire [11-1:0] node3062;
	wire [11-1:0] node3063;
	wire [11-1:0] node3064;
	wire [11-1:0] node3065;
	wire [11-1:0] node3069;
	wire [11-1:0] node3071;
	wire [11-1:0] node3074;
	wire [11-1:0] node3075;
	wire [11-1:0] node3076;
	wire [11-1:0] node3079;
	wire [11-1:0] node3082;
	wire [11-1:0] node3083;
	wire [11-1:0] node3087;
	wire [11-1:0] node3088;
	wire [11-1:0] node3089;
	wire [11-1:0] node3090;
	wire [11-1:0] node3091;
	wire [11-1:0] node3092;
	wire [11-1:0] node3093;
	wire [11-1:0] node3094;
	wire [11-1:0] node3098;
	wire [11-1:0] node3099;
	wire [11-1:0] node3102;
	wire [11-1:0] node3105;
	wire [11-1:0] node3106;
	wire [11-1:0] node3108;
	wire [11-1:0] node3111;
	wire [11-1:0] node3113;
	wire [11-1:0] node3116;
	wire [11-1:0] node3117;
	wire [11-1:0] node3118;
	wire [11-1:0] node3119;
	wire [11-1:0] node3122;
	wire [11-1:0] node3125;
	wire [11-1:0] node3126;
	wire [11-1:0] node3129;
	wire [11-1:0] node3132;
	wire [11-1:0] node3133;
	wire [11-1:0] node3136;
	wire [11-1:0] node3137;
	wire [11-1:0] node3140;
	wire [11-1:0] node3143;
	wire [11-1:0] node3144;
	wire [11-1:0] node3145;
	wire [11-1:0] node3146;
	wire [11-1:0] node3147;
	wire [11-1:0] node3150;
	wire [11-1:0] node3153;
	wire [11-1:0] node3154;
	wire [11-1:0] node3157;
	wire [11-1:0] node3160;
	wire [11-1:0] node3161;
	wire [11-1:0] node3162;
	wire [11-1:0] node3165;
	wire [11-1:0] node3168;
	wire [11-1:0] node3169;
	wire [11-1:0] node3172;
	wire [11-1:0] node3175;
	wire [11-1:0] node3176;
	wire [11-1:0] node3177;
	wire [11-1:0] node3178;
	wire [11-1:0] node3181;
	wire [11-1:0] node3184;
	wire [11-1:0] node3186;
	wire [11-1:0] node3189;
	wire [11-1:0] node3190;
	wire [11-1:0] node3191;
	wire [11-1:0] node3194;
	wire [11-1:0] node3197;
	wire [11-1:0] node3198;
	wire [11-1:0] node3201;
	wire [11-1:0] node3204;
	wire [11-1:0] node3205;
	wire [11-1:0] node3206;
	wire [11-1:0] node3207;
	wire [11-1:0] node3208;
	wire [11-1:0] node3209;
	wire [11-1:0] node3212;
	wire [11-1:0] node3215;
	wire [11-1:0] node3216;
	wire [11-1:0] node3219;
	wire [11-1:0] node3222;
	wire [11-1:0] node3223;
	wire [11-1:0] node3225;
	wire [11-1:0] node3228;
	wire [11-1:0] node3229;
	wire [11-1:0] node3232;
	wire [11-1:0] node3235;
	wire [11-1:0] node3236;
	wire [11-1:0] node3237;
	wire [11-1:0] node3239;
	wire [11-1:0] node3242;
	wire [11-1:0] node3243;
	wire [11-1:0] node3246;
	wire [11-1:0] node3249;
	wire [11-1:0] node3250;
	wire [11-1:0] node3252;
	wire [11-1:0] node3255;
	wire [11-1:0] node3256;
	wire [11-1:0] node3259;
	wire [11-1:0] node3262;
	wire [11-1:0] node3263;
	wire [11-1:0] node3264;
	wire [11-1:0] node3265;
	wire [11-1:0] node3266;
	wire [11-1:0] node3270;
	wire [11-1:0] node3272;
	wire [11-1:0] node3275;
	wire [11-1:0] node3276;
	wire [11-1:0] node3277;
	wire [11-1:0] node3281;
	wire [11-1:0] node3283;
	wire [11-1:0] node3286;
	wire [11-1:0] node3287;
	wire [11-1:0] node3288;
	wire [11-1:0] node3289;
	wire [11-1:0] node3292;
	wire [11-1:0] node3295;
	wire [11-1:0] node3296;
	wire [11-1:0] node3299;
	wire [11-1:0] node3302;
	wire [11-1:0] node3303;
	wire [11-1:0] node3305;
	wire [11-1:0] node3308;
	wire [11-1:0] node3309;
	wire [11-1:0] node3312;
	wire [11-1:0] node3315;
	wire [11-1:0] node3316;
	wire [11-1:0] node3317;
	wire [11-1:0] node3318;
	wire [11-1:0] node3319;
	wire [11-1:0] node3320;
	wire [11-1:0] node3321;
	wire [11-1:0] node3324;
	wire [11-1:0] node3327;
	wire [11-1:0] node3329;
	wire [11-1:0] node3332;
	wire [11-1:0] node3333;
	wire [11-1:0] node3336;
	wire [11-1:0] node3338;
	wire [11-1:0] node3341;
	wire [11-1:0] node3342;
	wire [11-1:0] node3343;
	wire [11-1:0] node3344;
	wire [11-1:0] node3347;
	wire [11-1:0] node3350;
	wire [11-1:0] node3352;
	wire [11-1:0] node3355;
	wire [11-1:0] node3356;
	wire [11-1:0] node3357;
	wire [11-1:0] node3360;
	wire [11-1:0] node3363;
	wire [11-1:0] node3366;
	wire [11-1:0] node3367;
	wire [11-1:0] node3368;
	wire [11-1:0] node3369;
	wire [11-1:0] node3370;
	wire [11-1:0] node3373;
	wire [11-1:0] node3376;
	wire [11-1:0] node3377;
	wire [11-1:0] node3381;
	wire [11-1:0] node3382;
	wire [11-1:0] node3383;
	wire [11-1:0] node3386;
	wire [11-1:0] node3389;
	wire [11-1:0] node3390;
	wire [11-1:0] node3393;
	wire [11-1:0] node3396;
	wire [11-1:0] node3397;
	wire [11-1:0] node3398;
	wire [11-1:0] node3399;
	wire [11-1:0] node3403;
	wire [11-1:0] node3404;
	wire [11-1:0] node3407;
	wire [11-1:0] node3410;
	wire [11-1:0] node3411;
	wire [11-1:0] node3414;
	wire [11-1:0] node3417;
	wire [11-1:0] node3418;
	wire [11-1:0] node3419;
	wire [11-1:0] node3420;
	wire [11-1:0] node3421;
	wire [11-1:0] node3424;
	wire [11-1:0] node3426;
	wire [11-1:0] node3429;
	wire [11-1:0] node3430;
	wire [11-1:0] node3432;
	wire [11-1:0] node3435;
	wire [11-1:0] node3437;
	wire [11-1:0] node3440;
	wire [11-1:0] node3441;
	wire [11-1:0] node3442;
	wire [11-1:0] node3443;
	wire [11-1:0] node3446;
	wire [11-1:0] node3449;
	wire [11-1:0] node3451;
	wire [11-1:0] node3454;
	wire [11-1:0] node3455;
	wire [11-1:0] node3456;
	wire [11-1:0] node3460;
	wire [11-1:0] node3461;
	wire [11-1:0] node3465;
	wire [11-1:0] node3466;
	wire [11-1:0] node3467;
	wire [11-1:0] node3468;
	wire [11-1:0] node3470;
	wire [11-1:0] node3473;
	wire [11-1:0] node3474;
	wire [11-1:0] node3478;
	wire [11-1:0] node3479;
	wire [11-1:0] node3480;
	wire [11-1:0] node3483;
	wire [11-1:0] node3486;
	wire [11-1:0] node3487;
	wire [11-1:0] node3490;
	wire [11-1:0] node3493;
	wire [11-1:0] node3494;
	wire [11-1:0] node3495;
	wire [11-1:0] node3496;
	wire [11-1:0] node3501;
	wire [11-1:0] node3502;
	wire [11-1:0] node3503;
	wire [11-1:0] node3506;
	wire [11-1:0] node3509;
	wire [11-1:0] node3510;
	wire [11-1:0] node3514;
	wire [11-1:0] node3515;
	wire [11-1:0] node3516;
	wire [11-1:0] node3517;
	wire [11-1:0] node3518;
	wire [11-1:0] node3519;
	wire [11-1:0] node3520;
	wire [11-1:0] node3521;
	wire [11-1:0] node3522;
	wire [11-1:0] node3523;
	wire [11-1:0] node3524;
	wire [11-1:0] node3527;
	wire [11-1:0] node3530;
	wire [11-1:0] node3531;
	wire [11-1:0] node3534;
	wire [11-1:0] node3537;
	wire [11-1:0] node3538;
	wire [11-1:0] node3541;
	wire [11-1:0] node3542;
	wire [11-1:0] node3545;
	wire [11-1:0] node3548;
	wire [11-1:0] node3549;
	wire [11-1:0] node3550;
	wire [11-1:0] node3551;
	wire [11-1:0] node3554;
	wire [11-1:0] node3557;
	wire [11-1:0] node3559;
	wire [11-1:0] node3562;
	wire [11-1:0] node3563;
	wire [11-1:0] node3564;
	wire [11-1:0] node3568;
	wire [11-1:0] node3569;
	wire [11-1:0] node3572;
	wire [11-1:0] node3575;
	wire [11-1:0] node3576;
	wire [11-1:0] node3577;
	wire [11-1:0] node3578;
	wire [11-1:0] node3579;
	wire [11-1:0] node3582;
	wire [11-1:0] node3585;
	wire [11-1:0] node3586;
	wire [11-1:0] node3589;
	wire [11-1:0] node3592;
	wire [11-1:0] node3593;
	wire [11-1:0] node3594;
	wire [11-1:0] node3597;
	wire [11-1:0] node3600;
	wire [11-1:0] node3601;
	wire [11-1:0] node3604;
	wire [11-1:0] node3607;
	wire [11-1:0] node3608;
	wire [11-1:0] node3609;
	wire [11-1:0] node3611;
	wire [11-1:0] node3614;
	wire [11-1:0] node3616;
	wire [11-1:0] node3619;
	wire [11-1:0] node3620;
	wire [11-1:0] node3621;
	wire [11-1:0] node3625;
	wire [11-1:0] node3626;
	wire [11-1:0] node3629;
	wire [11-1:0] node3632;
	wire [11-1:0] node3633;
	wire [11-1:0] node3634;
	wire [11-1:0] node3635;
	wire [11-1:0] node3636;
	wire [11-1:0] node3638;
	wire [11-1:0] node3641;
	wire [11-1:0] node3643;
	wire [11-1:0] node3646;
	wire [11-1:0] node3647;
	wire [11-1:0] node3648;
	wire [11-1:0] node3651;
	wire [11-1:0] node3654;
	wire [11-1:0] node3656;
	wire [11-1:0] node3659;
	wire [11-1:0] node3660;
	wire [11-1:0] node3661;
	wire [11-1:0] node3662;
	wire [11-1:0] node3665;
	wire [11-1:0] node3668;
	wire [11-1:0] node3670;
	wire [11-1:0] node3673;
	wire [11-1:0] node3674;
	wire [11-1:0] node3676;
	wire [11-1:0] node3679;
	wire [11-1:0] node3680;
	wire [11-1:0] node3683;
	wire [11-1:0] node3686;
	wire [11-1:0] node3687;
	wire [11-1:0] node3688;
	wire [11-1:0] node3689;
	wire [11-1:0] node3690;
	wire [11-1:0] node3694;
	wire [11-1:0] node3695;
	wire [11-1:0] node3698;
	wire [11-1:0] node3701;
	wire [11-1:0] node3702;
	wire [11-1:0] node3703;
	wire [11-1:0] node3706;
	wire [11-1:0] node3709;
	wire [11-1:0] node3710;
	wire [11-1:0] node3713;
	wire [11-1:0] node3716;
	wire [11-1:0] node3717;
	wire [11-1:0] node3718;
	wire [11-1:0] node3719;
	wire [11-1:0] node3722;
	wire [11-1:0] node3725;
	wire [11-1:0] node3726;
	wire [11-1:0] node3729;
	wire [11-1:0] node3732;
	wire [11-1:0] node3733;
	wire [11-1:0] node3736;
	wire [11-1:0] node3739;
	wire [11-1:0] node3740;
	wire [11-1:0] node3741;
	wire [11-1:0] node3742;
	wire [11-1:0] node3743;
	wire [11-1:0] node3744;
	wire [11-1:0] node3746;
	wire [11-1:0] node3749;
	wire [11-1:0] node3750;
	wire [11-1:0] node3753;
	wire [11-1:0] node3756;
	wire [11-1:0] node3757;
	wire [11-1:0] node3758;
	wire [11-1:0] node3761;
	wire [11-1:0] node3764;
	wire [11-1:0] node3765;
	wire [11-1:0] node3768;
	wire [11-1:0] node3771;
	wire [11-1:0] node3772;
	wire [11-1:0] node3773;
	wire [11-1:0] node3774;
	wire [11-1:0] node3777;
	wire [11-1:0] node3780;
	wire [11-1:0] node3781;
	wire [11-1:0] node3784;
	wire [11-1:0] node3787;
	wire [11-1:0] node3788;
	wire [11-1:0] node3789;
	wire [11-1:0] node3792;
	wire [11-1:0] node3795;
	wire [11-1:0] node3796;
	wire [11-1:0] node3799;
	wire [11-1:0] node3802;
	wire [11-1:0] node3803;
	wire [11-1:0] node3804;
	wire [11-1:0] node3805;
	wire [11-1:0] node3808;
	wire [11-1:0] node3809;
	wire [11-1:0] node3812;
	wire [11-1:0] node3815;
	wire [11-1:0] node3816;
	wire [11-1:0] node3817;
	wire [11-1:0] node3820;
	wire [11-1:0] node3823;
	wire [11-1:0] node3824;
	wire [11-1:0] node3827;
	wire [11-1:0] node3830;
	wire [11-1:0] node3831;
	wire [11-1:0] node3832;
	wire [11-1:0] node3833;
	wire [11-1:0] node3836;
	wire [11-1:0] node3839;
	wire [11-1:0] node3840;
	wire [11-1:0] node3843;
	wire [11-1:0] node3846;
	wire [11-1:0] node3847;
	wire [11-1:0] node3848;
	wire [11-1:0] node3851;
	wire [11-1:0] node3854;
	wire [11-1:0] node3856;
	wire [11-1:0] node3859;
	wire [11-1:0] node3860;
	wire [11-1:0] node3861;
	wire [11-1:0] node3862;
	wire [11-1:0] node3863;
	wire [11-1:0] node3866;
	wire [11-1:0] node3867;
	wire [11-1:0] node3870;
	wire [11-1:0] node3873;
	wire [11-1:0] node3874;
	wire [11-1:0] node3875;
	wire [11-1:0] node3879;
	wire [11-1:0] node3882;
	wire [11-1:0] node3883;
	wire [11-1:0] node3884;
	wire [11-1:0] node3885;
	wire [11-1:0] node3888;
	wire [11-1:0] node3891;
	wire [11-1:0] node3892;
	wire [11-1:0] node3895;
	wire [11-1:0] node3898;
	wire [11-1:0] node3899;
	wire [11-1:0] node3900;
	wire [11-1:0] node3903;
	wire [11-1:0] node3906;
	wire [11-1:0] node3907;
	wire [11-1:0] node3910;
	wire [11-1:0] node3913;
	wire [11-1:0] node3914;
	wire [11-1:0] node3915;
	wire [11-1:0] node3916;
	wire [11-1:0] node3919;
	wire [11-1:0] node3921;
	wire [11-1:0] node3924;
	wire [11-1:0] node3925;
	wire [11-1:0] node3928;
	wire [11-1:0] node3929;
	wire [11-1:0] node3933;
	wire [11-1:0] node3934;
	wire [11-1:0] node3935;
	wire [11-1:0] node3936;
	wire [11-1:0] node3939;
	wire [11-1:0] node3942;
	wire [11-1:0] node3943;
	wire [11-1:0] node3946;
	wire [11-1:0] node3949;
	wire [11-1:0] node3950;
	wire [11-1:0] node3953;
	wire [11-1:0] node3956;
	wire [11-1:0] node3957;
	wire [11-1:0] node3958;
	wire [11-1:0] node3959;
	wire [11-1:0] node3960;
	wire [11-1:0] node3961;
	wire [11-1:0] node3962;
	wire [11-1:0] node3963;
	wire [11-1:0] node3966;
	wire [11-1:0] node3969;
	wire [11-1:0] node3970;
	wire [11-1:0] node3973;
	wire [11-1:0] node3976;
	wire [11-1:0] node3977;
	wire [11-1:0] node3978;
	wire [11-1:0] node3981;
	wire [11-1:0] node3985;
	wire [11-1:0] node3986;
	wire [11-1:0] node3987;
	wire [11-1:0] node3988;
	wire [11-1:0] node3991;
	wire [11-1:0] node3994;
	wire [11-1:0] node3995;
	wire [11-1:0] node3998;
	wire [11-1:0] node4001;
	wire [11-1:0] node4002;
	wire [11-1:0] node4003;
	wire [11-1:0] node4007;
	wire [11-1:0] node4008;
	wire [11-1:0] node4011;
	wire [11-1:0] node4014;
	wire [11-1:0] node4015;
	wire [11-1:0] node4016;
	wire [11-1:0] node4017;
	wire [11-1:0] node4018;
	wire [11-1:0] node4021;
	wire [11-1:0] node4024;
	wire [11-1:0] node4025;
	wire [11-1:0] node4029;
	wire [11-1:0] node4030;
	wire [11-1:0] node4033;
	wire [11-1:0] node4034;
	wire [11-1:0] node4037;
	wire [11-1:0] node4040;
	wire [11-1:0] node4041;
	wire [11-1:0] node4042;
	wire [11-1:0] node4043;
	wire [11-1:0] node4046;
	wire [11-1:0] node4049;
	wire [11-1:0] node4050;
	wire [11-1:0] node4053;
	wire [11-1:0] node4056;
	wire [11-1:0] node4057;
	wire [11-1:0] node4059;
	wire [11-1:0] node4062;
	wire [11-1:0] node4063;
	wire [11-1:0] node4066;
	wire [11-1:0] node4069;
	wire [11-1:0] node4070;
	wire [11-1:0] node4071;
	wire [11-1:0] node4072;
	wire [11-1:0] node4073;
	wire [11-1:0] node4074;
	wire [11-1:0] node4078;
	wire [11-1:0] node4079;
	wire [11-1:0] node4083;
	wire [11-1:0] node4084;
	wire [11-1:0] node4085;
	wire [11-1:0] node4088;
	wire [11-1:0] node4091;
	wire [11-1:0] node4094;
	wire [11-1:0] node4095;
	wire [11-1:0] node4096;
	wire [11-1:0] node4097;
	wire [11-1:0] node4100;
	wire [11-1:0] node4103;
	wire [11-1:0] node4104;
	wire [11-1:0] node4108;
	wire [11-1:0] node4109;
	wire [11-1:0] node4110;
	wire [11-1:0] node4113;
	wire [11-1:0] node4116;
	wire [11-1:0] node4117;
	wire [11-1:0] node4120;
	wire [11-1:0] node4123;
	wire [11-1:0] node4124;
	wire [11-1:0] node4125;
	wire [11-1:0] node4126;
	wire [11-1:0] node4127;
	wire [11-1:0] node4131;
	wire [11-1:0] node4132;
	wire [11-1:0] node4135;
	wire [11-1:0] node4138;
	wire [11-1:0] node4139;
	wire [11-1:0] node4142;
	wire [11-1:0] node4143;
	wire [11-1:0] node4146;
	wire [11-1:0] node4149;
	wire [11-1:0] node4150;
	wire [11-1:0] node4151;
	wire [11-1:0] node4152;
	wire [11-1:0] node4155;
	wire [11-1:0] node4158;
	wire [11-1:0] node4159;
	wire [11-1:0] node4163;
	wire [11-1:0] node4164;
	wire [11-1:0] node4165;
	wire [11-1:0] node4168;
	wire [11-1:0] node4171;
	wire [11-1:0] node4172;
	wire [11-1:0] node4175;
	wire [11-1:0] node4178;
	wire [11-1:0] node4179;
	wire [11-1:0] node4180;
	wire [11-1:0] node4181;
	wire [11-1:0] node4182;
	wire [11-1:0] node4183;
	wire [11-1:0] node4184;
	wire [11-1:0] node4187;
	wire [11-1:0] node4190;
	wire [11-1:0] node4191;
	wire [11-1:0] node4194;
	wire [11-1:0] node4197;
	wire [11-1:0] node4198;
	wire [11-1:0] node4199;
	wire [11-1:0] node4202;
	wire [11-1:0] node4205;
	wire [11-1:0] node4206;
	wire [11-1:0] node4210;
	wire [11-1:0] node4211;
	wire [11-1:0] node4212;
	wire [11-1:0] node4213;
	wire [11-1:0] node4216;
	wire [11-1:0] node4219;
	wire [11-1:0] node4222;
	wire [11-1:0] node4223;
	wire [11-1:0] node4224;
	wire [11-1:0] node4227;
	wire [11-1:0] node4230;
	wire [11-1:0] node4231;
	wire [11-1:0] node4234;
	wire [11-1:0] node4237;
	wire [11-1:0] node4238;
	wire [11-1:0] node4239;
	wire [11-1:0] node4240;
	wire [11-1:0] node4242;
	wire [11-1:0] node4245;
	wire [11-1:0] node4246;
	wire [11-1:0] node4249;
	wire [11-1:0] node4252;
	wire [11-1:0] node4253;
	wire [11-1:0] node4254;
	wire [11-1:0] node4257;
	wire [11-1:0] node4260;
	wire [11-1:0] node4263;
	wire [11-1:0] node4264;
	wire [11-1:0] node4265;
	wire [11-1:0] node4266;
	wire [11-1:0] node4269;
	wire [11-1:0] node4272;
	wire [11-1:0] node4273;
	wire [11-1:0] node4277;
	wire [11-1:0] node4278;
	wire [11-1:0] node4279;
	wire [11-1:0] node4282;
	wire [11-1:0] node4285;
	wire [11-1:0] node4286;
	wire [11-1:0] node4290;
	wire [11-1:0] node4291;
	wire [11-1:0] node4292;
	wire [11-1:0] node4293;
	wire [11-1:0] node4294;
	wire [11-1:0] node4295;
	wire [11-1:0] node4299;
	wire [11-1:0] node4300;
	wire [11-1:0] node4304;
	wire [11-1:0] node4305;
	wire [11-1:0] node4306;
	wire [11-1:0] node4309;
	wire [11-1:0] node4312;
	wire [11-1:0] node4313;
	wire [11-1:0] node4316;
	wire [11-1:0] node4319;
	wire [11-1:0] node4320;
	wire [11-1:0] node4321;
	wire [11-1:0] node4322;
	wire [11-1:0] node4325;
	wire [11-1:0] node4328;
	wire [11-1:0] node4329;
	wire [11-1:0] node4332;
	wire [11-1:0] node4335;
	wire [11-1:0] node4336;
	wire [11-1:0] node4337;
	wire [11-1:0] node4340;
	wire [11-1:0] node4343;
	wire [11-1:0] node4344;
	wire [11-1:0] node4347;
	wire [11-1:0] node4350;
	wire [11-1:0] node4351;
	wire [11-1:0] node4352;
	wire [11-1:0] node4353;
	wire [11-1:0] node4354;
	wire [11-1:0] node4358;
	wire [11-1:0] node4359;
	wire [11-1:0] node4362;
	wire [11-1:0] node4365;
	wire [11-1:0] node4366;
	wire [11-1:0] node4367;
	wire [11-1:0] node4370;
	wire [11-1:0] node4373;
	wire [11-1:0] node4374;
	wire [11-1:0] node4377;
	wire [11-1:0] node4380;
	wire [11-1:0] node4381;
	wire [11-1:0] node4382;
	wire [11-1:0] node4383;
	wire [11-1:0] node4386;
	wire [11-1:0] node4389;
	wire [11-1:0] node4390;
	wire [11-1:0] node4393;
	wire [11-1:0] node4396;
	wire [11-1:0] node4397;
	wire [11-1:0] node4398;
	wire [11-1:0] node4401;
	wire [11-1:0] node4404;
	wire [11-1:0] node4407;
	wire [11-1:0] node4408;
	wire [11-1:0] node4409;
	wire [11-1:0] node4410;
	wire [11-1:0] node4411;
	wire [11-1:0] node4412;
	wire [11-1:0] node4413;
	wire [11-1:0] node4414;
	wire [11-1:0] node4415;
	wire [11-1:0] node4418;
	wire [11-1:0] node4421;
	wire [11-1:0] node4422;
	wire [11-1:0] node4426;
	wire [11-1:0] node4427;
	wire [11-1:0] node4428;
	wire [11-1:0] node4432;
	wire [11-1:0] node4434;
	wire [11-1:0] node4437;
	wire [11-1:0] node4438;
	wire [11-1:0] node4439;
	wire [11-1:0] node4442;
	wire [11-1:0] node4443;
	wire [11-1:0] node4446;
	wire [11-1:0] node4449;
	wire [11-1:0] node4450;
	wire [11-1:0] node4451;
	wire [11-1:0] node4454;
	wire [11-1:0] node4457;
	wire [11-1:0] node4458;
	wire [11-1:0] node4461;
	wire [11-1:0] node4464;
	wire [11-1:0] node4465;
	wire [11-1:0] node4466;
	wire [11-1:0] node4467;
	wire [11-1:0] node4468;
	wire [11-1:0] node4471;
	wire [11-1:0] node4474;
	wire [11-1:0] node4475;
	wire [11-1:0] node4478;
	wire [11-1:0] node4481;
	wire [11-1:0] node4482;
	wire [11-1:0] node4483;
	wire [11-1:0] node4486;
	wire [11-1:0] node4489;
	wire [11-1:0] node4490;
	wire [11-1:0] node4493;
	wire [11-1:0] node4496;
	wire [11-1:0] node4497;
	wire [11-1:0] node4498;
	wire [11-1:0] node4499;
	wire [11-1:0] node4502;
	wire [11-1:0] node4505;
	wire [11-1:0] node4506;
	wire [11-1:0] node4509;
	wire [11-1:0] node4512;
	wire [11-1:0] node4513;
	wire [11-1:0] node4516;
	wire [11-1:0] node4517;
	wire [11-1:0] node4520;
	wire [11-1:0] node4523;
	wire [11-1:0] node4524;
	wire [11-1:0] node4525;
	wire [11-1:0] node4526;
	wire [11-1:0] node4527;
	wire [11-1:0] node4529;
	wire [11-1:0] node4532;
	wire [11-1:0] node4533;
	wire [11-1:0] node4536;
	wire [11-1:0] node4539;
	wire [11-1:0] node4540;
	wire [11-1:0] node4541;
	wire [11-1:0] node4544;
	wire [11-1:0] node4547;
	wire [11-1:0] node4548;
	wire [11-1:0] node4551;
	wire [11-1:0] node4554;
	wire [11-1:0] node4555;
	wire [11-1:0] node4556;
	wire [11-1:0] node4557;
	wire [11-1:0] node4561;
	wire [11-1:0] node4562;
	wire [11-1:0] node4566;
	wire [11-1:0] node4567;
	wire [11-1:0] node4569;
	wire [11-1:0] node4572;
	wire [11-1:0] node4573;
	wire [11-1:0] node4577;
	wire [11-1:0] node4578;
	wire [11-1:0] node4579;
	wire [11-1:0] node4580;
	wire [11-1:0] node4582;
	wire [11-1:0] node4585;
	wire [11-1:0] node4586;
	wire [11-1:0] node4589;
	wire [11-1:0] node4592;
	wire [11-1:0] node4593;
	wire [11-1:0] node4594;
	wire [11-1:0] node4597;
	wire [11-1:0] node4600;
	wire [11-1:0] node4601;
	wire [11-1:0] node4605;
	wire [11-1:0] node4606;
	wire [11-1:0] node4607;
	wire [11-1:0] node4608;
	wire [11-1:0] node4611;
	wire [11-1:0] node4614;
	wire [11-1:0] node4616;
	wire [11-1:0] node4619;
	wire [11-1:0] node4620;
	wire [11-1:0] node4623;
	wire [11-1:0] node4625;
	wire [11-1:0] node4628;
	wire [11-1:0] node4629;
	wire [11-1:0] node4630;
	wire [11-1:0] node4631;
	wire [11-1:0] node4632;
	wire [11-1:0] node4633;
	wire [11-1:0] node4634;
	wire [11-1:0] node4638;
	wire [11-1:0] node4639;
	wire [11-1:0] node4642;
	wire [11-1:0] node4645;
	wire [11-1:0] node4646;
	wire [11-1:0] node4649;
	wire [11-1:0] node4650;
	wire [11-1:0] node4653;
	wire [11-1:0] node4656;
	wire [11-1:0] node4657;
	wire [11-1:0] node4658;
	wire [11-1:0] node4660;
	wire [11-1:0] node4663;
	wire [11-1:0] node4665;
	wire [11-1:0] node4668;
	wire [11-1:0] node4669;
	wire [11-1:0] node4670;
	wire [11-1:0] node4673;
	wire [11-1:0] node4676;
	wire [11-1:0] node4677;
	wire [11-1:0] node4680;
	wire [11-1:0] node4683;
	wire [11-1:0] node4684;
	wire [11-1:0] node4685;
	wire [11-1:0] node4686;
	wire [11-1:0] node4687;
	wire [11-1:0] node4690;
	wire [11-1:0] node4693;
	wire [11-1:0] node4695;
	wire [11-1:0] node4698;
	wire [11-1:0] node4699;
	wire [11-1:0] node4700;
	wire [11-1:0] node4703;
	wire [11-1:0] node4706;
	wire [11-1:0] node4707;
	wire [11-1:0] node4710;
	wire [11-1:0] node4713;
	wire [11-1:0] node4714;
	wire [11-1:0] node4715;
	wire [11-1:0] node4716;
	wire [11-1:0] node4719;
	wire [11-1:0] node4722;
	wire [11-1:0] node4723;
	wire [11-1:0] node4726;
	wire [11-1:0] node4729;
	wire [11-1:0] node4730;
	wire [11-1:0] node4731;
	wire [11-1:0] node4735;
	wire [11-1:0] node4736;
	wire [11-1:0] node4740;
	wire [11-1:0] node4741;
	wire [11-1:0] node4742;
	wire [11-1:0] node4743;
	wire [11-1:0] node4744;
	wire [11-1:0] node4745;
	wire [11-1:0] node4748;
	wire [11-1:0] node4751;
	wire [11-1:0] node4752;
	wire [11-1:0] node4755;
	wire [11-1:0] node4758;
	wire [11-1:0] node4759;
	wire [11-1:0] node4760;
	wire [11-1:0] node4763;
	wire [11-1:0] node4766;
	wire [11-1:0] node4768;
	wire [11-1:0] node4771;
	wire [11-1:0] node4772;
	wire [11-1:0] node4773;
	wire [11-1:0] node4774;
	wire [11-1:0] node4777;
	wire [11-1:0] node4780;
	wire [11-1:0] node4781;
	wire [11-1:0] node4784;
	wire [11-1:0] node4787;
	wire [11-1:0] node4788;
	wire [11-1:0] node4789;
	wire [11-1:0] node4793;
	wire [11-1:0] node4794;
	wire [11-1:0] node4797;
	wire [11-1:0] node4800;
	wire [11-1:0] node4801;
	wire [11-1:0] node4802;
	wire [11-1:0] node4803;
	wire [11-1:0] node4804;
	wire [11-1:0] node4807;
	wire [11-1:0] node4810;
	wire [11-1:0] node4811;
	wire [11-1:0] node4815;
	wire [11-1:0] node4816;
	wire [11-1:0] node4817;
	wire [11-1:0] node4820;
	wire [11-1:0] node4823;
	wire [11-1:0] node4824;
	wire [11-1:0] node4827;
	wire [11-1:0] node4830;
	wire [11-1:0] node4831;
	wire [11-1:0] node4832;
	wire [11-1:0] node4833;
	wire [11-1:0] node4836;
	wire [11-1:0] node4839;
	wire [11-1:0] node4840;
	wire [11-1:0] node4844;
	wire [11-1:0] node4845;
	wire [11-1:0] node4848;
	wire [11-1:0] node4849;
	wire [11-1:0] node4853;
	wire [11-1:0] node4854;
	wire [11-1:0] node4855;
	wire [11-1:0] node4856;
	wire [11-1:0] node4857;
	wire [11-1:0] node4858;
	wire [11-1:0] node4860;
	wire [11-1:0] node4862;
	wire [11-1:0] node4865;
	wire [11-1:0] node4866;
	wire [11-1:0] node4867;
	wire [11-1:0] node4871;
	wire [11-1:0] node4872;
	wire [11-1:0] node4876;
	wire [11-1:0] node4877;
	wire [11-1:0] node4878;
	wire [11-1:0] node4879;
	wire [11-1:0] node4882;
	wire [11-1:0] node4885;
	wire [11-1:0] node4886;
	wire [11-1:0] node4890;
	wire [11-1:0] node4891;
	wire [11-1:0] node4892;
	wire [11-1:0] node4895;
	wire [11-1:0] node4898;
	wire [11-1:0] node4900;
	wire [11-1:0] node4903;
	wire [11-1:0] node4904;
	wire [11-1:0] node4905;
	wire [11-1:0] node4906;
	wire [11-1:0] node4907;
	wire [11-1:0] node4910;
	wire [11-1:0] node4913;
	wire [11-1:0] node4914;
	wire [11-1:0] node4917;
	wire [11-1:0] node4920;
	wire [11-1:0] node4921;
	wire [11-1:0] node4922;
	wire [11-1:0] node4925;
	wire [11-1:0] node4928;
	wire [11-1:0] node4929;
	wire [11-1:0] node4932;
	wire [11-1:0] node4935;
	wire [11-1:0] node4936;
	wire [11-1:0] node4937;
	wire [11-1:0] node4938;
	wire [11-1:0] node4941;
	wire [11-1:0] node4944;
	wire [11-1:0] node4945;
	wire [11-1:0] node4948;
	wire [11-1:0] node4951;
	wire [11-1:0] node4952;
	wire [11-1:0] node4953;
	wire [11-1:0] node4956;
	wire [11-1:0] node4959;
	wire [11-1:0] node4960;
	wire [11-1:0] node4964;
	wire [11-1:0] node4965;
	wire [11-1:0] node4966;
	wire [11-1:0] node4967;
	wire [11-1:0] node4968;
	wire [11-1:0] node4970;
	wire [11-1:0] node4973;
	wire [11-1:0] node4974;
	wire [11-1:0] node4977;
	wire [11-1:0] node4980;
	wire [11-1:0] node4981;
	wire [11-1:0] node4982;
	wire [11-1:0] node4986;
	wire [11-1:0] node4987;
	wire [11-1:0] node4991;
	wire [11-1:0] node4992;
	wire [11-1:0] node4993;
	wire [11-1:0] node4994;
	wire [11-1:0] node4997;
	wire [11-1:0] node5000;
	wire [11-1:0] node5001;
	wire [11-1:0] node5004;
	wire [11-1:0] node5007;
	wire [11-1:0] node5008;
	wire [11-1:0] node5009;
	wire [11-1:0] node5012;
	wire [11-1:0] node5015;
	wire [11-1:0] node5016;
	wire [11-1:0] node5019;
	wire [11-1:0] node5022;
	wire [11-1:0] node5023;
	wire [11-1:0] node5024;
	wire [11-1:0] node5025;
	wire [11-1:0] node5026;
	wire [11-1:0] node5029;
	wire [11-1:0] node5032;
	wire [11-1:0] node5034;
	wire [11-1:0] node5037;
	wire [11-1:0] node5038;
	wire [11-1:0] node5039;
	wire [11-1:0] node5042;
	wire [11-1:0] node5045;
	wire [11-1:0] node5046;
	wire [11-1:0] node5049;
	wire [11-1:0] node5052;
	wire [11-1:0] node5053;
	wire [11-1:0] node5054;
	wire [11-1:0] node5056;
	wire [11-1:0] node5059;
	wire [11-1:0] node5060;
	wire [11-1:0] node5063;
	wire [11-1:0] node5066;
	wire [11-1:0] node5067;
	wire [11-1:0] node5069;
	wire [11-1:0] node5072;
	wire [11-1:0] node5073;
	wire [11-1:0] node5077;
	wire [11-1:0] node5078;
	wire [11-1:0] node5079;
	wire [11-1:0] node5080;
	wire [11-1:0] node5081;
	wire [11-1:0] node5082;
	wire [11-1:0] node5083;
	wire [11-1:0] node5086;
	wire [11-1:0] node5089;
	wire [11-1:0] node5090;
	wire [11-1:0] node5093;
	wire [11-1:0] node5096;
	wire [11-1:0] node5097;
	wire [11-1:0] node5098;
	wire [11-1:0] node5101;
	wire [11-1:0] node5104;
	wire [11-1:0] node5105;
	wire [11-1:0] node5108;
	wire [11-1:0] node5111;
	wire [11-1:0] node5112;
	wire [11-1:0] node5113;
	wire [11-1:0] node5115;
	wire [11-1:0] node5118;
	wire [11-1:0] node5119;
	wire [11-1:0] node5123;
	wire [11-1:0] node5124;
	wire [11-1:0] node5127;
	wire [11-1:0] node5129;
	wire [11-1:0] node5132;
	wire [11-1:0] node5133;
	wire [11-1:0] node5134;
	wire [11-1:0] node5135;
	wire [11-1:0] node5136;
	wire [11-1:0] node5140;
	wire [11-1:0] node5141;
	wire [11-1:0] node5144;
	wire [11-1:0] node5147;
	wire [11-1:0] node5148;
	wire [11-1:0] node5149;
	wire [11-1:0] node5152;
	wire [11-1:0] node5155;
	wire [11-1:0] node5156;
	wire [11-1:0] node5160;
	wire [11-1:0] node5161;
	wire [11-1:0] node5162;
	wire [11-1:0] node5165;
	wire [11-1:0] node5166;
	wire [11-1:0] node5169;
	wire [11-1:0] node5172;
	wire [11-1:0] node5173;
	wire [11-1:0] node5174;
	wire [11-1:0] node5177;
	wire [11-1:0] node5180;
	wire [11-1:0] node5181;
	wire [11-1:0] node5185;
	wire [11-1:0] node5186;
	wire [11-1:0] node5187;
	wire [11-1:0] node5188;
	wire [11-1:0] node5189;
	wire [11-1:0] node5191;
	wire [11-1:0] node5194;
	wire [11-1:0] node5195;
	wire [11-1:0] node5198;
	wire [11-1:0] node5201;
	wire [11-1:0] node5202;
	wire [11-1:0] node5204;
	wire [11-1:0] node5207;
	wire [11-1:0] node5209;
	wire [11-1:0] node5212;
	wire [11-1:0] node5213;
	wire [11-1:0] node5214;
	wire [11-1:0] node5215;
	wire [11-1:0] node5218;
	wire [11-1:0] node5221;
	wire [11-1:0] node5222;
	wire [11-1:0] node5226;
	wire [11-1:0] node5227;
	wire [11-1:0] node5229;
	wire [11-1:0] node5232;
	wire [11-1:0] node5235;
	wire [11-1:0] node5236;
	wire [11-1:0] node5237;
	wire [11-1:0] node5238;
	wire [11-1:0] node5240;
	wire [11-1:0] node5243;
	wire [11-1:0] node5245;
	wire [11-1:0] node5248;
	wire [11-1:0] node5249;
	wire [11-1:0] node5250;
	wire [11-1:0] node5253;
	wire [11-1:0] node5256;
	wire [11-1:0] node5257;
	wire [11-1:0] node5260;
	wire [11-1:0] node5263;
	wire [11-1:0] node5264;
	wire [11-1:0] node5265;
	wire [11-1:0] node5266;
	wire [11-1:0] node5269;
	wire [11-1:0] node5272;
	wire [11-1:0] node5273;
	wire [11-1:0] node5276;
	wire [11-1:0] node5279;
	wire [11-1:0] node5280;
	wire [11-1:0] node5281;
	wire [11-1:0] node5285;
	wire [11-1:0] node5286;
	wire [11-1:0] node5290;
	wire [11-1:0] node5291;
	wire [11-1:0] node5292;
	wire [11-1:0] node5293;
	wire [11-1:0] node5294;
	wire [11-1:0] node5295;
	wire [11-1:0] node5296;
	wire [11-1:0] node5297;
	wire [11-1:0] node5299;
	wire [11-1:0] node5300;
	wire [11-1:0] node5303;
	wire [11-1:0] node5306;
	wire [11-1:0] node5307;
	wire [11-1:0] node5310;
	wire [11-1:0] node5311;
	wire [11-1:0] node5314;
	wire [11-1:0] node5317;
	wire [11-1:0] node5318;
	wire [11-1:0] node5319;
	wire [11-1:0] node5320;
	wire [11-1:0] node5323;
	wire [11-1:0] node5326;
	wire [11-1:0] node5327;
	wire [11-1:0] node5330;
	wire [11-1:0] node5333;
	wire [11-1:0] node5334;
	wire [11-1:0] node5335;
	wire [11-1:0] node5338;
	wire [11-1:0] node5341;
	wire [11-1:0] node5342;
	wire [11-1:0] node5345;
	wire [11-1:0] node5348;
	wire [11-1:0] node5349;
	wire [11-1:0] node5350;
	wire [11-1:0] node5351;
	wire [11-1:0] node5353;
	wire [11-1:0] node5356;
	wire [11-1:0] node5359;
	wire [11-1:0] node5360;
	wire [11-1:0] node5361;
	wire [11-1:0] node5364;
	wire [11-1:0] node5367;
	wire [11-1:0] node5368;
	wire [11-1:0] node5371;
	wire [11-1:0] node5374;
	wire [11-1:0] node5375;
	wire [11-1:0] node5376;
	wire [11-1:0] node5378;
	wire [11-1:0] node5381;
	wire [11-1:0] node5382;
	wire [11-1:0] node5385;
	wire [11-1:0] node5388;
	wire [11-1:0] node5389;
	wire [11-1:0] node5390;
	wire [11-1:0] node5394;
	wire [11-1:0] node5395;
	wire [11-1:0] node5398;
	wire [11-1:0] node5401;
	wire [11-1:0] node5402;
	wire [11-1:0] node5403;
	wire [11-1:0] node5404;
	wire [11-1:0] node5405;
	wire [11-1:0] node5407;
	wire [11-1:0] node5410;
	wire [11-1:0] node5411;
	wire [11-1:0] node5414;
	wire [11-1:0] node5417;
	wire [11-1:0] node5418;
	wire [11-1:0] node5419;
	wire [11-1:0] node5422;
	wire [11-1:0] node5425;
	wire [11-1:0] node5428;
	wire [11-1:0] node5429;
	wire [11-1:0] node5430;
	wire [11-1:0] node5431;
	wire [11-1:0] node5435;
	wire [11-1:0] node5436;
	wire [11-1:0] node5439;
	wire [11-1:0] node5442;
	wire [11-1:0] node5443;
	wire [11-1:0] node5444;
	wire [11-1:0] node5447;
	wire [11-1:0] node5450;
	wire [11-1:0] node5452;
	wire [11-1:0] node5455;
	wire [11-1:0] node5456;
	wire [11-1:0] node5457;
	wire [11-1:0] node5458;
	wire [11-1:0] node5459;
	wire [11-1:0] node5463;
	wire [11-1:0] node5464;
	wire [11-1:0] node5467;
	wire [11-1:0] node5470;
	wire [11-1:0] node5471;
	wire [11-1:0] node5472;
	wire [11-1:0] node5475;
	wire [11-1:0] node5478;
	wire [11-1:0] node5480;
	wire [11-1:0] node5483;
	wire [11-1:0] node5484;
	wire [11-1:0] node5485;
	wire [11-1:0] node5488;
	wire [11-1:0] node5489;
	wire [11-1:0] node5492;
	wire [11-1:0] node5495;
	wire [11-1:0] node5496;
	wire [11-1:0] node5498;
	wire [11-1:0] node5501;
	wire [11-1:0] node5503;
	wire [11-1:0] node5506;
	wire [11-1:0] node5507;
	wire [11-1:0] node5508;
	wire [11-1:0] node5509;
	wire [11-1:0] node5510;
	wire [11-1:0] node5511;
	wire [11-1:0] node5512;
	wire [11-1:0] node5516;
	wire [11-1:0] node5517;
	wire [11-1:0] node5520;
	wire [11-1:0] node5523;
	wire [11-1:0] node5524;
	wire [11-1:0] node5525;
	wire [11-1:0] node5529;
	wire [11-1:0] node5531;
	wire [11-1:0] node5534;
	wire [11-1:0] node5535;
	wire [11-1:0] node5536;
	wire [11-1:0] node5537;
	wire [11-1:0] node5541;
	wire [11-1:0] node5542;
	wire [11-1:0] node5545;
	wire [11-1:0] node5548;
	wire [11-1:0] node5549;
	wire [11-1:0] node5550;
	wire [11-1:0] node5553;
	wire [11-1:0] node5556;
	wire [11-1:0] node5557;
	wire [11-1:0] node5561;
	wire [11-1:0] node5562;
	wire [11-1:0] node5563;
	wire [11-1:0] node5564;
	wire [11-1:0] node5565;
	wire [11-1:0] node5568;
	wire [11-1:0] node5571;
	wire [11-1:0] node5572;
	wire [11-1:0] node5576;
	wire [11-1:0] node5577;
	wire [11-1:0] node5578;
	wire [11-1:0] node5582;
	wire [11-1:0] node5583;
	wire [11-1:0] node5586;
	wire [11-1:0] node5589;
	wire [11-1:0] node5590;
	wire [11-1:0] node5591;
	wire [11-1:0] node5592;
	wire [11-1:0] node5595;
	wire [11-1:0] node5598;
	wire [11-1:0] node5599;
	wire [11-1:0] node5602;
	wire [11-1:0] node5605;
	wire [11-1:0] node5606;
	wire [11-1:0] node5607;
	wire [11-1:0] node5611;
	wire [11-1:0] node5613;
	wire [11-1:0] node5616;
	wire [11-1:0] node5617;
	wire [11-1:0] node5618;
	wire [11-1:0] node5619;
	wire [11-1:0] node5620;
	wire [11-1:0] node5623;
	wire [11-1:0] node5624;
	wire [11-1:0] node5627;
	wire [11-1:0] node5630;
	wire [11-1:0] node5631;
	wire [11-1:0] node5632;
	wire [11-1:0] node5636;
	wire [11-1:0] node5637;
	wire [11-1:0] node5640;
	wire [11-1:0] node5643;
	wire [11-1:0] node5644;
	wire [11-1:0] node5645;
	wire [11-1:0] node5646;
	wire [11-1:0] node5649;
	wire [11-1:0] node5652;
	wire [11-1:0] node5653;
	wire [11-1:0] node5656;
	wire [11-1:0] node5659;
	wire [11-1:0] node5660;
	wire [11-1:0] node5661;
	wire [11-1:0] node5664;
	wire [11-1:0] node5667;
	wire [11-1:0] node5669;
	wire [11-1:0] node5672;
	wire [11-1:0] node5673;
	wire [11-1:0] node5674;
	wire [11-1:0] node5675;
	wire [11-1:0] node5676;
	wire [11-1:0] node5679;
	wire [11-1:0] node5682;
	wire [11-1:0] node5683;
	wire [11-1:0] node5686;
	wire [11-1:0] node5689;
	wire [11-1:0] node5690;
	wire [11-1:0] node5691;
	wire [11-1:0] node5694;
	wire [11-1:0] node5697;
	wire [11-1:0] node5698;
	wire [11-1:0] node5701;
	wire [11-1:0] node5704;
	wire [11-1:0] node5705;
	wire [11-1:0] node5706;
	wire [11-1:0] node5707;
	wire [11-1:0] node5710;
	wire [11-1:0] node5713;
	wire [11-1:0] node5714;
	wire [11-1:0] node5718;
	wire [11-1:0] node5719;
	wire [11-1:0] node5721;
	wire [11-1:0] node5724;
	wire [11-1:0] node5725;
	wire [11-1:0] node5728;
	wire [11-1:0] node5731;
	wire [11-1:0] node5732;
	wire [11-1:0] node5733;
	wire [11-1:0] node5734;
	wire [11-1:0] node5735;
	wire [11-1:0] node5736;
	wire [11-1:0] node5737;
	wire [11-1:0] node5738;
	wire [11-1:0] node5742;
	wire [11-1:0] node5744;
	wire [11-1:0] node5747;
	wire [11-1:0] node5748;
	wire [11-1:0] node5750;
	wire [11-1:0] node5753;
	wire [11-1:0] node5754;
	wire [11-1:0] node5757;
	wire [11-1:0] node5760;
	wire [11-1:0] node5761;
	wire [11-1:0] node5762;
	wire [11-1:0] node5763;
	wire [11-1:0] node5767;
	wire [11-1:0] node5770;
	wire [11-1:0] node5771;
	wire [11-1:0] node5772;
	wire [11-1:0] node5775;
	wire [11-1:0] node5778;
	wire [11-1:0] node5780;
	wire [11-1:0] node5783;
	wire [11-1:0] node5784;
	wire [11-1:0] node5785;
	wire [11-1:0] node5786;
	wire [11-1:0] node5787;
	wire [11-1:0] node5790;
	wire [11-1:0] node5793;
	wire [11-1:0] node5794;
	wire [11-1:0] node5797;
	wire [11-1:0] node5800;
	wire [11-1:0] node5801;
	wire [11-1:0] node5803;
	wire [11-1:0] node5806;
	wire [11-1:0] node5807;
	wire [11-1:0] node5810;
	wire [11-1:0] node5813;
	wire [11-1:0] node5814;
	wire [11-1:0] node5815;
	wire [11-1:0] node5816;
	wire [11-1:0] node5820;
	wire [11-1:0] node5821;
	wire [11-1:0] node5825;
	wire [11-1:0] node5826;
	wire [11-1:0] node5828;
	wire [11-1:0] node5831;
	wire [11-1:0] node5832;
	wire [11-1:0] node5836;
	wire [11-1:0] node5837;
	wire [11-1:0] node5838;
	wire [11-1:0] node5839;
	wire [11-1:0] node5840;
	wire [11-1:0] node5841;
	wire [11-1:0] node5844;
	wire [11-1:0] node5847;
	wire [11-1:0] node5848;
	wire [11-1:0] node5851;
	wire [11-1:0] node5854;
	wire [11-1:0] node5855;
	wire [11-1:0] node5856;
	wire [11-1:0] node5859;
	wire [11-1:0] node5862;
	wire [11-1:0] node5863;
	wire [11-1:0] node5866;
	wire [11-1:0] node5869;
	wire [11-1:0] node5870;
	wire [11-1:0] node5871;
	wire [11-1:0] node5872;
	wire [11-1:0] node5875;
	wire [11-1:0] node5878;
	wire [11-1:0] node5879;
	wire [11-1:0] node5882;
	wire [11-1:0] node5885;
	wire [11-1:0] node5886;
	wire [11-1:0] node5889;
	wire [11-1:0] node5890;
	wire [11-1:0] node5893;
	wire [11-1:0] node5896;
	wire [11-1:0] node5897;
	wire [11-1:0] node5898;
	wire [11-1:0] node5899;
	wire [11-1:0] node5902;
	wire [11-1:0] node5903;
	wire [11-1:0] node5906;
	wire [11-1:0] node5909;
	wire [11-1:0] node5910;
	wire [11-1:0] node5913;
	wire [11-1:0] node5914;
	wire [11-1:0] node5918;
	wire [11-1:0] node5919;
	wire [11-1:0] node5920;
	wire [11-1:0] node5921;
	wire [11-1:0] node5924;
	wire [11-1:0] node5927;
	wire [11-1:0] node5928;
	wire [11-1:0] node5932;
	wire [11-1:0] node5933;
	wire [11-1:0] node5934;
	wire [11-1:0] node5937;
	wire [11-1:0] node5940;
	wire [11-1:0] node5942;
	wire [11-1:0] node5945;
	wire [11-1:0] node5946;
	wire [11-1:0] node5947;
	wire [11-1:0] node5948;
	wire [11-1:0] node5949;
	wire [11-1:0] node5950;
	wire [11-1:0] node5951;
	wire [11-1:0] node5954;
	wire [11-1:0] node5957;
	wire [11-1:0] node5958;
	wire [11-1:0] node5961;
	wire [11-1:0] node5964;
	wire [11-1:0] node5965;
	wire [11-1:0] node5966;
	wire [11-1:0] node5969;
	wire [11-1:0] node5972;
	wire [11-1:0] node5973;
	wire [11-1:0] node5976;
	wire [11-1:0] node5979;
	wire [11-1:0] node5980;
	wire [11-1:0] node5981;
	wire [11-1:0] node5982;
	wire [11-1:0] node5985;
	wire [11-1:0] node5988;
	wire [11-1:0] node5989;
	wire [11-1:0] node5992;
	wire [11-1:0] node5995;
	wire [11-1:0] node5996;
	wire [11-1:0] node5997;
	wire [11-1:0] node6000;
	wire [11-1:0] node6003;
	wire [11-1:0] node6005;
	wire [11-1:0] node6008;
	wire [11-1:0] node6009;
	wire [11-1:0] node6010;
	wire [11-1:0] node6011;
	wire [11-1:0] node6012;
	wire [11-1:0] node6015;
	wire [11-1:0] node6018;
	wire [11-1:0] node6019;
	wire [11-1:0] node6022;
	wire [11-1:0] node6025;
	wire [11-1:0] node6026;
	wire [11-1:0] node6029;
	wire [11-1:0] node6030;
	wire [11-1:0] node6034;
	wire [11-1:0] node6035;
	wire [11-1:0] node6036;
	wire [11-1:0] node6037;
	wire [11-1:0] node6040;
	wire [11-1:0] node6043;
	wire [11-1:0] node6044;
	wire [11-1:0] node6047;
	wire [11-1:0] node6050;
	wire [11-1:0] node6051;
	wire [11-1:0] node6053;
	wire [11-1:0] node6056;
	wire [11-1:0] node6057;
	wire [11-1:0] node6061;
	wire [11-1:0] node6062;
	wire [11-1:0] node6063;
	wire [11-1:0] node6064;
	wire [11-1:0] node6065;
	wire [11-1:0] node6066;
	wire [11-1:0] node6069;
	wire [11-1:0] node6072;
	wire [11-1:0] node6073;
	wire [11-1:0] node6077;
	wire [11-1:0] node6078;
	wire [11-1:0] node6081;
	wire [11-1:0] node6082;
	wire [11-1:0] node6085;
	wire [11-1:0] node6088;
	wire [11-1:0] node6089;
	wire [11-1:0] node6090;
	wire [11-1:0] node6091;
	wire [11-1:0] node6095;
	wire [11-1:0] node6096;
	wire [11-1:0] node6100;
	wire [11-1:0] node6101;
	wire [11-1:0] node6104;
	wire [11-1:0] node6105;
	wire [11-1:0] node6109;
	wire [11-1:0] node6110;
	wire [11-1:0] node6111;
	wire [11-1:0] node6112;
	wire [11-1:0] node6113;
	wire [11-1:0] node6117;
	wire [11-1:0] node6118;
	wire [11-1:0] node6121;
	wire [11-1:0] node6124;
	wire [11-1:0] node6125;
	wire [11-1:0] node6126;
	wire [11-1:0] node6129;
	wire [11-1:0] node6132;
	wire [11-1:0] node6133;
	wire [11-1:0] node6136;
	wire [11-1:0] node6139;
	wire [11-1:0] node6140;
	wire [11-1:0] node6141;
	wire [11-1:0] node6142;
	wire [11-1:0] node6146;
	wire [11-1:0] node6147;
	wire [11-1:0] node6150;
	wire [11-1:0] node6153;
	wire [11-1:0] node6154;
	wire [11-1:0] node6158;
	wire [11-1:0] node6159;
	wire [11-1:0] node6160;
	wire [11-1:0] node6161;
	wire [11-1:0] node6162;
	wire [11-1:0] node6163;
	wire [11-1:0] node6164;
	wire [11-1:0] node6165;
	wire [11-1:0] node6167;
	wire [11-1:0] node6170;
	wire [11-1:0] node6171;
	wire [11-1:0] node6174;
	wire [11-1:0] node6177;
	wire [11-1:0] node6178;
	wire [11-1:0] node6179;
	wire [11-1:0] node6182;
	wire [11-1:0] node6185;
	wire [11-1:0] node6186;
	wire [11-1:0] node6190;
	wire [11-1:0] node6191;
	wire [11-1:0] node6192;
	wire [11-1:0] node6193;
	wire [11-1:0] node6196;
	wire [11-1:0] node6199;
	wire [11-1:0] node6201;
	wire [11-1:0] node6204;
	wire [11-1:0] node6205;
	wire [11-1:0] node6206;
	wire [11-1:0] node6210;
	wire [11-1:0] node6212;
	wire [11-1:0] node6215;
	wire [11-1:0] node6216;
	wire [11-1:0] node6217;
	wire [11-1:0] node6218;
	wire [11-1:0] node6219;
	wire [11-1:0] node6223;
	wire [11-1:0] node6225;
	wire [11-1:0] node6228;
	wire [11-1:0] node6229;
	wire [11-1:0] node6230;
	wire [11-1:0] node6234;
	wire [11-1:0] node6235;
	wire [11-1:0] node6239;
	wire [11-1:0] node6240;
	wire [11-1:0] node6241;
	wire [11-1:0] node6242;
	wire [11-1:0] node6245;
	wire [11-1:0] node6248;
	wire [11-1:0] node6250;
	wire [11-1:0] node6253;
	wire [11-1:0] node6254;
	wire [11-1:0] node6255;
	wire [11-1:0] node6258;
	wire [11-1:0] node6261;
	wire [11-1:0] node6264;
	wire [11-1:0] node6265;
	wire [11-1:0] node6266;
	wire [11-1:0] node6267;
	wire [11-1:0] node6268;
	wire [11-1:0] node6270;
	wire [11-1:0] node6273;
	wire [11-1:0] node6276;
	wire [11-1:0] node6277;
	wire [11-1:0] node6278;
	wire [11-1:0] node6281;
	wire [11-1:0] node6284;
	wire [11-1:0] node6285;
	wire [11-1:0] node6288;
	wire [11-1:0] node6291;
	wire [11-1:0] node6292;
	wire [11-1:0] node6293;
	wire [11-1:0] node6294;
	wire [11-1:0] node6297;
	wire [11-1:0] node6300;
	wire [11-1:0] node6301;
	wire [11-1:0] node6304;
	wire [11-1:0] node6307;
	wire [11-1:0] node6308;
	wire [11-1:0] node6309;
	wire [11-1:0] node6312;
	wire [11-1:0] node6315;
	wire [11-1:0] node6316;
	wire [11-1:0] node6319;
	wire [11-1:0] node6322;
	wire [11-1:0] node6323;
	wire [11-1:0] node6324;
	wire [11-1:0] node6325;
	wire [11-1:0] node6326;
	wire [11-1:0] node6330;
	wire [11-1:0] node6331;
	wire [11-1:0] node6334;
	wire [11-1:0] node6337;
	wire [11-1:0] node6338;
	wire [11-1:0] node6340;
	wire [11-1:0] node6343;
	wire [11-1:0] node6344;
	wire [11-1:0] node6348;
	wire [11-1:0] node6349;
	wire [11-1:0] node6350;
	wire [11-1:0] node6353;
	wire [11-1:0] node6354;
	wire [11-1:0] node6357;
	wire [11-1:0] node6360;
	wire [11-1:0] node6361;
	wire [11-1:0] node6362;
	wire [11-1:0] node6366;
	wire [11-1:0] node6367;
	wire [11-1:0] node6371;
	wire [11-1:0] node6372;
	wire [11-1:0] node6373;
	wire [11-1:0] node6374;
	wire [11-1:0] node6375;
	wire [11-1:0] node6376;
	wire [11-1:0] node6378;
	wire [11-1:0] node6381;
	wire [11-1:0] node6383;
	wire [11-1:0] node6386;
	wire [11-1:0] node6387;
	wire [11-1:0] node6388;
	wire [11-1:0] node6392;
	wire [11-1:0] node6393;
	wire [11-1:0] node6396;
	wire [11-1:0] node6399;
	wire [11-1:0] node6400;
	wire [11-1:0] node6401;
	wire [11-1:0] node6402;
	wire [11-1:0] node6406;
	wire [11-1:0] node6408;
	wire [11-1:0] node6411;
	wire [11-1:0] node6412;
	wire [11-1:0] node6413;
	wire [11-1:0] node6416;
	wire [11-1:0] node6419;
	wire [11-1:0] node6420;
	wire [11-1:0] node6423;
	wire [11-1:0] node6426;
	wire [11-1:0] node6427;
	wire [11-1:0] node6428;
	wire [11-1:0] node6429;
	wire [11-1:0] node6430;
	wire [11-1:0] node6433;
	wire [11-1:0] node6436;
	wire [11-1:0] node6437;
	wire [11-1:0] node6441;
	wire [11-1:0] node6442;
	wire [11-1:0] node6443;
	wire [11-1:0] node6447;
	wire [11-1:0] node6449;
	wire [11-1:0] node6452;
	wire [11-1:0] node6453;
	wire [11-1:0] node6454;
	wire [11-1:0] node6455;
	wire [11-1:0] node6458;
	wire [11-1:0] node6461;
	wire [11-1:0] node6462;
	wire [11-1:0] node6466;
	wire [11-1:0] node6467;
	wire [11-1:0] node6468;
	wire [11-1:0] node6471;
	wire [11-1:0] node6474;
	wire [11-1:0] node6475;
	wire [11-1:0] node6479;
	wire [11-1:0] node6480;
	wire [11-1:0] node6481;
	wire [11-1:0] node6482;
	wire [11-1:0] node6483;
	wire [11-1:0] node6484;
	wire [11-1:0] node6487;
	wire [11-1:0] node6490;
	wire [11-1:0] node6491;
	wire [11-1:0] node6495;
	wire [11-1:0] node6496;
	wire [11-1:0] node6497;
	wire [11-1:0] node6500;
	wire [11-1:0] node6503;
	wire [11-1:0] node6504;
	wire [11-1:0] node6507;
	wire [11-1:0] node6510;
	wire [11-1:0] node6511;
	wire [11-1:0] node6512;
	wire [11-1:0] node6513;
	wire [11-1:0] node6517;
	wire [11-1:0] node6518;
	wire [11-1:0] node6522;
	wire [11-1:0] node6523;
	wire [11-1:0] node6524;
	wire [11-1:0] node6527;
	wire [11-1:0] node6530;
	wire [11-1:0] node6531;
	wire [11-1:0] node6535;
	wire [11-1:0] node6536;
	wire [11-1:0] node6537;
	wire [11-1:0] node6538;
	wire [11-1:0] node6540;
	wire [11-1:0] node6543;
	wire [11-1:0] node6545;
	wire [11-1:0] node6548;
	wire [11-1:0] node6549;
	wire [11-1:0] node6550;
	wire [11-1:0] node6553;
	wire [11-1:0] node6556;
	wire [11-1:0] node6559;
	wire [11-1:0] node6560;
	wire [11-1:0] node6561;
	wire [11-1:0] node6564;
	wire [11-1:0] node6565;
	wire [11-1:0] node6569;
	wire [11-1:0] node6570;
	wire [11-1:0] node6573;
	wire [11-1:0] node6574;
	wire [11-1:0] node6578;
	wire [11-1:0] node6579;
	wire [11-1:0] node6580;
	wire [11-1:0] node6581;
	wire [11-1:0] node6582;
	wire [11-1:0] node6583;
	wire [11-1:0] node6584;
	wire [11-1:0] node6585;
	wire [11-1:0] node6588;
	wire [11-1:0] node6591;
	wire [11-1:0] node6592;
	wire [11-1:0] node6595;
	wire [11-1:0] node6598;
	wire [11-1:0] node6599;
	wire [11-1:0] node6601;
	wire [11-1:0] node6604;
	wire [11-1:0] node6605;
	wire [11-1:0] node6608;
	wire [11-1:0] node6611;
	wire [11-1:0] node6612;
	wire [11-1:0] node6613;
	wire [11-1:0] node6616;
	wire [11-1:0] node6617;
	wire [11-1:0] node6621;
	wire [11-1:0] node6622;
	wire [11-1:0] node6623;
	wire [11-1:0] node6626;
	wire [11-1:0] node6629;
	wire [11-1:0] node6630;
	wire [11-1:0] node6634;
	wire [11-1:0] node6635;
	wire [11-1:0] node6636;
	wire [11-1:0] node6637;
	wire [11-1:0] node6638;
	wire [11-1:0] node6641;
	wire [11-1:0] node6644;
	wire [11-1:0] node6645;
	wire [11-1:0] node6648;
	wire [11-1:0] node6651;
	wire [11-1:0] node6652;
	wire [11-1:0] node6653;
	wire [11-1:0] node6656;
	wire [11-1:0] node6659;
	wire [11-1:0] node6660;
	wire [11-1:0] node6663;
	wire [11-1:0] node6666;
	wire [11-1:0] node6667;
	wire [11-1:0] node6668;
	wire [11-1:0] node6669;
	wire [11-1:0] node6672;
	wire [11-1:0] node6675;
	wire [11-1:0] node6676;
	wire [11-1:0] node6679;
	wire [11-1:0] node6682;
	wire [11-1:0] node6683;
	wire [11-1:0] node6684;
	wire [11-1:0] node6687;
	wire [11-1:0] node6690;
	wire [11-1:0] node6691;
	wire [11-1:0] node6694;
	wire [11-1:0] node6697;
	wire [11-1:0] node6698;
	wire [11-1:0] node6699;
	wire [11-1:0] node6700;
	wire [11-1:0] node6701;
	wire [11-1:0] node6703;
	wire [11-1:0] node6706;
	wire [11-1:0] node6707;
	wire [11-1:0] node6710;
	wire [11-1:0] node6713;
	wire [11-1:0] node6714;
	wire [11-1:0] node6715;
	wire [11-1:0] node6718;
	wire [11-1:0] node6721;
	wire [11-1:0] node6723;
	wire [11-1:0] node6726;
	wire [11-1:0] node6727;
	wire [11-1:0] node6728;
	wire [11-1:0] node6729;
	wire [11-1:0] node6732;
	wire [11-1:0] node6735;
	wire [11-1:0] node6736;
	wire [11-1:0] node6739;
	wire [11-1:0] node6742;
	wire [11-1:0] node6743;
	wire [11-1:0] node6745;
	wire [11-1:0] node6748;
	wire [11-1:0] node6751;
	wire [11-1:0] node6752;
	wire [11-1:0] node6753;
	wire [11-1:0] node6754;
	wire [11-1:0] node6756;
	wire [11-1:0] node6759;
	wire [11-1:0] node6760;
	wire [11-1:0] node6764;
	wire [11-1:0] node6766;
	wire [11-1:0] node6767;
	wire [11-1:0] node6771;
	wire [11-1:0] node6772;
	wire [11-1:0] node6773;
	wire [11-1:0] node6776;
	wire [11-1:0] node6777;
	wire [11-1:0] node6780;
	wire [11-1:0] node6783;
	wire [11-1:0] node6784;
	wire [11-1:0] node6786;
	wire [11-1:0] node6790;
	wire [11-1:0] node6791;
	wire [11-1:0] node6792;
	wire [11-1:0] node6793;
	wire [11-1:0] node6794;
	wire [11-1:0] node6795;
	wire [11-1:0] node6796;
	wire [11-1:0] node6800;
	wire [11-1:0] node6801;
	wire [11-1:0] node6804;
	wire [11-1:0] node6807;
	wire [11-1:0] node6808;
	wire [11-1:0] node6811;
	wire [11-1:0] node6814;
	wire [11-1:0] node6815;
	wire [11-1:0] node6816;
	wire [11-1:0] node6817;
	wire [11-1:0] node6820;
	wire [11-1:0] node6823;
	wire [11-1:0] node6824;
	wire [11-1:0] node6828;
	wire [11-1:0] node6829;
	wire [11-1:0] node6831;
	wire [11-1:0] node6834;
	wire [11-1:0] node6837;
	wire [11-1:0] node6838;
	wire [11-1:0] node6839;
	wire [11-1:0] node6840;
	wire [11-1:0] node6841;
	wire [11-1:0] node6844;
	wire [11-1:0] node6847;
	wire [11-1:0] node6848;
	wire [11-1:0] node6851;
	wire [11-1:0] node6854;
	wire [11-1:0] node6855;
	wire [11-1:0] node6856;
	wire [11-1:0] node6859;
	wire [11-1:0] node6862;
	wire [11-1:0] node6863;
	wire [11-1:0] node6866;
	wire [11-1:0] node6869;
	wire [11-1:0] node6870;
	wire [11-1:0] node6871;
	wire [11-1:0] node6873;
	wire [11-1:0] node6876;
	wire [11-1:0] node6877;
	wire [11-1:0] node6880;
	wire [11-1:0] node6883;
	wire [11-1:0] node6884;
	wire [11-1:0] node6885;
	wire [11-1:0] node6889;
	wire [11-1:0] node6890;
	wire [11-1:0] node6894;
	wire [11-1:0] node6895;
	wire [11-1:0] node6896;
	wire [11-1:0] node6897;
	wire [11-1:0] node6898;
	wire [11-1:0] node6900;
	wire [11-1:0] node6903;
	wire [11-1:0] node6904;
	wire [11-1:0] node6907;
	wire [11-1:0] node6910;
	wire [11-1:0] node6911;
	wire [11-1:0] node6913;
	wire [11-1:0] node6916;
	wire [11-1:0] node6917;
	wire [11-1:0] node6920;
	wire [11-1:0] node6923;
	wire [11-1:0] node6924;
	wire [11-1:0] node6925;
	wire [11-1:0] node6926;
	wire [11-1:0] node6930;
	wire [11-1:0] node6931;
	wire [11-1:0] node6934;
	wire [11-1:0] node6937;
	wire [11-1:0] node6938;
	wire [11-1:0] node6940;
	wire [11-1:0] node6943;
	wire [11-1:0] node6944;
	wire [11-1:0] node6948;
	wire [11-1:0] node6949;
	wire [11-1:0] node6950;
	wire [11-1:0] node6951;
	wire [11-1:0] node6952;
	wire [11-1:0] node6956;
	wire [11-1:0] node6957;
	wire [11-1:0] node6960;
	wire [11-1:0] node6963;
	wire [11-1:0] node6964;
	wire [11-1:0] node6965;
	wire [11-1:0] node6968;
	wire [11-1:0] node6971;
	wire [11-1:0] node6972;
	wire [11-1:0] node6976;
	wire [11-1:0] node6977;
	wire [11-1:0] node6978;
	wire [11-1:0] node6979;
	wire [11-1:0] node6983;
	wire [11-1:0] node6985;
	wire [11-1:0] node6988;
	wire [11-1:0] node6989;
	wire [11-1:0] node6991;

	assign outp = (inp[1]) ? node3514 : node1;
		assign node1 = (inp[7]) ? node1751 : node2;
			assign node2 = (inp[2]) ? node874 : node3;
				assign node3 = (inp[0]) ? node439 : node4;
					assign node4 = (inp[4]) ? node218 : node5;
						assign node5 = (inp[10]) ? node115 : node6;
							assign node6 = (inp[3]) ? node60 : node7;
								assign node7 = (inp[9]) ? node31 : node8;
									assign node8 = (inp[5]) ? node20 : node9;
										assign node9 = (inp[6]) ? node15 : node10;
											assign node10 = (inp[8]) ? node12 : 11'b01001101011;
												assign node12 = (inp[11]) ? 11'b01000001001 : 11'b01000001010;
											assign node15 = (inp[8]) ? 11'b01011101000 : node16;
												assign node16 = (inp[11]) ? 11'b01010000010 : 11'b01001100010;
										assign node20 = (inp[11]) ? node28 : node21;
											assign node21 = (inp[8]) ? node25 : node22;
												assign node22 = (inp[6]) ? 11'b01001011011 : 11'b01001111010;
												assign node25 = (inp[6]) ? 11'b01000111011 : 11'b01000011011;
											assign node28 = (inp[8]) ? 11'b01001011010 : 11'b01011011001;
									assign node31 = (inp[11]) ? node45 : node32;
										assign node32 = (inp[6]) ? node40 : node33;
											assign node33 = (inp[8]) ? node37 : node34;
												assign node34 = (inp[5]) ? 11'b01001111010 : 11'b01001101011;
												assign node37 = (inp[5]) ? 11'b01010111010 : 11'b01010101011;
											assign node40 = (inp[5]) ? 11'b01010011001 : node41;
												assign node41 = (inp[8]) ? 11'b01010001000 : 11'b01000100000;
										assign node45 = (inp[5]) ? node53 : node46;
											assign node46 = (inp[6]) ? node50 : node47;
												assign node47 = (inp[8]) ? 11'b01110111001 : 11'b01101111011;
												assign node50 = (inp[8]) ? 11'b01101011010 : 11'b01111111001;
											assign node53 = (inp[6]) ? node57 : node54;
												assign node54 = (inp[8]) ? 11'b01001101010 : 11'b01110101000;
												assign node57 = (inp[8]) ? 11'b01010101001 : 11'b01111001011;
								assign node60 = (inp[9]) ? node88 : node61;
									assign node61 = (inp[11]) ? node75 : node62;
										assign node62 = (inp[5]) ? node70 : node63;
											assign node63 = (inp[6]) ? node67 : node64;
												assign node64 = (inp[8]) ? 11'b11101101011 : 11'b11001101011;
												assign node67 = (inp[8]) ? 11'b11111001010 : 11'b11011100010;
											assign node70 = (inp[8]) ? 11'b11000111001 : node71;
												assign node71 = (inp[6]) ? 11'b11011011011 : 11'b11001111010;
										assign node75 = (inp[5]) ? node81 : node76;
											assign node76 = (inp[8]) ? 11'b11100011001 : node77;
												assign node77 = (inp[6]) ? 11'b11000010010 : 11'b11001111011;
											assign node81 = (inp[8]) ? node85 : node82;
												assign node82 = (inp[6]) ? 11'b11100001001 : 11'b11101101000;
												assign node85 = (inp[6]) ? 11'b11001101011 : 11'b11010001010;
									assign node88 = (inp[5]) ? node102 : node89;
										assign node89 = (inp[6]) ? node97 : node90;
											assign node90 = (inp[11]) ? node94 : node91;
												assign node91 = (inp[8]) ? 11'b11111101111 : 11'b11001101111;
												assign node94 = (inp[8]) ? 11'b11100101101 : 11'b11101101111;
											assign node97 = (inp[8]) ? node99 : 11'b11100101101;
												assign node99 = (inp[11]) ? 11'b11111001110 : 11'b11100001100;
										assign node102 = (inp[6]) ? node108 : node103;
											assign node103 = (inp[8]) ? 11'b11100111110 : node104;
												assign node104 = (inp[11]) ? 11'b11011111100 : 11'b11001111110;
											assign node108 = (inp[8]) ? node112 : node109;
												assign node109 = (inp[11]) ? 11'b11010011111 : 11'b11001111111;
												assign node112 = (inp[11]) ? 11'b11100111111 : 11'b11010111111;
							assign node115 = (inp[3]) ? node165 : node116;
								assign node116 = (inp[9]) ? node138 : node117;
									assign node117 = (inp[5]) ? node127 : node118;
										assign node118 = (inp[6]) ? node124 : node119;
											assign node119 = (inp[8]) ? node121 : 11'b11000101011;
												assign node121 = (inp[11]) ? 11'b11111101001 : 11'b11001101011;
											assign node124 = (inp[11]) ? 11'b11011101011 : 11'b11011001010;
										assign node127 = (inp[6]) ? node133 : node128;
											assign node128 = (inp[11]) ? 11'b11010011010 : node129;
												assign node129 = (inp[8]) ? 11'b11101111010 : 11'b11100111010;
											assign node133 = (inp[8]) ? node135 : 11'b11110011001;
												assign node135 = (inp[11]) ? 11'b11001111001 : 11'b11110111001;
									assign node138 = (inp[5]) ? node150 : node139;
										assign node139 = (inp[8]) ? node145 : node140;
											assign node140 = (inp[6]) ? 11'b11110111101 : node141;
												assign node141 = (inp[11]) ? 11'b11100111111 : 11'b11000111111;
											assign node145 = (inp[6]) ? 11'b11001011110 : node146;
												assign node146 = (inp[11]) ? 11'b11001111101 : 11'b11011111111;
										assign node150 = (inp[6]) ? node158 : node151;
											assign node151 = (inp[11]) ? node155 : node152;
												assign node152 = (inp[8]) ? 11'b11000101100 : 11'b11100101110;
												assign node155 = (inp[8]) ? 11'b11110101110 : 11'b11111101100;
											assign node158 = (inp[8]) ? node162 : node159;
												assign node159 = (inp[11]) ? 11'b11100001101 : 11'b11111101111;
												assign node162 = (inp[11]) ? 11'b11111101111 : 11'b11010101111;
								assign node165 = (inp[8]) ? node187 : node166;
									assign node166 = (inp[11]) ? node176 : node167;
										assign node167 = (inp[5]) ? node173 : node168;
											assign node168 = (inp[6]) ? node170 : 11'b01000101111;
												assign node170 = (inp[9]) ? 11'b01010110100 : 11'b01010100110;
											assign node173 = (inp[6]) ? 11'b01000101111 : 11'b01100111110;
										assign node176 = (inp[5]) ? node184 : node177;
											assign node177 = (inp[6]) ? node181 : node178;
												assign node178 = (inp[9]) ? 11'b01010111111 : 11'b01000111111;
												assign node181 = (inp[9]) ? 11'b01001111111 : 11'b01001111101;
											assign node184 = (inp[6]) ? 11'b01010001101 : 11'b01000101100;
									assign node187 = (inp[5]) ? node203 : node188;
										assign node188 = (inp[6]) ? node196 : node189;
											assign node189 = (inp[11]) ? node193 : node190;
												assign node190 = (inp[9]) ? 11'b01110111111 : 11'b01100101111;
												assign node193 = (inp[9]) ? 11'b01101111101 : 11'b01011111101;
											assign node196 = (inp[11]) ? node200 : node197;
												assign node197 = (inp[9]) ? 11'b01111011110 : 11'b01101001100;
												assign node200 = (inp[9]) ? 11'b01100011100 : 11'b01010111110;
										assign node203 = (inp[6]) ? node211 : node204;
											assign node204 = (inp[9]) ? node208 : node205;
												assign node205 = (inp[11]) ? 11'b01001101110 : 11'b01111111110;
												assign node208 = (inp[11]) ? 11'b01111101110 : 11'b01101101100;
											assign node211 = (inp[11]) ? node215 : node212;
												assign node212 = (inp[9]) ? 11'b01100101101 : 11'b01101111101;
												assign node215 = (inp[9]) ? 11'b01111101111 : 11'b01011101101;
						assign node218 = (inp[9]) ? node328 : node219;
							assign node219 = (inp[5]) ? node269 : node220;
								assign node220 = (inp[10]) ? node244 : node221;
									assign node221 = (inp[3]) ? node231 : node222;
										assign node222 = (inp[6]) ? node228 : node223;
											assign node223 = (inp[8]) ? 11'b01110101101 : node224;
												assign node224 = (inp[11]) ? 11'b01011001111 : 11'b01001001111;
											assign node228 = (inp[8]) ? 11'b01100001110 : 11'b01000100110;
										assign node231 = (inp[11]) ? node237 : node232;
											assign node232 = (inp[6]) ? node234 : 11'b11001001111;
												assign node234 = (inp[8]) ? 11'b11000001100 : 11'b11011000110;
											assign node237 = (inp[8]) ? node241 : node238;
												assign node238 = (inp[6]) ? 11'b11100101111 : 11'b11111001111;
												assign node241 = (inp[6]) ? 11'b11011001110 : 11'b11010101101;
									assign node244 = (inp[3]) ? node258 : node245;
										assign node245 = (inp[8]) ? node251 : node246;
											assign node246 = (inp[11]) ? node248 : 11'b11000011111;
												assign node248 = (inp[6]) ? 11'b11110111111 : 11'b11110011111;
											assign node251 = (inp[6]) ? node255 : node252;
												assign node252 = (inp[11]) ? 11'b11111011101 : 11'b11101011111;
												assign node255 = (inp[11]) ? 11'b11101011110 : 11'b11110011100;
										assign node258 = (inp[11]) ? node262 : node259;
											assign node259 = (inp[6]) ? 11'b01110000010 : 11'b01100001011;
											assign node262 = (inp[8]) ? node266 : node263;
												assign node263 = (inp[6]) ? 11'b01100111001 : 11'b01110011011;
												assign node266 = (inp[6]) ? 11'b01110011010 : 11'b01101011011;
								assign node269 = (inp[10]) ? node299 : node270;
									assign node270 = (inp[3]) ? node286 : node271;
										assign node271 = (inp[11]) ? node279 : node272;
											assign node272 = (inp[8]) ? node276 : node273;
												assign node273 = (inp[6]) ? 11'b01010111111 : 11'b01011011110;
												assign node276 = (inp[6]) ? 11'b01111011101 : 11'b01111111100;
											assign node279 = (inp[8]) ? node283 : node280;
												assign node280 = (inp[6]) ? 11'b01001111100 : 11'b01000111100;
												assign node283 = (inp[6]) ? 11'b01101111101 : 11'b01101111100;
										assign node286 = (inp[6]) ? node292 : node287;
											assign node287 = (inp[8]) ? 11'b11010111100 : node288;
												assign node288 = (inp[11]) ? 11'b11101011100 : 11'b11111011110;
											assign node292 = (inp[11]) ? node296 : node293;
												assign node293 = (inp[8]) ? 11'b11011011101 : 11'b11100111101;
												assign node296 = (inp[8]) ? 11'b11100111101 : 11'b11111111100;
									assign node299 = (inp[3]) ? node315 : node300;
										assign node300 = (inp[6]) ? node308 : node301;
											assign node301 = (inp[8]) ? node305 : node302;
												assign node302 = (inp[11]) ? 11'b11001001100 : 11'b11010001110;
												assign node305 = (inp[11]) ? 11'b11110101100 : 11'b11000101100;
											assign node308 = (inp[11]) ? node312 : node309;
												assign node309 = (inp[8]) ? 11'b11000001111 : 11'b11001101101;
												assign node312 = (inp[8]) ? 11'b11110101101 : 11'b11010101110;
										assign node315 = (inp[11]) ? node323 : node316;
											assign node316 = (inp[6]) ? node320 : node317;
												assign node317 = (inp[8]) ? 11'b01001011000 : 11'b01010011010;
												assign node320 = (inp[8]) ? 11'b01000011011 : 11'b01011111001;
											assign node323 = (inp[6]) ? node325 : 11'b01110101000;
												assign node325 = (inp[8]) ? 11'b01111001011 : 11'b01100101010;
							assign node328 = (inp[5]) ? node388 : node329;
								assign node329 = (inp[6]) ? node361 : node330;
									assign node330 = (inp[11]) ? node346 : node331;
										assign node331 = (inp[3]) ? node339 : node332;
											assign node332 = (inp[10]) ? node336 : node333;
												assign node333 = (inp[8]) ? 11'b01110001111 : 11'b01101001111;
												assign node336 = (inp[8]) ? 11'b11001001001 : 11'b11100001011;
											assign node339 = (inp[10]) ? node343 : node340;
												assign node340 = (inp[8]) ? 11'b11011011011 : 11'b11101011011;
												assign node343 = (inp[8]) ? 11'b01101011001 : 11'b01100011011;
										assign node346 = (inp[10]) ? node354 : node347;
											assign node347 = (inp[3]) ? node351 : node348;
												assign node348 = (inp[8]) ? 11'b01000011111 : 11'b01011011111;
												assign node351 = (inp[8]) ? 11'b11010011011 : 11'b11011011011;
											assign node354 = (inp[8]) ? node358 : node355;
												assign node355 = (inp[3]) ? 11'b01110011011 : 11'b11110011011;
												assign node358 = (inp[3]) ? 11'b01111011011 : 11'b11111011011;
									assign node361 = (inp[8]) ? node373 : node362;
										assign node362 = (inp[11]) ? node370 : node363;
											assign node363 = (inp[3]) ? node367 : node364;
												assign node364 = (inp[10]) ? 11'b11101000000 : 11'b01100000100;
												assign node367 = (inp[10]) ? 11'b01111010000 : 11'b11110010000;
											assign node370 = (inp[3]) ? 11'b11011011001 : 11'b11100011011;
										assign node373 = (inp[10]) ? node381 : node374;
											assign node374 = (inp[3]) ? node378 : node375;
												assign node375 = (inp[11]) ? 11'b01010011100 : 11'b01111101100;
												assign node378 = (inp[11]) ? 11'b11000011000 : 11'b11010111010;
											assign node381 = (inp[3]) ? node385 : node382;
												assign node382 = (inp[11]) ? 11'b11111111001 : 11'b11000101010;
												assign node385 = (inp[11]) ? 11'b01111111011 : 11'b01111111010;
								assign node388 = (inp[6]) ? node418 : node389;
									assign node389 = (inp[3]) ? node405 : node390;
										assign node390 = (inp[10]) ? node398 : node391;
											assign node391 = (inp[11]) ? node395 : node392;
												assign node392 = (inp[8]) ? 11'b01101011100 : 11'b01111011110;
												assign node395 = (inp[8]) ? 11'b01101001100 : 11'b01010001100;
											assign node398 = (inp[8]) ? node402 : node399;
												assign node399 = (inp[11]) ? 11'b11011001000 : 11'b11001011000;
												assign node402 = (inp[11]) ? 11'b11110001000 : 11'b11110011000;
										assign node405 = (inp[10]) ? node413 : node406;
											assign node406 = (inp[11]) ? node410 : node407;
												assign node407 = (inp[8]) ? 11'b11110001000 : 11'b11001001000;
												assign node410 = (inp[8]) ? 11'b11101001000 : 11'b11111001000;
											assign node413 = (inp[11]) ? 11'b01110001000 : node414;
												assign node414 = (inp[8]) ? 11'b01101001010 : 11'b01100001000;
									assign node418 = (inp[8]) ? node430 : node419;
										assign node419 = (inp[11]) ? node425 : node420;
											assign node420 = (inp[3]) ? node422 : 11'b11001011011;
												assign node422 = (inp[10]) ? 11'b01111001011 : 11'b11010101011;
											assign node425 = (inp[3]) ? node427 : 11'b11001101000;
												assign node427 = (inp[10]) ? 11'b01110101000 : 11'b11101101000;
										assign node430 = (inp[3]) ? node436 : node431;
											assign node431 = (inp[10]) ? 11'b11101011001 : node432;
												assign node432 = (inp[11]) ? 11'b01101001111 : 11'b01111011111;
											assign node436 = (inp[10]) ? 11'b01110001001 : 11'b11101001001;
					assign node439 = (inp[3]) ? node673 : node440;
						assign node440 = (inp[4]) ? node558 : node441;
							assign node441 = (inp[11]) ? node501 : node442;
								assign node442 = (inp[6]) ? node474 : node443;
									assign node443 = (inp[5]) ? node459 : node444;
										assign node444 = (inp[8]) ? node452 : node445;
											assign node445 = (inp[10]) ? node449 : node446;
												assign node446 = (inp[9]) ? 11'b01001101101 : 11'b01001101001;
												assign node449 = (inp[9]) ? 11'b01000111001 : 11'b01000101101;
											assign node452 = (inp[10]) ? node456 : node453;
												assign node453 = (inp[9]) ? 11'b01110101101 : 11'b01100001000;
												assign node456 = (inp[9]) ? 11'b01111111001 : 11'b01101101101;
										assign node459 = (inp[9]) ? node467 : node460;
											assign node460 = (inp[10]) ? node464 : node461;
												assign node461 = (inp[8]) ? 11'b01100001001 : 11'b01001101000;
												assign node464 = (inp[8]) ? 11'b01011101100 : 11'b01100101100;
											assign node467 = (inp[10]) ? node471 : node468;
												assign node468 = (inp[8]) ? 11'b01110101100 : 11'b01001101100;
												assign node471 = (inp[8]) ? 11'b01001111010 : 11'b01100111000;
									assign node474 = (inp[5]) ? node490 : node475;
										assign node475 = (inp[8]) ? node483 : node476;
											assign node476 = (inp[10]) ? node480 : node477;
												assign node477 = (inp[9]) ? 11'b01011100110 : 11'b01011100000;
												assign node480 = (inp[9]) ? 11'b01010110010 : 11'b01010100100;
											assign node483 = (inp[10]) ? node487 : node484;
												assign node484 = (inp[9]) ? 11'b01100001110 : 11'b01110101000;
												assign node487 = (inp[9]) ? 11'b01101011000 : 11'b01111001100;
										assign node490 = (inp[8]) ? node496 : node491;
											assign node491 = (inp[10]) ? 11'b01110001111 : node492;
												assign node492 = (inp[9]) ? 11'b01011101111 : 11'b01011001001;
											assign node496 = (inp[10]) ? node498 : 11'b01101101101;
												assign node498 = (inp[9]) ? 11'b01010111001 : 11'b01001101111;
								assign node501 = (inp[10]) ? node531 : node502;
									assign node502 = (inp[9]) ? node516 : node503;
										assign node503 = (inp[6]) ? node509 : node504;
											assign node504 = (inp[8]) ? node506 : 11'b01001111010;
												assign node506 = (inp[5]) ? 11'b01101011000 : 11'b01100011011;
											assign node509 = (inp[8]) ? node513 : node510;
												assign node510 = (inp[5]) ? 11'b01010011011 : 11'b01010010000;
												assign node513 = (inp[5]) ? 11'b01110011001 : 11'b01111111010;
										assign node516 = (inp[8]) ? node524 : node517;
											assign node517 = (inp[5]) ? node521 : node518;
												assign node518 = (inp[6]) ? 11'b01110111111 : 11'b01101111101;
												assign node521 = (inp[6]) ? 11'b01101011101 : 11'b01111111110;
											assign node524 = (inp[6]) ? node528 : node525;
												assign node525 = (inp[5]) ? 11'b01001111100 : 11'b01000111111;
												assign node528 = (inp[5]) ? 11'b01010111111 : 11'b01011011100;
									assign node531 = (inp[9]) ? node547 : node532;
										assign node532 = (inp[8]) ? node540 : node533;
											assign node533 = (inp[6]) ? node537 : node534;
												assign node534 = (inp[5]) ? 11'b01010111110 : 11'b01000111101;
												assign node537 = (inp[5]) ? 11'b01000011101 : 11'b01011111101;
											assign node540 = (inp[6]) ? node544 : node541;
												assign node541 = (inp[5]) ? 11'b01110011100 : 11'b01111111111;
												assign node544 = (inp[5]) ? 11'b01101111111 : 11'b01100111100;
										assign node547 = (inp[6]) ? node551 : node548;
											assign node548 = (inp[5]) ? 11'b01110101010 : 11'b01101101011;
											assign node551 = (inp[8]) ? node555 : node552;
												assign node552 = (inp[5]) ? 11'b01100001011 : 11'b01000101001;
												assign node555 = (inp[5]) ? 11'b01001101001 : 11'b01110001010;
							assign node558 = (inp[5]) ? node616 : node559;
								assign node559 = (inp[6]) ? node589 : node560;
									assign node560 = (inp[11]) ? node576 : node561;
										assign node561 = (inp[10]) ? node569 : node562;
											assign node562 = (inp[9]) ? node566 : node563;
												assign node563 = (inp[8]) ? 11'b01100101001 : 11'b01001001001;
												assign node566 = (inp[8]) ? 11'b01010011101 : 11'b01101011101;
											assign node569 = (inp[9]) ? node573 : node570;
												assign node570 = (inp[8]) ? 11'b01101011101 : 11'b01000011101;
												assign node573 = (inp[8]) ? 11'b01001011011 : 11'b01100011001;
										assign node576 = (inp[8]) ? node584 : node577;
											assign node577 = (inp[10]) ? node581 : node578;
												assign node578 = (inp[9]) ? 11'b01011001101 : 11'b01011011001;
												assign node581 = (inp[9]) ? 11'b01110001001 : 11'b01110001101;
											assign node584 = (inp[10]) ? 11'b01001001101 : node585;
												assign node585 = (inp[9]) ? 11'b01100001101 : 11'b01110111011;
									assign node589 = (inp[11]) ? node601 : node590;
										assign node590 = (inp[8]) ? node594 : node591;
											assign node591 = (inp[10]) ? 11'b01111010010 : 11'b01110010110;
											assign node594 = (inp[9]) ? node598 : node595;
												assign node595 = (inp[10]) ? 11'b01111111110 : 11'b01110001000;
												assign node598 = (inp[10]) ? 11'b01010111000 : 11'b01001111100;
										assign node601 = (inp[8]) ? node609 : node602;
											assign node602 = (inp[10]) ? node606 : node603;
												assign node603 = (inp[9]) ? 11'b01001001111 : 11'b01001111001;
												assign node606 = (inp[9]) ? 11'b01100001001 : 11'b01100101111;
											assign node609 = (inp[10]) ? node613 : node610;
												assign node610 = (inp[9]) ? 11'b01110001110 : 11'b01100011000;
												assign node613 = (inp[9]) ? 11'b01001101001 : 11'b01011001100;
								assign node616 = (inp[6]) ? node644 : node617;
									assign node617 = (inp[8]) ? node631 : node618;
										assign node618 = (inp[10]) ? node626 : node619;
											assign node619 = (inp[11]) ? node623 : node620;
												assign node620 = (inp[9]) ? 11'b01111011100 : 11'b01111001000;
												assign node623 = (inp[9]) ? 11'b01111001110 : 11'b01101011010;
											assign node626 = (inp[9]) ? node628 : 11'b01010011100;
												assign node628 = (inp[11]) ? 11'b01110001010 : 11'b01100011010;
										assign node631 = (inp[9]) ? node639 : node632;
											assign node632 = (inp[10]) ? node636 : node633;
												assign node633 = (inp[11]) ? 11'b01001111010 : 11'b01010101010;
												assign node636 = (inp[11]) ? 11'b01010101110 : 11'b01101011110;
											assign node639 = (inp[10]) ? 11'b01000011000 : node640;
												assign node640 = (inp[11]) ? 11'b01001001110 : 11'b01010011110;
									assign node644 = (inp[8]) ? node660 : node645;
										assign node645 = (inp[11]) ? node653 : node646;
											assign node646 = (inp[9]) ? node650 : node647;
												assign node647 = (inp[10]) ? 11'b01001111111 : 11'b01100101011;
												assign node650 = (inp[10]) ? 11'b01111011001 : 11'b01100111101;
											assign node653 = (inp[9]) ? node657 : node654;
												assign node654 = (inp[10]) ? 11'b01110101100 : 11'b01111111010;
												assign node657 = (inp[10]) ? 11'b01100101010 : 11'b01101101110;
										assign node660 = (inp[11]) ? node668 : node661;
											assign node661 = (inp[10]) ? node665 : node662;
												assign node662 = (inp[9]) ? 11'b01001011111 : 11'b01001001011;
												assign node665 = (inp[9]) ? 11'b01010011011 : 11'b01110011101;
											assign node668 = (inp[9]) ? 11'b01011001101 : node669;
												assign node669 = (inp[10]) ? 11'b01000101101 : 11'b01010111011;
						assign node673 = (inp[10]) ? node773 : node674;
							assign node674 = (inp[8]) ? node726 : node675;
								assign node675 = (inp[5]) ? node697 : node676;
									assign node676 = (inp[6]) ? node688 : node677;
										assign node677 = (inp[4]) ? node683 : node678;
											assign node678 = (inp[9]) ? node680 : 11'b01001101001;
												assign node680 = (inp[11]) ? 11'b01101111001 : 11'b01001111001;
											assign node683 = (inp[9]) ? 11'b01101001001 : node684;
												assign node684 = (inp[11]) ? 11'b01111011001 : 11'b01001011001;
										assign node688 = (inp[11]) ? node694 : node689;
											assign node689 = (inp[9]) ? node691 : 11'b01001010000;
												assign node691 = (inp[4]) ? 11'b01101000010 : 11'b01001110010;
											assign node694 = (inp[4]) ? 11'b01110111001 : 11'b01000000000;
									assign node697 = (inp[11]) ? node713 : node698;
										assign node698 = (inp[6]) ? node706 : node699;
											assign node699 = (inp[4]) ? node703 : node700;
												assign node700 = (inp[9]) ? 11'b01101111000 : 11'b01101101000;
												assign node703 = (inp[9]) ? 11'b01001001010 : 11'b01111011000;
											assign node706 = (inp[9]) ? node710 : node707;
												assign node707 = (inp[4]) ? 11'b01111111011 : 11'b01101001011;
												assign node710 = (inp[4]) ? 11'b01000101001 : 11'b01101111001;
										assign node713 = (inp[9]) ? node719 : node714;
											assign node714 = (inp[4]) ? node716 : 11'b01101101010;
												assign node716 = (inp[6]) ? 11'b01001111000 : 11'b01001011010;
											assign node719 = (inp[4]) ? node723 : node720;
												assign node720 = (inp[6]) ? 11'b01010011001 : 11'b01011111010;
												assign node723 = (inp[6]) ? 11'b01011101010 : 11'b01011001010;
								assign node726 = (inp[5]) ? node750 : node727;
									assign node727 = (inp[6]) ? node741 : node728;
										assign node728 = (inp[11]) ? node734 : node729;
											assign node729 = (inp[4]) ? 11'b01001011001 : node730;
												assign node730 = (inp[9]) ? 11'b01011111001 : 11'b01001101001;
											assign node734 = (inp[4]) ? node738 : node735;
												assign node735 = (inp[9]) ? 11'b01101111011 : 11'b01011101011;
												assign node738 = (inp[9]) ? 11'b01110001001 : 11'b01111011011;
										assign node741 = (inp[4]) ? 11'b01110101000 : node742;
											assign node742 = (inp[9]) ? node746 : node743;
												assign node743 = (inp[11]) ? 11'b01010101010 : 11'b01001001000;
												assign node746 = (inp[11]) ? 11'b01101011010 : 11'b01011011010;
									assign node750 = (inp[4]) ? node762 : node751;
										assign node751 = (inp[11]) ? node757 : node752;
											assign node752 = (inp[9]) ? 11'b01100111001 : node753;
												assign node753 = (inp[6]) ? 11'b01100101011 : 11'b01100001001;
											assign node757 = (inp[9]) ? node759 : 11'b01110001000;
												assign node759 = (inp[6]) ? 11'b01010111001 : 11'b01010111000;
										assign node762 = (inp[9]) ? node770 : node763;
											assign node763 = (inp[11]) ? node767 : node764;
												assign node764 = (inp[6]) ? 11'b01110011011 : 11'b01110111010;
												assign node767 = (inp[6]) ? 11'b01010111011 : 11'b01010111010;
											assign node770 = (inp[6]) ? 11'b01010001011 : 11'b01010001010;
							assign node773 = (inp[4]) ? node827 : node774;
								assign node774 = (inp[11]) ? node800 : node775;
									assign node775 = (inp[8]) ? node787 : node776;
										assign node776 = (inp[5]) ? node782 : node777;
											assign node777 = (inp[6]) ? node779 : 11'b01000101001;
												assign node779 = (inp[9]) ? 11'b01000100000 : 11'b01000100010;
											assign node782 = (inp[9]) ? node784 : 11'b01000001011;
												assign node784 = (inp[6]) ? 11'b01010101001 : 11'b01010101000;
										assign node787 = (inp[5]) ? node793 : node788;
											assign node788 = (inp[6]) ? node790 : 11'b01000101001;
												assign node790 = (inp[9]) ? 11'b01001001000 : 11'b01010001010;
											assign node793 = (inp[6]) ? node797 : node794;
												assign node794 = (inp[9]) ? 11'b01011101010 : 11'b01011101000;
												assign node797 = (inp[9]) ? 11'b01011001011 : 11'b01011101011;
									assign node800 = (inp[9]) ? node814 : node801;
										assign node801 = (inp[5]) ? node809 : node802;
											assign node802 = (inp[8]) ? node806 : node803;
												assign node803 = (inp[6]) ? 11'b01101101011 : 11'b01100101001;
												assign node806 = (inp[6]) ? 11'b01110101000 : 11'b01110101011;
											assign node809 = (inp[6]) ? 11'b01111001001 : node810;
												assign node810 = (inp[8]) ? 11'b01101101000 : 11'b01110101010;
										assign node814 = (inp[5]) ? node822 : node815;
											assign node815 = (inp[8]) ? node819 : node816;
												assign node816 = (inp[6]) ? 11'b01011101001 : 11'b01010101001;
												assign node819 = (inp[6]) ? 11'b01010001010 : 11'b01010101011;
											assign node822 = (inp[6]) ? 11'b01001101010 : node823;
												assign node823 = (inp[8]) ? 11'b01001101010 : 11'b01000101010;
								assign node827 = (inp[9]) ? node851 : node828;
									assign node828 = (inp[11]) ? node838 : node829;
										assign node829 = (inp[8]) ? node835 : node830;
											assign node830 = (inp[5]) ? 11'b01110101011 : node831;
												assign node831 = (inp[6]) ? 11'b01100000010 : 11'b01100001001;
											assign node835 = (inp[5]) ? 11'b01100001001 : 11'b01110001001;
										assign node838 = (inp[8]) ? node844 : node839;
											assign node839 = (inp[5]) ? node841 : 11'b01011001011;
												assign node841 = (inp[6]) ? 11'b01010101000 : 11'b01010001010;
											assign node844 = (inp[6]) ? node848 : node845;
												assign node845 = (inp[5]) ? 11'b01001001010 : 11'b01001001001;
												assign node848 = (inp[5]) ? 11'b01001001001 : 11'b01000001010;
									assign node851 = (inp[11]) ? node863 : node852;
										assign node852 = (inp[8]) ? node858 : node853;
											assign node853 = (inp[6]) ? 11'b01001000000 : node854;
												assign node854 = (inp[5]) ? 11'b01000001010 : 11'b01000001001;
											assign node858 = (inp[5]) ? node860 : 11'b01001101010;
												assign node860 = (inp[6]) ? 11'b01000001001 : 11'b01001001000;
										assign node863 = (inp[5]) ? node867 : node864;
											assign node864 = (inp[8]) ? 11'b01001101001 : 11'b01000001001;
											assign node867 = (inp[8]) ? node871 : node868;
												assign node868 = (inp[6]) ? 11'b01000101000 : 11'b01000001000;
												assign node871 = (inp[6]) ? 11'b01000001001 : 11'b01000001000;
				assign node874 = (inp[0]) ? node1300 : node875;
					assign node875 = (inp[8]) ? node1079 : node876;
						assign node876 = (inp[6]) ? node974 : node877;
							assign node877 = (inp[4]) ? node927 : node878;
								assign node878 = (inp[9]) ? node906 : node879;
									assign node879 = (inp[5]) ? node895 : node880;
										assign node880 = (inp[11]) ? node888 : node881;
											assign node881 = (inp[10]) ? node885 : node882;
												assign node882 = (inp[3]) ? 11'b11101001010 : 11'b01101001010;
												assign node885 = (inp[3]) ? 11'b01110001110 : 11'b11110001010;
											assign node888 = (inp[3]) ? node892 : node889;
												assign node889 = (inp[10]) ? 11'b11111000011 : 11'b01100000011;
												assign node892 = (inp[10]) ? 11'b01100010111 : 11'b11111010011;
										assign node895 = (inp[11]) ? node899 : node896;
											assign node896 = (inp[3]) ? 11'b11100010011 : 11'b11011010011;
											assign node899 = (inp[10]) ? node903 : node900;
												assign node900 = (inp[3]) ? 11'b11011000000 : 11'b01101010000;
												assign node903 = (inp[3]) ? 11'b01100000100 : 11'b11000010000;
									assign node906 = (inp[5]) ? node916 : node907;
										assign node907 = (inp[10]) ? node911 : node908;
											assign node908 = (inp[11]) ? 11'b11011100111 : 11'b11101100111;
											assign node911 = (inp[11]) ? node913 : 11'b11110110111;
												assign node913 = (inp[3]) ? 11'b01101110101 : 11'b11001110101;
										assign node916 = (inp[3]) ? node922 : node917;
											assign node917 = (inp[10]) ? node919 : 11'b01011000000;
												assign node919 = (inp[11]) ? 11'b11010000110 : 11'b11000000101;
											assign node922 = (inp[10]) ? 11'b01101100100 : node923;
												assign node923 = (inp[11]) ? 11'b11101010110 : 11'b11110010101;
								assign node927 = (inp[5]) ? node949 : node928;
									assign node928 = (inp[9]) ? node940 : node929;
										assign node929 = (inp[3]) ? node935 : node930;
											assign node930 = (inp[10]) ? node932 : 11'b01110100101;
												assign node932 = (inp[11]) ? 11'b11001110101 : 11'b11111110101;
											assign node935 = (inp[10]) ? 11'b01000100001 : node936;
												assign node936 = (inp[11]) ? 11'b11000100101 : 11'b11101100101;
										assign node940 = (inp[10]) ? node946 : node941;
											assign node941 = (inp[3]) ? node943 : 11'b01000100101;
												assign node943 = (inp[11]) ? 11'b11100110011 : 11'b11011010001;
											assign node946 = (inp[3]) ? 11'b01011010011 : 11'b11011010011;
									assign node949 = (inp[10]) ? node961 : node950;
										assign node950 = (inp[3]) ? node954 : node951;
											assign node951 = (inp[9]) ? 11'b01001110110 : 11'b01111110100;
											assign node954 = (inp[9]) ? node958 : node955;
												assign node955 = (inp[11]) ? 11'b11011110110 : 11'b11000110110;
												assign node958 = (inp[11]) ? 11'b11001100000 : 11'b11100100010;
										assign node961 = (inp[3]) ? node967 : node962;
											assign node962 = (inp[9]) ? node964 : 11'b11110100110;
												assign node964 = (inp[11]) ? 11'b11101100000 : 11'b11110110010;
											assign node967 = (inp[9]) ? node971 : node968;
												assign node968 = (inp[11]) ? 11'b01000100000 : 11'b01111110010;
												assign node971 = (inp[11]) ? 11'b01010100000 : 11'b01000100000;
							assign node974 = (inp[5]) ? node1030 : node975;
								assign node975 = (inp[4]) ? node1005 : node976;
									assign node976 = (inp[11]) ? node990 : node977;
										assign node977 = (inp[10]) ? node983 : node978;
											assign node978 = (inp[3]) ? 11'b11101101110 : node979;
												assign node979 = (inp[9]) ? 11'b01100001001 : 11'b01101001011;
											assign node983 = (inp[9]) ? node987 : node984;
												assign node984 = (inp[3]) ? 11'b01110001101 : 11'b11110001011;
												assign node987 = (inp[3]) ? 11'b01110111110 : 11'b11111111110;
										assign node990 = (inp[10]) ? node998 : node991;
											assign node991 = (inp[3]) ? node995 : node992;
												assign node992 = (inp[9]) ? 11'b01011011000 : 11'b01111001010;
												assign node995 = (inp[9]) ? 11'b11011001110 : 11'b11100011010;
											assign node998 = (inp[3]) ? node1002 : node999;
												assign node999 = (inp[9]) ? 11'b11000011110 : 11'b11100001000;
												assign node1002 = (inp[9]) ? 11'b01100011100 : 11'b01110011100;
									assign node1005 = (inp[10]) ? node1019 : node1006;
										assign node1006 = (inp[3]) ? node1014 : node1007;
											assign node1007 = (inp[9]) ? node1011 : node1008;
												assign node1008 = (inp[11]) ? 11'b01110001100 : 11'b01100101100;
												assign node1011 = (inp[11]) ? 11'b01100111100 : 11'b01010101110;
											assign node1014 = (inp[9]) ? node1016 : 11'b11011101100;
												assign node1016 = (inp[11]) ? 11'b11110111000 : 11'b11000111000;
										assign node1019 = (inp[3]) ? node1025 : node1020;
											assign node1020 = (inp[11]) ? node1022 : 11'b11000101000;
												assign node1022 = (inp[9]) ? 11'b11011111000 : 11'b11011111110;
											assign node1025 = (inp[9]) ? node1027 : 11'b01000111010;
												assign node1027 = (inp[11]) ? 11'b01011111010 : 11'b01011011000;
								assign node1030 = (inp[11]) ? node1058 : node1031;
									assign node1031 = (inp[4]) ? node1047 : node1032;
										assign node1032 = (inp[10]) ? node1040 : node1033;
											assign node1033 = (inp[9]) ? node1037 : node1034;
												assign node1034 = (inp[3]) ? 11'b11100111000 : 11'b01100111010;
												assign node1037 = (inp[3]) ? 11'b11100011110 : 11'b01111011010;
											assign node1040 = (inp[9]) ? node1044 : node1041;
												assign node1041 = (inp[3]) ? 11'b01011011100 : 11'b11000111000;
												assign node1044 = (inp[3]) ? 11'b01100001100 : 11'b11000001100;
										assign node1047 = (inp[9]) ? node1051 : node1048;
											assign node1048 = (inp[3]) ? 11'b01100011000 : 11'b11110001110;
											assign node1051 = (inp[3]) ? node1055 : node1052;
												assign node1052 = (inp[10]) ? 11'b11111110011 : 11'b01000011100;
												assign node1055 = (inp[10]) ? 11'b01010100011 : 11'b11101100011;
									assign node1058 = (inp[4]) ? node1068 : node1059;
										assign node1059 = (inp[10]) ? node1063 : node1060;
											assign node1060 = (inp[3]) ? 11'b11010100001 : 11'b01110110001;
											assign node1063 = (inp[9]) ? 11'b11010100101 : node1064;
												assign node1064 = (inp[3]) ? 11'b01101100111 : 11'b11001110011;
										assign node1068 = (inp[3]) ? node1072 : node1069;
											assign node1069 = (inp[10]) ? 11'b11111000001 : 11'b01111000111;
											assign node1072 = (inp[10]) ? node1076 : node1073;
												assign node1073 = (inp[9]) ? 11'b11011000011 : 11'b11001010101;
												assign node1076 = (inp[9]) ? 11'b01010000001 : 11'b01000000011;
						assign node1079 = (inp[5]) ? node1195 : node1080;
							assign node1080 = (inp[9]) ? node1138 : node1081;
								assign node1081 = (inp[11]) ? node1109 : node1082;
									assign node1082 = (inp[6]) ? node1094 : node1083;
										assign node1083 = (inp[4]) ? node1091 : node1084;
											assign node1084 = (inp[3]) ? node1088 : node1085;
												assign node1085 = (inp[10]) ? 11'b11111000010 : 11'b01100100010;
												assign node1088 = (inp[10]) ? 11'b01000000110 : 11'b11011000010;
											assign node1091 = (inp[3]) ? 11'b01101100011 : 11'b01000000100;
										assign node1094 = (inp[4]) ? node1102 : node1095;
											assign node1095 = (inp[10]) ? node1099 : node1096;
												assign node1096 = (inp[3]) ? 11'b11001100011 : 11'b01100000011;
												assign node1099 = (inp[3]) ? 11'b01001100101 : 11'b11101100001;
											assign node1102 = (inp[3]) ? node1106 : node1103;
												assign node1103 = (inp[10]) ? 11'b11000110111 : 11'b01011100101;
												assign node1106 = (inp[10]) ? 11'b01100100001 : 11'b11100100111;
									assign node1109 = (inp[4]) ? node1125 : node1110;
										assign node1110 = (inp[3]) ? node1118 : node1111;
											assign node1111 = (inp[6]) ? node1115 : node1112;
												assign node1112 = (inp[10]) ? 11'b11000100001 : 11'b01101100001;
												assign node1115 = (inp[10]) ? 11'b11011000011 : 11'b01110000001;
											assign node1118 = (inp[10]) ? node1122 : node1119;
												assign node1119 = (inp[6]) ? 11'b11011010001 : 11'b11010110001;
												assign node1122 = (inp[6]) ? 11'b01100010111 : 11'b01111010101;
										assign node1125 = (inp[6]) ? node1133 : node1126;
											assign node1126 = (inp[10]) ? node1130 : node1127;
												assign node1127 = (inp[3]) ? 11'b11101000101 : 11'b01011000111;
												assign node1130 = (inp[3]) ? 11'b01000010001 : 11'b11010010101;
											assign node1133 = (inp[10]) ? 11'b11010110100 : node1134;
												assign node1134 = (inp[3]) ? 11'b11110100100 : 11'b01001100100;
								assign node1138 = (inp[4]) ? node1168 : node1139;
									assign node1139 = (inp[10]) ? node1153 : node1140;
										assign node1140 = (inp[3]) ? node1148 : node1141;
											assign node1141 = (inp[11]) ? node1145 : node1142;
												assign node1142 = (inp[6]) ? 11'b01110100001 : 11'b01110000010;
												assign node1145 = (inp[6]) ? 11'b01000010001 : 11'b01001010011;
											assign node1148 = (inp[11]) ? node1150 : 11'b11000000100;
												assign node1150 = (inp[6]) ? 11'b11000000101 : 11'b11010000111;
										assign node1153 = (inp[3]) ? node1161 : node1154;
											assign node1154 = (inp[6]) ? node1158 : node1155;
												assign node1155 = (inp[11]) ? 11'b11110010111 : 11'b11101010100;
												assign node1158 = (inp[11]) ? 11'b11101110110 : 11'b11111110111;
											assign node1161 = (inp[11]) ? node1165 : node1162;
												assign node1162 = (inp[6]) ? 11'b01011110101 : 11'b01011010100;
												assign node1165 = (inp[6]) ? 11'b01001110110 : 11'b01001010111;
									assign node1168 = (inp[11]) ? node1184 : node1169;
										assign node1169 = (inp[3]) ? node1177 : node1170;
											assign node1170 = (inp[10]) ? node1174 : node1171;
												assign node1171 = (inp[6]) ? 11'b01001000101 : 11'b01010100111;
												assign node1174 = (inp[6]) ? 11'b11110000011 : 11'b11111100011;
											assign node1177 = (inp[6]) ? node1181 : node1178;
												assign node1178 = (inp[10]) ? 11'b01001110001 : 11'b11100110011;
												assign node1181 = (inp[10]) ? 11'b01010010011 : 11'b11111010001;
										assign node1184 = (inp[10]) ? node1192 : node1185;
											assign node1185 = (inp[3]) ? node1189 : node1186;
												assign node1186 = (inp[6]) ? 11'b01111110110 : 11'b01101110101;
												assign node1189 = (inp[6]) ? 11'b11111110000 : 11'b11111110001;
											assign node1192 = (inp[6]) ? 11'b11010110000 : 11'b11000110011;
							assign node1195 = (inp[11]) ? node1245 : node1196;
								assign node1196 = (inp[6]) ? node1220 : node1197;
									assign node1197 = (inp[10]) ? node1205 : node1198;
										assign node1198 = (inp[3]) ? node1202 : node1199;
											assign node1199 = (inp[4]) ? 11'b01010010101 : 11'b01101110011;
											assign node1202 = (inp[9]) ? 11'b11101010101 : 11'b11101010111;
										assign node1205 = (inp[3]) ? node1213 : node1206;
											assign node1206 = (inp[4]) ? node1210 : node1207;
												assign node1207 = (inp[9]) ? 11'b11111000101 : 11'b11001110001;
												assign node1210 = (inp[9]) ? 11'b11011110000 : 11'b11111000111;
											assign node1213 = (inp[9]) ? node1217 : node1214;
												assign node1214 = (inp[4]) ? 11'b01101010001 : 11'b01010110101;
												assign node1217 = (inp[4]) ? 11'b01001100010 : 11'b01000000111;
									assign node1220 = (inp[4]) ? node1234 : node1221;
										assign node1221 = (inp[10]) ? node1227 : node1222;
											assign node1222 = (inp[3]) ? node1224 : 11'b01100010010;
												assign node1224 = (inp[9]) ? 11'b11100010100 : 11'b11101010000;
											assign node1227 = (inp[3]) ? node1231 : node1228;
												assign node1228 = (inp[9]) ? 11'b11101000100 : 11'b11001010000;
												assign node1231 = (inp[9]) ? 11'b01001000110 : 11'b01000010110;
										assign node1234 = (inp[9]) ? node1240 : node1235;
											assign node1235 = (inp[3]) ? node1237 : 11'b11110000100;
												assign node1237 = (inp[10]) ? 11'b01111110000 : 11'b11110010110;
											assign node1240 = (inp[10]) ? node1242 : 11'b11010100010;
												assign node1242 = (inp[3]) ? 11'b01010100000 : 11'b11010110000;
								assign node1245 = (inp[4]) ? node1273 : node1246;
									assign node1246 = (inp[9]) ? node1260 : node1247;
										assign node1247 = (inp[3]) ? node1253 : node1248;
											assign node1248 = (inp[10]) ? 11'b11101110010 : node1249;
												assign node1249 = (inp[6]) ? 11'b01111110010 : 11'b01100110010;
											assign node1253 = (inp[10]) ? node1257 : node1254;
												assign node1254 = (inp[6]) ? 11'b11111100010 : 11'b11110100010;
												assign node1257 = (inp[6]) ? 11'b01110100100 : 11'b01111100110;
										assign node1260 = (inp[3]) ? node1268 : node1261;
											assign node1261 = (inp[10]) ? node1265 : node1262;
												assign node1262 = (inp[6]) ? 11'b01110100010 : 11'b01101100000;
												assign node1265 = (inp[6]) ? 11'b11011000100 : 11'b11000100100;
											assign node1268 = (inp[10]) ? 11'b01011000100 : node1269;
												assign node1269 = (inp[6]) ? 11'b11011010110 : 11'b11010110100;
									assign node1273 = (inp[10]) ? node1287 : node1274;
										assign node1274 = (inp[3]) ? node1282 : node1275;
											assign node1275 = (inp[6]) ? node1279 : node1276;
												assign node1276 = (inp[9]) ? 11'b01001000100 : 11'b01001010110;
												assign node1279 = (inp[9]) ? 11'b01011000110 : 11'b01010010110;
											assign node1282 = (inp[9]) ? node1284 : 11'b11010010110;
												assign node1284 = (inp[6]) ? 11'b11010000010 : 11'b11011000000;
										assign node1287 = (inp[3]) ? node1295 : node1288;
											assign node1288 = (inp[6]) ? node1292 : node1289;
												assign node1289 = (inp[9]) ? 11'b11000000000 : 11'b11000000110;
												assign node1292 = (inp[9]) ? 11'b11010000000 : 11'b11010000100;
											assign node1295 = (inp[9]) ? 11'b01010000000 : node1296;
												assign node1296 = (inp[6]) ? 11'b01011000000 : 11'b01011000010;
					assign node1300 = (inp[3]) ? node1530 : node1301;
						assign node1301 = (inp[6]) ? node1415 : node1302;
							assign node1302 = (inp[5]) ? node1360 : node1303;
								assign node1303 = (inp[4]) ? node1331 : node1304;
									assign node1304 = (inp[11]) ? node1318 : node1305;
										assign node1305 = (inp[8]) ? node1311 : node1306;
											assign node1306 = (inp[9]) ? 11'b01010110001 : node1307;
												assign node1307 = (inp[10]) ? 11'b01010001100 : 11'b01001001000;
											assign node1311 = (inp[10]) ? node1315 : node1312;
												assign node1312 = (inp[9]) ? 11'b01110000100 : 11'b01100100000;
												assign node1315 = (inp[9]) ? 11'b01111010010 : 11'b01101000100;
										assign node1318 = (inp[10]) ? node1326 : node1319;
											assign node1319 = (inp[9]) ? node1323 : node1320;
												assign node1320 = (inp[8]) ? 11'b01110110011 : 11'b01010010001;
												assign node1323 = (inp[8]) ? 11'b01001010101 : 11'b01110010101;
											assign node1326 = (inp[9]) ? node1328 : 11'b01101010111;
												assign node1328 = (inp[8]) ? 11'b01100000001 : 11'b01001100011;
									assign node1331 = (inp[11]) ? node1347 : node1332;
										assign node1332 = (inp[10]) ? node1340 : node1333;
											assign node1333 = (inp[9]) ? node1337 : node1334;
												assign node1334 = (inp[8]) ? 11'b01100000010 : 11'b01001100011;
												assign node1337 = (inp[8]) ? 11'b01000110101 : 11'b01101010111;
											assign node1340 = (inp[8]) ? node1344 : node1341;
												assign node1341 = (inp[9]) ? 11'b01110010011 : 11'b01010110111;
												assign node1344 = (inp[9]) ? 11'b01011110001 : 11'b01101110101;
										assign node1347 = (inp[9]) ? node1353 : node1348;
											assign node1348 = (inp[10]) ? 11'b01101100111 : node1349;
												assign node1349 = (inp[8]) ? 11'b01111010001 : 11'b01010110011;
											assign node1353 = (inp[10]) ? node1357 : node1354;
												assign node1354 = (inp[8]) ? 11'b01111100111 : 11'b01000100101;
												assign node1357 = (inp[8]) ? 11'b01010100001 : 11'b01111000001;
								assign node1360 = (inp[11]) ? node1384 : node1361;
									assign node1361 = (inp[4]) ? node1373 : node1362;
										assign node1362 = (inp[9]) ? node1368 : node1363;
											assign node1363 = (inp[10]) ? 11'b01111000101 : node1364;
												assign node1364 = (inp[8]) ? 11'b01101100001 : 11'b01000000001;
											assign node1368 = (inp[10]) ? 11'b01101110010 : node1369;
												assign node1369 = (inp[8]) ? 11'b01101000111 : 11'b01010000111;
										assign node1373 = (inp[8]) ? node1381 : node1374;
											assign node1374 = (inp[9]) ? node1378 : node1375;
												assign node1375 = (inp[10]) ? 11'b01010110100 : 11'b01110100010;
												assign node1378 = (inp[10]) ? 11'b01110110000 : 11'b01101110100;
											assign node1381 = (inp[10]) ? 11'b01011110010 : 11'b01000000001;
									assign node1384 = (inp[9]) ? node1400 : node1385;
										assign node1385 = (inp[10]) ? node1393 : node1386;
											assign node1386 = (inp[4]) ? node1390 : node1387;
												assign node1387 = (inp[8]) ? 11'b01110110000 : 11'b01011010010;
												assign node1390 = (inp[8]) ? 11'b01011010000 : 11'b01101110000;
											assign node1393 = (inp[8]) ? node1397 : node1394;
												assign node1394 = (inp[4]) ? 11'b01100100110 : 11'b01000010110;
												assign node1397 = (inp[4]) ? 11'b01010000100 : 11'b01111110100;
										assign node1400 = (inp[10]) ? node1408 : node1401;
											assign node1401 = (inp[4]) ? node1405 : node1402;
												assign node1402 = (inp[8]) ? 11'b01010110110 : 11'b01111010110;
												assign node1405 = (inp[8]) ? 11'b01011000110 : 11'b01111100110;
											assign node1408 = (inp[8]) ? node1412 : node1409;
												assign node1409 = (inp[4]) ? 11'b01110100010 : 11'b01110000000;
												assign node1412 = (inp[4]) ? 11'b01010000010 : 11'b01011000010;
							assign node1415 = (inp[8]) ? node1473 : node1416;
								assign node1416 = (inp[5]) ? node1448 : node1417;
									assign node1417 = (inp[4]) ? node1433 : node1418;
										assign node1418 = (inp[11]) ? node1426 : node1419;
											assign node1419 = (inp[9]) ? node1423 : node1420;
												assign node1420 = (inp[10]) ? 11'b01000001111 : 11'b01011001001;
												assign node1423 = (inp[10]) ? 11'b01001111000 : 11'b01011101110;
											assign node1426 = (inp[10]) ? node1430 : node1427;
												assign node1427 = (inp[9]) ? 11'b01101011100 : 11'b01001011000;
												assign node1430 = (inp[9]) ? 11'b01010001000 : 11'b01010011110;
										assign node1433 = (inp[10]) ? node1441 : node1434;
											assign node1434 = (inp[9]) ? node1438 : node1435;
												assign node1435 = (inp[11]) ? 11'b01001111010 : 11'b01010101010;
												assign node1438 = (inp[11]) ? 11'b01010101110 : 11'b01110111100;
											assign node1441 = (inp[9]) ? node1445 : node1442;
												assign node1442 = (inp[11]) ? 11'b01111101100 : 11'b01001111100;
												assign node1445 = (inp[11]) ? 11'b01101101000 : 11'b01101011010;
									assign node1448 = (inp[11]) ? node1460 : node1449;
										assign node1449 = (inp[4]) ? node1453 : node1450;
											assign node1450 = (inp[9]) ? 11'b01001001100 : 11'b01010101000;
											assign node1453 = (inp[9]) ? node1457 : node1454;
												assign node1454 = (inp[10]) ? 11'b01000011110 : 11'b01101001000;
												assign node1457 = (inp[10]) ? 11'b01101110001 : 11'b01111110111;
										assign node1460 = (inp[4]) ? node1468 : node1461;
											assign node1461 = (inp[9]) ? node1465 : node1462;
												assign node1462 = (inp[10]) ? 11'b01011110101 : 11'b01000110011;
												assign node1465 = (inp[10]) ? 11'b01100100001 : 11'b01100110111;
											assign node1468 = (inp[10]) ? 11'b01110000111 : node1469;
												assign node1469 = (inp[9]) ? 11'b01101000101 : 11'b01111010001;
								assign node1473 = (inp[5]) ? node1503 : node1474;
									assign node1474 = (inp[4]) ? node1488 : node1475;
										assign node1475 = (inp[11]) ? node1481 : node1476;
											assign node1476 = (inp[10]) ? node1478 : 11'b01100100101;
												assign node1478 = (inp[9]) ? 11'b01101110011 : 11'b01111100111;
											assign node1481 = (inp[10]) ? node1485 : node1482;
												assign node1482 = (inp[9]) ? 11'b01010010111 : 11'b01101010011;
												assign node1485 = (inp[9]) ? 11'b01111100000 : 11'b01111010101;
										assign node1488 = (inp[11]) ? node1496 : node1489;
											assign node1489 = (inp[9]) ? node1493 : node1490;
												assign node1490 = (inp[10]) ? 11'b01110110101 : 11'b01110100011;
												assign node1493 = (inp[10]) ? 11'b01000010001 : 11'b01011010111;
											assign node1496 = (inp[10]) ? node1500 : node1497;
												assign node1497 = (inp[9]) ? 11'b01101100110 : 11'b01100110010;
												assign node1500 = (inp[9]) ? 11'b01000100000 : 11'b01000100100;
									assign node1503 = (inp[10]) ? node1517 : node1504;
										assign node1504 = (inp[11]) ? node1510 : node1505;
											assign node1505 = (inp[4]) ? 11'b01010000000 : node1506;
												assign node1506 = (inp[9]) ? 11'b01110000100 : 11'b01111000000;
											assign node1510 = (inp[9]) ? node1514 : node1511;
												assign node1511 = (inp[4]) ? 11'b01000010000 : 11'b01101110000;
												assign node1514 = (inp[4]) ? 11'b01001000100 : 11'b01000110100;
										assign node1517 = (inp[9]) ? node1525 : node1518;
											assign node1518 = (inp[4]) ? node1522 : node1519;
												assign node1519 = (inp[11]) ? 11'b01100110110 : 11'b01010000110;
												assign node1522 = (inp[11]) ? 11'b01001000110 : 11'b01101110110;
											assign node1525 = (inp[4]) ? 11'b01000110010 : node1526;
												assign node1526 = (inp[11]) ? 11'b01001000010 : 11'b01011010010;
						assign node1530 = (inp[10]) ? node1640 : node1531;
							assign node1531 = (inp[8]) ? node1589 : node1532;
								assign node1532 = (inp[4]) ? node1562 : node1533;
									assign node1533 = (inp[9]) ? node1549 : node1534;
										assign node1534 = (inp[5]) ? node1542 : node1535;
											assign node1535 = (inp[11]) ? node1539 : node1536;
												assign node1536 = (inp[6]) ? 11'b01011001001 : 11'b01011001000;
												assign node1539 = (inp[6]) ? 11'b01010001000 : 11'b01011000001;
											assign node1542 = (inp[6]) ? node1546 : node1543;
												assign node1543 = (inp[11]) ? 11'b01110000010 : 11'b01110000001;
												assign node1546 = (inp[11]) ? 11'b01111100011 : 11'b01110101010;
										assign node1549 = (inp[5]) ? node1555 : node1550;
											assign node1550 = (inp[6]) ? 11'b01111011000 : node1551;
												assign node1551 = (inp[11]) ? 11'b01111110001 : 11'b01011110001;
											assign node1555 = (inp[11]) ? node1559 : node1556;
												assign node1556 = (inp[6]) ? 11'b01110011000 : 11'b01110010011;
												assign node1559 = (inp[6]) ? 11'b01000110011 : 11'b01001010000;
									assign node1562 = (inp[9]) ? node1576 : node1563;
										assign node1563 = (inp[6]) ? node1571 : node1564;
											assign node1564 = (inp[5]) ? node1568 : node1565;
												assign node1565 = (inp[11]) ? 11'b01101110011 : 11'b01011110011;
												assign node1568 = (inp[11]) ? 11'b01011110000 : 11'b01100110000;
											assign node1571 = (inp[5]) ? 11'b01101011000 : node1572;
												assign node1572 = (inp[11]) ? 11'b01101111000 : 11'b01011111010;
										assign node1576 = (inp[5]) ? node1582 : node1577;
											assign node1577 = (inp[6]) ? node1579 : 11'b01111000011;
												assign node1579 = (inp[11]) ? 11'b01101101010 : 11'b01110101010;
											assign node1582 = (inp[11]) ? node1586 : node1583;
												assign node1583 = (inp[6]) ? 11'b01011100001 : 11'b01010100000;
												assign node1586 = (inp[6]) ? 11'b01001000011 : 11'b01001100010;
								assign node1589 = (inp[5]) ? node1617 : node1590;
									assign node1590 = (inp[11]) ? node1602 : node1591;
										assign node1591 = (inp[6]) ? node1597 : node1592;
											assign node1592 = (inp[4]) ? 11'b01011110011 : node1593;
												assign node1593 = (inp[9]) ? 11'b01001010010 : 11'b01011000000;
											assign node1597 = (inp[4]) ? 11'b01101000001 : node1598;
												assign node1598 = (inp[9]) ? 11'b01000110001 : 11'b01011100001;
										assign node1602 = (inp[6]) ? node1610 : node1603;
											assign node1603 = (inp[9]) ? node1607 : node1604;
												assign node1604 = (inp[4]) ? 11'b01100010011 : 11'b01000100011;
												assign node1607 = (inp[4]) ? 11'b01101100001 : 11'b01110010001;
											assign node1610 = (inp[4]) ? node1614 : node1611;
												assign node1611 = (inp[9]) ? 11'b01111110010 : 11'b01001000001;
												assign node1614 = (inp[9]) ? 11'b01100100010 : 11'b01100110010;
									assign node1617 = (inp[4]) ? node1627 : node1618;
										assign node1618 = (inp[11]) ? node1624 : node1619;
											assign node1619 = (inp[6]) ? node1621 : 11'b01111010011;
												assign node1621 = (inp[9]) ? 11'b01111010010 : 11'b01111000010;
											assign node1624 = (inp[9]) ? 11'b01001010010 : 11'b01101100010;
										assign node1627 = (inp[9]) ? node1635 : node1628;
											assign node1628 = (inp[11]) ? node1632 : node1629;
												assign node1629 = (inp[6]) ? 11'b01100010010 : 11'b01101010001;
												assign node1632 = (inp[6]) ? 11'b01000010010 : 11'b01000010000;
											assign node1635 = (inp[11]) ? 11'b01000000010 : node1636;
												assign node1636 = (inp[6]) ? 11'b01000100010 : 11'b01001100010;
							assign node1640 = (inp[9]) ? node1698 : node1641;
								assign node1641 = (inp[6]) ? node1669 : node1642;
									assign node1642 = (inp[5]) ? node1654 : node1643;
										assign node1643 = (inp[4]) ? node1647 : node1644;
											assign node1644 = (inp[8]) ? 11'b01010000000 : 11'b01100000001;
											assign node1647 = (inp[11]) ? node1651 : node1648;
												assign node1648 = (inp[8]) ? 11'b01111100001 : 11'b01100100011;
												assign node1651 = (inp[8]) ? 11'b01001100011 : 11'b01010100011;
										assign node1654 = (inp[11]) ? node1662 : node1655;
											assign node1655 = (inp[4]) ? node1659 : node1656;
												assign node1656 = (inp[8]) ? 11'b01010100011 : 11'b01001000011;
												assign node1659 = (inp[8]) ? 11'b01100000011 : 11'b01111100000;
											assign node1662 = (inp[4]) ? node1666 : node1663;
												assign node1663 = (inp[8]) ? 11'b01101100010 : 11'b01111000010;
												assign node1666 = (inp[8]) ? 11'b01001000010 : 11'b01010100010;
									assign node1669 = (inp[8]) ? node1685 : node1670;
										assign node1670 = (inp[4]) ? node1678 : node1671;
											assign node1671 = (inp[11]) ? node1675 : node1672;
												assign node1672 = (inp[5]) ? 11'b01001001000 : 11'b01000001011;
												assign node1675 = (inp[5]) ? 11'b01111100001 : 11'b01101001010;
											assign node1678 = (inp[11]) ? node1682 : node1679;
												assign node1679 = (inp[5]) ? 11'b01110001010 : 11'b01101101000;
												assign node1682 = (inp[5]) ? 11'b01010000001 : 11'b01010101000;
										assign node1685 = (inp[4]) ? node1693 : node1686;
											assign node1686 = (inp[5]) ? node1690 : node1687;
												assign node1687 = (inp[11]) ? 11'b01110000001 : 11'b01010100011;
												assign node1690 = (inp[11]) ? 11'b01100100000 : 11'b01010000000;
											assign node1693 = (inp[11]) ? node1695 : 11'b01111000011;
												assign node1695 = (inp[5]) ? 11'b01001000000 : 11'b01001100000;
								assign node1698 = (inp[11]) ? node1726 : node1699;
									assign node1699 = (inp[4]) ? node1711 : node1700;
										assign node1700 = (inp[5]) ? node1708 : node1701;
											assign node1701 = (inp[8]) ? node1705 : node1702;
												assign node1702 = (inp[6]) ? 11'b01000101010 : 11'b01000100011;
												assign node1705 = (inp[6]) ? 11'b01001100011 : 11'b01000000010;
											assign node1708 = (inp[6]) ? 11'b01011001010 : 11'b01011100010;
										assign node1711 = (inp[5]) ? node1719 : node1712;
											assign node1712 = (inp[8]) ? node1716 : node1713;
												assign node1713 = (inp[6]) ? 11'b01001001000 : 11'b01000000001;
												assign node1716 = (inp[6]) ? 11'b01000000011 : 11'b01001100011;
											assign node1719 = (inp[8]) ? node1723 : node1720;
												assign node1720 = (inp[6]) ? 11'b01000100011 : 11'b01001000010;
												assign node1723 = (inp[6]) ? 11'b01000100000 : 11'b01001100000;
									assign node1726 = (inp[5]) ? node1742 : node1727;
										assign node1727 = (inp[4]) ? node1735 : node1728;
											assign node1728 = (inp[8]) ? node1732 : node1729;
												assign node1729 = (inp[6]) ? 11'b01010001010 : 11'b01010100011;
												assign node1732 = (inp[6]) ? 11'b01011100000 : 11'b01011000001;
											assign node1735 = (inp[8]) ? node1739 : node1736;
												assign node1736 = (inp[6]) ? 11'b01001101000 : 11'b01001000001;
												assign node1739 = (inp[6]) ? 11'b01000100000 : 11'b01000100001;
										assign node1742 = (inp[4]) ? node1748 : node1743;
											assign node1743 = (inp[6]) ? 11'b01001000001 : node1744;
												assign node1744 = (inp[8]) ? 11'b01001000000 : 11'b01000000000;
											assign node1748 = (inp[8]) ? 11'b01000000000 : 11'b01000100000;
			assign node1751 = (inp[6]) ? node2641 : node1752;
				assign node1752 = (inp[2]) ? node2200 : node1753;
					assign node1753 = (inp[8]) ? node1981 : node1754;
						assign node1754 = (inp[5]) ? node1866 : node1755;
							assign node1755 = (inp[0]) ? node1815 : node1756;
								assign node1756 = (inp[4]) ? node1788 : node1757;
									assign node1757 = (inp[10]) ? node1773 : node1758;
										assign node1758 = (inp[3]) ? node1766 : node1759;
											assign node1759 = (inp[11]) ? node1763 : node1760;
												assign node1760 = (inp[9]) ? 11'b01010100011 : 11'b01011100011;
												assign node1763 = (inp[9]) ? 11'b01110010011 : 11'b01011000011;
											assign node1766 = (inp[9]) ? node1770 : node1767;
												assign node1767 = (inp[11]) ? 11'b11011010011 : 11'b11011100011;
												assign node1770 = (inp[11]) ? 11'b11111100111 : 11'b11011100111;
										assign node1773 = (inp[3]) ? node1781 : node1774;
											assign node1774 = (inp[9]) ? node1778 : node1775;
												assign node1775 = (inp[11]) ? 11'b11011000001 : 11'b11011100001;
												assign node1778 = (inp[11]) ? 11'b11111110101 : 11'b11011110101;
											assign node1781 = (inp[9]) ? node1785 : node1782;
												assign node1782 = (inp[11]) ? 11'b01010010101 : 11'b01010100101;
												assign node1785 = (inp[11]) ? 11'b01001110111 : 11'b01011110101;
									assign node1788 = (inp[11]) ? node1800 : node1789;
										assign node1789 = (inp[9]) ? node1795 : node1790;
											assign node1790 = (inp[10]) ? node1792 : 11'b11010100111;
												assign node1792 = (inp[3]) ? 11'b01111000001 : 11'b11010110101;
											assign node1795 = (inp[10]) ? 11'b11110000001 : node1796;
												assign node1796 = (inp[3]) ? 11'b11110010011 : 11'b01111000111;
										assign node1800 = (inp[10]) ? node1808 : node1801;
											assign node1801 = (inp[3]) ? node1805 : node1802;
												assign node1802 = (inp[9]) ? 11'b01001110111 : 11'b01000100111;
												assign node1805 = (inp[9]) ? 11'b11001110001 : 11'b11100100101;
											assign node1808 = (inp[3]) ? node1812 : node1809;
												assign node1809 = (inp[9]) ? 11'b11100110001 : 11'b11100110101;
												assign node1812 = (inp[9]) ? 11'b01100110011 : 11'b01101110011;
								assign node1815 = (inp[11]) ? node1837 : node1816;
									assign node1816 = (inp[4]) ? node1826 : node1817;
										assign node1817 = (inp[3]) ? node1823 : node1818;
											assign node1818 = (inp[10]) ? 11'b01001110011 : node1819;
												assign node1819 = (inp[9]) ? 11'b01000100101 : 11'b01001100001;
											assign node1823 = (inp[9]) ? 11'b01001110011 : 11'b01001100011;
										assign node1826 = (inp[9]) ? node1834 : node1827;
											assign node1827 = (inp[10]) ? node1831 : node1828;
												assign node1828 = (inp[3]) ? 11'b01000110011 : 11'b01000100001;
												assign node1831 = (inp[3]) ? 11'b01101000001 : 11'b01001010111;
											assign node1834 = (inp[10]) ? 11'b01100010011 : 11'b01101010101;
									assign node1837 = (inp[4]) ? node1851 : node1838;
										assign node1838 = (inp[9]) ? node1846 : node1839;
											assign node1839 = (inp[10]) ? node1843 : node1840;
												assign node1840 = (inp[3]) ? 11'b01001000011 : 11'b01001010001;
												assign node1843 = (inp[3]) ? 11'b01100000001 : 11'b01000010111;
											assign node1846 = (inp[10]) ? node1848 : 11'b01100010101;
												assign node1848 = (inp[3]) ? 11'b01011100001 : 11'b01011100011;
										assign node1851 = (inp[3]) ? node1859 : node1852;
											assign node1852 = (inp[10]) ? node1856 : node1853;
												assign node1853 = (inp[9]) ? 11'b01011100101 : 11'b01010110001;
												assign node1856 = (inp[9]) ? 11'b01110100011 : 11'b01111100111;
											assign node1859 = (inp[10]) ? node1863 : node1860;
												assign node1860 = (inp[9]) ? 11'b01110100011 : 11'b01110110011;
												assign node1863 = (inp[9]) ? 11'b01000100001 : 11'b01011100001;
							assign node1866 = (inp[11]) ? node1924 : node1867;
								assign node1867 = (inp[4]) ? node1897 : node1868;
									assign node1868 = (inp[0]) ? node1884 : node1869;
										assign node1869 = (inp[10]) ? node1877 : node1870;
											assign node1870 = (inp[3]) ? node1874 : node1871;
												assign node1871 = (inp[9]) ? 11'b01010010011 : 11'b01011010011;
												assign node1874 = (inp[9]) ? 11'b11010010101 : 11'b11011010001;
											assign node1877 = (inp[3]) ? node1881 : node1878;
												assign node1878 = (inp[9]) ? 11'b11111000101 : 11'b11111010001;
												assign node1881 = (inp[9]) ? 11'b01001000111 : 11'b01110010111;
										assign node1884 = (inp[10]) ? node1892 : node1885;
											assign node1885 = (inp[3]) ? node1889 : node1886;
												assign node1886 = (inp[9]) ? 11'b01000000111 : 11'b01001000011;
												assign node1889 = (inp[9]) ? 11'b01101010011 : 11'b01101000011;
											assign node1892 = (inp[3]) ? node1894 : 11'b01101010001;
												assign node1894 = (inp[9]) ? 11'b01011000001 : 11'b01000000001;
									assign node1897 = (inp[9]) ? node1913 : node1898;
										assign node1898 = (inp[0]) ? node1906 : node1899;
											assign node1899 = (inp[10]) ? node1903 : node1900;
												assign node1900 = (inp[3]) ? 11'b11100010101 : 11'b01001010101;
												assign node1903 = (inp[3]) ? 11'b01001110010 : 11'b11000000111;
											assign node1906 = (inp[10]) ? node1910 : node1907;
												assign node1907 = (inp[3]) ? 11'b01110010011 : 11'b01110000011;
												assign node1910 = (inp[3]) ? 11'b01111100000 : 11'b01010010101;
										assign node1913 = (inp[10]) ? node1921 : node1914;
											assign node1914 = (inp[3]) ? node1918 : node1915;
												assign node1915 = (inp[0]) ? 11'b01111110110 : 11'b01101110100;
												assign node1918 = (inp[0]) ? 11'b01001100000 : 11'b11011100000;
											assign node1921 = (inp[3]) ? 11'b01110100010 : 11'b11010110010;
								assign node1924 = (inp[4]) ? node1952 : node1925;
									assign node1925 = (inp[0]) ? node1937 : node1926;
										assign node1926 = (inp[9]) ? node1932 : node1927;
											assign node1927 = (inp[3]) ? node1929 : 11'b11111110010;
												assign node1929 = (inp[10]) ? 11'b01001100100 : 11'b11111100000;
											assign node1932 = (inp[3]) ? 11'b11000110110 : node1933;
												assign node1933 = (inp[10]) ? 11'b11101000110 : 11'b01100100000;
										assign node1937 = (inp[3]) ? node1945 : node1938;
											assign node1938 = (inp[10]) ? node1942 : node1939;
												assign node1939 = (inp[9]) ? 11'b01110110110 : 11'b01001110010;
												assign node1942 = (inp[9]) ? 11'b01111000000 : 11'b01011110100;
											assign node1945 = (inp[10]) ? node1949 : node1946;
												assign node1946 = (inp[9]) ? 11'b01010110000 : 11'b01101100000;
												assign node1949 = (inp[9]) ? 11'b01001000010 : 11'b01110100010;
									assign node1952 = (inp[10]) ? node1968 : node1953;
										assign node1953 = (inp[9]) ? node1961 : node1954;
											assign node1954 = (inp[0]) ? node1958 : node1955;
												assign node1955 = (inp[3]) ? 11'b11110010110 : 11'b01011010100;
												assign node1958 = (inp[3]) ? 11'b01000010000 : 11'b01101010000;
											assign node1961 = (inp[0]) ? node1965 : node1962;
												assign node1962 = (inp[3]) ? 11'b11101000010 : 11'b01001000110;
												assign node1965 = (inp[3]) ? 11'b01011000000 : 11'b01111000100;
										assign node1968 = (inp[0]) ? node1974 : node1969;
											assign node1969 = (inp[3]) ? node1971 : 11'b11001000000;
												assign node1971 = (inp[9]) ? 11'b01100000000 : 11'b01110000000;
											assign node1974 = (inp[3]) ? node1978 : node1975;
												assign node1975 = (inp[9]) ? 11'b01110000010 : 11'b01100000110;
												assign node1978 = (inp[9]) ? 11'b01000000000 : 11'b01011000010;
						assign node1981 = (inp[5]) ? node2093 : node1982;
							assign node1982 = (inp[11]) ? node2038 : node1983;
								assign node1983 = (inp[0]) ? node2013 : node1984;
									assign node1984 = (inp[9]) ? node1998 : node1985;
										assign node1985 = (inp[10]) ? node1993 : node1986;
											assign node1986 = (inp[3]) ? node1990 : node1987;
												assign node1987 = (inp[4]) ? 11'b01111100110 : 11'b01010000010;
												assign node1990 = (inp[4]) ? 11'b11011100100 : 11'b11111100010;
											assign node1993 = (inp[3]) ? node1995 : 11'b11110110100;
												assign node1995 = (inp[4]) ? 11'b01000100010 : 11'b01111100100;
										assign node1998 = (inp[4]) ? node2006 : node1999;
											assign node1999 = (inp[10]) ? node2003 : node2000;
												assign node2000 = (inp[3]) ? 11'b11100100100 : 11'b01000100010;
												assign node2003 = (inp[3]) ? 11'b01101110110 : 11'b11000110100;
											assign node2006 = (inp[10]) ? node2010 : node2007;
												assign node2007 = (inp[3]) ? 11'b11001010000 : 11'b01100100100;
												assign node2010 = (inp[3]) ? 11'b01110010010 : 11'b11011000010;
									assign node2013 = (inp[3]) ? node2023 : node2014;
										assign node2014 = (inp[4]) ? node2020 : node2015;
											assign node2015 = (inp[10]) ? 11'b01101100110 : node2016;
												assign node2016 = (inp[9]) ? 11'b01110100100 : 11'b01100000000;
											assign node2020 = (inp[9]) ? 11'b01001010000 : 11'b01100110100;
										assign node2023 = (inp[10]) ? node2031 : node2024;
											assign node2024 = (inp[9]) ? node2028 : node2025;
												assign node2025 = (inp[4]) ? 11'b01000110010 : 11'b01001100010;
												assign node2028 = (inp[4]) ? 11'b01111000010 : 11'b01010110010;
											assign node2031 = (inp[9]) ? node2035 : node2032;
												assign node2032 = (inp[4]) ? 11'b01110100000 : 11'b01011100000;
												assign node2035 = (inp[4]) ? 11'b01000000010 : 11'b01001100000;
								assign node2038 = (inp[4]) ? node2068 : node2039;
									assign node2039 = (inp[0]) ? node2053 : node2040;
										assign node2040 = (inp[3]) ? node2046 : node2041;
											assign node2041 = (inp[10]) ? node2043 : 11'b01101010000;
												assign node2043 = (inp[9]) ? 11'b11010010110 : 11'b11101000010;
											assign node2046 = (inp[10]) ? node2050 : node2047;
												assign node2047 = (inp[9]) ? 11'b11110000110 : 11'b11110010000;
												assign node2050 = (inp[9]) ? 11'b01110010100 : 11'b01001010100;
										assign node2053 = (inp[10]) ? node2061 : node2054;
											assign node2054 = (inp[3]) ? node2058 : node2055;
												assign node2055 = (inp[9]) ? 11'b01001010100 : 11'b01100010010;
												assign node2058 = (inp[9]) ? 11'b01100010000 : 11'b01010000000;
											assign node2061 = (inp[9]) ? node2065 : node2062;
												assign node2062 = (inp[3]) ? 11'b01111000010 : 11'b01111010100;
												assign node2065 = (inp[3]) ? 11'b00011101011 : 11'b01100000010;
									assign node2068 = (inp[0]) ? node2084 : node2069;
										assign node2069 = (inp[10]) ? node2077 : node2070;
											assign node2070 = (inp[9]) ? node2074 : node2071;
												assign node2071 = (inp[3]) ? 11'b10001101111 : 11'b00101101111;
												assign node2074 = (inp[3]) ? 11'b10000111001 : 11'b00010111111;
											assign node2077 = (inp[3]) ? node2081 : node2078;
												assign node2078 = (inp[9]) ? 11'b10101111001 : 11'b10101111101;
												assign node2081 = (inp[9]) ? 11'b00101111011 : 11'b00110111001;
										assign node2084 = (inp[10]) ? node2088 : node2085;
											assign node2085 = (inp[3]) ? 11'b00111101011 : 11'b00111111001;
											assign node2088 = (inp[3]) ? node2090 : 11'b00000101111;
												assign node2090 = (inp[9]) ? 11'b00001101001 : 11'b00000101001;
							assign node2093 = (inp[4]) ? node2147 : node2094;
								assign node2094 = (inp[0]) ? node2126 : node2095;
									assign node2095 = (inp[10]) ? node2111 : node2096;
										assign node2096 = (inp[3]) ? node2104 : node2097;
											assign node2097 = (inp[9]) ? node2101 : node2098;
												assign node2098 = (inp[11]) ? 11'b00011111011 : 11'b00010111011;
												assign node2101 = (inp[11]) ? 11'b00011101011 : 11'b00001011001;
											assign node2104 = (inp[9]) ? node2108 : node2105;
												assign node2105 = (inp[11]) ? 11'b10001101001 : 11'b10010111001;
												assign node2108 = (inp[11]) ? 11'b10111111101 : 11'b10011011101;
										assign node2111 = (inp[3]) ? node2119 : node2112;
											assign node2112 = (inp[9]) ? node2116 : node2113;
												assign node2113 = (inp[11]) ? 11'b10000111001 : 11'b10110111001;
												assign node2116 = (inp[11]) ? 11'b10101101111 : 11'b10010001111;
											assign node2119 = (inp[11]) ? node2123 : node2120;
												assign node2120 = (inp[9]) ? 11'b00110001111 : 11'b00101011111;
												assign node2123 = (inp[9]) ? 11'b00100101111 : 11'b00010101111;
									assign node2126 = (inp[9]) ? node2138 : node2127;
										assign node2127 = (inp[10]) ? node2131 : node2128;
											assign node2128 = (inp[11]) ? 11'b00110101011 : 11'b00100101011;
											assign node2131 = (inp[11]) ? node2135 : node2132;
												assign node2132 = (inp[3]) ? 11'b00011001001 : 11'b00010101101;
												assign node2135 = (inp[3]) ? 11'b00100101001 : 11'b00110111111;
										assign node2138 = (inp[11]) ? node2140 : 11'b00101011001;
											assign node2140 = (inp[10]) ? node2144 : node2141;
												assign node2141 = (inp[3]) ? 11'b00011111011 : 11'b00001111111;
												assign node2144 = (inp[3]) ? 11'b00000101011 : 11'b00011101001;
								assign node2147 = (inp[0]) ? node2177 : node2148;
									assign node2148 = (inp[10]) ? node2164 : node2149;
										assign node2149 = (inp[3]) ? node2157 : node2150;
											assign node2150 = (inp[11]) ? node2154 : node2151;
												assign node2151 = (inp[9]) ? 11'b00110011101 : 11'b00100011101;
												assign node2154 = (inp[9]) ? 11'b00111001101 : 11'b00110111101;
											assign node2157 = (inp[9]) ? node2161 : node2158;
												assign node2158 = (inp[11]) ? 11'b10110111101 : 11'b10001011111;
												assign node2161 = (inp[11]) ? 11'b10110001011 : 11'b10100001011;
										assign node2164 = (inp[3]) ? node2170 : node2165;
											assign node2165 = (inp[9]) ? 11'b10100001001 : node2166;
												assign node2166 = (inp[11]) ? 11'b10101001111 : 11'b10011001111;
											assign node2170 = (inp[11]) ? node2174 : node2171;
												assign node2171 = (inp[9]) ? 11'b00111101001 : 11'b00011011001;
												assign node2174 = (inp[9]) ? 11'b00100001001 : 11'b00101001001;
									assign node2177 = (inp[3]) ? node2187 : node2178;
										assign node2178 = (inp[11]) ? node2184 : node2179;
											assign node2179 = (inp[9]) ? 11'b00010011101 : node2180;
												assign node2180 = (inp[10]) ? 11'b00101011111 : 11'b00011001011;
											assign node2184 = (inp[10]) ? 11'b00011001101 : 11'b00001001101;
										assign node2187 = (inp[10]) ? node2193 : node2188;
											assign node2188 = (inp[11]) ? 11'b00010111001 : node2189;
												assign node2189 = (inp[9]) ? 11'b00010001001 : 11'b00111011001;
											assign node2193 = (inp[9]) ? node2197 : node2194;
												assign node2194 = (inp[11]) ? 11'b00001001011 : 11'b00100001011;
												assign node2197 = (inp[11]) ? 11'b00000001001 : 11'b00001101001;
					assign node2200 = (inp[0]) ? node2424 : node2201;
						assign node2201 = (inp[8]) ? node2305 : node2202;
							assign node2202 = (inp[10]) ? node2254 : node2203;
								assign node2203 = (inp[3]) ? node2227 : node2204;
									assign node2204 = (inp[4]) ? node2216 : node2205;
										assign node2205 = (inp[5]) ? node2211 : node2206;
											assign node2206 = (inp[11]) ? 11'b00110101010 : node2207;
												assign node2207 = (inp[9]) ? 11'b00110001011 : 11'b00111001011;
											assign node2211 = (inp[11]) ? node2213 : 11'b00111111000;
												assign node2213 = (inp[9]) ? 11'b00000001010 : 11'b00111011000;
										assign node2216 = (inp[5]) ? node2222 : node2217;
											assign node2217 = (inp[9]) ? 11'b00100011110 : node2218;
												assign node2218 = (inp[11]) ? 11'b00101001100 : 11'b00111101100;
											assign node2222 = (inp[9]) ? 11'b00010011110 : node2223;
												assign node2223 = (inp[11]) ? 11'b00110111111 : 11'b00100111110;
									assign node2227 = (inp[11]) ? node2243 : node2228;
										assign node2228 = (inp[5]) ? node2236 : node2229;
											assign node2229 = (inp[4]) ? node2233 : node2230;
												assign node2230 = (inp[9]) ? 11'b10110001101 : 11'b10111001011;
												assign node2233 = (inp[9]) ? 11'b10001111010 : 11'b10110101100;
											assign node2236 = (inp[4]) ? node2240 : node2237;
												assign node2237 = (inp[9]) ? 11'b10101111110 : 11'b10110111000;
												assign node2240 = (inp[9]) ? 11'b10110001000 : 11'b10011011110;
										assign node2243 = (inp[5]) ? node2249 : node2244;
											assign node2244 = (inp[4]) ? node2246 : 11'b10000001100;
												assign node2246 = (inp[9]) ? 11'b10111111010 : 11'b10011001110;
											assign node2249 = (inp[9]) ? node2251 : 11'b10000111101;
												assign node2251 = (inp[4]) ? 11'b10011101011 : 11'b10111111111;
								assign node2254 = (inp[3]) ? node2280 : node2255;
									assign node2255 = (inp[5]) ? node2267 : node2256;
										assign node2256 = (inp[4]) ? node2262 : node2257;
											assign node2257 = (inp[9]) ? 11'b10101111110 : node2258;
												assign node2258 = (inp[11]) ? 11'b10101001000 : 11'b10101001001;
											assign node2262 = (inp[9]) ? node2264 : 11'b10100111110;
												assign node2264 = (inp[11]) ? 11'b10001111000 : 11'b10001101000;
										assign node2267 = (inp[11]) ? node2275 : node2268;
											assign node2268 = (inp[4]) ? node2272 : node2269;
												assign node2269 = (inp[9]) ? 11'b10010101110 : 11'b10000111010;
												assign node2272 = (inp[9]) ? 11'b10100011010 : 11'b10111001100;
											assign node2275 = (inp[4]) ? node2277 : 11'b10001101101;
												assign node2277 = (inp[9]) ? 11'b10110101011 : 11'b10100101111;
									assign node2280 = (inp[4]) ? node2294 : node2281;
										assign node2281 = (inp[9]) ? node2289 : node2282;
											assign node2282 = (inp[11]) ? node2286 : node2283;
												assign node2283 = (inp[5]) ? 11'b00011111110 : 11'b00100001111;
												assign node2286 = (inp[5]) ? 11'b00110001100 : 11'b00111011110;
											assign node2289 = (inp[5]) ? node2291 : 11'b00101111110;
												assign node2291 = (inp[11]) ? 11'b00101101111 : 11'b00110101100;
										assign node2294 = (inp[11]) ? node2300 : node2295;
											assign node2295 = (inp[5]) ? 11'b00011001010 : node2296;
												assign node2296 = (inp[9]) ? 11'b00010111000 : 11'b00010101000;
											assign node2300 = (inp[5]) ? 11'b00000101001 : node2301;
												assign node2301 = (inp[9]) ? 11'b00001111010 : 11'b00000011000;
							assign node2305 = (inp[5]) ? node2365 : node2306;
								assign node2306 = (inp[11]) ? node2338 : node2307;
									assign node2307 = (inp[9]) ? node2323 : node2308;
										assign node2308 = (inp[4]) ? node2316 : node2309;
											assign node2309 = (inp[10]) ? node2313 : node2310;
												assign node2310 = (inp[3]) ? 11'b10000101001 : 11'b00110101011;
												assign node2313 = (inp[3]) ? 11'b00011001111 : 11'b10101001001;
											assign node2316 = (inp[3]) ? node2320 : node2317;
												assign node2317 = (inp[10]) ? 11'b10011011101 : 11'b00011001101;
												assign node2320 = (inp[10]) ? 11'b00110001001 : 11'b10101001111;
										assign node2323 = (inp[3]) ? node2331 : node2324;
											assign node2324 = (inp[10]) ? node2328 : node2325;
												assign node2325 = (inp[4]) ? 11'b00000001111 : 11'b00101001001;
												assign node2328 = (inp[4]) ? 11'b10101101011 : 11'b10110011111;
											assign node2331 = (inp[10]) ? node2335 : node2332;
												assign node2332 = (inp[4]) ? 11'b10110011001 : 11'b10010001101;
												assign node2335 = (inp[4]) ? 11'b00011111011 : 11'b00000011101;
									assign node2338 = (inp[4]) ? node2352 : node2339;
										assign node2339 = (inp[10]) ? node2347 : node2340;
											assign node2340 = (inp[3]) ? node2344 : node2341;
												assign node2341 = (inp[9]) ? 11'b00011111011 : 11'b00111101001;
												assign node2344 = (inp[9]) ? 11'b10001101101 : 11'b10000111011;
											assign node2347 = (inp[3]) ? node2349 : 11'b10101111101;
												assign node2349 = (inp[9]) ? 11'b00010111111 : 11'b00100111101;
										assign node2352 = (inp[10]) ? node2358 : node2353;
											assign node2353 = (inp[9]) ? 11'b10100011011 : node2354;
												assign node2354 = (inp[3]) ? 11'b10110101101 : 11'b00000101101;
											assign node2358 = (inp[9]) ? node2362 : node2359;
												assign node2359 = (inp[3]) ? 11'b00011011001 : 11'b10001011111;
												assign node2362 = (inp[3]) ? 11'b00000011011 : 11'b10010011001;
								assign node2365 = (inp[11]) ? node2397 : node2366;
									assign node2366 = (inp[4]) ? node2382 : node2367;
										assign node2367 = (inp[10]) ? node2375 : node2368;
											assign node2368 = (inp[3]) ? node2372 : node2369;
												assign node2369 = (inp[9]) ? 11'b00100011001 : 11'b00111011011;
												assign node2372 = (inp[9]) ? 11'b10110011111 : 11'b10101011001;
											assign node2375 = (inp[9]) ? node2379 : node2376;
												assign node2376 = (inp[3]) ? 11'b00001011101 : 11'b10011011011;
												assign node2379 = (inp[3]) ? 11'b00011101100 : 11'b10100001101;
										assign node2382 = (inp[3]) ? node2390 : node2383;
											assign node2383 = (inp[9]) ? node2387 : node2384;
												assign node2384 = (inp[10]) ? 11'b10100101110 : 11'b00001111110;
												assign node2387 = (inp[10]) ? 11'b10001111000 : 11'b00000111100;
											assign node2390 = (inp[9]) ? node2394 : node2391;
												assign node2391 = (inp[10]) ? 11'b00110111010 : 11'b10111111100;
												assign node2394 = (inp[10]) ? 11'b00011101000 : 11'b10011101010;
									assign node2397 = (inp[3]) ? node2411 : node2398;
										assign node2398 = (inp[4]) ? node2406 : node2399;
											assign node2399 = (inp[9]) ? node2403 : node2400;
												assign node2400 = (inp[10]) ? 11'b10110111000 : 11'b00110111010;
												assign node2403 = (inp[10]) ? 11'b10010001110 : 11'b00111001000;
											assign node2406 = (inp[10]) ? 11'b10011001100 : node2407;
												assign node2407 = (inp[9]) ? 11'b00011001100 : 11'b00010011110;
										assign node2411 = (inp[10]) ? node2419 : node2412;
											assign node2412 = (inp[9]) ? node2416 : node2413;
												assign node2413 = (inp[4]) ? 11'b10000011100 : 11'b10100101000;
												assign node2416 = (inp[4]) ? 11'b10000001010 : 11'b10001011110;
											assign node2419 = (inp[9]) ? node2421 : 11'b00001001010;
												assign node2421 = (inp[4]) ? 11'b00000001000 : 11'b00000001100;
						assign node2424 = (inp[3]) ? node2530 : node2425;
							assign node2425 = (inp[5]) ? node2473 : node2426;
								assign node2426 = (inp[8]) ? node2450 : node2427;
									assign node2427 = (inp[11]) ? node2441 : node2428;
										assign node2428 = (inp[4]) ? node2436 : node2429;
											assign node2429 = (inp[10]) ? node2433 : node2430;
												assign node2430 = (inp[9]) ? 11'b00000001111 : 11'b00001001001;
												assign node2433 = (inp[9]) ? 11'b00011111000 : 11'b00010001111;
											assign node2436 = (inp[9]) ? 11'b00101111100 : node2437;
												assign node2437 = (inp[10]) ? 11'b00010111100 : 11'b00000101010;
										assign node2441 = (inp[10]) ? node2447 : node2442;
											assign node2442 = (inp[9]) ? node2444 : 11'b00011011010;
												assign node2444 = (inp[4]) ? 11'b00000001100 : 11'b00110011110;
											assign node2447 = (inp[9]) ? 11'b00000001000 : 11'b00100001110;
									assign node2450 = (inp[11]) ? node2464 : node2451;
										assign node2451 = (inp[9]) ? node2457 : node2452;
											assign node2452 = (inp[10]) ? node2454 : 11'b00101001001;
												assign node2454 = (inp[4]) ? 11'b00100011111 : 11'b00101001101;
											assign node2457 = (inp[10]) ? node2461 : node2458;
												assign node2458 = (inp[4]) ? 11'b00000011111 : 11'b00110001111;
												assign node2461 = (inp[4]) ? 11'b00011111001 : 11'b00110011001;
										assign node2464 = (inp[9]) ? node2468 : node2465;
											assign node2465 = (inp[10]) ? 11'b00100111111 : 11'b00110111011;
											assign node2468 = (inp[4]) ? 11'b00111001101 : node2469;
												assign node2469 = (inp[10]) ? 11'b00101101001 : 11'b00001111101;
								assign node2473 = (inp[11]) ? node2503 : node2474;
									assign node2474 = (inp[4]) ? node2490 : node2475;
										assign node2475 = (inp[8]) ? node2483 : node2476;
											assign node2476 = (inp[10]) ? node2480 : node2477;
												assign node2477 = (inp[9]) ? 11'b00011101110 : 11'b00000101010;
												assign node2480 = (inp[9]) ? 11'b00100111010 : 11'b00110101100;
											assign node2483 = (inp[10]) ? node2487 : node2484;
												assign node2484 = (inp[9]) ? 11'b00100001101 : 11'b00101001011;
												assign node2487 = (inp[9]) ? 11'b00001111010 : 11'b00001001101;
										assign node2490 = (inp[8]) ? node2496 : node2491;
											assign node2491 = (inp[10]) ? node2493 : 11'b00110101000;
												assign node2493 = (inp[9]) ? 11'b00110011000 : 11'b00011011110;
											assign node2496 = (inp[10]) ? node2500 : node2497;
												assign node2497 = (inp[9]) ? 11'b00011111110 : 11'b00001101010;
												assign node2500 = (inp[9]) ? 11'b00011111010 : 11'b00110111100;
									assign node2503 = (inp[8]) ? node2517 : node2504;
										assign node2504 = (inp[4]) ? node2512 : node2505;
											assign node2505 = (inp[9]) ? node2509 : node2506;
												assign node2506 = (inp[10]) ? 11'b00000011110 : 11'b00011011010;
												assign node2509 = (inp[10]) ? 11'b00111101011 : 11'b00110011100;
											assign node2512 = (inp[9]) ? node2514 : 11'b00100101101;
												assign node2514 = (inp[10]) ? 11'b00110101011 : 11'b00111101111;
										assign node2517 = (inp[9]) ? node2525 : node2518;
											assign node2518 = (inp[4]) ? node2522 : node2519;
												assign node2519 = (inp[10]) ? 11'b00110111100 : 11'b00110111000;
												assign node2522 = (inp[10]) ? 11'b00011001100 : 11'b00010011000;
											assign node2525 = (inp[4]) ? node2527 : 11'b00011011110;
												assign node2527 = (inp[10]) ? 11'b00010001010 : 11'b00010001110;
							assign node2530 = (inp[10]) ? node2586 : node2531;
								assign node2531 = (inp[8]) ? node2559 : node2532;
									assign node2532 = (inp[11]) ? node2544 : node2533;
										assign node2533 = (inp[4]) ? node2539 : node2534;
											assign node2534 = (inp[9]) ? node2536 : 11'b00110101010;
												assign node2536 = (inp[5]) ? 11'b00111111000 : 11'b00011111010;
											assign node2539 = (inp[5]) ? 11'b00010001010 : node2540;
												assign node2540 = (inp[9]) ? 11'b00111101000 : 11'b00010111000;
										assign node2544 = (inp[5]) ? node2552 : node2545;
											assign node2545 = (inp[4]) ? node2549 : node2546;
												assign node2546 = (inp[9]) ? 11'b00110011010 : 11'b00011001010;
												assign node2549 = (inp[9]) ? 11'b00101101010 : 11'b00101011000;
											assign node2552 = (inp[9]) ? node2556 : node2553;
												assign node2553 = (inp[4]) ? 11'b00010111011 : 11'b00111001000;
												assign node2556 = (inp[4]) ? 11'b00001101001 : 11'b00001111011;
									assign node2559 = (inp[5]) ? node2573 : node2560;
										assign node2560 = (inp[4]) ? node2568 : node2561;
											assign node2561 = (inp[9]) ? node2565 : node2562;
												assign node2562 = (inp[11]) ? 11'b00000101001 : 11'b00011001011;
												assign node2565 = (inp[11]) ? 11'b00111111011 : 11'b00000011001;
											assign node2568 = (inp[9]) ? node2570 : 11'b00100111001;
												assign node2570 = (inp[11]) ? 11'b00100001011 : 11'b00101101011;
										assign node2573 = (inp[9]) ? node2581 : node2574;
											assign node2574 = (inp[4]) ? node2578 : node2575;
												assign node2575 = (inp[11]) ? 11'b00100101010 : 11'b00111001011;
												assign node2578 = (inp[11]) ? 11'b00001011010 : 11'b00100111010;
											assign node2581 = (inp[4]) ? 11'b00001101000 : node2582;
												assign node2582 = (inp[11]) ? 11'b00001011000 : 11'b00110011001;
								assign node2586 = (inp[9]) ? node2616 : node2587;
									assign node2587 = (inp[8]) ? node2601 : node2588;
										assign node2588 = (inp[11]) ? node2594 : node2589;
											assign node2589 = (inp[4]) ? node2591 : 11'b00001101010;
												assign node2591 = (inp[5]) ? 11'b00111001000 : 11'b00101101010;
											assign node2594 = (inp[4]) ? node2598 : node2595;
												assign node2595 = (inp[5]) ? 11'b00110001010 : 11'b00101001000;
												assign node2598 = (inp[5]) ? 11'b00011101011 : 11'b00010001010;
										assign node2601 = (inp[11]) ? node2609 : node2602;
											assign node2602 = (inp[4]) ? node2606 : node2603;
												assign node2603 = (inp[5]) ? 11'b00010001011 : 11'b00011001001;
												assign node2606 = (inp[5]) ? 11'b00100101010 : 11'b00110001001;
											assign node2609 = (inp[4]) ? node2613 : node2610;
												assign node2610 = (inp[5]) ? 11'b00101001010 : 11'b00111101011;
												assign node2613 = (inp[5]) ? 11'b00001001010 : 11'b00001001011;
									assign node2616 = (inp[11]) ? node2628 : node2617;
										assign node2617 = (inp[8]) ? node2625 : node2618;
											assign node2618 = (inp[5]) ? node2622 : node2619;
												assign node2619 = (inp[4]) ? 11'b00000101000 : 11'b00001101010;
												assign node2622 = (inp[4]) ? 11'b00001001010 : 11'b00010101010;
											assign node2625 = (inp[4]) ? 11'b00001101011 : 11'b00001001011;
										assign node2628 = (inp[8]) ? node2636 : node2629;
											assign node2629 = (inp[5]) ? node2633 : node2630;
												assign node2630 = (inp[4]) ? 11'b00001101000 : 11'b00011001010;
												assign node2633 = (inp[4]) ? 11'b00000101001 : 11'b00001101001;
											assign node2636 = (inp[5]) ? 11'b00000001000 : node2637;
												assign node2637 = (inp[4]) ? 11'b00000001001 : 11'b00010101001;
				assign node2641 = (inp[8]) ? node3087 : node2642;
					assign node2642 = (inp[5]) ? node2866 : node2643;
						assign node2643 = (inp[2]) ? node2753 : node2644;
							assign node2644 = (inp[11]) ? node2700 : node2645;
								assign node2645 = (inp[3]) ? node2673 : node2646;
									assign node2646 = (inp[9]) ? node2658 : node2647;
										assign node2647 = (inp[10]) ? node2651 : node2648;
											assign node2648 = (inp[0]) ? 11'b00011101000 : 11'b00011101010;
											assign node2651 = (inp[4]) ? node2655 : node2652;
												assign node2652 = (inp[0]) ? 11'b00011101100 : 11'b10011101000;
												assign node2655 = (inp[0]) ? 11'b00010111100 : 11'b10010111100;
										assign node2658 = (inp[4]) ? node2666 : node2659;
											assign node2659 = (inp[10]) ? node2663 : node2660;
												assign node2660 = (inp[0]) ? 11'b00010101110 : 11'b00010101000;
												assign node2663 = (inp[0]) ? 11'b00011111010 : 11'b10011111110;
											assign node2666 = (inp[10]) ? node2670 : node2667;
												assign node2667 = (inp[0]) ? 11'b00111011110 : 11'b00110101100;
												assign node2670 = (inp[0]) ? 11'b00111011010 : 11'b10111001010;
									assign node2673 = (inp[9]) ? node2687 : node2674;
										assign node2674 = (inp[10]) ? node2682 : node2675;
											assign node2675 = (inp[0]) ? node2679 : node2676;
												assign node2676 = (inp[4]) ? 11'b10001101100 : 11'b10001101000;
												assign node2679 = (inp[4]) ? 11'b00000111010 : 11'b00001101010;
											assign node2682 = (inp[4]) ? 11'b00100101010 : node2683;
												assign node2683 = (inp[0]) ? 11'b00000101010 : 11'b00000101110;
										assign node2687 = (inp[4]) ? node2693 : node2688;
											assign node2688 = (inp[10]) ? node2690 : 11'b00000111000;
												assign node2690 = (inp[0]) ? 11'b00001101000 : 11'b00001111100;
											assign node2693 = (inp[0]) ? node2697 : node2694;
												assign node2694 = (inp[10]) ? 11'b00101011000 : 11'b10101011010;
												assign node2697 = (inp[10]) ? 11'b00001001000 : 11'b00101001000;
								assign node2700 = (inp[4]) ? node2724 : node2701;
									assign node2701 = (inp[9]) ? node2713 : node2702;
										assign node2702 = (inp[0]) ? node2706 : node2703;
											assign node2703 = (inp[10]) ? 11'b10000001010 : 11'b10010011000;
											assign node2706 = (inp[3]) ? node2710 : node2707;
												assign node2707 = (inp[10]) ? 11'b00010011100 : 11'b00010011000;
												assign node2710 = (inp[10]) ? 11'b00101001010 : 11'b00000001010;
										assign node2713 = (inp[3]) ? node2719 : node2714;
											assign node2714 = (inp[0]) ? 11'b00111011110 : node2715;
												assign node2715 = (inp[10]) ? 11'b10101011100 : 11'b00101011000;
											assign node2719 = (inp[10]) ? node2721 : 11'b00101011000;
												assign node2721 = (inp[0]) ? 11'b00010001000 : 11'b00010011100;
									assign node2724 = (inp[9]) ? node2738 : node2725;
										assign node2725 = (inp[10]) ? node2733 : node2726;
											assign node2726 = (inp[0]) ? node2730 : node2727;
												assign node2727 = (inp[3]) ? 11'b10110001100 : 11'b00000001110;
												assign node2730 = (inp[3]) ? 11'b00111110011 : 11'b00000011010;
											assign node2733 = (inp[0]) ? 11'b00101100101 : node2734;
												assign node2734 = (inp[3]) ? 11'b00111110011 : 11'b10101110111;
										assign node2738 = (inp[0]) ? node2746 : node2739;
											assign node2739 = (inp[3]) ? node2743 : node2740;
												assign node2740 = (inp[10]) ? 11'b10110110001 : 11'b00011110101;
												assign node2743 = (inp[10]) ? 11'b00100110011 : 11'b10000110011;
											assign node2746 = (inp[10]) ? node2750 : node2747;
												assign node2747 = (inp[3]) ? 11'b00110100001 : 11'b00001100101;
												assign node2750 = (inp[3]) ? 11'b00000100001 : 11'b00100100011;
							assign node2753 = (inp[0]) ? node2811 : node2754;
								assign node2754 = (inp[11]) ? node2782 : node2755;
									assign node2755 = (inp[4]) ? node2769 : node2756;
										assign node2756 = (inp[10]) ? node2762 : node2757;
											assign node2757 = (inp[3]) ? 11'b10110000110 : node2758;
												assign node2758 = (inp[9]) ? 11'b00110000000 : 11'b00111000010;
											assign node2762 = (inp[9]) ? node2766 : node2763;
												assign node2763 = (inp[3]) ? 11'b00101000100 : 11'b10101000010;
												assign node2766 = (inp[3]) ? 11'b00101110111 : 11'b10100010100;
										assign node2769 = (inp[9]) ? node2777 : node2770;
											assign node2770 = (inp[10]) ? node2774 : node2771;
												assign node2771 = (inp[3]) ? 11'b10111100111 : 11'b00111100101;
												assign node2774 = (inp[3]) ? 11'b00000100011 : 11'b10101110101;
											assign node2777 = (inp[10]) ? 11'b10011100011 : node2778;
												assign node2778 = (inp[3]) ? 11'b10010110001 : 11'b00000100101;
									assign node2782 = (inp[4]) ? node2798 : node2783;
										assign node2783 = (inp[9]) ? node2791 : node2784;
											assign node2784 = (inp[3]) ? node2788 : node2785;
												assign node2785 = (inp[10]) ? 11'b10110100011 : 11'b00101100011;
												assign node2788 = (inp[10]) ? 11'b00100110101 : 11'b10111110001;
											assign node2791 = (inp[10]) ? node2795 : node2792;
												assign node2792 = (inp[3]) ? 11'b10000100101 : 11'b00000110011;
												assign node2795 = (inp[3]) ? 11'b00111010111 : 11'b10011010101;
										assign node2798 = (inp[3]) ? node2806 : node2799;
											assign node2799 = (inp[10]) ? node2803 : node2800;
												assign node2800 = (inp[9]) ? 11'b00110010101 : 11'b00101000101;
												assign node2803 = (inp[9]) ? 11'b10001010001 : 11'b10000010101;
											assign node2806 = (inp[10]) ? 11'b00010010011 : node2807;
												assign node2807 = (inp[9]) ? 11'b10101010011 : 11'b10000000111;
								assign node2811 = (inp[3]) ? node2837 : node2812;
									assign node2812 = (inp[4]) ? node2824 : node2813;
										assign node2813 = (inp[11]) ? node2817 : node2814;
											assign node2814 = (inp[9]) ? 11'b00010000100 : 11'b00011000000;
											assign node2817 = (inp[10]) ? node2821 : node2818;
												assign node2818 = (inp[9]) ? 11'b00100110101 : 11'b00001110011;
												assign node2821 = (inp[9]) ? 11'b00011000001 : 11'b00010110101;
										assign node2824 = (inp[11]) ? node2830 : node2825;
											assign node2825 = (inp[9]) ? node2827 : 11'b00011100011;
												assign node2827 = (inp[10]) ? 11'b00101110011 : 11'b00110110111;
											assign node2830 = (inp[10]) ? node2834 : node2831;
												assign node2831 = (inp[9]) ? 11'b00011000111 : 11'b00001010001;
												assign node2834 = (inp[9]) ? 11'b00101000011 : 11'b00110000111;
									assign node2837 = (inp[4]) ? node2853 : node2838;
										assign node2838 = (inp[10]) ? node2846 : node2839;
											assign node2839 = (inp[11]) ? node2843 : node2840;
												assign node2840 = (inp[9]) ? 11'b00010010010 : 11'b00011000010;
												assign node2843 = (inp[9]) ? 11'b00111010011 : 11'b00010100011;
											assign node2846 = (inp[9]) ? node2850 : node2847;
												assign node2847 = (inp[11]) ? 11'b00100100011 : 11'b00000000010;
												assign node2850 = (inp[11]) ? 11'b00011000011 : 11'b00001100011;
										assign node2853 = (inp[11]) ? node2859 : node2854;
											assign node2854 = (inp[10]) ? node2856 : 11'b00110100001;
												assign node2856 = (inp[9]) ? 11'b00001100001 : 11'b00100100001;
											assign node2859 = (inp[10]) ? node2863 : node2860;
												assign node2860 = (inp[9]) ? 11'b00101000001 : 11'b00100010011;
												assign node2863 = (inp[9]) ? 11'b00001000001 : 11'b00010000001;
						assign node2866 = (inp[0]) ? node2978 : node2867;
							assign node2867 = (inp[9]) ? node2921 : node2868;
								assign node2868 = (inp[4]) ? node2896 : node2869;
									assign node2869 = (inp[3]) ? node2885 : node2870;
										assign node2870 = (inp[11]) ? node2878 : node2871;
											assign node2871 = (inp[2]) ? node2875 : node2872;
												assign node2872 = (inp[10]) ? 11'b10111110011 : 11'b00011110011;
												assign node2875 = (inp[10]) ? 11'b10010010011 : 11'b00110010011;
											assign node2878 = (inp[10]) ? node2882 : node2879;
												assign node2879 = (inp[2]) ? 11'b00100110001 : 11'b00001010001;
												assign node2882 = (inp[2]) ? 11'b10010110001 : 11'b10100010001;
										assign node2885 = (inp[10]) ? node2893 : node2886;
											assign node2886 = (inp[11]) ? node2890 : node2887;
												assign node2887 = (inp[2]) ? 11'b10110010001 : 11'b10001110001;
												assign node2890 = (inp[2]) ? 11'b10000100011 : 11'b10110000011;
											assign node2893 = (inp[11]) ? 11'b00010000101 : 11'b00000010101;
									assign node2896 = (inp[10]) ? node2908 : node2897;
										assign node2897 = (inp[3]) ? node2905 : node2898;
											assign node2898 = (inp[2]) ? node2902 : node2899;
												assign node2899 = (inp[11]) ? 11'b00010110101 : 11'b00001010101;
												assign node2902 = (inp[11]) ? 11'b00110010111 : 11'b00100110111;
											assign node2905 = (inp[11]) ? 11'b10010010101 : 11'b10000110101;
										assign node2908 = (inp[3]) ? node2916 : node2909;
											assign node2909 = (inp[2]) ? node2913 : node2910;
												assign node2910 = (inp[11]) ? 11'b10000100101 : 11'b10010000111;
												assign node2913 = (inp[11]) ? 11'b10111000111 : 11'b10100100111;
											assign node2916 = (inp[11]) ? 11'b00111100011 : node2917;
												assign node2917 = (inp[2]) ? 11'b00111110011 : 11'b00000010001;
								assign node2921 = (inp[11]) ? node2949 : node2922;
									assign node2922 = (inp[2]) ? node2936 : node2923;
										assign node2923 = (inp[4]) ? node2931 : node2924;
											assign node2924 = (inp[10]) ? node2928 : node2925;
												assign node2925 = (inp[3]) ? 11'b10010110111 : 11'b00000110011;
												assign node2928 = (inp[3]) ? 11'b00011000111 : 11'b10100100101;
											assign node2931 = (inp[3]) ? 11'b10000000001 : node2932;
												assign node2932 = (inp[10]) ? 11'b10011010001 : 11'b00110010111;
										assign node2936 = (inp[10]) ? node2942 : node2937;
											assign node2937 = (inp[3]) ? 11'b10111110101 : node2938;
												assign node2938 = (inp[4]) ? 11'b00011110101 : 11'b00101110011;
											assign node2942 = (inp[4]) ? node2946 : node2943;
												assign node2943 = (inp[3]) ? 11'b00111100101 : 11'b10011100111;
												assign node2946 = (inp[3]) ? 11'b00000100011 : 11'b10101110001;
									assign node2949 = (inp[2]) ? node2963 : node2950;
										assign node2950 = (inp[3]) ? node2958 : node2951;
											assign node2951 = (inp[10]) ? node2955 : node2952;
												assign node2952 = (inp[4]) ? 11'b00001100101 : 11'b00101100011;
												assign node2955 = (inp[4]) ? 11'b10010100011 : 11'b10111100111;
											assign node2958 = (inp[4]) ? node2960 : 11'b00001100101;
												assign node2960 = (inp[10]) ? 11'b00100100001 : 11'b10111100001;
										assign node2963 = (inp[10]) ? node2971 : node2964;
											assign node2964 = (inp[3]) ? node2968 : node2965;
												assign node2965 = (inp[4]) ? 11'b00101000111 : 11'b00011000001;
												assign node2968 = (inp[4]) ? 11'b10001000001 : 11'b10101010111;
											assign node2971 = (inp[3]) ? node2975 : node2972;
												assign node2972 = (inp[4]) ? 11'b10100000011 : 11'b10001000101;
												assign node2975 = (inp[4]) ? 11'b00000000001 : 11'b00100000111;
							assign node2978 = (inp[3]) ? node3034 : node2979;
								assign node2979 = (inp[9]) ? node3007 : node2980;
									assign node2980 = (inp[10]) ? node2992 : node2981;
										assign node2981 = (inp[4]) ? node2987 : node2982;
											assign node2982 = (inp[11]) ? node2984 : 11'b00010000011;
												assign node2984 = (inp[2]) ? 11'b00000110001 : 11'b00010010011;
											assign node2987 = (inp[11]) ? node2989 : 11'b00100100001;
												assign node2989 = (inp[2]) ? 11'b00110010011 : 11'b00110110001;
										assign node2992 = (inp[11]) ? node3000 : node2993;
											assign node2993 = (inp[4]) ? node2997 : node2994;
												assign node2994 = (inp[2]) ? 11'b00100000111 : 11'b00111100101;
												assign node2997 = (inp[2]) ? 11'b00000110101 : 11'b00000010111;
											assign node3000 = (inp[4]) ? node3004 : node3001;
												assign node3001 = (inp[2]) ? 11'b00011010111 : 11'b00000010111;
												assign node3004 = (inp[2]) ? 11'b00111000111 : 11'b00111100111;
									assign node3007 = (inp[10]) ? node3021 : node3008;
										assign node3008 = (inp[11]) ? node3016 : node3009;
											assign node3009 = (inp[4]) ? node3013 : node3010;
												assign node3010 = (inp[2]) ? 11'b00001100111 : 11'b00010100101;
												assign node3013 = (inp[2]) ? 11'b00111110101 : 11'b00100010101;
											assign node3016 = (inp[4]) ? 11'b00101000111 : node3017;
												assign node3017 = (inp[2]) ? 11'b00101010111 : 11'b00101110111;
										assign node3021 = (inp[11]) ? node3029 : node3022;
											assign node3022 = (inp[2]) ? node3026 : node3023;
												assign node3023 = (inp[4]) ? 11'b00111010001 : 11'b00111010011;
												assign node3026 = (inp[4]) ? 11'b00101110001 : 11'b00111110001;
											assign node3029 = (inp[2]) ? 11'b00100000011 : node3030;
												assign node3030 = (inp[4]) ? 11'b00100100011 : 11'b00101100001;
								assign node3034 = (inp[10]) ? node3062 : node3035;
									assign node3035 = (inp[11]) ? node3049 : node3036;
										assign node3036 = (inp[9]) ? node3042 : node3037;
											assign node3037 = (inp[2]) ? 11'b00100110011 : node3038;
												assign node3038 = (inp[4]) ? 11'b00111010001 : 11'b00101100001;
											assign node3042 = (inp[4]) ? node3046 : node3043;
												assign node3043 = (inp[2]) ? 11'b00111110011 : 11'b00100110011;
												assign node3046 = (inp[2]) ? 11'b00011100011 : 11'b00001000011;
										assign node3049 = (inp[9]) ? node3055 : node3050;
											assign node3050 = (inp[4]) ? node3052 : 11'b00100000001;
												assign node3052 = (inp[2]) ? 11'b00010010001 : 11'b00000110011;
											assign node3055 = (inp[2]) ? node3059 : node3056;
												assign node3056 = (inp[4]) ? 11'b00011100001 : 11'b00011110011;
												assign node3059 = (inp[4]) ? 11'b00001000001 : 11'b00001010001;
									assign node3062 = (inp[9]) ? node3074 : node3063;
										assign node3063 = (inp[11]) ? node3069 : node3064;
											assign node3064 = (inp[4]) ? 11'b00110000011 : node3065;
												assign node3065 = (inp[2]) ? 11'b00000000001 : 11'b00000100011;
											assign node3069 = (inp[2]) ? node3071 : 11'b00011100001;
												assign node3071 = (inp[4]) ? 11'b00011000001 : 11'b00111000001;
										assign node3074 = (inp[11]) ? node3082 : node3075;
											assign node3075 = (inp[2]) ? node3079 : node3076;
												assign node3076 = (inp[4]) ? 11'b00001000011 : 11'b00011000001;
												assign node3079 = (inp[4]) ? 11'b00000100011 : 11'b00010100011;
											assign node3082 = (inp[2]) ? 11'b00000000001 : node3083;
												assign node3083 = (inp[4]) ? 11'b00000100001 : 11'b00000100011;
					assign node3087 = (inp[0]) ? node3315 : node3088;
						assign node3088 = (inp[11]) ? node3204 : node3089;
							assign node3089 = (inp[2]) ? node3143 : node3090;
								assign node3090 = (inp[5]) ? node3116 : node3091;
									assign node3091 = (inp[9]) ? node3105 : node3092;
										assign node3092 = (inp[4]) ? node3098 : node3093;
											assign node3093 = (inp[3]) ? 11'b10100100001 : node3094;
												assign node3094 = (inp[10]) ? 11'b10001000011 : 11'b00010100011;
											assign node3098 = (inp[3]) ? node3102 : node3099;
												assign node3099 = (inp[10]) ? 11'b10101010111 : 11'b00111000111;
												assign node3102 = (inp[10]) ? 11'b00011000001 : 11'b10011000101;
										assign node3105 = (inp[3]) ? node3111 : node3106;
											assign node3106 = (inp[10]) ? node3108 : 11'b00001000001;
												assign node3108 = (inp[4]) ? 11'b10010000001 : 11'b10010010101;
											assign node3111 = (inp[10]) ? node3113 : 11'b10000010001;
												assign node3113 = (inp[4]) ? 11'b00101110010 : 11'b00100010111;
									assign node3116 = (inp[9]) ? node3132 : node3117;
										assign node3117 = (inp[4]) ? node3125 : node3118;
											assign node3118 = (inp[3]) ? node3122 : node3119;
												assign node3119 = (inp[10]) ? 11'b10100010010 : 11'b00010010010;
												assign node3122 = (inp[10]) ? 11'b00110010100 : 11'b10010010000;
											assign node3125 = (inp[10]) ? node3129 : node3126;
												assign node3126 = (inp[3]) ? 11'b10000010110 : 11'b00100010100;
												assign node3129 = (inp[3]) ? 11'b00011110010 : 11'b10010000100;
										assign node3132 = (inp[4]) ? node3136 : node3133;
											assign node3133 = (inp[10]) ? 11'b10001000110 : 11'b00011010010;
											assign node3136 = (inp[3]) ? node3140 : node3137;
												assign node3137 = (inp[10]) ? 11'b10110110010 : 11'b00101110100;
												assign node3140 = (inp[10]) ? 11'b00100100000 : 11'b10111100000;
								assign node3143 = (inp[9]) ? node3175 : node3144;
									assign node3144 = (inp[5]) ? node3160 : node3145;
										assign node3145 = (inp[10]) ? node3153 : node3146;
											assign node3146 = (inp[4]) ? node3150 : node3147;
												assign node3147 = (inp[3]) ? 11'b10010000001 : 11'b00110000011;
												assign node3150 = (inp[3]) ? 11'b10111100110 : 11'b00000100110;
											assign node3153 = (inp[3]) ? node3157 : node3154;
												assign node3154 = (inp[4]) ? 11'b10011110100 : 11'b10111100010;
												assign node3157 = (inp[4]) ? 11'b00111100010 : 11'b00011100100;
										assign node3160 = (inp[3]) ? node3168 : node3161;
											assign node3161 = (inp[4]) ? node3165 : node3162;
												assign node3162 = (inp[10]) ? 11'b10011110010 : 11'b00111110010;
												assign node3165 = (inp[10]) ? 11'b10101100110 : 11'b00011110110;
											assign node3168 = (inp[10]) ? node3172 : node3169;
												assign node3169 = (inp[4]) ? 11'b10101110100 : 11'b10111110000;
												assign node3172 = (inp[4]) ? 11'b00101110000 : 11'b00011110100;
									assign node3175 = (inp[4]) ? node3189 : node3176;
										assign node3176 = (inp[3]) ? node3184 : node3177;
											assign node3177 = (inp[10]) ? node3181 : node3178;
												assign node3178 = (inp[5]) ? 11'b00110110010 : 11'b00101100010;
												assign node3181 = (inp[5]) ? 11'b10110100110 : 11'b10100110110;
											assign node3184 = (inp[10]) ? node3186 : 11'b10110110100;
												assign node3186 = (inp[5]) ? 11'b00010100100 : 11'b00000110100;
										assign node3189 = (inp[3]) ? node3197 : node3190;
											assign node3190 = (inp[10]) ? node3194 : node3191;
												assign node3191 = (inp[5]) ? 11'b00000110110 : 11'b00011100100;
												assign node3194 = (inp[5]) ? 11'b10000110010 : 11'b10100100000;
											assign node3197 = (inp[5]) ? node3201 : node3198;
												assign node3198 = (inp[10]) ? 11'b00000110010 : 11'b10100110010;
												assign node3201 = (inp[10]) ? 11'b00000100000 : 11'b10000100000;
							assign node3204 = (inp[2]) ? node3262 : node3205;
								assign node3205 = (inp[4]) ? node3235 : node3206;
									assign node3206 = (inp[9]) ? node3222 : node3207;
										assign node3207 = (inp[3]) ? node3215 : node3208;
											assign node3208 = (inp[5]) ? node3212 : node3209;
												assign node3209 = (inp[10]) ? 11'b10101100000 : 11'b00001100000;
												assign node3212 = (inp[10]) ? 11'b10011110010 : 11'b00000110010;
											assign node3215 = (inp[10]) ? node3219 : node3216;
												assign node3216 = (inp[5]) ? 11'b10010100000 : 11'b10111110010;
												assign node3219 = (inp[5]) ? 11'b00001100100 : 11'b00000110110;
										assign node3222 = (inp[3]) ? node3228 : node3223;
											assign node3223 = (inp[10]) ? node3225 : 11'b00001100010;
												assign node3225 = (inp[5]) ? 11'b10100100100 : 11'b10001110110;
											assign node3228 = (inp[10]) ? node3232 : node3229;
												assign node3229 = (inp[5]) ? 11'b10110110110 : 11'b10100100100;
												assign node3232 = (inp[5]) ? 11'b00100100110 : 11'b00111110100;
									assign node3235 = (inp[10]) ? node3249 : node3236;
										assign node3236 = (inp[3]) ? node3242 : node3237;
											assign node3237 = (inp[5]) ? node3239 : 11'b00000110100;
												assign node3239 = (inp[9]) ? 11'b00110000110 : 11'b00110110100;
											assign node3242 = (inp[9]) ? node3246 : node3243;
												assign node3243 = (inp[5]) ? 11'b10111010110 : 11'b10001100100;
												assign node3246 = (inp[5]) ? 11'b10110000000 : 11'b10011010010;
										assign node3249 = (inp[3]) ? node3255 : node3250;
											assign node3250 = (inp[5]) ? node3252 : 11'b10101010000;
												assign node3252 = (inp[9]) ? 11'b10100000010 : 11'b10101000100;
											assign node3255 = (inp[5]) ? node3259 : node3256;
												assign node3256 = (inp[9]) ? 11'b00101010010 : 11'b00100110010;
												assign node3259 = (inp[9]) ? 11'b00100000000 : 11'b00101000010;
								assign node3262 = (inp[9]) ? node3286 : node3263;
									assign node3263 = (inp[4]) ? node3275 : node3264;
										assign node3264 = (inp[5]) ? node3270 : node3265;
											assign node3265 = (inp[3]) ? 11'b10001010010 : node3266;
												assign node3266 = (inp[10]) ? 11'b10001000000 : 11'b00100100000;
											assign node3270 = (inp[3]) ? node3272 : 11'b10101010010;
												assign node3272 = (inp[10]) ? 11'b00101000100 : 11'b10101000000;
										assign node3275 = (inp[3]) ? node3281 : node3276;
											assign node3276 = (inp[5]) ? 11'b00001010110 : node3277;
												assign node3277 = (inp[10]) ? 11'b10001010100 : 11'b00010000100;
											assign node3281 = (inp[10]) ? node3283 : 11'b10001010100;
												assign node3283 = (inp[5]) ? 11'b00001000000 : 11'b00001010010;
									assign node3286 = (inp[5]) ? node3302 : node3287;
										assign node3287 = (inp[3]) ? node3295 : node3288;
											assign node3288 = (inp[10]) ? node3292 : node3289;
												assign node3289 = (inp[4]) ? 11'b00101010100 : 11'b00011010000;
												assign node3292 = (inp[4]) ? 11'b10000010000 : 11'b10110010100;
											assign node3295 = (inp[4]) ? node3299 : node3296;
												assign node3296 = (inp[10]) ? 11'b00010010110 : 11'b10010000110;
												assign node3299 = (inp[10]) ? 11'b00000010010 : 11'b10100010010;
										assign node3302 = (inp[3]) ? node3308 : node3303;
											assign node3303 = (inp[10]) ? node3305 : 11'b00000000110;
												assign node3305 = (inp[4]) ? 11'b10000000010 : 11'b10000000110;
											assign node3308 = (inp[10]) ? node3312 : node3309;
												assign node3309 = (inp[4]) ? 11'b10000000000 : 11'b10000010100;
												assign node3312 = (inp[4]) ? 11'b00000000000 : 11'b00000000100;
						assign node3315 = (inp[3]) ? node3417 : node3316;
							assign node3316 = (inp[5]) ? node3366 : node3317;
								assign node3317 = (inp[11]) ? node3341 : node3318;
									assign node3318 = (inp[2]) ? node3332 : node3319;
										assign node3319 = (inp[9]) ? node3327 : node3320;
											assign node3320 = (inp[10]) ? node3324 : node3321;
												assign node3321 = (inp[4]) ? 11'b00111000011 : 11'b00110100001;
												assign node3324 = (inp[4]) ? 11'b00111010101 : 11'b00111000101;
											assign node3327 = (inp[10]) ? node3329 : 11'b00101000101;
												assign node3329 = (inp[4]) ? 11'b00010010001 : 11'b00100010011;
										assign node3332 = (inp[9]) ? node3336 : node3333;
											assign node3333 = (inp[10]) ? 11'b00111110100 : 11'b00110100000;
											assign node3336 = (inp[10]) ? node3338 : 11'b00011110100;
												assign node3338 = (inp[4]) ? 11'b00000110000 : 11'b00100110000;
									assign node3341 = (inp[9]) ? node3355 : node3342;
										assign node3342 = (inp[10]) ? node3350 : node3343;
											assign node3343 = (inp[2]) ? node3347 : node3344;
												assign node3344 = (inp[4]) ? 11'b00101110000 : 11'b00111110010;
												assign node3347 = (inp[4]) ? 11'b00101010010 : 11'b00100110000;
											assign node3350 = (inp[4]) ? node3352 : 11'b00100110110;
												assign node3352 = (inp[2]) ? 11'b00001000110 : 11'b00010100100;
										assign node3355 = (inp[10]) ? node3363 : node3356;
											assign node3356 = (inp[4]) ? node3360 : node3357;
												assign node3357 = (inp[2]) ? 11'b00010010110 : 11'b00010110110;
												assign node3360 = (inp[2]) ? 11'b00100000110 : 11'b00111000110;
											assign node3363 = (inp[4]) ? 11'b00000000010 : 11'b00110000010;
								assign node3366 = (inp[4]) ? node3396 : node3367;
									assign node3367 = (inp[11]) ? node3381 : node3368;
										assign node3368 = (inp[2]) ? node3376 : node3369;
											assign node3369 = (inp[9]) ? node3373 : node3370;
												assign node3370 = (inp[10]) ? 11'b00000000110 : 11'b00110000010;
												assign node3373 = (inp[10]) ? 11'b00011010000 : 11'b00101000100;
											assign node3376 = (inp[9]) ? 11'b00110100110 : node3377;
												assign node3377 = (inp[10]) ? 11'b00011100110 : 11'b00111100010;
										assign node3381 = (inp[2]) ? node3389 : node3382;
											assign node3382 = (inp[10]) ? node3386 : node3383;
												assign node3383 = (inp[9]) ? 11'b00011110100 : 11'b00110110000;
												assign node3386 = (inp[9]) ? 11'b00000100000 : 11'b00101110100;
											assign node3389 = (inp[9]) ? node3393 : node3390;
												assign node3390 = (inp[10]) ? 11'b00101010110 : 11'b00101010010;
												assign node3393 = (inp[10]) ? 11'b00000000010 : 11'b00000010110;
									assign node3396 = (inp[11]) ? node3410 : node3397;
										assign node3397 = (inp[9]) ? node3403 : node3398;
											assign node3398 = (inp[10]) ? 11'b00111110110 : node3399;
												assign node3399 = (inp[2]) ? 11'b00011100010 : 11'b00000000000;
											assign node3403 = (inp[10]) ? node3407 : node3404;
												assign node3404 = (inp[2]) ? 11'b00000110110 : 11'b00001110110;
												assign node3407 = (inp[2]) ? 11'b00000110010 : 11'b00010110010;
										assign node3410 = (inp[9]) ? node3414 : node3411;
											assign node3411 = (inp[10]) ? 11'b00001000110 : 11'b00001010010;
											assign node3414 = (inp[10]) ? 11'b00000000010 : 11'b00010000110;
							assign node3417 = (inp[9]) ? node3465 : node3418;
								assign node3418 = (inp[4]) ? node3440 : node3419;
									assign node3419 = (inp[11]) ? node3429 : node3420;
										assign node3420 = (inp[2]) ? node3424 : node3421;
											assign node3421 = (inp[10]) ? 11'b00011000010 : 11'b00001000011;
											assign node3424 = (inp[5]) ? node3426 : 11'b00011100010;
												assign node3426 = (inp[10]) ? 11'b00011100000 : 11'b00111100000;
										assign node3429 = (inp[2]) ? node3435 : node3430;
											assign node3430 = (inp[5]) ? node3432 : 11'b00110100000;
												assign node3432 = (inp[10]) ? 11'b00101100010 : 11'b00111100010;
											assign node3435 = (inp[10]) ? node3437 : 11'b00001000010;
												assign node3437 = (inp[5]) ? 11'b00101000000 : 11'b00111000000;
									assign node3440 = (inp[10]) ? node3454 : node3441;
										assign node3441 = (inp[5]) ? node3449 : node3442;
											assign node3442 = (inp[11]) ? node3446 : node3443;
												assign node3443 = (inp[2]) ? 11'b00011110010 : 11'b00001010001;
												assign node3446 = (inp[2]) ? 11'b00101010000 : 11'b00110110010;
											assign node3449 = (inp[11]) ? node3451 : 11'b00110010000;
												assign node3451 = (inp[2]) ? 11'b00001010000 : 11'b00011010000;
										assign node3454 = (inp[11]) ? node3460 : node3455;
											assign node3455 = (inp[5]) ? 11'b00101100000 : node3456;
												assign node3456 = (inp[2]) ? 11'b00111100010 : 11'b00110000011;
											assign node3460 = (inp[2]) ? 11'b00001000000 : node3461;
												assign node3461 = (inp[5]) ? 11'b00001000000 : 11'b00000100010;
								assign node3465 = (inp[10]) ? node3493 : node3466;
									assign node3466 = (inp[4]) ? node3478 : node3467;
										assign node3467 = (inp[2]) ? node3473 : node3468;
											assign node3468 = (inp[5]) ? node3470 : 11'b00010010001;
												assign node3470 = (inp[11]) ? 11'b00010110010 : 11'b00101010010;
											assign node3473 = (inp[11]) ? 11'b00000010000 : node3474;
												assign node3474 = (inp[5]) ? 11'b00110110000 : 11'b00000110010;
										assign node3478 = (inp[2]) ? node3486 : node3479;
											assign node3479 = (inp[5]) ? node3483 : node3480;
												assign node3480 = (inp[11]) ? 11'b00111000000 : 11'b00110000011;
												assign node3483 = (inp[11]) ? 11'b00010000000 : 11'b00011100000;
											assign node3486 = (inp[11]) ? node3490 : node3487;
												assign node3487 = (inp[5]) ? 11'b00000100000 : 11'b00100100010;
												assign node3490 = (inp[5]) ? 11'b00000000000 : 11'b00100000000;
									assign node3493 = (inp[11]) ? node3501 : node3494;
										assign node3494 = (inp[5]) ? 11'b00000100000 : node3495;
											assign node3495 = (inp[2]) ? 11'b00000100010 : node3496;
												assign node3496 = (inp[4]) ? 11'b00001100010 : 11'b00000000001;
										assign node3501 = (inp[2]) ? node3509 : node3502;
											assign node3502 = (inp[4]) ? node3506 : node3503;
												assign node3503 = (inp[5]) ? 11'b00000100010 : 11'b00011100010;
												assign node3506 = (inp[5]) ? 11'b00000000000 : 11'b00001000000;
											assign node3509 = (inp[5]) ? 11'b00000000000 : node3510;
												assign node3510 = (inp[4]) ? 11'b00000000000 : 11'b00010000000;
		assign node3514 = (inp[7]) ? node5290 : node3515;
			assign node3515 = (inp[6]) ? node4407 : node3516;
				assign node3516 = (inp[8]) ? node3956 : node3517;
					assign node3517 = (inp[0]) ? node3739 : node3518;
						assign node3518 = (inp[9]) ? node3632 : node3519;
							assign node3519 = (inp[4]) ? node3575 : node3520;
								assign node3520 = (inp[2]) ? node3548 : node3521;
									assign node3521 = (inp[10]) ? node3537 : node3522;
										assign node3522 = (inp[3]) ? node3530 : node3523;
											assign node3523 = (inp[5]) ? node3527 : node3524;
												assign node3524 = (inp[11]) ? 11'b00001001011 : 11'b00001101011;
												assign node3527 = (inp[11]) ? 11'b00000111001 : 11'b00000011001;
											assign node3530 = (inp[11]) ? node3534 : node3531;
												assign node3531 = (inp[5]) ? 11'b10001111011 : 11'b10001101001;
												assign node3534 = (inp[5]) ? 11'b10101001011 : 11'b10001011001;
										assign node3537 = (inp[3]) ? node3541 : node3538;
											assign node3538 = (inp[5]) ? 11'b10101011001 : 11'b10001101011;
											assign node3541 = (inp[5]) ? node3545 : node3542;
												assign node3542 = (inp[11]) ? 11'b00001011101 : 11'b00001101101;
												assign node3545 = (inp[11]) ? 11'b00011001111 : 11'b00101111111;
									assign node3548 = (inp[11]) ? node3562 : node3549;
										assign node3549 = (inp[5]) ? node3557 : node3550;
											assign node3550 = (inp[10]) ? node3554 : node3551;
												assign node3551 = (inp[3]) ? 11'b10101001000 : 11'b00101001010;
												assign node3554 = (inp[3]) ? 11'b00111001100 : 11'b10111001010;
											assign node3557 = (inp[3]) ? node3559 : 11'b10010011001;
												assign node3559 = (inp[10]) ? 11'b00000011111 : 11'b10100011011;
										assign node3562 = (inp[10]) ? node3568 : node3563;
											assign node3563 = (inp[3]) ? 11'b10110111001 : node3564;
												assign node3564 = (inp[5]) ? 11'b00101111001 : 11'b00100101011;
											assign node3568 = (inp[3]) ? node3572 : node3569;
												assign node3569 = (inp[5]) ? 11'b10001111011 : 11'b10111101011;
												assign node3572 = (inp[5]) ? 11'b00101101101 : 11'b00101111111;
								assign node3575 = (inp[3]) ? node3607 : node3576;
									assign node3576 = (inp[10]) ? node3592 : node3577;
										assign node3577 = (inp[2]) ? node3585 : node3578;
											assign node3578 = (inp[5]) ? node3582 : node3579;
												assign node3579 = (inp[11]) ? 11'b00011001111 : 11'b00001101111;
												assign node3582 = (inp[11]) ? 11'b00000011111 : 11'b00010111101;
											assign node3585 = (inp[11]) ? node3589 : node3586;
												assign node3586 = (inp[5]) ? 11'b00111011111 : 11'b00100001100;
												assign node3589 = (inp[5]) ? 11'b00100111101 : 11'b00110101101;
										assign node3592 = (inp[5]) ? node3600 : node3593;
											assign node3593 = (inp[11]) ? node3597 : node3594;
												assign node3594 = (inp[2]) ? 11'b10111111101 : 11'b10001111111;
												assign node3597 = (inp[2]) ? 11'b10000111111 : 11'b10111011111;
											assign node3600 = (inp[2]) ? node3604 : node3601;
												assign node3601 = (inp[11]) ? 11'b10001001111 : 11'b10011101101;
												assign node3604 = (inp[11]) ? 11'b10111101101 : 11'b10100001111;
									assign node3607 = (inp[10]) ? node3619 : node3608;
										assign node3608 = (inp[2]) ? node3614 : node3609;
											assign node3609 = (inp[11]) ? node3611 : 11'b10111111111;
												assign node3611 = (inp[5]) ? 11'b10100011101 : 11'b10111001101;
											assign node3614 = (inp[5]) ? node3616 : 11'b10000101101;
												assign node3616 = (inp[11]) ? 11'b10011111111 : 11'b10001011101;
										assign node3619 = (inp[5]) ? node3625 : node3620;
											assign node3620 = (inp[11]) ? 11'b00111011001 : node3621;
												assign node3621 = (inp[2]) ? 11'b00001101001 : 11'b00101101001;
											assign node3625 = (inp[11]) ? node3629 : node3626;
												assign node3626 = (inp[2]) ? 11'b00110011001 : 11'b00011111011;
												assign node3629 = (inp[2]) ? 11'b00001101011 : 11'b00101001001;
							assign node3632 = (inp[4]) ? node3686 : node3633;
								assign node3633 = (inp[3]) ? node3659 : node3634;
									assign node3634 = (inp[10]) ? node3646 : node3635;
										assign node3635 = (inp[11]) ? node3641 : node3636;
											assign node3636 = (inp[5]) ? node3638 : 11'b00000101011;
												assign node3638 = (inp[2]) ? 11'b00100011001 : 11'b00001111001;
											assign node3641 = (inp[2]) ? node3643 : 11'b00111001001;
												assign node3643 = (inp[5]) ? 11'b00010101011 : 11'b00011111001;
										assign node3646 = (inp[5]) ? node3654 : node3647;
											assign node3647 = (inp[2]) ? node3651 : node3648;
												assign node3648 = (inp[11]) ? 11'b10100011111 : 11'b10000111111;
												assign node3651 = (inp[11]) ? 11'b10001111101 : 11'b10110011100;
											assign node3654 = (inp[2]) ? node3656 : 11'b10100101101;
												assign node3656 = (inp[11]) ? 11'b10010101111 : 11'b10001001111;
									assign node3659 = (inp[10]) ? node3673 : node3660;
										assign node3660 = (inp[5]) ? node3668 : node3661;
											assign node3661 = (inp[2]) ? node3665 : node3662;
												assign node3662 = (inp[11]) ? 11'b10100001101 : 11'b10000101101;
												assign node3665 = (inp[11]) ? 11'b10011101111 : 11'b10100001110;
											assign node3668 = (inp[2]) ? node3670 : 11'b10010011111;
												assign node3670 = (inp[11]) ? 11'b10100111101 : 11'b10111011111;
										assign node3673 = (inp[5]) ? node3679 : node3674;
											assign node3674 = (inp[2]) ? node3676 : 11'b00010011101;
												assign node3676 = (inp[11]) ? 11'b00100111111 : 11'b00110011110;
											assign node3679 = (inp[2]) ? node3683 : node3680;
												assign node3680 = (inp[11]) ? 11'b00000001101 : 11'b00010101111;
												assign node3683 = (inp[11]) ? 11'b00110101101 : 11'b00101001101;
								assign node3686 = (inp[11]) ? node3716 : node3687;
									assign node3687 = (inp[2]) ? node3701 : node3688;
										assign node3688 = (inp[3]) ? node3694 : node3689;
											assign node3689 = (inp[5]) ? 11'b00111111101 : node3690;
												assign node3690 = (inp[10]) ? 11'b10100101011 : 11'b00100101111;
											assign node3694 = (inp[5]) ? node3698 : node3695;
												assign node3695 = (inp[10]) ? 11'b00100111001 : 11'b10100111001;
												assign node3698 = (inp[10]) ? 11'b00100101011 : 11'b10000101011;
										assign node3701 = (inp[5]) ? node3709 : node3702;
											assign node3702 = (inp[3]) ? node3706 : node3703;
												assign node3703 = (inp[10]) ? 11'b10010101011 : 11'b00001101111;
												assign node3706 = (inp[10]) ? 11'b00000111001 : 11'b10011111001;
											assign node3709 = (inp[3]) ? node3713 : node3710;
												assign node3710 = (inp[10]) ? 11'b10110011001 : 11'b00000011101;
												assign node3713 = (inp[10]) ? 11'b00001101011 : 11'b10100001011;
									assign node3716 = (inp[5]) ? node3732 : node3717;
										assign node3717 = (inp[3]) ? node3725 : node3718;
											assign node3718 = (inp[10]) ? node3722 : node3719;
												assign node3719 = (inp[2]) ? 11'b00111011111 : 11'b00010011111;
												assign node3722 = (inp[2]) ? 11'b10011011011 : 11'b10110011011;
											assign node3725 = (inp[10]) ? node3729 : node3726;
												assign node3726 = (inp[2]) ? 11'b10101011001 : 11'b10010011001;
												assign node3729 = (inp[2]) ? 11'b00011011001 : 11'b00110011001;
										assign node3732 = (inp[10]) ? node3736 : node3733;
											assign node3733 = (inp[3]) ? 11'b10111001001 : 11'b00111101101;
											assign node3736 = (inp[3]) ? 11'b00110001001 : 11'b10100101011;
						assign node3739 = (inp[3]) ? node3859 : node3740;
							assign node3740 = (inp[9]) ? node3802 : node3741;
								assign node3741 = (inp[10]) ? node3771 : node3742;
									assign node3742 = (inp[11]) ? node3756 : node3743;
										assign node3743 = (inp[2]) ? node3749 : node3744;
											assign node3744 = (inp[4]) ? node3746 : 11'b00001101011;
												assign node3746 = (inp[5]) ? 11'b00111101011 : 11'b00001101011;
											assign node3749 = (inp[4]) ? node3753 : node3750;
												assign node3750 = (inp[5]) ? 11'b00000001011 : 11'b00001001010;
												assign node3753 = (inp[5]) ? 11'b00111001001 : 11'b00000001000;
										assign node3756 = (inp[5]) ? node3764 : node3757;
											assign node3757 = (inp[2]) ? node3761 : node3758;
												assign node3758 = (inp[4]) ? 11'b00011011011 : 11'b00001011011;
												assign node3761 = (inp[4]) ? 11'b00010111001 : 11'b00010111011;
											assign node3764 = (inp[4]) ? node3768 : node3765;
												assign node3765 = (inp[2]) ? 11'b00011111001 : 11'b00000111001;
												assign node3768 = (inp[2]) ? 11'b00101111011 : 11'b00100011001;
									assign node3771 = (inp[11]) ? node3787 : node3772;
										assign node3772 = (inp[2]) ? node3780 : node3773;
											assign node3773 = (inp[4]) ? node3777 : node3774;
												assign node3774 = (inp[5]) ? 11'b00101101111 : 11'b00001101111;
												assign node3777 = (inp[5]) ? 11'b00011111111 : 11'b00001111111;
											assign node3780 = (inp[5]) ? node3784 : node3781;
												assign node3781 = (inp[4]) ? 11'b00011111101 : 11'b00011001110;
												assign node3784 = (inp[4]) ? 11'b00010011111 : 11'b00110001111;
										assign node3787 = (inp[4]) ? node3795 : node3788;
											assign node3788 = (inp[5]) ? node3792 : node3789;
												assign node3789 = (inp[2]) ? 11'b00001111111 : 11'b00001011111;
												assign node3792 = (inp[2]) ? 11'b00001111101 : 11'b00011011101;
											assign node3795 = (inp[2]) ? node3799 : node3796;
												assign node3796 = (inp[5]) ? 11'b00101001101 : 11'b00111001111;
												assign node3799 = (inp[5]) ? 11'b00101101101 : 11'b00100101101;
								assign node3802 = (inp[10]) ? node3830 : node3803;
									assign node3803 = (inp[11]) ? node3815 : node3804;
										assign node3804 = (inp[4]) ? node3808 : node3805;
											assign node3805 = (inp[2]) ? 11'b00010001101 : 11'b00000101111;
											assign node3808 = (inp[5]) ? node3812 : node3809;
												assign node3809 = (inp[2]) ? 11'b00101111101 : 11'b00100111111;
												assign node3812 = (inp[2]) ? 11'b00100011111 : 11'b00110111111;
										assign node3815 = (inp[5]) ? node3823 : node3816;
											assign node3816 = (inp[4]) ? node3820 : node3817;
												assign node3817 = (inp[2]) ? 11'b00111111111 : 11'b00100011111;
												assign node3820 = (inp[2]) ? 11'b00001001111 : 11'b00010001111;
											assign node3823 = (inp[2]) ? node3827 : node3824;
												assign node3824 = (inp[4]) ? 11'b00111001101 : 11'b00111011101;
												assign node3827 = (inp[4]) ? 11'b00111101101 : 11'b00110111101;
									assign node3830 = (inp[11]) ? node3846 : node3831;
										assign node3831 = (inp[2]) ? node3839 : node3832;
											assign node3832 = (inp[4]) ? node3836 : node3833;
												assign node3833 = (inp[5]) ? 11'b00100111011 : 11'b00000111011;
												assign node3836 = (inp[5]) ? 11'b00100111001 : 11'b00100111011;
											assign node3839 = (inp[4]) ? node3843 : node3840;
												assign node3840 = (inp[5]) ? 11'b00101011001 : 11'b00010011010;
												assign node3843 = (inp[5]) ? 11'b00111111011 : 11'b00110111001;
										assign node3846 = (inp[5]) ? node3854 : node3847;
											assign node3847 = (inp[2]) ? node3851 : node3848;
												assign node3848 = (inp[4]) ? 11'b00110001011 : 11'b00010001011;
												assign node3851 = (inp[4]) ? 11'b00111001011 : 11'b00001101001;
											assign node3854 = (inp[2]) ? node3856 : 11'b00110001001;
												assign node3856 = (inp[4]) ? 11'b00110101001 : 11'b00110101011;
							assign node3859 = (inp[9]) ? node3913 : node3860;
								assign node3860 = (inp[4]) ? node3882 : node3861;
									assign node3861 = (inp[5]) ? node3873 : node3862;
										assign node3862 = (inp[2]) ? node3866 : node3863;
											assign node3863 = (inp[11]) ? 11'b00001001001 : 11'b00001101001;
											assign node3866 = (inp[11]) ? node3870 : node3867;
												assign node3867 = (inp[10]) ? 11'b00001001000 : 11'b00011001000;
												assign node3870 = (inp[10]) ? 11'b00101101001 : 11'b00010101001;
										assign node3873 = (inp[2]) ? node3879 : node3874;
											assign node3874 = (inp[11]) ? 11'b00111001011 : node3875;
												assign node3875 = (inp[10]) ? 11'b00001101001 : 11'b00101101001;
											assign node3879 = (inp[11]) ? 11'b00110101011 : 11'b00110001001;
									assign node3882 = (inp[10]) ? node3898 : node3883;
										assign node3883 = (inp[5]) ? node3891 : node3884;
											assign node3884 = (inp[2]) ? node3888 : node3885;
												assign node3885 = (inp[11]) ? 11'b00111011001 : 11'b00001111001;
												assign node3888 = (inp[11]) ? 11'b00100111011 : 11'b00011111011;
											assign node3891 = (inp[11]) ? node3895 : node3892;
												assign node3892 = (inp[2]) ? 11'b00101011001 : 11'b00111111001;
												assign node3895 = (inp[2]) ? 11'b00011111001 : 11'b00001011011;
										assign node3898 = (inp[11]) ? node3906 : node3899;
											assign node3899 = (inp[5]) ? node3903 : node3900;
												assign node3900 = (inp[2]) ? 11'b00101101011 : 11'b00101101001;
												assign node3903 = (inp[2]) ? 11'b00110001001 : 11'b00111101001;
											assign node3906 = (inp[5]) ? node3910 : node3907;
												assign node3907 = (inp[2]) ? 11'b00011001011 : 11'b00011001001;
												assign node3910 = (inp[2]) ? 11'b00011101011 : 11'b00011001011;
								assign node3913 = (inp[10]) ? node3933 : node3914;
									assign node3914 = (inp[4]) ? node3924 : node3915;
										assign node3915 = (inp[2]) ? node3919 : node3916;
											assign node3916 = (inp[11]) ? 11'b00010011011 : 11'b00000111001;
											assign node3919 = (inp[11]) ? node3921 : 11'b00111011011;
												assign node3921 = (inp[5]) ? 11'b00000111001 : 11'b00111111001;
										assign node3924 = (inp[5]) ? node3928 : node3925;
											assign node3925 = (inp[11]) ? 11'b00110001001 : 11'b00100101001;
											assign node3928 = (inp[11]) ? 11'b00000101011 : node3929;
												assign node3929 = (inp[2]) ? 11'b00010001001 : 11'b00000101011;
									assign node3933 = (inp[4]) ? node3949 : node3934;
										assign node3934 = (inp[2]) ? node3942 : node3935;
											assign node3935 = (inp[11]) ? node3939 : node3936;
												assign node3936 = (inp[5]) ? 11'b00010101001 : 11'b00000101001;
												assign node3939 = (inp[5]) ? 11'b00000001011 : 11'b00010001001;
											assign node3942 = (inp[11]) ? node3946 : node3943;
												assign node3943 = (inp[5]) ? 11'b00011001011 : 11'b00000001010;
												assign node3946 = (inp[5]) ? 11'b00000101001 : 11'b00010101011;
										assign node3949 = (inp[11]) ? node3953 : node3950;
											assign node3950 = (inp[5]) ? 11'b00000101011 : 11'b00000101001;
											assign node3953 = (inp[2]) ? 11'b00001001001 : 11'b00000001001;
					assign node3956 = (inp[0]) ? node4178 : node3957;
						assign node3957 = (inp[2]) ? node4069 : node3958;
							assign node3958 = (inp[11]) ? node4014 : node3959;
								assign node3959 = (inp[9]) ? node3985 : node3960;
									assign node3960 = (inp[4]) ? node3976 : node3961;
										assign node3961 = (inp[5]) ? node3969 : node3962;
											assign node3962 = (inp[10]) ? node3966 : node3963;
												assign node3963 = (inp[3]) ? 11'b10100001001 : 11'b00000001011;
												assign node3966 = (inp[3]) ? 11'b00101101100 : 11'b10001101010;
											assign node3969 = (inp[3]) ? node3973 : node3970;
												assign node3970 = (inp[10]) ? 11'b10100011000 : 11'b00001011000;
												assign node3973 = (inp[10]) ? 11'b00110011110 : 11'b10000011010;
										assign node3976 = (inp[3]) ? 11'b10010111110 : node3977;
											assign node3977 = (inp[10]) ? node3981 : node3978;
												assign node3978 = (inp[5]) ? 11'b00111111100 : 11'b00100101100;
												assign node3981 = (inp[5]) ? 11'b10000101110 : 11'b10100111100;
									assign node3985 = (inp[4]) ? node4001 : node3986;
										assign node3986 = (inp[3]) ? node3994 : node3987;
											assign node3987 = (inp[10]) ? node3991 : node3988;
												assign node3988 = (inp[5]) ? 11'b00010011000 : 11'b00011101010;
												assign node3991 = (inp[5]) ? 11'b10001101100 : 11'b10010111110;
											assign node3994 = (inp[5]) ? node3998 : node3995;
												assign node3995 = (inp[10]) ? 11'b00110111100 : 11'b10111101100;
												assign node3998 = (inp[10]) ? 11'b00101101110 : 11'b10001111110;
										assign node4001 = (inp[10]) ? node4007 : node4002;
											assign node4002 = (inp[3]) ? 11'b10011111010 : node4003;
												assign node4003 = (inp[5]) ? 11'b00100111110 : 11'b00111101100;
											assign node4007 = (inp[3]) ? node4011 : node4008;
												assign node4008 = (inp[5]) ? 11'b10111111010 : 11'b10001101000;
												assign node4011 = (inp[5]) ? 11'b00101101000 : 11'b00100111010;
								assign node4014 = (inp[4]) ? node4040 : node4015;
									assign node4015 = (inp[9]) ? node4029 : node4016;
										assign node4016 = (inp[10]) ? node4024 : node4017;
											assign node4017 = (inp[3]) ? node4021 : node4018;
												assign node4018 = (inp[5]) ? 11'b00001111010 : 11'b00000101000;
												assign node4021 = (inp[5]) ? 11'b10011101000 : 11'b10100111010;
											assign node4024 = (inp[3]) ? 11'b00011011110 : node4025;
												assign node4025 = (inp[5]) ? 11'b10010111010 : 11'b10110101000;
										assign node4029 = (inp[5]) ? node4033 : node4030;
											assign node4030 = (inp[3]) ? 11'b10101001100 : 11'b10001011110;
											assign node4033 = (inp[10]) ? node4037 : node4034;
												assign node4034 = (inp[3]) ? 11'b10100111110 : 11'b00000101000;
												assign node4037 = (inp[3]) ? 11'b00111001110 : 11'b10110101100;
									assign node4040 = (inp[10]) ? node4056 : node4041;
										assign node4041 = (inp[3]) ? node4049 : node4042;
											assign node4042 = (inp[5]) ? node4046 : node4043;
												assign node4043 = (inp[9]) ? 11'b00001011110 : 11'b00110001110;
												assign node4046 = (inp[9]) ? 11'b00100001110 : 11'b00101011100;
											assign node4049 = (inp[5]) ? node4053 : node4050;
												assign node4050 = (inp[9]) ? 11'b10011011000 : 11'b10010001100;
												assign node4053 = (inp[9]) ? 11'b10100001000 : 11'b10101011110;
										assign node4056 = (inp[3]) ? node4062 : node4057;
											assign node4057 = (inp[9]) ? node4059 : 11'b10111001100;
												assign node4059 = (inp[5]) ? 11'b10110001010 : 11'b10111011010;
											assign node4062 = (inp[5]) ? node4066 : node4063;
												assign node4063 = (inp[9]) ? 11'b00111011000 : 11'b00100011000;
												assign node4066 = (inp[9]) ? 11'b00110001000 : 11'b00110001010;
							assign node4069 = (inp[5]) ? node4123 : node4070;
								assign node4070 = (inp[11]) ? node4094 : node4071;
									assign node4071 = (inp[9]) ? node4083 : node4072;
										assign node4072 = (inp[4]) ? node4078 : node4073;
											assign node4073 = (inp[10]) ? 11'b00001001111 : node4074;
												assign node4074 = (inp[3]) ? 11'b10010101001 : 11'b00100101011;
											assign node4078 = (inp[3]) ? 11'b00100001001 : node4079;
												assign node4079 = (inp[10]) ? 11'b10000011111 : 11'b00000001111;
										assign node4083 = (inp[3]) ? node4091 : node4084;
											assign node4084 = (inp[10]) ? node4088 : node4085;
												assign node4085 = (inp[4]) ? 11'b00011001111 : 11'b00111001001;
												assign node4088 = (inp[4]) ? 11'b10111001001 : 11'b10101011101;
											assign node4091 = (inp[10]) ? 11'b00010011111 : 11'b10101011011;
									assign node4094 = (inp[4]) ? node4108 : node4095;
										assign node4095 = (inp[3]) ? node4103 : node4096;
											assign node4096 = (inp[10]) ? node4100 : node4097;
												assign node4097 = (inp[9]) ? 11'b00000011011 : 11'b00101001001;
												assign node4100 = (inp[9]) ? 11'b10111111110 : 11'b10000001011;
											assign node4103 = (inp[10]) ? 11'b00110011101 : node4104;
												assign node4104 = (inp[9]) ? 11'b10010001101 : 11'b10010011011;
										assign node4108 = (inp[9]) ? node4116 : node4109;
											assign node4109 = (inp[10]) ? node4113 : node4110;
												assign node4110 = (inp[3]) ? 11'b10101101110 : 11'b00011101100;
												assign node4113 = (inp[3]) ? 11'b00001111000 : 11'b10011111100;
											assign node4116 = (inp[3]) ? node4120 : node4117;
												assign node4117 = (inp[10]) ? 11'b10000111010 : 11'b00100111110;
												assign node4120 = (inp[10]) ? 11'b00010111000 : 11'b10110111000;
								assign node4123 = (inp[11]) ? node4149 : node4124;
									assign node4124 = (inp[4]) ? node4138 : node4125;
										assign node4125 = (inp[10]) ? node4131 : node4126;
											assign node4126 = (inp[3]) ? 11'b10101111100 : node4127;
												assign node4127 = (inp[9]) ? 11'b00111111000 : 11'b00100111000;
											assign node4131 = (inp[9]) ? node4135 : node4132;
												assign node4132 = (inp[3]) ? 11'b00011111110 : 11'b10001111000;
												assign node4135 = (inp[3]) ? 11'b00000101100 : 11'b10110101110;
										assign node4138 = (inp[9]) ? node4142 : node4139;
											assign node4139 = (inp[10]) ? 11'b10110101100 : 11'b00010111110;
											assign node4142 = (inp[3]) ? node4146 : node4143;
												assign node4143 = (inp[10]) ? 11'b10011011010 : 11'b00011011100;
												assign node4146 = (inp[10]) ? 11'b00001001000 : 11'b10001001000;
									assign node4149 = (inp[3]) ? node4163 : node4150;
										assign node4150 = (inp[4]) ? node4158 : node4151;
											assign node4151 = (inp[10]) ? node4155 : node4152;
												assign node4152 = (inp[9]) ? 11'b00100001000 : 11'b00100011010;
												assign node4155 = (inp[9]) ? 11'b10001001110 : 11'b10100011000;
											assign node4158 = (inp[10]) ? 11'b10001001100 : node4159;
												assign node4159 = (inp[9]) ? 11'b00000001100 : 11'b00001011110;
										assign node4163 = (inp[10]) ? node4171 : node4164;
											assign node4164 = (inp[9]) ? node4168 : node4165;
												assign node4165 = (inp[4]) ? 11'b10011011100 : 11'b10110001000;
												assign node4168 = (inp[4]) ? 11'b10010001010 : 11'b10011011110;
											assign node4171 = (inp[4]) ? node4175 : node4172;
												assign node4172 = (inp[9]) ? 11'b00011001100 : 11'b00110001110;
												assign node4175 = (inp[9]) ? 11'b00010001000 : 11'b00010001010;
						assign node4178 = (inp[3]) ? node4290 : node4179;
							assign node4179 = (inp[5]) ? node4237 : node4180;
								assign node4180 = (inp[2]) ? node4210 : node4181;
									assign node4181 = (inp[11]) ? node4197 : node4182;
										assign node4182 = (inp[9]) ? node4190 : node4183;
											assign node4183 = (inp[10]) ? node4187 : node4184;
												assign node4184 = (inp[4]) ? 11'b00100101010 : 11'b00100001011;
												assign node4187 = (inp[4]) ? 11'b00101111110 : 11'b00101101110;
											assign node4190 = (inp[4]) ? node4194 : node4191;
												assign node4191 = (inp[10]) ? 11'b00110111010 : 11'b00111101110;
												assign node4194 = (inp[10]) ? 11'b00001111000 : 11'b00011111110;
										assign node4197 = (inp[9]) ? node4205 : node4198;
											assign node4198 = (inp[10]) ? node4202 : node4199;
												assign node4199 = (inp[4]) ? 11'b00110011000 : 11'b00100111000;
												assign node4202 = (inp[4]) ? 11'b00000001110 : 11'b00110111100;
											assign node4205 = (inp[4]) ? 11'b00101001110 : node4206;
												assign node4206 = (inp[10]) ? 11'b00101001000 : 11'b00001011100;
									assign node4210 = (inp[11]) ? node4222 : node4211;
										assign node4211 = (inp[9]) ? node4219 : node4212;
											assign node4212 = (inp[10]) ? node4216 : node4213;
												assign node4213 = (inp[4]) ? 11'b00100001001 : 11'b00100101011;
												assign node4216 = (inp[4]) ? 11'b00100011111 : 11'b00101001111;
											assign node4219 = (inp[10]) ? 11'b00011011011 : 11'b00001011111;
										assign node4222 = (inp[4]) ? node4230 : node4223;
											assign node4223 = (inp[9]) ? node4227 : node4224;
												assign node4224 = (inp[10]) ? 11'b00100011101 : 11'b00111011001;
												assign node4227 = (inp[10]) ? 11'b00101101010 : 11'b00000011111;
											assign node4230 = (inp[9]) ? node4234 : node4231;
												assign node4231 = (inp[10]) ? 11'b00011101100 : 11'b00111111010;
												assign node4234 = (inp[10]) ? 11'b00010101010 : 11'b00110101100;
								assign node4237 = (inp[11]) ? node4263 : node4238;
									assign node4238 = (inp[4]) ? node4252 : node4239;
										assign node4239 = (inp[10]) ? node4245 : node4240;
											assign node4240 = (inp[9]) ? node4242 : 11'b00101101010;
												assign node4242 = (inp[2]) ? 11'b00101101100 : 11'b00111101110;
											assign node4245 = (inp[9]) ? node4249 : node4246;
												assign node4246 = (inp[2]) ? 11'b00001101100 : 11'b00010001110;
												assign node4249 = (inp[2]) ? 11'b00000111010 : 11'b00001111000;
										assign node4252 = (inp[10]) ? node4260 : node4253;
											assign node4253 = (inp[9]) ? node4257 : node4254;
												assign node4254 = (inp[2]) ? 11'b00000101010 : 11'b00011101000;
												assign node4257 = (inp[2]) ? 11'b00011011100 : 11'b00010111100;
											assign node4260 = (inp[9]) ? 11'b00001111010 : 11'b00111011110;
									assign node4263 = (inp[9]) ? node4277 : node4264;
										assign node4264 = (inp[4]) ? node4272 : node4265;
											assign node4265 = (inp[10]) ? node4269 : node4266;
												assign node4266 = (inp[2]) ? 11'b00110011010 : 11'b00101111010;
												assign node4269 = (inp[2]) ? 11'b00110011110 : 11'b00110111110;
											assign node4272 = (inp[10]) ? 11'b00011001100 : node4273;
												assign node4273 = (inp[2]) ? 11'b00011011010 : 11'b00001011000;
										assign node4277 = (inp[10]) ? node4285 : node4278;
											assign node4278 = (inp[4]) ? node4282 : node4279;
												assign node4279 = (inp[2]) ? 11'b00010011100 : 11'b00000111110;
												assign node4282 = (inp[2]) ? 11'b00010001100 : 11'b00000001100;
											assign node4285 = (inp[4]) ? 11'b00010001000 : node4286;
												assign node4286 = (inp[2]) ? 11'b00011001000 : 11'b00011001010;
							assign node4290 = (inp[10]) ? node4350 : node4291;
								assign node4291 = (inp[2]) ? node4319 : node4292;
									assign node4292 = (inp[11]) ? node4304 : node4293;
										assign node4293 = (inp[9]) ? node4299 : node4294;
											assign node4294 = (inp[4]) ? 11'b00000111000 : node4295;
												assign node4295 = (inp[5]) ? 11'b00100001000 : 11'b00000001001;
											assign node4299 = (inp[5]) ? 11'b00101111010 : node4300;
												assign node4300 = (inp[4]) ? 11'b00111101000 : 11'b00011111000;
										assign node4304 = (inp[4]) ? node4312 : node4305;
											assign node4305 = (inp[5]) ? node4309 : node4306;
												assign node4306 = (inp[9]) ? 11'b00101011010 : 11'b00010101010;
												assign node4309 = (inp[9]) ? 11'b00010111000 : 11'b00111101000;
											assign node4312 = (inp[9]) ? node4316 : node4313;
												assign node4313 = (inp[5]) ? 11'b00011011010 : 11'b00110011010;
												assign node4316 = (inp[5]) ? 11'b00010001010 : 11'b00111001000;
									assign node4319 = (inp[5]) ? node4335 : node4320;
										assign node4320 = (inp[9]) ? node4328 : node4321;
											assign node4321 = (inp[11]) ? node4325 : node4322;
												assign node4322 = (inp[4]) ? 11'b00010011011 : 11'b00010101001;
												assign node4325 = (inp[4]) ? 11'b00101111010 : 11'b00000001011;
											assign node4328 = (inp[4]) ? node4332 : node4329;
												assign node4329 = (inp[11]) ? 11'b00110011001 : 11'b00001011011;
												assign node4332 = (inp[11]) ? 11'b00100101000 : 11'b00101001001;
										assign node4335 = (inp[9]) ? node4343 : node4336;
											assign node4336 = (inp[11]) ? node4340 : node4337;
												assign node4337 = (inp[4]) ? 11'b00100111000 : 11'b00111101000;
												assign node4340 = (inp[4]) ? 11'b00001011000 : 11'b00100001000;
											assign node4343 = (inp[4]) ? node4347 : node4344;
												assign node4344 = (inp[11]) ? 11'b00001011010 : 11'b00110111010;
												assign node4347 = (inp[11]) ? 11'b00000001010 : 11'b00001001010;
								assign node4350 = (inp[9]) ? node4380 : node4351;
									assign node4351 = (inp[5]) ? node4365 : node4352;
										assign node4352 = (inp[2]) ? node4358 : node4353;
											assign node4353 = (inp[11]) ? 11'b00111001010 : node4354;
												assign node4354 = (inp[4]) ? 11'b00111101000 : 11'b00011101000;
											assign node4358 = (inp[11]) ? node4362 : node4359;
												assign node4359 = (inp[4]) ? 11'b00110001001 : 11'b00011001001;
												assign node4362 = (inp[4]) ? 11'b00000101010 : 11'b00110001011;
										assign node4365 = (inp[2]) ? node4373 : node4366;
											assign node4366 = (inp[4]) ? node4370 : node4367;
												assign node4367 = (inp[11]) ? 11'b00100101000 : 11'b00010001000;
												assign node4370 = (inp[11]) ? 11'b00000001010 : 11'b00100101010;
											assign node4373 = (inp[11]) ? node4377 : node4374;
												assign node4374 = (inp[4]) ? 11'b00101001010 : 11'b00011101010;
												assign node4377 = (inp[4]) ? 11'b00000001010 : 11'b00100001010;
									assign node4380 = (inp[11]) ? node4396 : node4381;
										assign node4381 = (inp[5]) ? node4389 : node4382;
											assign node4382 = (inp[2]) ? node4386 : node4383;
												assign node4383 = (inp[4]) ? 11'b00000101010 : 11'b00000101000;
												assign node4386 = (inp[4]) ? 11'b00001001011 : 11'b00000001011;
											assign node4389 = (inp[4]) ? node4393 : node4390;
												assign node4390 = (inp[2]) ? 11'b00010101000 : 11'b00011101010;
												assign node4393 = (inp[2]) ? 11'b00001001000 : 11'b00001101000;
										assign node4396 = (inp[4]) ? node4404 : node4397;
											assign node4397 = (inp[5]) ? node4401 : node4398;
												assign node4398 = (inp[2]) ? 11'b00011101000 : 11'b00010001010;
												assign node4401 = (inp[2]) ? 11'b00001001000 : 11'b00001001010;
											assign node4404 = (inp[5]) ? 11'b00000001000 : 11'b00001001000;
				assign node4407 = (inp[2]) ? node4853 : node4408;
					assign node4408 = (inp[8]) ? node4628 : node4409;
						assign node4409 = (inp[5]) ? node4523 : node4410;
							assign node4410 = (inp[11]) ? node4464 : node4411;
								assign node4411 = (inp[4]) ? node4437 : node4412;
									assign node4412 = (inp[9]) ? node4426 : node4413;
										assign node4413 = (inp[0]) ? node4421 : node4414;
											assign node4414 = (inp[3]) ? node4418 : node4415;
												assign node4415 = (inp[10]) ? 11'b10001101000 : 11'b00001101010;
												assign node4418 = (inp[10]) ? 11'b00011101110 : 11'b10011101000;
											assign node4421 = (inp[3]) ? 11'b00001101010 : node4422;
												assign node4422 = (inp[10]) ? 11'b00011101110 : 11'b00011101010;
										assign node4426 = (inp[3]) ? node4432 : node4427;
											assign node4427 = (inp[10]) ? 11'b00010111000 : node4428;
												assign node4428 = (inp[0]) ? 11'b00011101100 : 11'b00001101000;
											assign node4432 = (inp[0]) ? node4434 : 11'b00010111100;
												assign node4434 = (inp[10]) ? 11'b00000101000 : 11'b00000111010;
									assign node4437 = (inp[9]) ? node4449 : node4438;
										assign node4438 = (inp[0]) ? node4442 : node4439;
											assign node4439 = (inp[3]) ? 11'b10010101100 : 11'b10000111100;
											assign node4442 = (inp[3]) ? node4446 : node4443;
												assign node4443 = (inp[10]) ? 11'b00011111110 : 11'b00010101010;
												assign node4446 = (inp[10]) ? 11'b00101101010 : 11'b00000111000;
										assign node4449 = (inp[0]) ? node4457 : node4450;
											assign node4450 = (inp[3]) ? node4454 : node4451;
												assign node4451 = (inp[10]) ? 11'b10101101010 : 11'b00101101100;
												assign node4454 = (inp[10]) ? 11'b00111111000 : 11'b10111111010;
											assign node4457 = (inp[3]) ? node4461 : node4458;
												assign node4458 = (inp[10]) ? 11'b00111111000 : 11'b00111111100;
												assign node4461 = (inp[10]) ? 11'b00001101000 : 11'b00101101010;
								assign node4464 = (inp[0]) ? node4496 : node4465;
									assign node4465 = (inp[4]) ? node4481 : node4466;
										assign node4466 = (inp[9]) ? node4474 : node4467;
											assign node4467 = (inp[3]) ? node4471 : node4468;
												assign node4468 = (inp[10]) ? 11'b10010101000 : 11'b00010101010;
												assign node4471 = (inp[10]) ? 11'b00000111110 : 11'b10000111010;
											assign node4474 = (inp[10]) ? node4478 : node4475;
												assign node4475 = (inp[3]) ? 11'b10100101100 : 11'b00110111000;
												assign node4478 = (inp[3]) ? 11'b00001011100 : 11'b10111011110;
										assign node4481 = (inp[10]) ? node4489 : node4482;
											assign node4482 = (inp[9]) ? node4486 : node4483;
												assign node4483 = (inp[3]) ? 11'b10101001110 : 11'b00011001110;
												assign node4486 = (inp[3]) ? 11'b10010011000 : 11'b00000011110;
											assign node4489 = (inp[3]) ? node4493 : node4490;
												assign node4490 = (inp[9]) ? 11'b10100011010 : 11'b10111011100;
												assign node4493 = (inp[9]) ? 11'b00110011000 : 11'b00100011010;
									assign node4496 = (inp[10]) ? node4512 : node4497;
										assign node4497 = (inp[4]) ? node4505 : node4498;
											assign node4498 = (inp[9]) ? node4502 : node4499;
												assign node4499 = (inp[3]) ? 11'b00000101000 : 11'b00010111010;
												assign node4502 = (inp[3]) ? 11'b00101011010 : 11'b00110111100;
											assign node4505 = (inp[3]) ? node4509 : node4506;
												assign node4506 = (inp[9]) ? 11'b00000001100 : 11'b00001011010;
												assign node4509 = (inp[9]) ? 11'b00110001010 : 11'b00111011000;
										assign node4512 = (inp[9]) ? node4516 : node4513;
											assign node4513 = (inp[4]) ? 11'b00010001010 : 11'b00100101010;
											assign node4516 = (inp[4]) ? node4520 : node4517;
												assign node4517 = (inp[3]) ? 11'b00011001000 : 11'b00001001010;
												assign node4520 = (inp[3]) ? 11'b00000001000 : 11'b00100001010;
							assign node4523 = (inp[11]) ? node4577 : node4524;
								assign node4524 = (inp[4]) ? node4554 : node4525;
									assign node4525 = (inp[0]) ? node4539 : node4526;
										assign node4526 = (inp[10]) ? node4532 : node4527;
											assign node4527 = (inp[3]) ? node4529 : 11'b00011011010;
												assign node4529 = (inp[9]) ? 11'b10001011100 : 11'b10011011010;
											assign node4532 = (inp[9]) ? node4536 : node4533;
												assign node4533 = (inp[3]) ? 11'b00111011110 : 11'b10101011000;
												assign node4536 = (inp[3]) ? 11'b00000001110 : 11'b10110001110;
										assign node4539 = (inp[9]) ? node4547 : node4540;
											assign node4540 = (inp[3]) ? node4544 : node4541;
												assign node4541 = (inp[10]) ? 11'b00111001100 : 11'b00011001010;
												assign node4544 = (inp[10]) ? 11'b00001001010 : 11'b00101001010;
											assign node4547 = (inp[10]) ? node4551 : node4548;
												assign node4548 = (inp[3]) ? 11'b00101011000 : 11'b00011001100;
												assign node4551 = (inp[3]) ? 11'b00010001000 : 11'b00110011010;
									assign node4554 = (inp[9]) ? node4566 : node4555;
										assign node4555 = (inp[0]) ? node4561 : node4556;
											assign node4556 = (inp[10]) ? 11'b10000001110 : node4557;
												assign node4557 = (inp[3]) ? 11'b10100011110 : 11'b00010011100;
											assign node4561 = (inp[10]) ? 11'b00111100011 : node4562;
												assign node4562 = (inp[3]) ? 11'b00110011010 : 11'b00100001000;
										assign node4566 = (inp[3]) ? node4572 : node4567;
											assign node4567 = (inp[10]) ? node4569 : 11'b00101110111;
												assign node4569 = (inp[0]) ? 11'b00111110011 : 11'b10001110001;
											assign node4572 = (inp[10]) ? 11'b00111100011 : node4573;
												assign node4573 = (inp[0]) ? 11'b00001100001 : 11'b10011100001;
								assign node4577 = (inp[3]) ? node4605 : node4578;
									assign node4578 = (inp[9]) ? node4592 : node4579;
										assign node4579 = (inp[10]) ? node4585 : node4580;
											assign node4580 = (inp[4]) ? node4582 : 11'b00011110001;
												assign node4582 = (inp[0]) ? 11'b00111110001 : 11'b00001110111;
											assign node4585 = (inp[4]) ? node4589 : node4586;
												assign node4586 = (inp[0]) ? 11'b00000110111 : 11'b10110110011;
												assign node4589 = (inp[0]) ? 11'b00111100111 : 11'b10011100111;
										assign node4592 = (inp[10]) ? node4600 : node4593;
											assign node4593 = (inp[4]) ? node4597 : node4594;
												assign node4594 = (inp[0]) ? 11'b00100110111 : 11'b00110100011;
												assign node4597 = (inp[0]) ? 11'b00101100101 : 11'b00011100101;
											assign node4600 = (inp[0]) ? 11'b00100100001 : node4601;
												assign node4601 = (inp[4]) ? 11'b10000100011 : 11'b10100100101;
									assign node4605 = (inp[9]) ? node4619 : node4606;
										assign node4606 = (inp[4]) ? node4614 : node4607;
											assign node4607 = (inp[0]) ? node4611 : node4608;
												assign node4608 = (inp[10]) ? 11'b00000100101 : 11'b10101100001;
												assign node4611 = (inp[10]) ? 11'b00110100001 : 11'b00100100011;
											assign node4614 = (inp[0]) ? node4616 : 11'b00101100011;
												assign node4616 = (inp[10]) ? 11'b00011100001 : 11'b00001110001;
										assign node4619 = (inp[4]) ? node4623 : node4620;
											assign node4620 = (inp[0]) ? 11'b00010110001 : 11'b00011100111;
											assign node4623 = (inp[10]) ? node4625 : 11'b00010100011;
												assign node4625 = (inp[0]) ? 11'b00000100001 : 11'b00110100001;
						assign node4628 = (inp[0]) ? node4740 : node4629;
							assign node4629 = (inp[5]) ? node4683 : node4630;
								assign node4630 = (inp[11]) ? node4656 : node4631;
									assign node4631 = (inp[9]) ? node4645 : node4632;
										assign node4632 = (inp[4]) ? node4638 : node4633;
											assign node4633 = (inp[10]) ? 11'b00101000111 : node4634;
												assign node4634 = (inp[3]) ? 11'b10110100001 : 11'b00000100011;
											assign node4638 = (inp[3]) ? node4642 : node4639;
												assign node4639 = (inp[10]) ? 11'b10110010101 : 11'b00101000101;
												assign node4642 = (inp[10]) ? 11'b00000000001 : 11'b10000000111;
										assign node4645 = (inp[4]) ? node4649 : node4646;
											assign node4646 = (inp[10]) ? 11'b00111010101 : 11'b10101000101;
											assign node4649 = (inp[3]) ? node4653 : node4650;
												assign node4650 = (inp[10]) ? 11'b10000000001 : 11'b00110000111;
												assign node4653 = (inp[10]) ? 11'b00111010011 : 11'b10010010001;
									assign node4656 = (inp[4]) ? node4668 : node4657;
										assign node4657 = (inp[10]) ? node4663 : node4658;
											assign node4658 = (inp[3]) ? node4660 : 11'b00101010001;
												assign node4660 = (inp[9]) ? 11'b10110000111 : 11'b10101010001;
											assign node4663 = (inp[9]) ? node4665 : 11'b00011010101;
												assign node4665 = (inp[3]) ? 11'b00100010101 : 11'b10010010101;
										assign node4668 = (inp[9]) ? node4676 : node4669;
											assign node4669 = (inp[10]) ? node4673 : node4670;
												assign node4670 = (inp[3]) ? 11'b10010000101 : 11'b00110000111;
												assign node4673 = (inp[3]) ? 11'b00111110011 : 11'b10100010101;
											assign node4676 = (inp[10]) ? node4680 : node4677;
												assign node4677 = (inp[3]) ? 11'b10001110001 : 11'b00011110101;
												assign node4680 = (inp[3]) ? 11'b00111110001 : 11'b10111110011;
								assign node4683 = (inp[11]) ? node4713 : node4684;
									assign node4684 = (inp[9]) ? node4698 : node4685;
										assign node4685 = (inp[4]) ? node4693 : node4686;
											assign node4686 = (inp[10]) ? node4690 : node4687;
												assign node4687 = (inp[3]) ? 11'b10000110011 : 11'b00001110001;
												assign node4690 = (inp[3]) ? 11'b00100110101 : 11'b10110110001;
											assign node4693 = (inp[10]) ? node4695 : 11'b00111110101;
												assign node4695 = (inp[3]) ? 11'b00001110011 : 11'b10001100111;
										assign node4698 = (inp[4]) ? node4706 : node4699;
											assign node4699 = (inp[10]) ? node4703 : node4700;
												assign node4700 = (inp[3]) ? 11'b10010110101 : 11'b00000110011;
												assign node4703 = (inp[3]) ? 11'b00101100111 : 11'b10010100101;
											assign node4706 = (inp[3]) ? node4710 : node4707;
												assign node4707 = (inp[10]) ? 11'b10100110011 : 11'b00111110101;
												assign node4710 = (inp[10]) ? 11'b00110100001 : 11'b10100100011;
									assign node4713 = (inp[4]) ? node4729 : node4714;
										assign node4714 = (inp[9]) ? node4722 : node4715;
											assign node4715 = (inp[3]) ? node4719 : node4716;
												assign node4716 = (inp[10]) ? 11'b10000110001 : 11'b00010110011;
												assign node4719 = (inp[10]) ? 11'b00011000111 : 11'b10000100011;
											assign node4722 = (inp[3]) ? node4726 : node4723;
												assign node4723 = (inp[10]) ? 11'b10111000111 : 11'b00011000011;
												assign node4726 = (inp[10]) ? 11'b00111000111 : 11'b10101010101;
										assign node4729 = (inp[10]) ? node4735 : node4730;
											assign node4730 = (inp[3]) ? 11'b10100000011 : node4731;
												assign node4731 = (inp[9]) ? 11'b00100000101 : 11'b00101010101;
											assign node4735 = (inp[3]) ? 11'b00110000001 : node4736;
												assign node4736 = (inp[9]) ? 11'b10110000001 : 11'b10110000111;
							assign node4740 = (inp[3]) ? node4800 : node4741;
								assign node4741 = (inp[5]) ? node4771 : node4742;
									assign node4742 = (inp[4]) ? node4758 : node4743;
										assign node4743 = (inp[11]) ? node4751 : node4744;
											assign node4744 = (inp[9]) ? node4748 : node4745;
												assign node4745 = (inp[10]) ? 11'b00111000111 : 11'b00110100011;
												assign node4748 = (inp[10]) ? 11'b00101010011 : 11'b00101000101;
											assign node4751 = (inp[9]) ? node4755 : node4752;
												assign node4752 = (inp[10]) ? 11'b00101010111 : 11'b00111010001;
												assign node4755 = (inp[10]) ? 11'b00110000001 : 11'b00010010111;
										assign node4758 = (inp[10]) ? node4766 : node4759;
											assign node4759 = (inp[9]) ? node4763 : node4760;
												assign node4760 = (inp[11]) ? 11'b00100010011 : 11'b00110000011;
												assign node4763 = (inp[11]) ? 11'b00111100101 : 11'b00000010111;
											assign node4766 = (inp[11]) ? node4768 : 11'b00011010011;
												assign node4768 = (inp[9]) ? 11'b00001100011 : 11'b00011100111;
									assign node4771 = (inp[11]) ? node4787 : node4772;
										assign node4772 = (inp[4]) ? node4780 : node4773;
											assign node4773 = (inp[10]) ? node4777 : node4774;
												assign node4774 = (inp[9]) ? 11'b00100100111 : 11'b00110100011;
												assign node4777 = (inp[9]) ? 11'b00011110011 : 11'b00000100101;
											assign node4780 = (inp[10]) ? node4784 : node4781;
												assign node4781 = (inp[9]) ? 11'b00001110101 : 11'b00001100001;
												assign node4784 = (inp[9]) ? 11'b00010110001 : 11'b00111110111;
										assign node4787 = (inp[10]) ? node4793 : node4788;
											assign node4788 = (inp[9]) ? 11'b00011010101 : node4789;
												assign node4789 = (inp[4]) ? 11'b00011010001 : 11'b00110110011;
											assign node4793 = (inp[9]) ? node4797 : node4794;
												assign node4794 = (inp[4]) ? 11'b00000000111 : 11'b00100110101;
												assign node4797 = (inp[4]) ? 11'b00000000001 : 11'b00001000011;
								assign node4800 = (inp[10]) ? node4830 : node4801;
									assign node4801 = (inp[11]) ? node4815 : node4802;
										assign node4802 = (inp[5]) ? node4810 : node4803;
											assign node4803 = (inp[9]) ? node4807 : node4804;
												assign node4804 = (inp[4]) ? 11'b00000010011 : 11'b00000100001;
												assign node4807 = (inp[4]) ? 11'b00110000001 : 11'b00011010011;
											assign node4810 = (inp[4]) ? 11'b00111110011 : node4811;
												assign node4811 = (inp[9]) ? 11'b00100110001 : 11'b00100100011;
										assign node4815 = (inp[5]) ? node4823 : node4816;
											assign node4816 = (inp[9]) ? node4820 : node4817;
												assign node4817 = (inp[4]) ? 11'b00110010001 : 11'b00011000011;
												assign node4820 = (inp[4]) ? 11'b00111100011 : 11'b00100010011;
											assign node4823 = (inp[4]) ? node4827 : node4824;
												assign node4824 = (inp[9]) ? 11'b00011010001 : 11'b00110100001;
												assign node4827 = (inp[9]) ? 11'b00010000011 : 11'b00010010011;
									assign node4830 = (inp[5]) ? node4844 : node4831;
										assign node4831 = (inp[4]) ? node4839 : node4832;
											assign node4832 = (inp[9]) ? node4836 : node4833;
												assign node4833 = (inp[11]) ? 11'b00111000001 : 11'b00011000011;
												assign node4836 = (inp[11]) ? 11'b00010000011 : 11'b00001000001;
											assign node4839 = (inp[11]) ? 11'b00001100011 : node4840;
												assign node4840 = (inp[9]) ? 11'b00001000011 : 11'b00110000011;
										assign node4844 = (inp[4]) ? node4848 : node4845;
											assign node4845 = (inp[9]) ? 11'b00001000011 : 11'b00101000011;
											assign node4848 = (inp[11]) ? 11'b00000000001 : node4849;
												assign node4849 = (inp[9]) ? 11'b00000100001 : 11'b00101100001;
					assign node4853 = (inp[5]) ? node5077 : node4854;
						assign node4854 = (inp[0]) ? node4964 : node4855;
							assign node4855 = (inp[11]) ? node4903 : node4856;
								assign node4856 = (inp[8]) ? node4876 : node4857;
									assign node4857 = (inp[10]) ? node4865 : node4858;
										assign node4858 = (inp[3]) ? node4860 : 11'b00101000011;
											assign node4860 = (inp[9]) ? node4862 : 11'b10100000101;
												assign node4862 = (inp[4]) ? 11'b10001110010 : 11'b10101000101;
										assign node4865 = (inp[3]) ? node4871 : node4866;
											assign node4866 = (inp[4]) ? 11'b10110010111 : node4867;
												assign node4867 = (inp[9]) ? 11'b10110010111 : 11'b10111000001;
											assign node4871 = (inp[4]) ? 11'b00011110000 : node4872;
												assign node4872 = (inp[9]) ? 11'b00110010111 : 11'b00111000111;
									assign node4876 = (inp[9]) ? node4890 : node4877;
										assign node4877 = (inp[4]) ? node4885 : node4878;
											assign node4878 = (inp[3]) ? node4882 : node4879;
												assign node4879 = (inp[10]) ? 11'b10100000000 : 11'b00100000010;
												assign node4882 = (inp[10]) ? 11'b00000000100 : 11'b10000000010;
											assign node4885 = (inp[3]) ? 11'b10101100100 : node4886;
												assign node4886 = (inp[10]) ? 11'b10001110100 : 11'b00011100110;
										assign node4890 = (inp[4]) ? node4898 : node4891;
											assign node4891 = (inp[10]) ? node4895 : node4892;
												assign node4892 = (inp[3]) ? 11'b10011100100 : 11'b00111100010;
												assign node4895 = (inp[3]) ? 11'b00011110110 : 11'b10111110100;
											assign node4898 = (inp[10]) ? node4900 : 11'b00000100110;
												assign node4900 = (inp[3]) ? 11'b00010110010 : 11'b10110100010;
								assign node4903 = (inp[10]) ? node4935 : node4904;
									assign node4904 = (inp[3]) ? node4920 : node4905;
										assign node4905 = (inp[4]) ? node4913 : node4906;
											assign node4906 = (inp[9]) ? node4910 : node4907;
												assign node4907 = (inp[8]) ? 11'b00110100000 : 11'b00111100010;
												assign node4910 = (inp[8]) ? 11'b00001110000 : 11'b00010110010;
											assign node4913 = (inp[9]) ? node4917 : node4914;
												assign node4914 = (inp[8]) ? 11'b00001100100 : 11'b00110100100;
												assign node4917 = (inp[8]) ? 11'b00110110100 : 11'b00101110100;
										assign node4920 = (inp[4]) ? node4928 : node4921;
											assign node4921 = (inp[9]) ? node4925 : node4922;
												assign node4922 = (inp[8]) ? 11'b10010110000 : 11'b10101110010;
												assign node4925 = (inp[8]) ? 11'b10001100100 : 11'b10010100100;
											assign node4928 = (inp[9]) ? node4932 : node4929;
												assign node4929 = (inp[8]) ? 11'b10110100110 : 11'b10010100100;
												assign node4932 = (inp[8]) ? 11'b10110110010 : 11'b10111110010;
									assign node4935 = (inp[3]) ? node4951 : node4936;
										assign node4936 = (inp[4]) ? node4944 : node4937;
											assign node4937 = (inp[9]) ? node4941 : node4938;
												assign node4938 = (inp[8]) ? 11'b10011100010 : 11'b10101100000;
												assign node4941 = (inp[8]) ? 11'b10101110110 : 11'b10000110100;
											assign node4944 = (inp[8]) ? node4948 : node4945;
												assign node4945 = (inp[9]) ? 11'b10011110010 : 11'b10011110110;
												assign node4948 = (inp[9]) ? 11'b10010110010 : 11'b10010110110;
										assign node4951 = (inp[4]) ? node4959 : node4952;
											assign node4952 = (inp[8]) ? node4956 : node4953;
												assign node4953 = (inp[9]) ? 11'b00100110110 : 11'b00110110110;
												assign node4956 = (inp[9]) ? 11'b00001110110 : 11'b00101110110;
											assign node4959 = (inp[8]) ? 11'b00010110000 : node4960;
												assign node4960 = (inp[9]) ? 11'b00011110000 : 11'b00001110010;
							assign node4964 = (inp[11]) ? node5022 : node4965;
								assign node4965 = (inp[8]) ? node4991 : node4966;
									assign node4966 = (inp[10]) ? node4980 : node4967;
										assign node4967 = (inp[4]) ? node4973 : node4968;
											assign node4968 = (inp[3]) ? node4970 : 11'b00011000101;
												assign node4970 = (inp[9]) ? 11'b00011010001 : 11'b00011000001;
											assign node4973 = (inp[9]) ? node4977 : node4974;
												assign node4974 = (inp[3]) ? 11'b00010010011 : 11'b00010000001;
												assign node4977 = (inp[3]) ? 11'b00111100010 : 11'b00111110110;
										assign node4980 = (inp[3]) ? node4986 : node4981;
											assign node4981 = (inp[9]) ? 11'b00000010011 : node4982;
												assign node4982 = (inp[4]) ? 11'b00000010111 : 11'b00001000101;
											assign node4986 = (inp[4]) ? 11'b00100000001 : node4987;
												assign node4987 = (inp[9]) ? 11'b00000000011 : 11'b00001000011;
									assign node4991 = (inp[9]) ? node5007 : node4992;
										assign node4992 = (inp[4]) ? node5000 : node4993;
											assign node4993 = (inp[3]) ? node4997 : node4994;
												assign node4994 = (inp[10]) ? 11'b00110000100 : 11'b00110000010;
												assign node4997 = (inp[10]) ? 11'b00011100010 : 11'b00010000000;
											assign node5000 = (inp[10]) ? node5004 : node5001;
												assign node5001 = (inp[3]) ? 11'b00011110000 : 11'b00111100000;
												assign node5004 = (inp[3]) ? 11'b00110100010 : 11'b00110110110;
										assign node5007 = (inp[4]) ? node5015 : node5008;
											assign node5008 = (inp[3]) ? node5012 : node5009;
												assign node5009 = (inp[10]) ? 11'b00101110000 : 11'b00101100110;
												assign node5012 = (inp[10]) ? 11'b00001100010 : 11'b00001110000;
											assign node5015 = (inp[3]) ? node5019 : node5016;
												assign node5016 = (inp[10]) ? 11'b00000110010 : 11'b00010110100;
												assign node5019 = (inp[10]) ? 11'b00000100010 : 11'b00100100000;
								assign node5022 = (inp[10]) ? node5052 : node5023;
									assign node5023 = (inp[9]) ? node5037 : node5024;
										assign node5024 = (inp[4]) ? node5032 : node5025;
											assign node5025 = (inp[8]) ? node5029 : node5026;
												assign node5026 = (inp[3]) ? 11'b00011100000 : 11'b00001110010;
												assign node5029 = (inp[3]) ? 11'b00000100000 : 11'b00100110000;
											assign node5032 = (inp[3]) ? node5034 : 11'b00101110000;
												assign node5034 = (inp[8]) ? 11'b00100110010 : 11'b00100110000;
										assign node5037 = (inp[3]) ? node5045 : node5038;
											assign node5038 = (inp[4]) ? node5042 : node5039;
												assign node5039 = (inp[8]) ? 11'b00011110100 : 11'b00100110110;
												assign node5042 = (inp[8]) ? 11'b00100100100 : 11'b00011100100;
											assign node5045 = (inp[4]) ? node5049 : node5046;
												assign node5046 = (inp[8]) ? 11'b00111110010 : 11'b00110110000;
												assign node5049 = (inp[8]) ? 11'b00100100010 : 11'b00101100010;
									assign node5052 = (inp[3]) ? node5066 : node5053;
										assign node5053 = (inp[9]) ? node5059 : node5054;
											assign node5054 = (inp[4]) ? node5056 : 11'b00111110110;
												assign node5056 = (inp[8]) ? 11'b00000100110 : 11'b00111100110;
											assign node5059 = (inp[4]) ? node5063 : node5060;
												assign node5060 = (inp[8]) ? 11'b00111100010 : 11'b00010100010;
												assign node5063 = (inp[8]) ? 11'b00000100010 : 11'b00101100010;
										assign node5066 = (inp[4]) ? node5072 : node5067;
											assign node5067 = (inp[9]) ? node5069 : 11'b00100100010;
												assign node5069 = (inp[8]) ? 11'b00011100000 : 11'b00010100010;
											assign node5072 = (inp[8]) ? 11'b00000100000 : node5073;
												assign node5073 = (inp[9]) ? 11'b00001100000 : 11'b00011100000;
						assign node5077 = (inp[0]) ? node5185 : node5078;
							assign node5078 = (inp[11]) ? node5132 : node5079;
								assign node5079 = (inp[4]) ? node5111 : node5080;
									assign node5080 = (inp[8]) ? node5096 : node5081;
										assign node5081 = (inp[10]) ? node5089 : node5082;
											assign node5082 = (inp[3]) ? node5086 : node5083;
												assign node5083 = (inp[9]) ? 11'b00110110010 : 11'b00101110000;
												assign node5086 = (inp[9]) ? 11'b10100110110 : 11'b10100110010;
											assign node5089 = (inp[3]) ? node5093 : node5090;
												assign node5090 = (inp[9]) ? 11'b10000100100 : 11'b10000110010;
												assign node5093 = (inp[9]) ? 11'b00100100100 : 11'b00010110100;
										assign node5096 = (inp[10]) ? node5104 : node5097;
											assign node5097 = (inp[3]) ? node5101 : node5098;
												assign node5098 = (inp[9]) ? 11'b00101010000 : 11'b00100110000;
												assign node5101 = (inp[9]) ? 11'b10101010110 : 11'b10101010010;
											assign node5104 = (inp[3]) ? node5108 : node5105;
												assign node5105 = (inp[9]) ? 11'b10101000110 : 11'b10001010010;
												assign node5108 = (inp[9]) ? 11'b00001000100 : 11'b00001010100;
									assign node5111 = (inp[10]) ? node5123 : node5112;
										assign node5112 = (inp[3]) ? node5118 : node5113;
											assign node5113 = (inp[9]) ? node5115 : 11'b00111010110;
												assign node5115 = (inp[8]) ? 11'b00010010110 : 11'b00001010110;
											assign node5118 = (inp[8]) ? 11'b10010000010 : node5119;
												assign node5119 = (inp[9]) ? 11'b10101000000 : 11'b10011010100;
										assign node5123 = (inp[3]) ? node5127 : node5124;
											assign node5124 = (inp[8]) ? 11'b10110000100 : 11'b10110010010;
											assign node5127 = (inp[9]) ? node5129 : 11'b00110010000;
												assign node5129 = (inp[8]) ? 11'b00010000000 : 11'b00010000010;
								assign node5132 = (inp[10]) ? node5160 : node5133;
									assign node5133 = (inp[3]) ? node5147 : node5134;
										assign node5134 = (inp[8]) ? node5140 : node5135;
											assign node5135 = (inp[9]) ? 11'b00000000000 : node5136;
												assign node5136 = (inp[4]) ? 11'b00101010100 : 11'b00110010000;
											assign node5140 = (inp[4]) ? node5144 : node5141;
												assign node5141 = (inp[9]) ? 11'b00111000010 : 11'b00111010010;
												assign node5144 = (inp[9]) ? 11'b00010000110 : 11'b00010010110;
										assign node5147 = (inp[4]) ? node5155 : node5148;
											assign node5148 = (inp[9]) ? node5152 : node5149;
												assign node5149 = (inp[8]) ? 11'b10111000010 : 11'b10010000000;
												assign node5152 = (inp[8]) ? 11'b10011010110 : 11'b10111010110;
											assign node5155 = (inp[9]) ? 11'b10010000010 : node5156;
												assign node5156 = (inp[8]) ? 11'b10010010110 : 11'b10001010110;
									assign node5160 = (inp[3]) ? node5172 : node5161;
										assign node5161 = (inp[8]) ? node5165 : node5162;
											assign node5162 = (inp[9]) ? 11'b10011000110 : 11'b10101000110;
											assign node5165 = (inp[4]) ? node5169 : node5166;
												assign node5166 = (inp[9]) ? 11'b10011000100 : 11'b10111010000;
												assign node5169 = (inp[9]) ? 11'b10010000000 : 11'b10010000100;
										assign node5172 = (inp[4]) ? node5180 : node5173;
											assign node5173 = (inp[8]) ? node5177 : node5174;
												assign node5174 = (inp[9]) ? 11'b00111000100 : 11'b00100000110;
												assign node5177 = (inp[9]) ? 11'b00011000100 : 11'b00111000100;
											assign node5180 = (inp[9]) ? 11'b00010000000 : node5181;
												assign node5181 = (inp[8]) ? 11'b00010000000 : 11'b00001000000;
							assign node5185 = (inp[10]) ? node5235 : node5186;
								assign node5186 = (inp[11]) ? node5212 : node5187;
									assign node5187 = (inp[8]) ? node5201 : node5188;
										assign node5188 = (inp[4]) ? node5194 : node5189;
											assign node5189 = (inp[3]) ? node5191 : 11'b00000100110;
												assign node5191 = (inp[9]) ? 11'b00110110000 : 11'b00110100010;
											assign node5194 = (inp[9]) ? node5198 : node5195;
												assign node5195 = (inp[3]) ? 11'b00101010000 : 11'b00101000010;
												assign node5198 = (inp[3]) ? 11'b00011000000 : 11'b00111010100;
										assign node5201 = (inp[4]) ? node5207 : node5202;
											assign node5202 = (inp[9]) ? node5204 : 11'b00111000010;
												assign node5204 = (inp[3]) ? 11'b00111010010 : 11'b00111000110;
											assign node5207 = (inp[3]) ? node5209 : 11'b00010000010;
												assign node5209 = (inp[9]) ? 11'b00000000010 : 11'b00100010010;
									assign node5212 = (inp[9]) ? node5226 : node5213;
										assign node5213 = (inp[4]) ? node5221 : node5214;
											assign node5214 = (inp[3]) ? node5218 : node5215;
												assign node5215 = (inp[8]) ? 11'b00101010010 : 11'b00000010000;
												assign node5218 = (inp[8]) ? 11'b00101000010 : 11'b00110000010;
											assign node5221 = (inp[8]) ? 11'b00000010010 : node5222;
												assign node5222 = (inp[3]) ? 11'b00011010010 : 11'b00111010010;
										assign node5226 = (inp[3]) ? node5232 : node5227;
											assign node5227 = (inp[4]) ? node5229 : 11'b00100010100;
												assign node5229 = (inp[8]) ? 11'b00000000110 : 11'b00100000110;
											assign node5232 = (inp[4]) ? 11'b00000000010 : 11'b00001010010;
								assign node5235 = (inp[3]) ? node5263 : node5236;
									assign node5236 = (inp[9]) ? node5248 : node5237;
										assign node5237 = (inp[11]) ? node5243 : node5238;
											assign node5238 = (inp[4]) ? node5240 : 11'b00100100100;
												assign node5240 = (inp[8]) ? 11'b00100010100 : 11'b00001010100;
											assign node5243 = (inp[8]) ? node5245 : 11'b00010010110;
												assign node5245 = (inp[4]) ? 11'b00000000100 : 11'b00101010100;
										assign node5248 = (inp[11]) ? node5256 : node5249;
											assign node5249 = (inp[8]) ? node5253 : node5250;
												assign node5250 = (inp[4]) ? 11'b00100010010 : 11'b00110110000;
												assign node5253 = (inp[4]) ? 11'b00000010000 : 11'b00011010000;
											assign node5256 = (inp[4]) ? node5260 : node5257;
												assign node5257 = (inp[8]) ? 11'b00001000000 : 11'b00101000010;
												assign node5260 = (inp[8]) ? 11'b00000000000 : 11'b00100000000;
									assign node5263 = (inp[9]) ? node5279 : node5264;
										assign node5264 = (inp[8]) ? node5272 : node5265;
											assign node5265 = (inp[4]) ? node5269 : node5266;
												assign node5266 = (inp[11]) ? 11'b00110000000 : 11'b00000100000;
												assign node5269 = (inp[11]) ? 11'b00011000000 : 11'b00111000010;
											assign node5272 = (inp[4]) ? node5276 : node5273;
												assign node5273 = (inp[11]) ? 11'b00101000000 : 11'b00011000000;
												assign node5276 = (inp[11]) ? 11'b00000000000 : 11'b00100000000;
										assign node5279 = (inp[4]) ? node5285 : node5280;
											assign node5280 = (inp[11]) ? 11'b00001000000 : node5281;
												assign node5281 = (inp[8]) ? 11'b00011000000 : 11'b00011000010;
											assign node5285 = (inp[11]) ? 11'b00000000000 : node5286;
												assign node5286 = (inp[8]) ? 11'b00000000000 : 11'b00000000010;
			assign node5290 = (inp[6]) ? node6158 : node5291;
				assign node5291 = (inp[2]) ? node5731 : node5292;
					assign node5292 = (inp[5]) ? node5506 : node5293;
						assign node5293 = (inp[0]) ? node5401 : node5294;
							assign node5294 = (inp[10]) ? node5348 : node5295;
								assign node5295 = (inp[3]) ? node5317 : node5296;
									assign node5296 = (inp[4]) ? node5306 : node5297;
										assign node5297 = (inp[8]) ? node5299 : 11'b00011100011;
											assign node5299 = (inp[11]) ? node5303 : node5300;
												assign node5300 = (inp[9]) ? 11'b00000000001 : 11'b00010000011;
												assign node5303 = (inp[9]) ? 11'b00100110011 : 11'b00010100001;
										assign node5306 = (inp[8]) ? node5310 : node5307;
											assign node5307 = (inp[11]) ? 11'b00000110101 : 11'b00010100111;
											assign node5310 = (inp[11]) ? node5314 : node5311;
												assign node5311 = (inp[9]) ? 11'b00101100101 : 11'b00111100101;
												assign node5314 = (inp[9]) ? 11'b00011110111 : 11'b00101100111;
									assign node5317 = (inp[4]) ? node5333 : node5318;
										assign node5318 = (inp[8]) ? node5326 : node5319;
											assign node5319 = (inp[9]) ? node5323 : node5320;
												assign node5320 = (inp[11]) ? 11'b10011110011 : 11'b10011100011;
												assign node5323 = (inp[11]) ? 11'b10111100111 : 11'b10011100111;
											assign node5326 = (inp[9]) ? node5330 : node5327;
												assign node5327 = (inp[11]) ? 11'b10110110001 : 11'b10110000011;
												assign node5330 = (inp[11]) ? 11'b10110100101 : 11'b10101100111;
										assign node5333 = (inp[9]) ? node5341 : node5334;
											assign node5334 = (inp[8]) ? node5338 : node5335;
												assign node5335 = (inp[11]) ? 11'b10100100111 : 11'b10010100111;
												assign node5338 = (inp[11]) ? 11'b10001100111 : 11'b10011100111;
											assign node5341 = (inp[8]) ? node5345 : node5342;
												assign node5342 = (inp[11]) ? 11'b10000110011 : 11'b10110110011;
												assign node5345 = (inp[11]) ? 11'b10001110011 : 11'b10001110001;
								assign node5348 = (inp[3]) ? node5374 : node5349;
									assign node5349 = (inp[8]) ? node5359 : node5350;
										assign node5350 = (inp[4]) ? node5356 : node5351;
											assign node5351 = (inp[9]) ? node5353 : 11'b10011100001;
												assign node5353 = (inp[11]) ? 11'b10111110101 : 11'b10011110101;
											assign node5356 = (inp[9]) ? 11'b10110100001 : 11'b10010110101;
										assign node5359 = (inp[11]) ? node5367 : node5360;
											assign node5360 = (inp[9]) ? node5364 : node5361;
												assign node5361 = (inp[4]) ? 11'b10111110111 : 11'b10010000001;
												assign node5364 = (inp[4]) ? 11'b10010100011 : 11'b10001110111;
											assign node5367 = (inp[4]) ? node5371 : node5368;
												assign node5368 = (inp[9]) ? 11'b10010110101 : 11'b10100100001;
												assign node5371 = (inp[9]) ? 11'b10101110011 : 11'b10101110101;
									assign node5374 = (inp[4]) ? node5388 : node5375;
										assign node5375 = (inp[8]) ? node5381 : node5376;
											assign node5376 = (inp[9]) ? node5378 : 11'b00011100101;
												assign node5378 = (inp[11]) ? 11'b00001110101 : 11'b00011110101;
											assign node5381 = (inp[9]) ? node5385 : node5382;
												assign node5382 = (inp[11]) ? 11'b00000110111 : 11'b00110000101;
												assign node5385 = (inp[11]) ? 11'b00111110111 : 11'b00101110101;
										assign node5388 = (inp[8]) ? node5394 : node5389;
											assign node5389 = (inp[11]) ? 11'b00100110001 : node5390;
												assign node5390 = (inp[9]) ? 11'b00110110001 : 11'b00110100001;
											assign node5394 = (inp[11]) ? node5398 : node5395;
												assign node5395 = (inp[9]) ? 11'b00110110011 : 11'b00001100011;
												assign node5398 = (inp[9]) ? 11'b00101110001 : 11'b00111110001;
							assign node5401 = (inp[10]) ? node5455 : node5402;
								assign node5402 = (inp[8]) ? node5428 : node5403;
									assign node5403 = (inp[4]) ? node5417 : node5404;
										assign node5404 = (inp[9]) ? node5410 : node5405;
											assign node5405 = (inp[11]) ? node5407 : 11'b00001100011;
												assign node5407 = (inp[3]) ? 11'b00001100011 : 11'b00001110011;
											assign node5410 = (inp[3]) ? node5414 : node5411;
												assign node5411 = (inp[11]) ? 11'b00101110111 : 11'b00001100111;
												assign node5414 = (inp[11]) ? 11'b00101110011 : 11'b00001110011;
										assign node5417 = (inp[11]) ? node5425 : node5418;
											assign node5418 = (inp[9]) ? node5422 : node5419;
												assign node5419 = (inp[3]) ? 11'b00000110011 : 11'b00000100011;
												assign node5422 = (inp[3]) ? 11'b00100100011 : 11'b00100110111;
											assign node5425 = (inp[9]) ? 11'b00010100111 : 11'b00010110011;
									assign node5428 = (inp[4]) ? node5442 : node5429;
										assign node5429 = (inp[11]) ? node5435 : node5430;
											assign node5430 = (inp[9]) ? 11'b00111100111 : node5431;
												assign node5431 = (inp[3]) ? 11'b00000000011 : 11'b00100000011;
											assign node5435 = (inp[3]) ? node5439 : node5436;
												assign node5436 = (inp[9]) ? 11'b00000110111 : 11'b00100110001;
												assign node5439 = (inp[9]) ? 11'b00100110001 : 11'b00010100001;
										assign node5442 = (inp[9]) ? node5450 : node5443;
											assign node5443 = (inp[11]) ? node5447 : node5444;
												assign node5444 = (inp[3]) ? 11'b00001110011 : 11'b00101100001;
												assign node5447 = (inp[3]) ? 11'b00111110001 : 11'b00111110011;
											assign node5450 = (inp[3]) ? node5452 : 11'b00011110101;
												assign node5452 = (inp[11]) ? 11'b00111100011 : 11'b00110100011;
								assign node5455 = (inp[3]) ? node5483 : node5456;
									assign node5456 = (inp[9]) ? node5470 : node5457;
										assign node5457 = (inp[8]) ? node5463 : node5458;
											assign node5458 = (inp[4]) ? 11'b00000110101 : node5459;
												assign node5459 = (inp[11]) ? 11'b00001110101 : 11'b00001100101;
											assign node5463 = (inp[4]) ? node5467 : node5464;
												assign node5464 = (inp[11]) ? 11'b00110110111 : 11'b00100000101;
												assign node5467 = (inp[11]) ? 11'b00001100101 : 11'b00101110111;
										assign node5470 = (inp[11]) ? node5478 : node5471;
											assign node5471 = (inp[4]) ? node5475 : node5472;
												assign node5472 = (inp[8]) ? 11'b00111110001 : 11'b00001110001;
												assign node5475 = (inp[8]) ? 11'b00000110011 : 11'b00100110001;
											assign node5478 = (inp[8]) ? node5480 : 11'b00011100001;
												assign node5480 = (inp[4]) ? 11'b00011100001 : 11'b00100100001;
									assign node5483 = (inp[9]) ? node5495 : node5484;
										assign node5484 = (inp[8]) ? node5488 : node5485;
											assign node5485 = (inp[11]) ? 11'b00101100001 : 11'b00001100001;
											assign node5488 = (inp[4]) ? node5492 : node5489;
												assign node5489 = (inp[11]) ? 11'b00110100011 : 11'b00010000001;
												assign node5492 = (inp[11]) ? 11'b00001100001 : 11'b00111100001;
										assign node5495 = (inp[4]) ? node5501 : node5496;
											assign node5496 = (inp[11]) ? node5498 : 11'b00001100001;
												assign node5498 = (inp[8]) ? 11'b00011100011 : 11'b00011100001;
											assign node5501 = (inp[8]) ? node5503 : 11'b00000100001;
												assign node5503 = (inp[11]) ? 11'b00001100001 : 11'b00000100011;
						assign node5506 = (inp[0]) ? node5616 : node5507;
							assign node5507 = (inp[11]) ? node5561 : node5508;
								assign node5508 = (inp[8]) ? node5534 : node5509;
									assign node5509 = (inp[10]) ? node5523 : node5510;
										assign node5510 = (inp[3]) ? node5516 : node5511;
											assign node5511 = (inp[4]) ? 11'b00001010101 : node5512;
												assign node5512 = (inp[9]) ? 11'b00011010001 : 11'b00010110001;
											assign node5516 = (inp[4]) ? node5520 : node5517;
												assign node5517 = (inp[9]) ? 11'b10011010111 : 11'b10011010011;
												assign node5520 = (inp[9]) ? 11'b10010000001 : 11'b10101010101;
										assign node5523 = (inp[4]) ? node5529 : node5524;
											assign node5524 = (inp[9]) ? 11'b00001000111 : node5525;
												assign node5525 = (inp[3]) ? 11'b00111010101 : 11'b10111010011;
											assign node5529 = (inp[3]) ? node5531 : 11'b10010010011;
												assign node5531 = (inp[9]) ? 11'b00110000011 : 11'b00000010011;
									assign node5534 = (inp[4]) ? node5548 : node5535;
										assign node5535 = (inp[10]) ? node5541 : node5536;
											assign node5536 = (inp[3]) ? 11'b10010110011 : node5537;
												assign node5537 = (inp[9]) ? 11'b00000110001 : 11'b00011110001;
											assign node5541 = (inp[3]) ? node5545 : node5542;
												assign node5542 = (inp[9]) ? 11'b10010100111 : 11'b10110110011;
												assign node5545 = (inp[9]) ? 11'b00110100111 : 11'b00100110111;
										assign node5548 = (inp[9]) ? node5556 : node5549;
											assign node5549 = (inp[10]) ? node5553 : node5550;
												assign node5550 = (inp[3]) ? 11'b10000110101 : 11'b00100110111;
												assign node5553 = (inp[3]) ? 11'b00011010011 : 11'b10010100101;
											assign node5556 = (inp[10]) ? 11'b10101010001 : node5557;
												assign node5557 = (inp[3]) ? 11'b10101000011 : 11'b00111010111;
								assign node5561 = (inp[4]) ? node5589 : node5562;
									assign node5562 = (inp[9]) ? node5576 : node5563;
										assign node5563 = (inp[3]) ? node5571 : node5564;
											assign node5564 = (inp[10]) ? node5568 : node5565;
												assign node5565 = (inp[8]) ? 11'b00011010011 : 11'b00010010001;
												assign node5568 = (inp[8]) ? 11'b10001010011 : 11'b10111010011;
											assign node5571 = (inp[10]) ? 11'b00001000111 : node5572;
												assign node5572 = (inp[8]) ? 11'b10001000011 : 11'b10110000001;
										assign node5576 = (inp[3]) ? node5582 : node5577;
											assign node5577 = (inp[10]) ? 11'b10101000101 : node5578;
												assign node5578 = (inp[8]) ? 11'b00011000001 : 11'b00101000011;
											assign node5582 = (inp[10]) ? node5586 : node5583;
												assign node5583 = (inp[8]) ? 11'b10110010111 : 11'b10001010101;
												assign node5586 = (inp[8]) ? 11'b00100000111 : 11'b00011000111;
									assign node5589 = (inp[9]) ? node5605 : node5590;
										assign node5590 = (inp[10]) ? node5598 : node5591;
											assign node5591 = (inp[8]) ? node5595 : node5592;
												assign node5592 = (inp[3]) ? 11'b10111010101 : 11'b00011010111;
												assign node5595 = (inp[3]) ? 11'b10110010101 : 11'b00110010101;
											assign node5598 = (inp[3]) ? node5602 : node5599;
												assign node5599 = (inp[8]) ? 11'b10100000101 : 11'b10011000101;
												assign node5602 = (inp[8]) ? 11'b00100000011 : 11'b00110000011;
										assign node5605 = (inp[8]) ? node5611 : node5606;
											assign node5606 = (inp[3]) ? 11'b10100000011 : node5607;
												assign node5607 = (inp[10]) ? 11'b10000000001 : 11'b00000000111;
											assign node5611 = (inp[3]) ? node5613 : 11'b00110000111;
												assign node5613 = (inp[10]) ? 11'b00100000001 : 11'b10110000001;
							assign node5616 = (inp[3]) ? node5672 : node5617;
								assign node5617 = (inp[8]) ? node5643 : node5618;
									assign node5618 = (inp[4]) ? node5630 : node5619;
										assign node5619 = (inp[10]) ? node5623 : node5620;
											assign node5620 = (inp[9]) ? 11'b00001000101 : 11'b00000100001;
											assign node5623 = (inp[9]) ? node5627 : node5624;
												assign node5624 = (inp[11]) ? 11'b00011010111 : 11'b00101000111;
												assign node5627 = (inp[11]) ? 11'b00111000011 : 11'b00101010011;
										assign node5630 = (inp[9]) ? node5636 : node5631;
											assign node5631 = (inp[10]) ? 11'b00010010111 : node5632;
												assign node5632 = (inp[11]) ? 11'b00101010011 : 11'b00111000001;
											assign node5636 = (inp[11]) ? node5640 : node5637;
												assign node5637 = (inp[10]) ? 11'b00100010011 : 11'b00110010101;
												assign node5640 = (inp[10]) ? 11'b00110000001 : 11'b00110000111;
									assign node5643 = (inp[11]) ? node5659 : node5644;
										assign node5644 = (inp[10]) ? node5652 : node5645;
											assign node5645 = (inp[4]) ? node5649 : node5646;
												assign node5646 = (inp[9]) ? 11'b00110100101 : 11'b00101100001;
												assign node5649 = (inp[9]) ? 11'b00011010111 : 11'b00010100001;
											assign node5652 = (inp[9]) ? node5656 : node5653;
												assign node5653 = (inp[4]) ? 11'b00100110101 : 11'b00010100111;
												assign node5656 = (inp[4]) ? 11'b00001010001 : 11'b00000110011;
										assign node5659 = (inp[10]) ? node5667 : node5660;
											assign node5660 = (inp[9]) ? node5664 : node5661;
												assign node5661 = (inp[4]) ? 11'b00000010001 : 11'b00101010011;
												assign node5664 = (inp[4]) ? 11'b00000000111 : 11'b00001010101;
											assign node5667 = (inp[9]) ? node5669 : 11'b00010000111;
												assign node5669 = (inp[4]) ? 11'b00010000001 : 11'b00010000011;
								assign node5672 = (inp[10]) ? node5704 : node5673;
									assign node5673 = (inp[4]) ? node5689 : node5674;
										assign node5674 = (inp[9]) ? node5682 : node5675;
											assign node5675 = (inp[11]) ? node5679 : node5676;
												assign node5676 = (inp[8]) ? 11'b00100100011 : 11'b00101000011;
												assign node5679 = (inp[8]) ? 11'b00111000011 : 11'b00100000001;
											assign node5682 = (inp[11]) ? node5686 : node5683;
												assign node5683 = (inp[8]) ? 11'b00100110001 : 11'b00101010011;
												assign node5686 = (inp[8]) ? 11'b00010010011 : 11'b00011010001;
										assign node5689 = (inp[9]) ? node5697 : node5690;
											assign node5690 = (inp[11]) ? node5694 : node5691;
												assign node5691 = (inp[8]) ? 11'b00110110001 : 11'b00110010011;
												assign node5694 = (inp[8]) ? 11'b00010010001 : 11'b00001010001;
											assign node5697 = (inp[8]) ? node5701 : node5698;
												assign node5698 = (inp[11]) ? 11'b00010000001 : 11'b00000000001;
												assign node5701 = (inp[11]) ? 11'b00010000001 : 11'b00011000001;
									assign node5704 = (inp[4]) ? node5718 : node5705;
										assign node5705 = (inp[11]) ? node5713 : node5706;
											assign node5706 = (inp[8]) ? node5710 : node5707;
												assign node5707 = (inp[9]) ? 11'b00011000001 : 11'b00001000001;
												assign node5710 = (inp[9]) ? 11'b00010100011 : 11'b00010100001;
											assign node5713 = (inp[9]) ? 11'b00001000011 : node5714;
												assign node5714 = (inp[8]) ? 11'b00101000001 : 11'b00111000011;
										assign node5718 = (inp[9]) ? node5724 : node5719;
											assign node5719 = (inp[11]) ? node5721 : 11'b00101000011;
												assign node5721 = (inp[8]) ? 11'b00000000011 : 11'b00010000011;
											assign node5724 = (inp[8]) ? node5728 : node5725;
												assign node5725 = (inp[11]) ? 11'b00000000001 : 11'b00000000011;
												assign node5728 = (inp[11]) ? 11'b00000000001 : 11'b00001000001;
					assign node5731 = (inp[8]) ? node5945 : node5732;
						assign node5732 = (inp[5]) ? node5836 : node5733;
							assign node5733 = (inp[11]) ? node5783 : node5734;
								assign node5734 = (inp[4]) ? node5760 : node5735;
									assign node5735 = (inp[0]) ? node5747 : node5736;
										assign node5736 = (inp[10]) ? node5742 : node5737;
											assign node5737 = (inp[3]) ? 11'b10111000011 : node5738;
												assign node5738 = (inp[9]) ? 11'b00111000001 : 11'b00111000011;
											assign node5742 = (inp[9]) ? node5744 : 11'b00101000101;
												assign node5744 = (inp[3]) ? 11'b00101010111 : 11'b10101010111;
										assign node5747 = (inp[3]) ? node5753 : node5748;
											assign node5748 = (inp[10]) ? node5750 : 11'b00001000101;
												assign node5750 = (inp[9]) ? 11'b00011010011 : 11'b00011000101;
											assign node5753 = (inp[10]) ? node5757 : node5754;
												assign node5754 = (inp[9]) ? 11'b00011010011 : 11'b00011000011;
												assign node5757 = (inp[9]) ? 11'b00001000011 : 11'b00001000001;
									assign node5760 = (inp[9]) ? node5770 : node5761;
										assign node5761 = (inp[10]) ? node5767 : node5762;
											assign node5762 = (inp[0]) ? 11'b00001000001 : node5763;
												assign node5763 = (inp[3]) ? 11'b10111000101 : 11'b00111000101;
											assign node5767 = (inp[0]) ? 11'b00100000011 : 11'b00010000011;
										assign node5770 = (inp[10]) ? node5778 : node5771;
											assign node5771 = (inp[0]) ? node5775 : node5772;
												assign node5772 = (inp[3]) ? 11'b10000010011 : 11'b00010000111;
												assign node5775 = (inp[3]) ? 11'b00110000001 : 11'b00100010111;
											assign node5778 = (inp[3]) ? node5780 : 11'b00110010001;
												assign node5780 = (inp[0]) ? 11'b00000000001 : 11'b00010010001;
								assign node5783 = (inp[4]) ? node5813 : node5784;
									assign node5784 = (inp[9]) ? node5800 : node5785;
										assign node5785 = (inp[0]) ? node5793 : node5786;
											assign node5786 = (inp[3]) ? node5790 : node5787;
												assign node5787 = (inp[10]) ? 11'b10100000011 : 11'b00110000011;
												assign node5790 = (inp[10]) ? 11'b00110010101 : 11'b10100010011;
											assign node5793 = (inp[3]) ? node5797 : node5794;
												assign node5794 = (inp[10]) ? 11'b00000010111 : 11'b00010010011;
												assign node5797 = (inp[10]) ? 11'b00100000001 : 11'b00010000011;
										assign node5800 = (inp[10]) ? node5806 : node5801;
											assign node5801 = (inp[0]) ? node5803 : 11'b10000000101;
												assign node5803 = (inp[3]) ? 11'b00111110010 : 11'b00110010101;
											assign node5806 = (inp[0]) ? node5810 : node5807;
												assign node5807 = (inp[3]) ? 11'b00111110110 : 11'b10011110110;
												assign node5810 = (inp[3]) ? 11'b00011100010 : 11'b00001100010;
									assign node5813 = (inp[0]) ? node5825 : node5814;
										assign node5814 = (inp[10]) ? node5820 : node5815;
											assign node5815 = (inp[3]) ? 11'b10111110010 : node5816;
												assign node5816 = (inp[9]) ? 11'b00101110110 : 11'b00101100110;
											assign node5820 = (inp[3]) ? 11'b00001110000 : node5821;
												assign node5821 = (inp[9]) ? 11'b10001110010 : 11'b10011110100;
										assign node5825 = (inp[3]) ? node5831 : node5826;
											assign node5826 = (inp[10]) ? node5828 : 11'b00001100110;
												assign node5828 = (inp[9]) ? 11'b00111100000 : 11'b00101100100;
											assign node5831 = (inp[10]) ? 11'b00011100010 : node5832;
												assign node5832 = (inp[9]) ? 11'b00101100010 : 11'b00101110000;
							assign node5836 = (inp[0]) ? node5896 : node5837;
								assign node5837 = (inp[11]) ? node5869 : node5838;
									assign node5838 = (inp[10]) ? node5854 : node5839;
										assign node5839 = (inp[3]) ? node5847 : node5840;
											assign node5840 = (inp[4]) ? node5844 : node5841;
												assign node5841 = (inp[9]) ? 11'b00110110000 : 11'b00111110000;
												assign node5844 = (inp[9]) ? 11'b00010110100 : 11'b00100110110;
											assign node5847 = (inp[4]) ? node5851 : node5848;
												assign node5848 = (inp[9]) ? 11'b10100110100 : 11'b10110110010;
												assign node5851 = (inp[9]) ? 11'b10111100010 : 11'b10010110110;
										assign node5854 = (inp[3]) ? node5862 : node5855;
											assign node5855 = (inp[4]) ? node5859 : node5856;
												assign node5856 = (inp[9]) ? 11'b10010100100 : 11'b10000110010;
												assign node5859 = (inp[9]) ? 11'b10101110010 : 11'b10110100100;
											assign node5862 = (inp[9]) ? node5866 : node5863;
												assign node5863 = (inp[4]) ? 11'b00100110000 : 11'b00010110110;
												assign node5866 = (inp[4]) ? 11'b00011100010 : 11'b00110100110;
									assign node5869 = (inp[4]) ? node5885 : node5870;
										assign node5870 = (inp[9]) ? node5878 : node5871;
											assign node5871 = (inp[3]) ? node5875 : node5872;
												assign node5872 = (inp[10]) ? 11'b10011110000 : 11'b00111110000;
												assign node5875 = (inp[10]) ? 11'b00111100110 : 11'b10001100000;
											assign node5878 = (inp[3]) ? node5882 : node5879;
												assign node5879 = (inp[10]) ? 11'b10001100110 : 11'b00001100010;
												assign node5882 = (inp[10]) ? 11'b00101100100 : 11'b10111110110;
										assign node5885 = (inp[3]) ? node5889 : node5886;
											assign node5886 = (inp[9]) ? 11'b10110100000 : 11'b10100100110;
											assign node5889 = (inp[10]) ? node5893 : node5890;
												assign node5890 = (inp[9]) ? 11'b10010100000 : 11'b10001110100;
												assign node5893 = (inp[9]) ? 11'b00000100000 : 11'b00010100010;
								assign node5896 = (inp[3]) ? node5918 : node5897;
									assign node5897 = (inp[9]) ? node5909 : node5898;
										assign node5898 = (inp[10]) ? node5902 : node5899;
											assign node5899 = (inp[4]) ? 11'b00110100010 : 11'b00001100000;
											assign node5902 = (inp[11]) ? node5906 : node5903;
												assign node5903 = (inp[4]) ? 11'b00010110100 : 11'b00110100110;
												assign node5906 = (inp[4]) ? 11'b00100100110 : 11'b00001110100;
										assign node5909 = (inp[10]) ? node5913 : node5910;
											assign node5910 = (inp[11]) ? 11'b00110100100 : 11'b00100110100;
											assign node5913 = (inp[11]) ? 11'b00111100000 : node5914;
												assign node5914 = (inp[4]) ? 11'b00111110010 : 11'b00100110000;
									assign node5918 = (inp[9]) ? node5932 : node5919;
										assign node5919 = (inp[11]) ? node5927 : node5920;
											assign node5920 = (inp[4]) ? node5924 : node5921;
												assign node5921 = (inp[10]) ? 11'b00000100010 : 11'b00110100010;
												assign node5924 = (inp[10]) ? 11'b00110100000 : 11'b00100110010;
											assign node5927 = (inp[4]) ? 11'b00010100010 : node5928;
												assign node5928 = (inp[10]) ? 11'b00111100010 : 11'b00111100000;
										assign node5932 = (inp[11]) ? node5940 : node5933;
											assign node5933 = (inp[4]) ? node5937 : node5934;
												assign node5934 = (inp[10]) ? 11'b00010100010 : 11'b00110110000;
												assign node5937 = (inp[10]) ? 11'b00001100010 : 11'b00011100010;
											assign node5940 = (inp[10]) ? node5942 : 11'b00001110010;
												assign node5942 = (inp[4]) ? 11'b00000100000 : 11'b00001100000;
						assign node5945 = (inp[11]) ? node6061 : node5946;
							assign node5946 = (inp[4]) ? node6008 : node5947;
								assign node5947 = (inp[5]) ? node5979 : node5948;
									assign node5948 = (inp[3]) ? node5964 : node5949;
										assign node5949 = (inp[10]) ? node5957 : node5950;
											assign node5950 = (inp[9]) ? node5954 : node5951;
												assign node5951 = (inp[0]) ? 11'b00100100010 : 11'b00110100010;
												assign node5954 = (inp[0]) ? 11'b00110100100 : 11'b00100100000;
											assign node5957 = (inp[9]) ? node5961 : node5958;
												assign node5958 = (inp[0]) ? 11'b00100100110 : 11'b10100100010;
												assign node5961 = (inp[0]) ? 11'b00111010010 : 11'b10111010110;
										assign node5964 = (inp[9]) ? node5972 : node5965;
											assign node5965 = (inp[10]) ? node5969 : node5966;
												assign node5966 = (inp[0]) ? 11'b00010100010 : 11'b10000100010;
												assign node5969 = (inp[0]) ? 11'b00010100000 : 11'b00010100100;
											assign node5972 = (inp[10]) ? node5976 : node5973;
												assign node5973 = (inp[0]) ? 11'b00000110000 : 11'b10010100100;
												assign node5976 = (inp[0]) ? 11'b00001000010 : 11'b00001010110;
									assign node5979 = (inp[10]) ? node5995 : node5980;
										assign node5980 = (inp[9]) ? node5988 : node5981;
											assign node5981 = (inp[0]) ? node5985 : node5982;
												assign node5982 = (inp[3]) ? 11'b10100010000 : 11'b00110010000;
												assign node5985 = (inp[3]) ? 11'b00111000010 : 11'b00100000000;
											assign node5988 = (inp[3]) ? node5992 : node5989;
												assign node5989 = (inp[0]) ? 11'b00101000110 : 11'b00101010010;
												assign node5992 = (inp[0]) ? 11'b00111010000 : 11'b10111010100;
										assign node5995 = (inp[9]) ? node6003 : node5996;
											assign node5996 = (inp[0]) ? node6000 : node5997;
												assign node5997 = (inp[3]) ? 11'b00001010110 : 11'b10011010010;
												assign node6000 = (inp[3]) ? 11'b00011000010 : 11'b00001000110;
											assign node6003 = (inp[3]) ? node6005 : 11'b00001010000;
												assign node6005 = (inp[0]) ? 11'b00011000000 : 11'b00011000100;
								assign node6008 = (inp[9]) ? node6034 : node6009;
									assign node6009 = (inp[0]) ? node6025 : node6010;
										assign node6010 = (inp[3]) ? node6018 : node6011;
											assign node6011 = (inp[10]) ? node6015 : node6012;
												assign node6012 = (inp[5]) ? 11'b00001010100 : 11'b00011000110;
												assign node6015 = (inp[5]) ? 11'b10101000110 : 11'b10011010100;
											assign node6018 = (inp[10]) ? node6022 : node6019;
												assign node6019 = (inp[5]) ? 11'b10111010110 : 11'b10101000110;
												assign node6022 = (inp[5]) ? 11'b00111010010 : 11'b00111000000;
										assign node6025 = (inp[10]) ? node6029 : node6026;
											assign node6026 = (inp[3]) ? 11'b00011010000 : 11'b00101000010;
											assign node6029 = (inp[3]) ? 11'b00101000010 : node6030;
												assign node6030 = (inp[5]) ? 11'b00111010110 : 11'b00101010100;
									assign node6034 = (inp[3]) ? node6050 : node6035;
										assign node6035 = (inp[10]) ? node6043 : node6036;
											assign node6036 = (inp[5]) ? node6040 : node6037;
												assign node6037 = (inp[0]) ? 11'b00001010100 : 11'b00001000100;
												assign node6040 = (inp[0]) ? 11'b00011010100 : 11'b00001010110;
											assign node6043 = (inp[0]) ? node6047 : node6044;
												assign node6044 = (inp[5]) ? 11'b10001010000 : 11'b10101000010;
												assign node6047 = (inp[5]) ? 11'b00011010000 : 11'b00011010010;
										assign node6050 = (inp[0]) ? node6056 : node6051;
											assign node6051 = (inp[5]) ? node6053 : 11'b00011010010;
												assign node6053 = (inp[10]) ? 11'b00011000000 : 11'b10011000000;
											assign node6056 = (inp[5]) ? 11'b00001000000 : node6057;
												assign node6057 = (inp[10]) ? 11'b00001000010 : 11'b00101000010;
							assign node6061 = (inp[3]) ? node6109 : node6062;
								assign node6062 = (inp[4]) ? node6088 : node6063;
									assign node6063 = (inp[9]) ? node6077 : node6064;
										assign node6064 = (inp[5]) ? node6072 : node6065;
											assign node6065 = (inp[0]) ? node6069 : node6066;
												assign node6066 = (inp[10]) ? 11'b10011000000 : 11'b00111000000;
												assign node6069 = (inp[10]) ? 11'b00101010100 : 11'b00111010000;
											assign node6072 = (inp[0]) ? 11'b00110010110 : node6073;
												assign node6073 = (inp[10]) ? 11'b10110010010 : 11'b00110010010;
										assign node6077 = (inp[5]) ? node6081 : node6078;
											assign node6078 = (inp[10]) ? 11'b00100000010 : 11'b00000010110;
											assign node6081 = (inp[0]) ? node6085 : node6082;
												assign node6082 = (inp[10]) ? 11'b10010000100 : 11'b00110000000;
												assign node6085 = (inp[10]) ? 11'b00010000000 : 11'b00010010100;
									assign node6088 = (inp[10]) ? node6100 : node6089;
										assign node6089 = (inp[5]) ? node6095 : node6090;
											assign node6090 = (inp[0]) ? 11'b00110010000 : node6091;
												assign node6091 = (inp[9]) ? 11'b00110010110 : 11'b00000000100;
											assign node6095 = (inp[9]) ? 11'b00010000100 : node6096;
												assign node6096 = (inp[0]) ? 11'b00010010010 : 11'b00010010110;
										assign node6100 = (inp[9]) ? node6104 : node6101;
											assign node6101 = (inp[0]) ? 11'b00010000110 : 11'b10010000110;
											assign node6104 = (inp[0]) ? 11'b00010000000 : node6105;
												assign node6105 = (inp[5]) ? 11'b10010000000 : 11'b10010010000;
								assign node6109 = (inp[0]) ? node6139 : node6110;
									assign node6110 = (inp[10]) ? node6124 : node6111;
										assign node6111 = (inp[9]) ? node6117 : node6112;
											assign node6112 = (inp[4]) ? 11'b10110000100 : node6113;
												assign node6113 = (inp[5]) ? 11'b10100000010 : 11'b10001010000;
											assign node6117 = (inp[5]) ? node6121 : node6118;
												assign node6118 = (inp[4]) ? 11'b10100010010 : 11'b10000000110;
												assign node6121 = (inp[4]) ? 11'b10000000000 : 11'b10000010100;
										assign node6124 = (inp[5]) ? node6132 : node6125;
											assign node6125 = (inp[4]) ? node6129 : node6126;
												assign node6126 = (inp[9]) ? 11'b00010010100 : 11'b00101010100;
												assign node6129 = (inp[9]) ? 11'b00000010000 : 11'b00010010010;
											assign node6132 = (inp[9]) ? node6136 : node6133;
												assign node6133 = (inp[4]) ? 11'b00000000010 : 11'b00100000110;
												assign node6136 = (inp[4]) ? 11'b00000000000 : 11'b00000000100;
									assign node6139 = (inp[5]) ? node6153 : node6140;
										assign node6140 = (inp[4]) ? node6146 : node6141;
											assign node6141 = (inp[9]) ? 11'b00110010010 : node6142;
												assign node6142 = (inp[10]) ? 11'b00110000010 : 11'b00001000000;
											assign node6146 = (inp[10]) ? node6150 : node6147;
												assign node6147 = (inp[9]) ? 11'b00100000010 : 11'b00100010000;
												assign node6150 = (inp[9]) ? 11'b00000000000 : 11'b00000000010;
										assign node6153 = (inp[9]) ? 11'b00000000000 : node6154;
											assign node6154 = (inp[10]) ? 11'b00000000010 : 11'b00000010010;
				assign node6158 = (inp[2]) ? node6578 : node6159;
					assign node6159 = (inp[8]) ? node6371 : node6160;
						assign node6160 = (inp[11]) ? node6264 : node6161;
							assign node6161 = (inp[3]) ? node6215 : node6162;
								assign node6162 = (inp[9]) ? node6190 : node6163;
									assign node6163 = (inp[5]) ? node6177 : node6164;
										assign node6164 = (inp[10]) ? node6170 : node6165;
											assign node6165 = (inp[4]) ? node6167 : 11'b00011100010;
												assign node6167 = (inp[0]) ? 11'b00011100010 : 11'b00011100110;
											assign node6170 = (inp[0]) ? node6174 : node6171;
												assign node6171 = (inp[4]) ? 11'b10011110110 : 11'b10011100010;
												assign node6174 = (inp[4]) ? 11'b00011110110 : 11'b00011100110;
										assign node6177 = (inp[10]) ? node6185 : node6178;
											assign node6178 = (inp[4]) ? node6182 : node6179;
												assign node6179 = (inp[0]) ? 11'b00010100000 : 11'b00010110000;
												assign node6182 = (inp[0]) ? 11'b00101100000 : 11'b00001110100;
											assign node6185 = (inp[4]) ? 11'b10011100100 : node6186;
												assign node6186 = (inp[0]) ? 11'b00111100110 : 11'b10111110010;
									assign node6190 = (inp[5]) ? node6204 : node6191;
										assign node6191 = (inp[4]) ? node6199 : node6192;
											assign node6192 = (inp[10]) ? node6196 : node6193;
												assign node6193 = (inp[0]) ? 11'b00011100100 : 11'b00011100000;
												assign node6196 = (inp[0]) ? 11'b00011110000 : 11'b10011110100;
											assign node6199 = (inp[0]) ? node6201 : 11'b00111100100;
												assign node6201 = (inp[10]) ? 11'b00111110000 : 11'b00111110100;
										assign node6204 = (inp[0]) ? node6210 : node6205;
											assign node6205 = (inp[10]) ? 11'b10101100110 : node6206;
												assign node6206 = (inp[4]) ? 11'b00111110110 : 11'b00001110010;
											assign node6210 = (inp[10]) ? node6212 : 11'b00101110110;
												assign node6212 = (inp[4]) ? 11'b00111110010 : 11'b00111110000;
								assign node6215 = (inp[0]) ? node6239 : node6216;
									assign node6216 = (inp[10]) ? node6228 : node6217;
										assign node6217 = (inp[5]) ? node6223 : node6218;
											assign node6218 = (inp[9]) ? 11'b10001100100 : node6219;
												assign node6219 = (inp[4]) ? 11'b10001100110 : 11'b10001100010;
											assign node6223 = (inp[9]) ? node6225 : 11'b10111110100;
												assign node6225 = (inp[4]) ? 11'b10001100010 : 11'b10011110110;
										assign node6228 = (inp[4]) ? node6234 : node6229;
											assign node6229 = (inp[9]) ? 11'b00011100100 : node6230;
												assign node6230 = (inp[5]) ? 11'b00101110110 : 11'b00001100110;
											assign node6234 = (inp[5]) ? 11'b00101100010 : node6235;
												assign node6235 = (inp[9]) ? 11'b00101110000 : 11'b00101100010;
									assign node6239 = (inp[9]) ? node6253 : node6240;
										assign node6240 = (inp[5]) ? node6248 : node6241;
											assign node6241 = (inp[10]) ? node6245 : node6242;
												assign node6242 = (inp[4]) ? 11'b00001110010 : 11'b00001100010;
												assign node6245 = (inp[4]) ? 11'b00101100010 : 11'b00001100010;
											assign node6248 = (inp[10]) ? node6250 : 11'b00100100000;
												assign node6250 = (inp[4]) ? 11'b00111100010 : 11'b00001100010;
										assign node6253 = (inp[10]) ? node6261 : node6254;
											assign node6254 = (inp[4]) ? node6258 : node6255;
												assign node6255 = (inp[5]) ? 11'b00101110010 : 11'b00001110000;
												assign node6258 = (inp[5]) ? 11'b00001100010 : 11'b00101100000;
											assign node6261 = (inp[5]) ? 11'b00011100000 : 11'b00001100000;
							assign node6264 = (inp[0]) ? node6322 : node6265;
								assign node6265 = (inp[5]) ? node6291 : node6266;
									assign node6266 = (inp[10]) ? node6276 : node6267;
										assign node6267 = (inp[3]) ? node6273 : node6268;
											assign node6268 = (inp[9]) ? node6270 : 11'b00001100000;
												assign node6270 = (inp[4]) ? 11'b00010110110 : 11'b00100110010;
											assign node6273 = (inp[9]) ? 11'b10000110010 : 11'b10010110010;
										assign node6276 = (inp[3]) ? node6284 : node6277;
											assign node6277 = (inp[9]) ? node6281 : node6278;
												assign node6278 = (inp[4]) ? 11'b10100110110 : 11'b10000100010;
												assign node6281 = (inp[4]) ? 11'b10110110000 : 11'b10100110100;
											assign node6284 = (inp[4]) ? node6288 : node6285;
												assign node6285 = (inp[9]) ? 11'b00010110100 : 11'b00010110110;
												assign node6288 = (inp[9]) ? 11'b00100110000 : 11'b00110110010;
									assign node6291 = (inp[4]) ? node6307 : node6292;
										assign node6292 = (inp[3]) ? node6300 : node6293;
											assign node6293 = (inp[10]) ? node6297 : node6294;
												assign node6294 = (inp[9]) ? 11'b00101100000 : 11'b00001110010;
												assign node6297 = (inp[9]) ? 11'b10110100110 : 11'b10101110000;
											assign node6300 = (inp[10]) ? node6304 : node6301;
												assign node6301 = (inp[9]) ? 11'b10001110100 : 11'b10111100000;
												assign node6304 = (inp[9]) ? 11'b00000100110 : 11'b00011100100;
										assign node6307 = (inp[3]) ? node6315 : node6308;
											assign node6308 = (inp[10]) ? node6312 : node6309;
												assign node6309 = (inp[9]) ? 11'b00000100100 : 11'b00010110110;
												assign node6312 = (inp[9]) ? 11'b10010100000 : 11'b10000100110;
											assign node6315 = (inp[10]) ? node6319 : node6316;
												assign node6316 = (inp[9]) ? 11'b10110100000 : 11'b10100110110;
												assign node6319 = (inp[9]) ? 11'b00100100000 : 11'b00110100000;
								assign node6322 = (inp[10]) ? node6348 : node6323;
									assign node6323 = (inp[9]) ? node6337 : node6324;
										assign node6324 = (inp[4]) ? node6330 : node6325;
											assign node6325 = (inp[3]) ? 11'b00101100000 : node6326;
												assign node6326 = (inp[5]) ? 11'b00011110000 : 11'b00010110010;
											assign node6330 = (inp[5]) ? node6334 : node6331;
												assign node6331 = (inp[3]) ? 11'b00110110010 : 11'b00000110000;
												assign node6334 = (inp[3]) ? 11'b00000110010 : 11'b00110110010;
										assign node6337 = (inp[3]) ? node6343 : node6338;
											assign node6338 = (inp[5]) ? node6340 : 11'b00110110100;
												assign node6340 = (inp[4]) ? 11'b00100100100 : 11'b00101110100;
											assign node6343 = (inp[5]) ? 11'b00010110010 : node6344;
												assign node6344 = (inp[4]) ? 11'b00110100000 : 11'b00100110000;
									assign node6348 = (inp[9]) ? node6360 : node6349;
										assign node6349 = (inp[3]) ? node6353 : node6350;
											assign node6350 = (inp[5]) ? 11'b00001110100 : 11'b00010110110;
											assign node6353 = (inp[4]) ? node6357 : node6354;
												assign node6354 = (inp[5]) ? 11'b00111100000 : 11'b00100100010;
												assign node6357 = (inp[5]) ? 11'b00010100000 : 11'b00010100010;
										assign node6360 = (inp[3]) ? node6366 : node6361;
											assign node6361 = (inp[4]) ? 11'b00100100000 : node6362;
												assign node6362 = (inp[5]) ? 11'b00100100010 : 11'b00000100000;
											assign node6366 = (inp[4]) ? 11'b00000100000 : node6367;
												assign node6367 = (inp[5]) ? 11'b00000100010 : 11'b00010100000;
						assign node6371 = (inp[5]) ? node6479 : node6372;
							assign node6372 = (inp[11]) ? node6426 : node6373;
								assign node6373 = (inp[4]) ? node6399 : node6374;
									assign node6374 = (inp[9]) ? node6386 : node6375;
										assign node6375 = (inp[10]) ? node6381 : node6376;
											assign node6376 = (inp[3]) ? node6378 : 11'b00110100010;
												assign node6378 = (inp[0]) ? 11'b00000100010 : 11'b10100100010;
											assign node6381 = (inp[3]) ? node6383 : 11'b00110100110;
												assign node6383 = (inp[0]) ? 11'b00010100010 : 11'b00110100110;
										assign node6386 = (inp[3]) ? node6392 : node6387;
											assign node6387 = (inp[10]) ? 11'b10010110100 : node6388;
												assign node6388 = (inp[0]) ? 11'b00100100110 : 11'b00000100010;
											assign node6392 = (inp[0]) ? node6396 : node6393;
												assign node6393 = (inp[10]) ? 11'b00100110100 : 11'b10110100100;
												assign node6396 = (inp[10]) ? 11'b00000100000 : 11'b00010110000;
									assign node6399 = (inp[9]) ? node6411 : node6400;
										assign node6400 = (inp[10]) ? node6406 : node6401;
											assign node6401 = (inp[3]) ? 11'b00000110000 : node6402;
												assign node6402 = (inp[0]) ? 11'b00110100000 : 11'b00110100100;
											assign node6406 = (inp[3]) ? node6408 : 11'b00111010110;
												assign node6408 = (inp[0]) ? 11'b00111000010 : 11'b00011000010;
										assign node6411 = (inp[10]) ? node6419 : node6412;
											assign node6412 = (inp[3]) ? node6416 : node6413;
												assign node6413 = (inp[0]) ? 11'b00001010110 : 11'b00101000110;
												assign node6416 = (inp[0]) ? 11'b00111000010 : 11'b10001010010;
											assign node6419 = (inp[3]) ? node6423 : node6420;
												assign node6420 = (inp[0]) ? 11'b00011010010 : 11'b10011000010;
												assign node6423 = (inp[0]) ? 11'b00001000010 : 11'b00101010010;
								assign node6426 = (inp[0]) ? node6452 : node6427;
									assign node6427 = (inp[4]) ? node6441 : node6428;
										assign node6428 = (inp[10]) ? node6436 : node6429;
											assign node6429 = (inp[3]) ? node6433 : node6430;
												assign node6430 = (inp[9]) ? 11'b00111010000 : 11'b00001000010;
												assign node6433 = (inp[9]) ? 11'b10101000100 : 11'b10111010000;
											assign node6436 = (inp[3]) ? 11'b00001010100 : node6437;
												assign node6437 = (inp[9]) ? 11'b10001010100 : 11'b10101000000;
										assign node6441 = (inp[10]) ? node6447 : node6442;
											assign node6442 = (inp[3]) ? 11'b10001000110 : node6443;
												assign node6443 = (inp[9]) ? 11'b00001010110 : 11'b00101000110;
											assign node6447 = (inp[3]) ? node6449 : 11'b10111010110;
												assign node6449 = (inp[9]) ? 11'b00101010000 : 11'b00101010010;
									assign node6452 = (inp[10]) ? node6466 : node6453;
										assign node6453 = (inp[4]) ? node6461 : node6454;
											assign node6454 = (inp[3]) ? node6458 : node6455;
												assign node6455 = (inp[9]) ? 11'b00011010100 : 11'b00111010000;
												assign node6458 = (inp[9]) ? 11'b00101010000 : 11'b00011000000;
											assign node6461 = (inp[9]) ? 11'b00111000000 : node6462;
												assign node6462 = (inp[3]) ? 11'b00111010010 : 11'b00101010010;
										assign node6466 = (inp[4]) ? node6474 : node6467;
											assign node6467 = (inp[9]) ? node6471 : node6468;
												assign node6468 = (inp[3]) ? 11'b00111000000 : 11'b00101010100;
												assign node6471 = (inp[3]) ? 11'b00011000010 : 11'b00111000010;
											assign node6474 = (inp[9]) ? 11'b00001000000 : node6475;
												assign node6475 = (inp[3]) ? 11'b00001000010 : 11'b00011000110;
							assign node6479 = (inp[4]) ? node6535 : node6480;
								assign node6480 = (inp[9]) ? node6510 : node6481;
									assign node6481 = (inp[0]) ? node6495 : node6482;
										assign node6482 = (inp[11]) ? node6490 : node6483;
											assign node6483 = (inp[10]) ? node6487 : node6484;
												assign node6484 = (inp[3]) ? 11'b10011010000 : 11'b00011010000;
												assign node6487 = (inp[3]) ? 11'b00110010110 : 11'b10101010000;
											assign node6490 = (inp[3]) ? 11'b10010000010 : node6491;
												assign node6491 = (inp[10]) ? 11'b10010010010 : 11'b00000010000;
										assign node6495 = (inp[11]) ? node6503 : node6496;
											assign node6496 = (inp[10]) ? node6500 : node6497;
												assign node6497 = (inp[3]) ? 11'b00101000000 : 11'b00111000000;
												assign node6500 = (inp[3]) ? 11'b00010000010 : 11'b00001000100;
											assign node6503 = (inp[10]) ? node6507 : node6504;
												assign node6504 = (inp[3]) ? 11'b00110000010 : 11'b00110010010;
												assign node6507 = (inp[3]) ? 11'b00100000010 : 11'b00100010110;
									assign node6510 = (inp[0]) ? node6522 : node6511;
										assign node6511 = (inp[3]) ? node6517 : node6512;
											assign node6512 = (inp[10]) ? 11'b10000000110 : node6513;
												assign node6513 = (inp[11]) ? 11'b00000000010 : 11'b00010010010;
											assign node6517 = (inp[10]) ? 11'b00110000110 : node6518;
												assign node6518 = (inp[11]) ? 11'b10110010110 : 11'b10000010110;
										assign node6522 = (inp[10]) ? node6530 : node6523;
											assign node6523 = (inp[11]) ? node6527 : node6524;
												assign node6524 = (inp[3]) ? 11'b00100010010 : 11'b00100000110;
												assign node6527 = (inp[3]) ? 11'b00010010010 : 11'b00010010110;
											assign node6530 = (inp[11]) ? 11'b00000000010 : node6531;
												assign node6531 = (inp[3]) ? 11'b00010000010 : 11'b00010010010;
								assign node6535 = (inp[0]) ? node6559 : node6536;
									assign node6536 = (inp[9]) ? node6548 : node6537;
										assign node6537 = (inp[11]) ? node6543 : node6538;
											assign node6538 = (inp[10]) ? node6540 : 11'b10000010110;
												assign node6540 = (inp[3]) ? 11'b00010010000 : 11'b10010000100;
											assign node6543 = (inp[10]) ? node6545 : 11'b00110010100;
												assign node6545 = (inp[3]) ? 11'b00100000000 : 11'b10100000100;
										assign node6548 = (inp[3]) ? node6556 : node6549;
											assign node6549 = (inp[10]) ? node6553 : node6550;
												assign node6550 = (inp[11]) ? 11'b00110000100 : 11'b00100010100;
												assign node6553 = (inp[11]) ? 11'b10100000000 : 11'b10110010000;
											assign node6556 = (inp[10]) ? 11'b00100000000 : 11'b10110000000;
									assign node6559 = (inp[3]) ? node6569 : node6560;
										assign node6560 = (inp[11]) ? node6564 : node6561;
											assign node6561 = (inp[10]) ? 11'b00010010000 : 11'b00000010100;
											assign node6564 = (inp[10]) ? 11'b00000000100 : node6565;
												assign node6565 = (inp[9]) ? 11'b00010000100 : 11'b00010010000;
										assign node6569 = (inp[10]) ? node6573 : node6570;
											assign node6570 = (inp[9]) ? 11'b00010000000 : 11'b00110010000;
											assign node6573 = (inp[9]) ? 11'b00000000000 : node6574;
												assign node6574 = (inp[11]) ? 11'b00000000000 : 11'b00100000000;
					assign node6578 = (inp[0]) ? node6790 : node6579;
						assign node6579 = (inp[8]) ? node6697 : node6580;
							assign node6580 = (inp[5]) ? node6634 : node6581;
								assign node6581 = (inp[4]) ? node6611 : node6582;
									assign node6582 = (inp[9]) ? node6598 : node6583;
										assign node6583 = (inp[10]) ? node6591 : node6584;
											assign node6584 = (inp[3]) ? node6588 : node6585;
												assign node6585 = (inp[11]) ? 11'b00101000000 : 11'b00111000010;
												assign node6588 = (inp[11]) ? 11'b10111010010 : 11'b10111000010;
											assign node6591 = (inp[3]) ? node6595 : node6592;
												assign node6592 = (inp[11]) ? 11'b10111000010 : 11'b10101000010;
												assign node6595 = (inp[11]) ? 11'b00101010110 : 11'b00101000110;
										assign node6598 = (inp[10]) ? node6604 : node6599;
											assign node6599 = (inp[3]) ? node6601 : 11'b00001010010;
												assign node6601 = (inp[11]) ? 11'b10001000110 : 11'b10111000110;
											assign node6604 = (inp[3]) ? node6608 : node6605;
												assign node6605 = (inp[11]) ? 11'b10011010110 : 11'b10101010110;
												assign node6608 = (inp[11]) ? 11'b00111010110 : 11'b00101010110;
									assign node6611 = (inp[9]) ? node6621 : node6612;
										assign node6612 = (inp[11]) ? node6616 : node6613;
											assign node6613 = (inp[3]) ? 11'b10111000100 : 11'b00111000100;
											assign node6616 = (inp[10]) ? 11'b10001010110 : node6617;
												assign node6617 = (inp[3]) ? 11'b10001000110 : 11'b00101000110;
										assign node6621 = (inp[11]) ? node6629 : node6622;
											assign node6622 = (inp[3]) ? node6626 : node6623;
												assign node6623 = (inp[10]) ? 11'b10011000000 : 11'b00001000100;
												assign node6626 = (inp[10]) ? 11'b00001010000 : 11'b10011010000;
											assign node6629 = (inp[10]) ? 11'b10001010000 : node6630;
												assign node6630 = (inp[3]) ? 11'b10101010000 : 11'b00111010100;
								assign node6634 = (inp[11]) ? node6666 : node6635;
									assign node6635 = (inp[4]) ? node6651 : node6636;
										assign node6636 = (inp[9]) ? node6644 : node6637;
											assign node6637 = (inp[10]) ? node6641 : node6638;
												assign node6638 = (inp[3]) ? 11'b10111010000 : 11'b00111010000;
												assign node6641 = (inp[3]) ? 11'b00001010100 : 11'b10011010000;
											assign node6644 = (inp[10]) ? node6648 : node6645;
												assign node6645 = (inp[3]) ? 11'b10110010110 : 11'b00101010000;
												assign node6648 = (inp[3]) ? 11'b00110000110 : 11'b10010000110;
										assign node6651 = (inp[10]) ? node6659 : node6652;
											assign node6652 = (inp[9]) ? node6656 : node6653;
												assign node6653 = (inp[3]) ? 11'b10000010110 : 11'b00100010110;
												assign node6656 = (inp[3]) ? 11'b10110000010 : 11'b00010010110;
											assign node6659 = (inp[3]) ? node6663 : node6660;
												assign node6660 = (inp[9]) ? 11'b10100010010 : 11'b10100000110;
												assign node6663 = (inp[9]) ? 11'b00000000010 : 11'b00110010010;
									assign node6666 = (inp[9]) ? node6682 : node6667;
										assign node6667 = (inp[10]) ? node6675 : node6668;
											assign node6668 = (inp[4]) ? node6672 : node6669;
												assign node6669 = (inp[3]) ? 11'b10000000010 : 11'b00100010010;
												assign node6672 = (inp[3]) ? 11'b10010010100 : 11'b00110010100;
											assign node6675 = (inp[3]) ? node6679 : node6676;
												assign node6676 = (inp[4]) ? 11'b10110000100 : 11'b10010010000;
												assign node6679 = (inp[4]) ? 11'b00010000000 : 11'b00110000100;
										assign node6682 = (inp[4]) ? node6690 : node6683;
											assign node6683 = (inp[3]) ? node6687 : node6684;
												assign node6684 = (inp[10]) ? 11'b10000000100 : 11'b00010000000;
												assign node6687 = (inp[10]) ? 11'b00100000100 : 11'b10100010100;
											assign node6690 = (inp[3]) ? node6694 : node6691;
												assign node6691 = (inp[10]) ? 11'b10100000000 : 11'b00100000100;
												assign node6694 = (inp[10]) ? 11'b00000000000 : 11'b10000000000;
							assign node6697 = (inp[5]) ? node6751 : node6698;
								assign node6698 = (inp[11]) ? node6726 : node6699;
									assign node6699 = (inp[9]) ? node6713 : node6700;
										assign node6700 = (inp[4]) ? node6706 : node6701;
											assign node6701 = (inp[3]) ? node6703 : 11'b10110000010;
												assign node6703 = (inp[10]) ? 11'b00010000110 : 11'b10010000010;
											assign node6706 = (inp[3]) ? node6710 : node6707;
												assign node6707 = (inp[10]) ? 11'b10010010110 : 11'b00000000110;
												assign node6710 = (inp[10]) ? 11'b00110000010 : 11'b10110000110;
										assign node6713 = (inp[3]) ? node6721 : node6714;
											assign node6714 = (inp[10]) ? node6718 : node6715;
												assign node6715 = (inp[4]) ? 11'b00010000110 : 11'b00100000010;
												assign node6718 = (inp[4]) ? 11'b10100000010 : 11'b10100010110;
											assign node6721 = (inp[4]) ? node6723 : 11'b10000000110;
												assign node6723 = (inp[10]) ? 11'b00000010010 : 11'b10100010010;
									assign node6726 = (inp[4]) ? node6742 : node6727;
										assign node6727 = (inp[9]) ? node6735 : node6728;
											assign node6728 = (inp[3]) ? node6732 : node6729;
												assign node6729 = (inp[10]) ? 11'b10000000010 : 11'b00100000010;
												assign node6732 = (inp[10]) ? 11'b00110010100 : 11'b10000010010;
											assign node6735 = (inp[10]) ? node6739 : node6736;
												assign node6736 = (inp[3]) ? 11'b10010000100 : 11'b00010010000;
												assign node6739 = (inp[3]) ? 11'b00010010100 : 11'b10110010100;
										assign node6742 = (inp[10]) ? node6748 : node6743;
											assign node6743 = (inp[9]) ? node6745 : 11'b10100000100;
												assign node6745 = (inp[3]) ? 11'b10100010000 : 11'b00100010100;
											assign node6748 = (inp[3]) ? 11'b00000010000 : 11'b10000010000;
								assign node6751 = (inp[10]) ? node6771 : node6752;
									assign node6752 = (inp[4]) ? node6764 : node6753;
										assign node6753 = (inp[11]) ? node6759 : node6754;
											assign node6754 = (inp[3]) ? node6756 : 11'b00110010000;
												assign node6756 = (inp[9]) ? 11'b10110010100 : 11'b10110010000;
											assign node6759 = (inp[3]) ? 11'b10100000000 : node6760;
												assign node6760 = (inp[9]) ? 11'b00100000000 : 11'b00100010000;
										assign node6764 = (inp[3]) ? node6766 : 11'b00000010100;
											assign node6766 = (inp[9]) ? 11'b10000000000 : node6767;
												assign node6767 = (inp[11]) ? 11'b10000010100 : 11'b10100010100;
									assign node6771 = (inp[3]) ? node6783 : node6772;
										assign node6772 = (inp[11]) ? node6776 : node6773;
											assign node6773 = (inp[4]) ? 11'b10100000100 : 11'b10110000100;
											assign node6776 = (inp[4]) ? node6780 : node6777;
												assign node6777 = (inp[9]) ? 11'b10000000100 : 11'b10100010000;
												assign node6780 = (inp[9]) ? 11'b10000000000 : 11'b10000000100;
										assign node6783 = (inp[4]) ? 11'b00000000000 : node6784;
											assign node6784 = (inp[11]) ? node6786 : 11'b00010000100;
												assign node6786 = (inp[9]) ? 11'b00000000100 : 11'b00100000100;
						assign node6790 = (inp[8]) ? node6894 : node6791;
							assign node6791 = (inp[5]) ? node6837 : node6792;
								assign node6792 = (inp[4]) ? node6814 : node6793;
									assign node6793 = (inp[10]) ? node6807 : node6794;
										assign node6794 = (inp[9]) ? node6800 : node6795;
											assign node6795 = (inp[3]) ? 11'b00011000010 : node6796;
												assign node6796 = (inp[11]) ? 11'b00001010000 : 11'b00011000010;
											assign node6800 = (inp[3]) ? node6804 : node6801;
												assign node6801 = (inp[11]) ? 11'b00101010110 : 11'b00011000110;
												assign node6804 = (inp[11]) ? 11'b00111010010 : 11'b00011010010;
										assign node6807 = (inp[11]) ? node6811 : node6808;
											assign node6808 = (inp[3]) ? 11'b00001000010 : 11'b00001010010;
											assign node6811 = (inp[9]) ? 11'b00011000010 : 11'b00101000010;
									assign node6814 = (inp[10]) ? node6828 : node6815;
										assign node6815 = (inp[9]) ? node6823 : node6816;
											assign node6816 = (inp[11]) ? node6820 : node6817;
												assign node6817 = (inp[3]) ? 11'b00011010000 : 11'b00011000000;
												assign node6820 = (inp[3]) ? 11'b00101010010 : 11'b00001010010;
											assign node6823 = (inp[11]) ? 11'b00011000100 : node6824;
												assign node6824 = (inp[3]) ? 11'b00111000000 : 11'b00111010100;
										assign node6828 = (inp[9]) ? node6834 : node6829;
											assign node6829 = (inp[11]) ? node6831 : 11'b00001010100;
												assign node6831 = (inp[3]) ? 11'b00011000000 : 11'b00111000100;
											assign node6834 = (inp[3]) ? 11'b00001000000 : 11'b00101000000;
								assign node6837 = (inp[11]) ? node6869 : node6838;
									assign node6838 = (inp[4]) ? node6854 : node6839;
										assign node6839 = (inp[9]) ? node6847 : node6840;
											assign node6840 = (inp[10]) ? node6844 : node6841;
												assign node6841 = (inp[3]) ? 11'b00111000000 : 11'b00011000000;
												assign node6844 = (inp[3]) ? 11'b00001000000 : 11'b00101000100;
											assign node6847 = (inp[10]) ? node6851 : node6848;
												assign node6848 = (inp[3]) ? 11'b00110010010 : 11'b00001000100;
												assign node6851 = (inp[3]) ? 11'b00010000010 : 11'b00110010010;
										assign node6854 = (inp[3]) ? node6862 : node6855;
											assign node6855 = (inp[9]) ? node6859 : node6856;
												assign node6856 = (inp[10]) ? 11'b00000010110 : 11'b00100000010;
												assign node6859 = (inp[10]) ? 11'b00100010010 : 11'b00110010110;
											assign node6862 = (inp[9]) ? node6866 : node6863;
												assign node6863 = (inp[10]) ? 11'b00110000010 : 11'b00100010010;
												assign node6866 = (inp[10]) ? 11'b00000000010 : 11'b00010000010;
									assign node6869 = (inp[9]) ? node6883 : node6870;
										assign node6870 = (inp[10]) ? node6876 : node6871;
											assign node6871 = (inp[4]) ? node6873 : 11'b00000010010;
												assign node6873 = (inp[3]) ? 11'b00010010000 : 11'b00110010000;
											assign node6876 = (inp[3]) ? node6880 : node6877;
												assign node6877 = (inp[4]) ? 11'b00110000100 : 11'b00010010100;
												assign node6880 = (inp[4]) ? 11'b00010000000 : 11'b00110000000;
										assign node6883 = (inp[3]) ? node6889 : node6884;
											assign node6884 = (inp[10]) ? 11'b00100000000 : node6885;
												assign node6885 = (inp[4]) ? 11'b00100000100 : 11'b00100010100;
											assign node6889 = (inp[10]) ? 11'b00000000000 : node6890;
												assign node6890 = (inp[4]) ? 11'b00000000000 : 11'b00000010000;
							assign node6894 = (inp[5]) ? node6948 : node6895;
								assign node6895 = (inp[11]) ? node6923 : node6896;
									assign node6896 = (inp[9]) ? node6910 : node6897;
										assign node6897 = (inp[3]) ? node6903 : node6898;
											assign node6898 = (inp[10]) ? node6900 : 11'b00110000010;
												assign node6900 = (inp[4]) ? 11'b00110010110 : 11'b00110000110;
											assign node6903 = (inp[10]) ? node6907 : node6904;
												assign node6904 = (inp[4]) ? 11'b00010010010 : 11'b00010000010;
												assign node6907 = (inp[4]) ? 11'b00110000010 : 11'b00010000010;
										assign node6910 = (inp[3]) ? node6916 : node6911;
											assign node6911 = (inp[10]) ? node6913 : 11'b00010010110;
												assign node6913 = (inp[4]) ? 11'b00000010010 : 11'b00100010010;
											assign node6916 = (inp[4]) ? node6920 : node6917;
												assign node6917 = (inp[10]) ? 11'b00000000010 : 11'b00000010010;
												assign node6920 = (inp[10]) ? 11'b00000000010 : 11'b00100000010;
									assign node6923 = (inp[4]) ? node6937 : node6924;
										assign node6924 = (inp[3]) ? node6930 : node6925;
											assign node6925 = (inp[9]) ? 11'b00010010100 : node6926;
												assign node6926 = (inp[10]) ? 11'b00110010100 : 11'b00100010010;
											assign node6930 = (inp[9]) ? node6934 : node6931;
												assign node6931 = (inp[10]) ? 11'b00110000000 : 11'b00000000010;
												assign node6934 = (inp[10]) ? 11'b00010000000 : 11'b00110010000;
										assign node6937 = (inp[10]) ? node6943 : node6938;
											assign node6938 = (inp[9]) ? node6940 : 11'b00100010000;
												assign node6940 = (inp[3]) ? 11'b00100000000 : 11'b00100000100;
											assign node6943 = (inp[9]) ? 11'b00000000000 : node6944;
												assign node6944 = (inp[3]) ? 11'b00000000000 : 11'b00000000100;
								assign node6948 = (inp[11]) ? node6976 : node6949;
									assign node6949 = (inp[4]) ? node6963 : node6950;
										assign node6950 = (inp[10]) ? node6956 : node6951;
											assign node6951 = (inp[3]) ? 11'b00110010000 : node6952;
												assign node6952 = (inp[9]) ? 11'b00110000100 : 11'b00110000000;
											assign node6956 = (inp[9]) ? node6960 : node6957;
												assign node6957 = (inp[3]) ? 11'b00010000000 : 11'b00010000100;
												assign node6960 = (inp[3]) ? 11'b00010000000 : 11'b00010010000;
										assign node6963 = (inp[3]) ? node6971 : node6964;
											assign node6964 = (inp[10]) ? node6968 : node6965;
												assign node6965 = (inp[9]) ? 11'b00000010100 : 11'b00010000000;
												assign node6968 = (inp[9]) ? 11'b00000010000 : 11'b00100010100;
											assign node6971 = (inp[9]) ? 11'b00000000000 : node6972;
												assign node6972 = (inp[10]) ? 11'b00100000000 : 11'b00100010000;
									assign node6976 = (inp[9]) ? node6988 : node6977;
										assign node6977 = (inp[4]) ? node6983 : node6978;
											assign node6978 = (inp[3]) ? 11'b00100000000 : node6979;
												assign node6979 = (inp[10]) ? 11'b00100010100 : 11'b00100010000;
											assign node6983 = (inp[10]) ? node6985 : 11'b00000010000;
												assign node6985 = (inp[3]) ? 11'b00000000000 : 11'b00000000100;
										assign node6988 = (inp[10]) ? 11'b00000000000 : node6989;
											assign node6989 = (inp[4]) ? node6991 : 11'b00000010000;
												assign node6991 = (inp[3]) ? 11'b00000000000 : 11'b00000000100;

endmodule