module dtc_split66_bm15 (
	input  wire [15-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node14;
	wire [1-1:0] node17;
	wire [1-1:0] node18;
	wire [1-1:0] node20;
	wire [1-1:0] node22;
	wire [1-1:0] node24;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node30;
	wire [1-1:0] node32;
	wire [1-1:0] node35;
	wire [1-1:0] node36;
	wire [1-1:0] node38;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node45;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node50;
	wire [1-1:0] node52;
	wire [1-1:0] node54;
	wire [1-1:0] node56;
	wire [1-1:0] node59;
	wire [1-1:0] node60;
	wire [1-1:0] node62;
	wire [1-1:0] node64;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node70;
	wire [1-1:0] node73;
	wire [1-1:0] node74;
	wire [1-1:0] node77;
	wire [1-1:0] node80;
	wire [1-1:0] node81;
	wire [1-1:0] node82;
	wire [1-1:0] node84;
	wire [1-1:0] node86;
	wire [1-1:0] node89;
	wire [1-1:0] node90;
	wire [1-1:0] node92;
	wire [1-1:0] node95;
	wire [1-1:0] node96;
	wire [1-1:0] node99;
	wire [1-1:0] node102;
	wire [1-1:0] node103;
	wire [1-1:0] node104;
	wire [1-1:0] node106;
	wire [1-1:0] node109;
	wire [1-1:0] node110;
	wire [1-1:0] node113;
	wire [1-1:0] node116;
	wire [1-1:0] node117;
	wire [1-1:0] node118;
	wire [1-1:0] node121;
	wire [1-1:0] node124;
	wire [1-1:0] node125;
	wire [1-1:0] node128;
	wire [1-1:0] node131;
	wire [1-1:0] node132;
	wire [1-1:0] node133;
	wire [1-1:0] node134;
	wire [1-1:0] node136;
	wire [1-1:0] node138;
	wire [1-1:0] node140;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node146;
	wire [1-1:0] node148;
	wire [1-1:0] node151;
	wire [1-1:0] node152;
	wire [1-1:0] node154;
	wire [1-1:0] node157;
	wire [1-1:0] node158;
	wire [1-1:0] node161;
	wire [1-1:0] node164;
	wire [1-1:0] node165;
	wire [1-1:0] node166;
	wire [1-1:0] node168;
	wire [1-1:0] node170;
	wire [1-1:0] node173;
	wire [1-1:0] node174;
	wire [1-1:0] node176;
	wire [1-1:0] node179;
	wire [1-1:0] node180;
	wire [1-1:0] node183;
	wire [1-1:0] node186;
	wire [1-1:0] node187;
	wire [1-1:0] node188;
	wire [1-1:0] node190;
	wire [1-1:0] node193;
	wire [1-1:0] node194;
	wire [1-1:0] node197;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node205;
	wire [1-1:0] node208;
	wire [1-1:0] node209;
	wire [1-1:0] node212;
	wire [1-1:0] node215;
	wire [1-1:0] node216;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node220;
	wire [1-1:0] node222;
	wire [1-1:0] node225;
	wire [1-1:0] node226;
	wire [1-1:0] node228;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node235;
	wire [1-1:0] node238;
	wire [1-1:0] node239;
	wire [1-1:0] node240;
	wire [1-1:0] node242;
	wire [1-1:0] node245;
	wire [1-1:0] node246;
	wire [1-1:0] node249;
	wire [1-1:0] node252;
	wire [1-1:0] node253;
	wire [1-1:0] node254;
	wire [1-1:0] node257;
	wire [1-1:0] node260;
	wire [1-1:0] node261;
	wire [1-1:0] node264;
	wire [1-1:0] node267;
	wire [1-1:0] node268;
	wire [1-1:0] node269;
	wire [1-1:0] node270;
	wire [1-1:0] node272;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node279;
	wire [1-1:0] node282;
	wire [1-1:0] node283;
	wire [1-1:0] node284;
	wire [1-1:0] node287;
	wire [1-1:0] node290;
	wire [1-1:0] node291;
	wire [1-1:0] node294;
	wire [1-1:0] node297;
	wire [1-1:0] node298;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node303;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node310;
	wire [1-1:0] node313;
	wire [1-1:0] node314;
	wire [1-1:0] node315;
	wire [1-1:0] node318;
	wire [1-1:0] node321;
	wire [1-1:0] node322;
	wire [1-1:0] node326;
	wire [1-1:0] node327;
	wire [1-1:0] node328;
	wire [1-1:0] node329;
	wire [1-1:0] node330;
	wire [1-1:0] node332;
	wire [1-1:0] node334;
	wire [1-1:0] node336;
	wire [1-1:0] node339;
	wire [1-1:0] node340;
	wire [1-1:0] node342;
	wire [1-1:0] node344;
	wire [1-1:0] node347;
	wire [1-1:0] node348;
	wire [1-1:0] node350;
	wire [1-1:0] node353;
	wire [1-1:0] node354;
	wire [1-1:0] node357;
	wire [1-1:0] node360;
	wire [1-1:0] node361;
	wire [1-1:0] node362;
	wire [1-1:0] node364;
	wire [1-1:0] node366;
	wire [1-1:0] node369;
	wire [1-1:0] node370;
	wire [1-1:0] node372;
	wire [1-1:0] node375;
	wire [1-1:0] node376;
	wire [1-1:0] node379;
	wire [1-1:0] node382;
	wire [1-1:0] node383;
	wire [1-1:0] node384;
	wire [1-1:0] node386;
	wire [1-1:0] node389;
	wire [1-1:0] node390;
	wire [1-1:0] node393;
	wire [1-1:0] node396;
	wire [1-1:0] node397;
	wire [1-1:0] node398;
	wire [1-1:0] node401;
	wire [1-1:0] node404;
	wire [1-1:0] node405;
	wire [1-1:0] node408;
	wire [1-1:0] node411;
	wire [1-1:0] node412;
	wire [1-1:0] node413;
	wire [1-1:0] node414;
	wire [1-1:0] node416;
	wire [1-1:0] node418;
	wire [1-1:0] node421;
	wire [1-1:0] node422;
	wire [1-1:0] node424;
	wire [1-1:0] node427;
	wire [1-1:0] node428;
	wire [1-1:0] node431;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node438;
	wire [1-1:0] node441;
	wire [1-1:0] node442;
	wire [1-1:0] node445;
	wire [1-1:0] node448;
	wire [1-1:0] node449;
	wire [1-1:0] node450;
	wire [1-1:0] node453;
	wire [1-1:0] node456;
	wire [1-1:0] node457;
	wire [1-1:0] node460;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node465;
	wire [1-1:0] node466;
	wire [1-1:0] node468;
	wire [1-1:0] node471;
	wire [1-1:0] node472;
	wire [1-1:0] node475;
	wire [1-1:0] node478;
	wire [1-1:0] node479;
	wire [1-1:0] node480;
	wire [1-1:0] node483;
	wire [1-1:0] node486;
	wire [1-1:0] node487;
	wire [1-1:0] node490;
	wire [1-1:0] node493;
	wire [1-1:0] node494;
	wire [1-1:0] node495;
	wire [1-1:0] node496;
	wire [1-1:0] node499;
	wire [1-1:0] node502;
	wire [1-1:0] node503;
	wire [1-1:0] node506;
	wire [1-1:0] node509;
	wire [1-1:0] node510;
	wire [1-1:0] node511;
	wire [1-1:0] node514;
	wire [1-1:0] node517;
	wire [1-1:0] node518;
	wire [1-1:0] node522;
	wire [1-1:0] node523;
	wire [1-1:0] node524;
	wire [1-1:0] node525;
	wire [1-1:0] node526;
	wire [1-1:0] node528;
	wire [1-1:0] node530;
	wire [1-1:0] node533;
	wire [1-1:0] node534;
	wire [1-1:0] node536;
	wire [1-1:0] node539;
	wire [1-1:0] node540;
	wire [1-1:0] node543;
	wire [1-1:0] node546;
	wire [1-1:0] node547;
	wire [1-1:0] node548;
	wire [1-1:0] node550;
	wire [1-1:0] node553;
	wire [1-1:0] node554;
	wire [1-1:0] node557;
	wire [1-1:0] node560;
	wire [1-1:0] node561;
	wire [1-1:0] node562;
	wire [1-1:0] node565;
	wire [1-1:0] node568;
	wire [1-1:0] node569;
	wire [1-1:0] node572;
	wire [1-1:0] node575;
	wire [1-1:0] node576;
	wire [1-1:0] node577;
	wire [1-1:0] node578;
	wire [1-1:0] node580;
	wire [1-1:0] node583;
	wire [1-1:0] node584;
	wire [1-1:0] node587;
	wire [1-1:0] node590;
	wire [1-1:0] node591;
	wire [1-1:0] node592;
	wire [1-1:0] node595;
	wire [1-1:0] node598;
	wire [1-1:0] node599;
	wire [1-1:0] node602;
	wire [1-1:0] node605;
	wire [1-1:0] node606;
	wire [1-1:0] node607;
	wire [1-1:0] node608;
	wire [1-1:0] node611;
	wire [1-1:0] node614;
	wire [1-1:0] node615;
	wire [1-1:0] node618;
	wire [1-1:0] node621;
	wire [1-1:0] node622;
	wire [1-1:0] node623;
	wire [1-1:0] node626;
	wire [1-1:0] node629;
	wire [1-1:0] node630;
	wire [1-1:0] node634;
	wire [1-1:0] node635;
	wire [1-1:0] node636;
	wire [1-1:0] node637;
	wire [1-1:0] node638;
	wire [1-1:0] node640;
	wire [1-1:0] node643;
	wire [1-1:0] node644;
	wire [1-1:0] node647;
	wire [1-1:0] node650;
	wire [1-1:0] node651;
	wire [1-1:0] node652;
	wire [1-1:0] node655;
	wire [1-1:0] node658;
	wire [1-1:0] node659;
	wire [1-1:0] node662;
	wire [1-1:0] node665;
	wire [1-1:0] node666;
	wire [1-1:0] node667;
	wire [1-1:0] node668;
	wire [1-1:0] node671;
	wire [1-1:0] node674;
	wire [1-1:0] node675;
	wire [1-1:0] node678;
	wire [1-1:0] node681;
	wire [1-1:0] node682;
	wire [1-1:0] node683;
	wire [1-1:0] node686;
	wire [1-1:0] node689;
	wire [1-1:0] node690;
	wire [1-1:0] node694;
	wire [1-1:0] node695;
	wire [1-1:0] node696;
	wire [1-1:0] node697;
	wire [1-1:0] node698;
	wire [1-1:0] node701;
	wire [1-1:0] node704;
	wire [1-1:0] node705;
	wire [1-1:0] node708;
	wire [1-1:0] node711;
	wire [1-1:0] node712;
	wire [1-1:0] node713;
	wire [1-1:0] node716;
	wire [1-1:0] node719;
	wire [1-1:0] node720;
	wire [1-1:0] node724;
	wire [1-1:0] node725;
	wire [1-1:0] node726;
	wire [1-1:0] node727;
	wire [1-1:0] node730;
	wire [1-1:0] node733;
	wire [1-1:0] node734;
	wire [1-1:0] node738;
	wire [1-1:0] node739;
	wire [1-1:0] node740;
	wire [1-1:0] node745;
	wire [1-1:0] node746;
	wire [1-1:0] node747;
	wire [1-1:0] node748;
	wire [1-1:0] node749;
	wire [1-1:0] node750;
	wire [1-1:0] node752;
	wire [1-1:0] node754;
	wire [1-1:0] node756;
	wire [1-1:0] node759;
	wire [1-1:0] node760;
	wire [1-1:0] node762;
	wire [1-1:0] node764;
	wire [1-1:0] node767;
	wire [1-1:0] node768;
	wire [1-1:0] node770;
	wire [1-1:0] node773;
	wire [1-1:0] node774;
	wire [1-1:0] node777;
	wire [1-1:0] node780;
	wire [1-1:0] node781;
	wire [1-1:0] node782;
	wire [1-1:0] node784;
	wire [1-1:0] node786;
	wire [1-1:0] node789;
	wire [1-1:0] node790;
	wire [1-1:0] node792;
	wire [1-1:0] node795;
	wire [1-1:0] node796;
	wire [1-1:0] node799;
	wire [1-1:0] node802;
	wire [1-1:0] node803;
	wire [1-1:0] node804;
	wire [1-1:0] node806;
	wire [1-1:0] node809;
	wire [1-1:0] node810;
	wire [1-1:0] node813;
	wire [1-1:0] node816;
	wire [1-1:0] node817;
	wire [1-1:0] node818;
	wire [1-1:0] node821;
	wire [1-1:0] node824;
	wire [1-1:0] node825;
	wire [1-1:0] node828;
	wire [1-1:0] node831;
	wire [1-1:0] node832;
	wire [1-1:0] node833;
	wire [1-1:0] node834;
	wire [1-1:0] node836;
	wire [1-1:0] node838;
	wire [1-1:0] node841;
	wire [1-1:0] node842;
	wire [1-1:0] node844;
	wire [1-1:0] node847;
	wire [1-1:0] node848;
	wire [1-1:0] node851;
	wire [1-1:0] node854;
	wire [1-1:0] node855;
	wire [1-1:0] node856;
	wire [1-1:0] node858;
	wire [1-1:0] node861;
	wire [1-1:0] node862;
	wire [1-1:0] node865;
	wire [1-1:0] node868;
	wire [1-1:0] node869;
	wire [1-1:0] node870;
	wire [1-1:0] node873;
	wire [1-1:0] node876;
	wire [1-1:0] node877;
	wire [1-1:0] node880;
	wire [1-1:0] node883;
	wire [1-1:0] node884;
	wire [1-1:0] node885;
	wire [1-1:0] node886;
	wire [1-1:0] node888;
	wire [1-1:0] node891;
	wire [1-1:0] node892;
	wire [1-1:0] node895;
	wire [1-1:0] node898;
	wire [1-1:0] node899;
	wire [1-1:0] node900;
	wire [1-1:0] node903;
	wire [1-1:0] node906;
	wire [1-1:0] node907;
	wire [1-1:0] node910;
	wire [1-1:0] node913;
	wire [1-1:0] node914;
	wire [1-1:0] node915;
	wire [1-1:0] node916;
	wire [1-1:0] node919;
	wire [1-1:0] node922;
	wire [1-1:0] node923;
	wire [1-1:0] node926;
	wire [1-1:0] node929;
	wire [1-1:0] node930;
	wire [1-1:0] node931;
	wire [1-1:0] node934;
	wire [1-1:0] node937;
	wire [1-1:0] node938;
	wire [1-1:0] node942;
	wire [1-1:0] node943;
	wire [1-1:0] node944;
	wire [1-1:0] node945;
	wire [1-1:0] node946;
	wire [1-1:0] node948;
	wire [1-1:0] node950;
	wire [1-1:0] node953;
	wire [1-1:0] node954;
	wire [1-1:0] node956;
	wire [1-1:0] node959;
	wire [1-1:0] node960;
	wire [1-1:0] node963;
	wire [1-1:0] node966;
	wire [1-1:0] node967;
	wire [1-1:0] node968;
	wire [1-1:0] node970;
	wire [1-1:0] node973;
	wire [1-1:0] node974;
	wire [1-1:0] node977;
	wire [1-1:0] node980;
	wire [1-1:0] node981;
	wire [1-1:0] node982;
	wire [1-1:0] node985;
	wire [1-1:0] node988;
	wire [1-1:0] node989;
	wire [1-1:0] node992;
	wire [1-1:0] node995;
	wire [1-1:0] node996;
	wire [1-1:0] node997;
	wire [1-1:0] node998;
	wire [1-1:0] node1000;
	wire [1-1:0] node1003;
	wire [1-1:0] node1004;
	wire [1-1:0] node1007;
	wire [1-1:0] node1010;
	wire [1-1:0] node1011;
	wire [1-1:0] node1012;
	wire [1-1:0] node1015;
	wire [1-1:0] node1018;
	wire [1-1:0] node1019;
	wire [1-1:0] node1022;
	wire [1-1:0] node1025;
	wire [1-1:0] node1026;
	wire [1-1:0] node1027;
	wire [1-1:0] node1028;
	wire [1-1:0] node1031;
	wire [1-1:0] node1034;
	wire [1-1:0] node1035;
	wire [1-1:0] node1038;
	wire [1-1:0] node1041;
	wire [1-1:0] node1042;
	wire [1-1:0] node1043;
	wire [1-1:0] node1046;
	wire [1-1:0] node1049;
	wire [1-1:0] node1050;
	wire [1-1:0] node1054;
	wire [1-1:0] node1055;
	wire [1-1:0] node1056;
	wire [1-1:0] node1057;
	wire [1-1:0] node1058;
	wire [1-1:0] node1060;
	wire [1-1:0] node1063;
	wire [1-1:0] node1064;
	wire [1-1:0] node1067;
	wire [1-1:0] node1070;
	wire [1-1:0] node1071;
	wire [1-1:0] node1072;
	wire [1-1:0] node1075;
	wire [1-1:0] node1078;
	wire [1-1:0] node1079;
	wire [1-1:0] node1082;
	wire [1-1:0] node1085;
	wire [1-1:0] node1086;
	wire [1-1:0] node1087;
	wire [1-1:0] node1088;
	wire [1-1:0] node1091;
	wire [1-1:0] node1094;
	wire [1-1:0] node1095;
	wire [1-1:0] node1098;
	wire [1-1:0] node1101;
	wire [1-1:0] node1102;
	wire [1-1:0] node1103;
	wire [1-1:0] node1106;
	wire [1-1:0] node1109;
	wire [1-1:0] node1110;
	wire [1-1:0] node1114;
	wire [1-1:0] node1115;
	wire [1-1:0] node1116;
	wire [1-1:0] node1117;
	wire [1-1:0] node1118;
	wire [1-1:0] node1121;
	wire [1-1:0] node1124;
	wire [1-1:0] node1125;
	wire [1-1:0] node1128;
	wire [1-1:0] node1131;
	wire [1-1:0] node1132;
	wire [1-1:0] node1133;
	wire [1-1:0] node1136;
	wire [1-1:0] node1139;
	wire [1-1:0] node1140;
	wire [1-1:0] node1144;
	wire [1-1:0] node1145;
	wire [1-1:0] node1146;
	wire [1-1:0] node1147;
	wire [1-1:0] node1150;
	wire [1-1:0] node1153;
	wire [1-1:0] node1154;
	wire [1-1:0] node1158;
	wire [1-1:0] node1159;
	wire [1-1:0] node1160;
	wire [1-1:0] node1165;
	wire [1-1:0] node1166;
	wire [1-1:0] node1167;
	wire [1-1:0] node1168;
	wire [1-1:0] node1169;
	wire [1-1:0] node1170;
	wire [1-1:0] node1172;
	wire [1-1:0] node1174;
	wire [1-1:0] node1177;
	wire [1-1:0] node1178;
	wire [1-1:0] node1180;
	wire [1-1:0] node1183;
	wire [1-1:0] node1184;
	wire [1-1:0] node1187;
	wire [1-1:0] node1190;
	wire [1-1:0] node1191;
	wire [1-1:0] node1192;
	wire [1-1:0] node1194;
	wire [1-1:0] node1197;
	wire [1-1:0] node1198;
	wire [1-1:0] node1201;
	wire [1-1:0] node1204;
	wire [1-1:0] node1205;
	wire [1-1:0] node1206;
	wire [1-1:0] node1209;
	wire [1-1:0] node1212;
	wire [1-1:0] node1213;
	wire [1-1:0] node1216;
	wire [1-1:0] node1219;
	wire [1-1:0] node1220;
	wire [1-1:0] node1221;
	wire [1-1:0] node1222;
	wire [1-1:0] node1224;
	wire [1-1:0] node1227;
	wire [1-1:0] node1228;
	wire [1-1:0] node1231;
	wire [1-1:0] node1234;
	wire [1-1:0] node1235;
	wire [1-1:0] node1236;
	wire [1-1:0] node1239;
	wire [1-1:0] node1242;
	wire [1-1:0] node1243;
	wire [1-1:0] node1246;
	wire [1-1:0] node1249;
	wire [1-1:0] node1250;
	wire [1-1:0] node1251;
	wire [1-1:0] node1252;
	wire [1-1:0] node1255;
	wire [1-1:0] node1258;
	wire [1-1:0] node1259;
	wire [1-1:0] node1262;
	wire [1-1:0] node1265;
	wire [1-1:0] node1266;
	wire [1-1:0] node1267;
	wire [1-1:0] node1270;
	wire [1-1:0] node1273;
	wire [1-1:0] node1274;
	wire [1-1:0] node1278;
	wire [1-1:0] node1279;
	wire [1-1:0] node1280;
	wire [1-1:0] node1281;
	wire [1-1:0] node1282;
	wire [1-1:0] node1284;
	wire [1-1:0] node1287;
	wire [1-1:0] node1288;
	wire [1-1:0] node1291;
	wire [1-1:0] node1294;
	wire [1-1:0] node1295;
	wire [1-1:0] node1296;
	wire [1-1:0] node1299;
	wire [1-1:0] node1302;
	wire [1-1:0] node1303;
	wire [1-1:0] node1306;
	wire [1-1:0] node1309;
	wire [1-1:0] node1310;
	wire [1-1:0] node1311;
	wire [1-1:0] node1312;
	wire [1-1:0] node1315;
	wire [1-1:0] node1318;
	wire [1-1:0] node1319;
	wire [1-1:0] node1322;
	wire [1-1:0] node1325;
	wire [1-1:0] node1326;
	wire [1-1:0] node1327;
	wire [1-1:0] node1330;
	wire [1-1:0] node1333;
	wire [1-1:0] node1334;
	wire [1-1:0] node1338;
	wire [1-1:0] node1339;
	wire [1-1:0] node1340;
	wire [1-1:0] node1341;
	wire [1-1:0] node1342;
	wire [1-1:0] node1345;
	wire [1-1:0] node1348;
	wire [1-1:0] node1349;
	wire [1-1:0] node1352;
	wire [1-1:0] node1355;
	wire [1-1:0] node1356;
	wire [1-1:0] node1357;
	wire [1-1:0] node1360;
	wire [1-1:0] node1363;
	wire [1-1:0] node1364;
	wire [1-1:0] node1368;
	wire [1-1:0] node1369;
	wire [1-1:0] node1370;
	wire [1-1:0] node1371;
	wire [1-1:0] node1374;
	wire [1-1:0] node1377;
	wire [1-1:0] node1378;
	wire [1-1:0] node1382;
	wire [1-1:0] node1383;
	wire [1-1:0] node1384;
	wire [1-1:0] node1389;
	wire [1-1:0] node1390;
	wire [1-1:0] node1391;
	wire [1-1:0] node1392;
	wire [1-1:0] node1393;
	wire [1-1:0] node1394;
	wire [1-1:0] node1396;
	wire [1-1:0] node1399;
	wire [1-1:0] node1400;
	wire [1-1:0] node1403;
	wire [1-1:0] node1406;
	wire [1-1:0] node1407;
	wire [1-1:0] node1408;
	wire [1-1:0] node1411;
	wire [1-1:0] node1414;
	wire [1-1:0] node1415;
	wire [1-1:0] node1418;
	wire [1-1:0] node1421;
	wire [1-1:0] node1422;
	wire [1-1:0] node1423;
	wire [1-1:0] node1424;
	wire [1-1:0] node1427;
	wire [1-1:0] node1430;
	wire [1-1:0] node1431;
	wire [1-1:0] node1434;
	wire [1-1:0] node1437;
	wire [1-1:0] node1438;
	wire [1-1:0] node1439;
	wire [1-1:0] node1442;
	wire [1-1:0] node1445;
	wire [1-1:0] node1446;
	wire [1-1:0] node1450;
	wire [1-1:0] node1451;
	wire [1-1:0] node1452;
	wire [1-1:0] node1453;
	wire [1-1:0] node1454;
	wire [1-1:0] node1457;
	wire [1-1:0] node1460;
	wire [1-1:0] node1461;
	wire [1-1:0] node1464;
	wire [1-1:0] node1467;
	wire [1-1:0] node1468;
	wire [1-1:0] node1469;
	wire [1-1:0] node1472;
	wire [1-1:0] node1475;
	wire [1-1:0] node1476;
	wire [1-1:0] node1480;
	wire [1-1:0] node1481;
	wire [1-1:0] node1482;
	wire [1-1:0] node1483;
	wire [1-1:0] node1486;
	wire [1-1:0] node1490;
	wire [1-1:0] node1491;
	wire [1-1:0] node1492;
	wire [1-1:0] node1497;
	wire [1-1:0] node1498;
	wire [1-1:0] node1499;
	wire [1-1:0] node1500;
	wire [1-1:0] node1501;
	wire [1-1:0] node1502;
	wire [1-1:0] node1505;
	wire [1-1:0] node1508;
	wire [1-1:0] node1509;
	wire [1-1:0] node1512;
	wire [1-1:0] node1515;
	wire [1-1:0] node1516;
	wire [1-1:0] node1517;
	wire [1-1:0] node1520;
	wire [1-1:0] node1523;
	wire [1-1:0] node1524;
	wire [1-1:0] node1528;
	wire [1-1:0] node1529;
	wire [1-1:0] node1530;
	wire [1-1:0] node1531;
	wire [1-1:0] node1534;
	wire [1-1:0] node1537;
	wire [1-1:0] node1538;
	wire [1-1:0] node1542;
	wire [1-1:0] node1543;
	wire [1-1:0] node1544;
	wire [1-1:0] node1549;
	wire [1-1:0] node1550;
	wire [1-1:0] node1551;
	wire [1-1:0] node1552;
	wire [1-1:0] node1553;
	wire [1-1:0] node1556;
	wire [1-1:0] node1559;
	wire [1-1:0] node1560;
	wire [1-1:0] node1564;
	wire [1-1:0] node1565;
	wire [1-1:0] node1566;
	wire [1-1:0] node1571;
	wire [1-1:0] node1572;
	wire [1-1:0] node1573;
	wire [1-1:0] node1574;
	wire [1-1:0] node1580;
	wire [1-1:0] node1581;
	wire [1-1:0] node1582;
	wire [1-1:0] node1583;
	wire [1-1:0] node1584;
	wire [1-1:0] node1585;
	wire [1-1:0] node1586;
	wire [1-1:0] node1588;
	wire [1-1:0] node1590;
	wire [1-1:0] node1592;
	wire [1-1:0] node1595;
	wire [1-1:0] node1596;
	wire [1-1:0] node1598;
	wire [1-1:0] node1600;
	wire [1-1:0] node1603;
	wire [1-1:0] node1604;
	wire [1-1:0] node1606;
	wire [1-1:0] node1609;
	wire [1-1:0] node1610;
	wire [1-1:0] node1613;
	wire [1-1:0] node1616;
	wire [1-1:0] node1617;
	wire [1-1:0] node1618;
	wire [1-1:0] node1620;
	wire [1-1:0] node1622;
	wire [1-1:0] node1625;
	wire [1-1:0] node1626;
	wire [1-1:0] node1628;
	wire [1-1:0] node1631;
	wire [1-1:0] node1632;
	wire [1-1:0] node1635;
	wire [1-1:0] node1638;
	wire [1-1:0] node1639;
	wire [1-1:0] node1640;
	wire [1-1:0] node1642;
	wire [1-1:0] node1645;
	wire [1-1:0] node1646;
	wire [1-1:0] node1649;
	wire [1-1:0] node1652;
	wire [1-1:0] node1653;
	wire [1-1:0] node1654;
	wire [1-1:0] node1657;
	wire [1-1:0] node1660;
	wire [1-1:0] node1661;
	wire [1-1:0] node1664;
	wire [1-1:0] node1667;
	wire [1-1:0] node1668;
	wire [1-1:0] node1669;
	wire [1-1:0] node1670;
	wire [1-1:0] node1672;
	wire [1-1:0] node1674;
	wire [1-1:0] node1677;
	wire [1-1:0] node1678;
	wire [1-1:0] node1680;
	wire [1-1:0] node1683;
	wire [1-1:0] node1684;
	wire [1-1:0] node1687;
	wire [1-1:0] node1690;
	wire [1-1:0] node1691;
	wire [1-1:0] node1692;
	wire [1-1:0] node1694;
	wire [1-1:0] node1697;
	wire [1-1:0] node1698;
	wire [1-1:0] node1701;
	wire [1-1:0] node1704;
	wire [1-1:0] node1705;
	wire [1-1:0] node1706;
	wire [1-1:0] node1709;
	wire [1-1:0] node1712;
	wire [1-1:0] node1713;
	wire [1-1:0] node1717;
	wire [1-1:0] node1718;
	wire [1-1:0] node1719;
	wire [1-1:0] node1720;
	wire [1-1:0] node1722;
	wire [1-1:0] node1725;
	wire [1-1:0] node1726;
	wire [1-1:0] node1729;
	wire [1-1:0] node1732;
	wire [1-1:0] node1733;
	wire [1-1:0] node1734;
	wire [1-1:0] node1737;
	wire [1-1:0] node1740;
	wire [1-1:0] node1741;
	wire [1-1:0] node1744;
	wire [1-1:0] node1747;
	wire [1-1:0] node1748;
	wire [1-1:0] node1749;
	wire [1-1:0] node1750;
	wire [1-1:0] node1753;
	wire [1-1:0] node1756;
	wire [1-1:0] node1757;
	wire [1-1:0] node1760;
	wire [1-1:0] node1763;
	wire [1-1:0] node1764;
	wire [1-1:0] node1765;
	wire [1-1:0] node1768;
	wire [1-1:0] node1771;
	wire [1-1:0] node1772;
	wire [1-1:0] node1776;
	wire [1-1:0] node1777;
	wire [1-1:0] node1778;
	wire [1-1:0] node1779;
	wire [1-1:0] node1780;
	wire [1-1:0] node1782;
	wire [1-1:0] node1784;
	wire [1-1:0] node1787;
	wire [1-1:0] node1788;
	wire [1-1:0] node1790;
	wire [1-1:0] node1793;
	wire [1-1:0] node1794;
	wire [1-1:0] node1797;
	wire [1-1:0] node1800;
	wire [1-1:0] node1801;
	wire [1-1:0] node1802;
	wire [1-1:0] node1804;
	wire [1-1:0] node1807;
	wire [1-1:0] node1808;
	wire [1-1:0] node1811;
	wire [1-1:0] node1814;
	wire [1-1:0] node1815;
	wire [1-1:0] node1816;
	wire [1-1:0] node1819;
	wire [1-1:0] node1822;
	wire [1-1:0] node1823;
	wire [1-1:0] node1826;
	wire [1-1:0] node1829;
	wire [1-1:0] node1830;
	wire [1-1:0] node1831;
	wire [1-1:0] node1832;
	wire [1-1:0] node1834;
	wire [1-1:0] node1837;
	wire [1-1:0] node1838;
	wire [1-1:0] node1841;
	wire [1-1:0] node1844;
	wire [1-1:0] node1845;
	wire [1-1:0] node1846;
	wire [1-1:0] node1849;
	wire [1-1:0] node1852;
	wire [1-1:0] node1853;
	wire [1-1:0] node1856;
	wire [1-1:0] node1859;
	wire [1-1:0] node1860;
	wire [1-1:0] node1861;
	wire [1-1:0] node1862;
	wire [1-1:0] node1865;
	wire [1-1:0] node1868;
	wire [1-1:0] node1869;
	wire [1-1:0] node1872;
	wire [1-1:0] node1875;
	wire [1-1:0] node1876;
	wire [1-1:0] node1877;
	wire [1-1:0] node1880;
	wire [1-1:0] node1883;
	wire [1-1:0] node1884;
	wire [1-1:0] node1888;
	wire [1-1:0] node1889;
	wire [1-1:0] node1890;
	wire [1-1:0] node1891;
	wire [1-1:0] node1892;
	wire [1-1:0] node1894;
	wire [1-1:0] node1897;
	wire [1-1:0] node1898;
	wire [1-1:0] node1901;
	wire [1-1:0] node1904;
	wire [1-1:0] node1905;
	wire [1-1:0] node1906;
	wire [1-1:0] node1909;
	wire [1-1:0] node1912;
	wire [1-1:0] node1913;
	wire [1-1:0] node1916;
	wire [1-1:0] node1919;
	wire [1-1:0] node1920;
	wire [1-1:0] node1921;
	wire [1-1:0] node1922;
	wire [1-1:0] node1925;
	wire [1-1:0] node1928;
	wire [1-1:0] node1929;
	wire [1-1:0] node1932;
	wire [1-1:0] node1935;
	wire [1-1:0] node1936;
	wire [1-1:0] node1937;
	wire [1-1:0] node1940;
	wire [1-1:0] node1943;
	wire [1-1:0] node1944;
	wire [1-1:0] node1948;
	wire [1-1:0] node1949;
	wire [1-1:0] node1950;
	wire [1-1:0] node1951;
	wire [1-1:0] node1952;
	wire [1-1:0] node1955;
	wire [1-1:0] node1958;
	wire [1-1:0] node1959;
	wire [1-1:0] node1962;
	wire [1-1:0] node1965;
	wire [1-1:0] node1966;
	wire [1-1:0] node1967;
	wire [1-1:0] node1970;
	wire [1-1:0] node1973;
	wire [1-1:0] node1974;
	wire [1-1:0] node1978;
	wire [1-1:0] node1979;
	wire [1-1:0] node1980;
	wire [1-1:0] node1981;
	wire [1-1:0] node1984;
	wire [1-1:0] node1987;
	wire [1-1:0] node1988;
	wire [1-1:0] node1992;
	wire [1-1:0] node1993;
	wire [1-1:0] node1994;
	wire [1-1:0] node1999;
	wire [1-1:0] node2000;
	wire [1-1:0] node2001;
	wire [1-1:0] node2002;
	wire [1-1:0] node2003;
	wire [1-1:0] node2004;
	wire [1-1:0] node2006;
	wire [1-1:0] node2008;
	wire [1-1:0] node2011;
	wire [1-1:0] node2012;
	wire [1-1:0] node2014;
	wire [1-1:0] node2017;
	wire [1-1:0] node2018;
	wire [1-1:0] node2021;
	wire [1-1:0] node2024;
	wire [1-1:0] node2025;
	wire [1-1:0] node2026;
	wire [1-1:0] node2028;
	wire [1-1:0] node2031;
	wire [1-1:0] node2032;
	wire [1-1:0] node2035;
	wire [1-1:0] node2038;
	wire [1-1:0] node2039;
	wire [1-1:0] node2040;
	wire [1-1:0] node2043;
	wire [1-1:0] node2046;
	wire [1-1:0] node2047;
	wire [1-1:0] node2050;
	wire [1-1:0] node2053;
	wire [1-1:0] node2054;
	wire [1-1:0] node2055;
	wire [1-1:0] node2056;
	wire [1-1:0] node2058;
	wire [1-1:0] node2061;
	wire [1-1:0] node2062;
	wire [1-1:0] node2065;
	wire [1-1:0] node2068;
	wire [1-1:0] node2069;
	wire [1-1:0] node2070;
	wire [1-1:0] node2073;
	wire [1-1:0] node2076;
	wire [1-1:0] node2077;
	wire [1-1:0] node2080;
	wire [1-1:0] node2083;
	wire [1-1:0] node2084;
	wire [1-1:0] node2085;
	wire [1-1:0] node2086;
	wire [1-1:0] node2089;
	wire [1-1:0] node2092;
	wire [1-1:0] node2093;
	wire [1-1:0] node2096;
	wire [1-1:0] node2099;
	wire [1-1:0] node2100;
	wire [1-1:0] node2101;
	wire [1-1:0] node2104;
	wire [1-1:0] node2107;
	wire [1-1:0] node2108;
	wire [1-1:0] node2112;
	wire [1-1:0] node2113;
	wire [1-1:0] node2114;
	wire [1-1:0] node2115;
	wire [1-1:0] node2116;
	wire [1-1:0] node2118;
	wire [1-1:0] node2121;
	wire [1-1:0] node2122;
	wire [1-1:0] node2125;
	wire [1-1:0] node2128;
	wire [1-1:0] node2129;
	wire [1-1:0] node2130;
	wire [1-1:0] node2133;
	wire [1-1:0] node2136;
	wire [1-1:0] node2137;
	wire [1-1:0] node2140;
	wire [1-1:0] node2143;
	wire [1-1:0] node2144;
	wire [1-1:0] node2145;
	wire [1-1:0] node2146;
	wire [1-1:0] node2149;
	wire [1-1:0] node2152;
	wire [1-1:0] node2153;
	wire [1-1:0] node2156;
	wire [1-1:0] node2159;
	wire [1-1:0] node2160;
	wire [1-1:0] node2161;
	wire [1-1:0] node2164;
	wire [1-1:0] node2167;
	wire [1-1:0] node2168;
	wire [1-1:0] node2172;
	wire [1-1:0] node2173;
	wire [1-1:0] node2174;
	wire [1-1:0] node2175;
	wire [1-1:0] node2176;
	wire [1-1:0] node2179;
	wire [1-1:0] node2182;
	wire [1-1:0] node2183;
	wire [1-1:0] node2186;
	wire [1-1:0] node2189;
	wire [1-1:0] node2190;
	wire [1-1:0] node2191;
	wire [1-1:0] node2194;
	wire [1-1:0] node2197;
	wire [1-1:0] node2198;
	wire [1-1:0] node2202;
	wire [1-1:0] node2203;
	wire [1-1:0] node2204;
	wire [1-1:0] node2205;
	wire [1-1:0] node2208;
	wire [1-1:0] node2211;
	wire [1-1:0] node2212;
	wire [1-1:0] node2216;
	wire [1-1:0] node2217;
	wire [1-1:0] node2218;
	wire [1-1:0] node2223;
	wire [1-1:0] node2224;
	wire [1-1:0] node2225;
	wire [1-1:0] node2226;
	wire [1-1:0] node2227;
	wire [1-1:0] node2228;
	wire [1-1:0] node2230;
	wire [1-1:0] node2233;
	wire [1-1:0] node2234;
	wire [1-1:0] node2237;
	wire [1-1:0] node2240;
	wire [1-1:0] node2241;
	wire [1-1:0] node2242;
	wire [1-1:0] node2245;
	wire [1-1:0] node2248;
	wire [1-1:0] node2249;
	wire [1-1:0] node2252;
	wire [1-1:0] node2255;
	wire [1-1:0] node2256;
	wire [1-1:0] node2257;
	wire [1-1:0] node2258;
	wire [1-1:0] node2261;
	wire [1-1:0] node2264;
	wire [1-1:0] node2265;
	wire [1-1:0] node2268;
	wire [1-1:0] node2271;
	wire [1-1:0] node2272;
	wire [1-1:0] node2273;
	wire [1-1:0] node2276;
	wire [1-1:0] node2279;
	wire [1-1:0] node2280;
	wire [1-1:0] node2284;
	wire [1-1:0] node2285;
	wire [1-1:0] node2286;
	wire [1-1:0] node2287;
	wire [1-1:0] node2288;
	wire [1-1:0] node2291;
	wire [1-1:0] node2294;
	wire [1-1:0] node2295;
	wire [1-1:0] node2298;
	wire [1-1:0] node2301;
	wire [1-1:0] node2302;
	wire [1-1:0] node2303;
	wire [1-1:0] node2306;
	wire [1-1:0] node2309;
	wire [1-1:0] node2310;
	wire [1-1:0] node2314;
	wire [1-1:0] node2315;
	wire [1-1:0] node2316;
	wire [1-1:0] node2317;
	wire [1-1:0] node2320;
	wire [1-1:0] node2323;
	wire [1-1:0] node2324;
	wire [1-1:0] node2328;
	wire [1-1:0] node2329;
	wire [1-1:0] node2330;
	wire [1-1:0] node2335;
	wire [1-1:0] node2336;
	wire [1-1:0] node2337;
	wire [1-1:0] node2338;
	wire [1-1:0] node2339;
	wire [1-1:0] node2340;
	wire [1-1:0] node2343;
	wire [1-1:0] node2346;
	wire [1-1:0] node2347;
	wire [1-1:0] node2350;
	wire [1-1:0] node2353;
	wire [1-1:0] node2354;
	wire [1-1:0] node2355;
	wire [1-1:0] node2358;
	wire [1-1:0] node2361;
	wire [1-1:0] node2362;
	wire [1-1:0] node2366;
	wire [1-1:0] node2367;
	wire [1-1:0] node2368;
	wire [1-1:0] node2369;
	wire [1-1:0] node2372;
	wire [1-1:0] node2375;
	wire [1-1:0] node2376;
	wire [1-1:0] node2380;
	wire [1-1:0] node2381;
	wire [1-1:0] node2382;
	wire [1-1:0] node2387;
	wire [1-1:0] node2388;
	wire [1-1:0] node2389;
	wire [1-1:0] node2390;
	wire [1-1:0] node2391;
	wire [1-1:0] node2394;
	wire [1-1:0] node2397;
	wire [1-1:0] node2398;
	wire [1-1:0] node2402;
	wire [1-1:0] node2403;
	wire [1-1:0] node2404;
	wire [1-1:0] node2409;
	wire [1-1:0] node2410;
	wire [1-1:0] node2411;
	wire [1-1:0] node2412;
	wire [1-1:0] node2418;
	wire [1-1:0] node2419;
	wire [1-1:0] node2420;
	wire [1-1:0] node2421;
	wire [1-1:0] node2422;
	wire [1-1:0] node2423;
	wire [1-1:0] node2424;
	wire [1-1:0] node2426;
	wire [1-1:0] node2428;
	wire [1-1:0] node2431;
	wire [1-1:0] node2432;
	wire [1-1:0] node2434;
	wire [1-1:0] node2437;
	wire [1-1:0] node2438;
	wire [1-1:0] node2441;
	wire [1-1:0] node2444;
	wire [1-1:0] node2445;
	wire [1-1:0] node2446;
	wire [1-1:0] node2448;
	wire [1-1:0] node2451;
	wire [1-1:0] node2452;
	wire [1-1:0] node2455;
	wire [1-1:0] node2458;
	wire [1-1:0] node2459;
	wire [1-1:0] node2460;
	wire [1-1:0] node2463;
	wire [1-1:0] node2466;
	wire [1-1:0] node2467;
	wire [1-1:0] node2470;
	wire [1-1:0] node2473;
	wire [1-1:0] node2474;
	wire [1-1:0] node2475;
	wire [1-1:0] node2476;
	wire [1-1:0] node2478;
	wire [1-1:0] node2481;
	wire [1-1:0] node2482;
	wire [1-1:0] node2485;
	wire [1-1:0] node2488;
	wire [1-1:0] node2489;
	wire [1-1:0] node2490;
	wire [1-1:0] node2493;
	wire [1-1:0] node2496;
	wire [1-1:0] node2497;
	wire [1-1:0] node2500;
	wire [1-1:0] node2503;
	wire [1-1:0] node2504;
	wire [1-1:0] node2505;
	wire [1-1:0] node2506;
	wire [1-1:0] node2509;
	wire [1-1:0] node2512;
	wire [1-1:0] node2513;
	wire [1-1:0] node2516;
	wire [1-1:0] node2519;
	wire [1-1:0] node2520;
	wire [1-1:0] node2521;
	wire [1-1:0] node2524;
	wire [1-1:0] node2527;
	wire [1-1:0] node2528;
	wire [1-1:0] node2532;
	wire [1-1:0] node2533;
	wire [1-1:0] node2534;
	wire [1-1:0] node2535;
	wire [1-1:0] node2536;
	wire [1-1:0] node2538;
	wire [1-1:0] node2541;
	wire [1-1:0] node2542;
	wire [1-1:0] node2545;
	wire [1-1:0] node2548;
	wire [1-1:0] node2549;
	wire [1-1:0] node2550;
	wire [1-1:0] node2553;
	wire [1-1:0] node2556;
	wire [1-1:0] node2557;
	wire [1-1:0] node2560;
	wire [1-1:0] node2563;
	wire [1-1:0] node2564;
	wire [1-1:0] node2565;
	wire [1-1:0] node2566;
	wire [1-1:0] node2569;
	wire [1-1:0] node2572;
	wire [1-1:0] node2573;
	wire [1-1:0] node2576;
	wire [1-1:0] node2579;
	wire [1-1:0] node2580;
	wire [1-1:0] node2581;
	wire [1-1:0] node2584;
	wire [1-1:0] node2587;
	wire [1-1:0] node2588;
	wire [1-1:0] node2592;
	wire [1-1:0] node2593;
	wire [1-1:0] node2594;
	wire [1-1:0] node2595;
	wire [1-1:0] node2596;
	wire [1-1:0] node2599;
	wire [1-1:0] node2602;
	wire [1-1:0] node2603;
	wire [1-1:0] node2606;
	wire [1-1:0] node2609;
	wire [1-1:0] node2610;
	wire [1-1:0] node2611;
	wire [1-1:0] node2614;
	wire [1-1:0] node2617;
	wire [1-1:0] node2618;
	wire [1-1:0] node2622;
	wire [1-1:0] node2623;
	wire [1-1:0] node2624;
	wire [1-1:0] node2625;
	wire [1-1:0] node2628;
	wire [1-1:0] node2631;
	wire [1-1:0] node2632;
	wire [1-1:0] node2636;
	wire [1-1:0] node2637;
	wire [1-1:0] node2638;
	wire [1-1:0] node2643;
	wire [1-1:0] node2644;
	wire [1-1:0] node2645;
	wire [1-1:0] node2646;
	wire [1-1:0] node2647;
	wire [1-1:0] node2648;
	wire [1-1:0] node2650;
	wire [1-1:0] node2653;
	wire [1-1:0] node2654;
	wire [1-1:0] node2657;
	wire [1-1:0] node2660;
	wire [1-1:0] node2661;
	wire [1-1:0] node2662;
	wire [1-1:0] node2665;
	wire [1-1:0] node2668;
	wire [1-1:0] node2669;
	wire [1-1:0] node2672;
	wire [1-1:0] node2675;
	wire [1-1:0] node2676;
	wire [1-1:0] node2677;
	wire [1-1:0] node2678;
	wire [1-1:0] node2681;
	wire [1-1:0] node2684;
	wire [1-1:0] node2685;
	wire [1-1:0] node2688;
	wire [1-1:0] node2691;
	wire [1-1:0] node2692;
	wire [1-1:0] node2693;
	wire [1-1:0] node2696;
	wire [1-1:0] node2699;
	wire [1-1:0] node2700;
	wire [1-1:0] node2704;
	wire [1-1:0] node2705;
	wire [1-1:0] node2706;
	wire [1-1:0] node2707;
	wire [1-1:0] node2708;
	wire [1-1:0] node2711;
	wire [1-1:0] node2714;
	wire [1-1:0] node2715;
	wire [1-1:0] node2718;
	wire [1-1:0] node2721;
	wire [1-1:0] node2722;
	wire [1-1:0] node2723;
	wire [1-1:0] node2726;
	wire [1-1:0] node2729;
	wire [1-1:0] node2730;
	wire [1-1:0] node2734;
	wire [1-1:0] node2735;
	wire [1-1:0] node2736;
	wire [1-1:0] node2737;
	wire [1-1:0] node2740;
	wire [1-1:0] node2743;
	wire [1-1:0] node2744;
	wire [1-1:0] node2748;
	wire [1-1:0] node2749;
	wire [1-1:0] node2750;
	wire [1-1:0] node2755;
	wire [1-1:0] node2756;
	wire [1-1:0] node2757;
	wire [1-1:0] node2758;
	wire [1-1:0] node2759;
	wire [1-1:0] node2760;
	wire [1-1:0] node2763;
	wire [1-1:0] node2766;
	wire [1-1:0] node2767;
	wire [1-1:0] node2770;
	wire [1-1:0] node2773;
	wire [1-1:0] node2774;
	wire [1-1:0] node2775;
	wire [1-1:0] node2778;
	wire [1-1:0] node2781;
	wire [1-1:0] node2782;
	wire [1-1:0] node2786;
	wire [1-1:0] node2787;
	wire [1-1:0] node2788;
	wire [1-1:0] node2789;
	wire [1-1:0] node2792;
	wire [1-1:0] node2795;
	wire [1-1:0] node2796;
	wire [1-1:0] node2800;
	wire [1-1:0] node2801;
	wire [1-1:0] node2802;
	wire [1-1:0] node2807;
	wire [1-1:0] node2808;
	wire [1-1:0] node2809;
	wire [1-1:0] node2810;
	wire [1-1:0] node2811;
	wire [1-1:0] node2814;
	wire [1-1:0] node2817;
	wire [1-1:0] node2818;
	wire [1-1:0] node2822;
	wire [1-1:0] node2823;
	wire [1-1:0] node2824;
	wire [1-1:0] node2829;
	wire [1-1:0] node2830;
	wire [1-1:0] node2831;
	wire [1-1:0] node2832;
	wire [1-1:0] node2838;
	wire [1-1:0] node2839;
	wire [1-1:0] node2840;
	wire [1-1:0] node2841;
	wire [1-1:0] node2842;
	wire [1-1:0] node2843;
	wire [1-1:0] node2844;
	wire [1-1:0] node2846;
	wire [1-1:0] node2849;
	wire [1-1:0] node2850;
	wire [1-1:0] node2853;
	wire [1-1:0] node2856;
	wire [1-1:0] node2857;
	wire [1-1:0] node2858;
	wire [1-1:0] node2861;
	wire [1-1:0] node2864;
	wire [1-1:0] node2865;
	wire [1-1:0] node2868;
	wire [1-1:0] node2871;
	wire [1-1:0] node2872;
	wire [1-1:0] node2873;
	wire [1-1:0] node2874;
	wire [1-1:0] node2877;
	wire [1-1:0] node2880;
	wire [1-1:0] node2881;
	wire [1-1:0] node2884;
	wire [1-1:0] node2887;
	wire [1-1:0] node2888;
	wire [1-1:0] node2889;
	wire [1-1:0] node2892;
	wire [1-1:0] node2895;
	wire [1-1:0] node2896;
	wire [1-1:0] node2900;
	wire [1-1:0] node2901;
	wire [1-1:0] node2902;
	wire [1-1:0] node2903;
	wire [1-1:0] node2904;
	wire [1-1:0] node2907;
	wire [1-1:0] node2910;
	wire [1-1:0] node2911;
	wire [1-1:0] node2914;
	wire [1-1:0] node2917;
	wire [1-1:0] node2918;
	wire [1-1:0] node2919;
	wire [1-1:0] node2922;
	wire [1-1:0] node2925;
	wire [1-1:0] node2926;
	wire [1-1:0] node2930;
	wire [1-1:0] node2931;
	wire [1-1:0] node2932;
	wire [1-1:0] node2933;
	wire [1-1:0] node2936;
	wire [1-1:0] node2939;
	wire [1-1:0] node2940;
	wire [1-1:0] node2944;
	wire [1-1:0] node2945;
	wire [1-1:0] node2946;
	wire [1-1:0] node2951;
	wire [1-1:0] node2952;
	wire [1-1:0] node2953;
	wire [1-1:0] node2954;
	wire [1-1:0] node2955;
	wire [1-1:0] node2956;
	wire [1-1:0] node2959;
	wire [1-1:0] node2962;
	wire [1-1:0] node2963;
	wire [1-1:0] node2966;
	wire [1-1:0] node2969;
	wire [1-1:0] node2970;
	wire [1-1:0] node2971;
	wire [1-1:0] node2974;
	wire [1-1:0] node2977;
	wire [1-1:0] node2978;
	wire [1-1:0] node2982;
	wire [1-1:0] node2983;
	wire [1-1:0] node2984;
	wire [1-1:0] node2985;
	wire [1-1:0] node2988;
	wire [1-1:0] node2991;
	wire [1-1:0] node2992;
	wire [1-1:0] node2996;
	wire [1-1:0] node2997;
	wire [1-1:0] node2998;
	wire [1-1:0] node3003;
	wire [1-1:0] node3004;
	wire [1-1:0] node3005;
	wire [1-1:0] node3006;
	wire [1-1:0] node3007;
	wire [1-1:0] node3010;
	wire [1-1:0] node3013;
	wire [1-1:0] node3014;
	wire [1-1:0] node3018;
	wire [1-1:0] node3019;
	wire [1-1:0] node3020;
	wire [1-1:0] node3025;
	wire [1-1:0] node3026;
	wire [1-1:0] node3027;
	wire [1-1:0] node3028;
	wire [1-1:0] node3034;
	wire [1-1:0] node3035;
	wire [1-1:0] node3036;
	wire [1-1:0] node3037;
	wire [1-1:0] node3038;
	wire [1-1:0] node3039;
	wire [1-1:0] node3040;
	wire [1-1:0] node3043;
	wire [1-1:0] node3046;
	wire [1-1:0] node3047;
	wire [1-1:0] node3050;
	wire [1-1:0] node3053;
	wire [1-1:0] node3054;
	wire [1-1:0] node3055;
	wire [1-1:0] node3058;
	wire [1-1:0] node3061;
	wire [1-1:0] node3062;
	wire [1-1:0] node3066;
	wire [1-1:0] node3067;
	wire [1-1:0] node3068;
	wire [1-1:0] node3069;
	wire [1-1:0] node3072;
	wire [1-1:0] node3075;
	wire [1-1:0] node3076;
	wire [1-1:0] node3080;
	wire [1-1:0] node3081;
	wire [1-1:0] node3082;
	wire [1-1:0] node3087;
	wire [1-1:0] node3088;
	wire [1-1:0] node3089;
	wire [1-1:0] node3090;
	wire [1-1:0] node3091;
	wire [1-1:0] node3094;
	wire [1-1:0] node3097;
	wire [1-1:0] node3098;
	wire [1-1:0] node3102;
	wire [1-1:0] node3103;
	wire [1-1:0] node3104;
	wire [1-1:0] node3109;
	wire [1-1:0] node3110;
	wire [1-1:0] node3111;
	wire [1-1:0] node3112;
	wire [1-1:0] node3118;
	wire [1-1:0] node3119;
	wire [1-1:0] node3120;
	wire [1-1:0] node3121;
	wire [1-1:0] node3122;
	wire [1-1:0] node3123;
	wire [1-1:0] node3126;
	wire [1-1:0] node3129;
	wire [1-1:0] node3130;
	wire [1-1:0] node3134;
	wire [1-1:0] node3135;
	wire [1-1:0] node3136;
	wire [1-1:0] node3141;
	wire [1-1:0] node3142;
	wire [1-1:0] node3143;
	wire [1-1:0] node3144;
	wire [1-1:0] node3150;
	wire [1-1:0] node3151;
	wire [1-1:0] node3152;
	wire [1-1:0] node3153;
	wire [1-1:0] node3154;

	assign outp = (inp[13]) ? node1580 : node1;
		assign node1 = (inp[9]) ? node745 : node2;
			assign node2 = (inp[6]) ? node326 : node3;
				assign node3 = (inp[10]) ? node131 : node4;
					assign node4 = (inp[0]) ? node48 : node5;
						assign node5 = (inp[7]) ? node17 : node6;
							assign node6 = (inp[8]) ? node8 : 1'b1;
								assign node8 = (inp[4]) ? node10 : 1'b1;
									assign node10 = (inp[5]) ? node12 : 1'b1;
										assign node12 = (inp[14]) ? node14 : 1'b1;
											assign node14 = (inp[12]) ? 1'b1 : 1'b1;
							assign node17 = (inp[2]) ? node27 : node18;
								assign node18 = (inp[1]) ? node20 : 1'b1;
									assign node20 = (inp[4]) ? node22 : 1'b1;
										assign node22 = (inp[3]) ? node24 : 1'b1;
											assign node24 = (inp[5]) ? 1'b1 : 1'b1;
								assign node27 = (inp[5]) ? node35 : node28;
									assign node28 = (inp[14]) ? node30 : 1'b1;
										assign node30 = (inp[12]) ? node32 : 1'b1;
											assign node32 = (inp[1]) ? 1'b1 : 1'b1;
									assign node35 = (inp[3]) ? node41 : node36;
										assign node36 = (inp[8]) ? node38 : 1'b1;
											assign node38 = (inp[4]) ? 1'b1 : 1'b1;
										assign node41 = (inp[12]) ? node45 : node42;
											assign node42 = (inp[4]) ? 1'b1 : 1'b1;
											assign node45 = (inp[14]) ? 1'b0 : 1'b1;
						assign node48 = (inp[14]) ? node80 : node49;
							assign node49 = (inp[3]) ? node59 : node50;
								assign node50 = (inp[8]) ? node52 : 1'b1;
									assign node52 = (inp[11]) ? node54 : 1'b1;
										assign node54 = (inp[1]) ? node56 : 1'b1;
											assign node56 = (inp[5]) ? 1'b1 : 1'b1;
								assign node59 = (inp[12]) ? node67 : node60;
									assign node60 = (inp[2]) ? node62 : 1'b1;
										assign node62 = (inp[5]) ? node64 : 1'b1;
											assign node64 = (inp[11]) ? 1'b1 : 1'b1;
									assign node67 = (inp[11]) ? node73 : node68;
										assign node68 = (inp[4]) ? node70 : 1'b1;
											assign node70 = (inp[5]) ? 1'b1 : 1'b1;
										assign node73 = (inp[7]) ? node77 : node74;
											assign node74 = (inp[4]) ? 1'b1 : 1'b1;
											assign node77 = (inp[1]) ? 1'b0 : 1'b1;
							assign node80 = (inp[2]) ? node102 : node81;
								assign node81 = (inp[1]) ? node89 : node82;
									assign node82 = (inp[4]) ? node84 : 1'b1;
										assign node84 = (inp[11]) ? node86 : 1'b1;
											assign node86 = (inp[3]) ? 1'b1 : 1'b1;
									assign node89 = (inp[7]) ? node95 : node90;
										assign node90 = (inp[8]) ? node92 : 1'b1;
											assign node92 = (inp[11]) ? 1'b1 : 1'b1;
										assign node95 = (inp[3]) ? node99 : node96;
											assign node96 = (inp[8]) ? 1'b1 : 1'b1;
											assign node99 = (inp[12]) ? 1'b0 : 1'b1;
								assign node102 = (inp[5]) ? node116 : node103;
									assign node103 = (inp[3]) ? node109 : node104;
										assign node104 = (inp[8]) ? node106 : 1'b1;
											assign node106 = (inp[7]) ? 1'b1 : 1'b1;
										assign node109 = (inp[11]) ? node113 : node110;
											assign node110 = (inp[1]) ? 1'b1 : 1'b1;
											assign node113 = (inp[4]) ? 1'b0 : 1'b1;
									assign node116 = (inp[4]) ? node124 : node117;
										assign node117 = (inp[12]) ? node121 : node118;
											assign node118 = (inp[8]) ? 1'b1 : 1'b1;
											assign node121 = (inp[8]) ? 1'b0 : 1'b1;
										assign node124 = (inp[11]) ? node128 : node125;
											assign node125 = (inp[1]) ? 1'b0 : 1'b1;
											assign node128 = (inp[3]) ? 1'b0 : 1'b0;
					assign node131 = (inp[4]) ? node215 : node132;
						assign node132 = (inp[11]) ? node164 : node133;
							assign node133 = (inp[2]) ? node143 : node134;
								assign node134 = (inp[1]) ? node136 : 1'b1;
									assign node136 = (inp[7]) ? node138 : 1'b1;
										assign node138 = (inp[8]) ? node140 : 1'b1;
											assign node140 = (inp[0]) ? 1'b1 : 1'b1;
								assign node143 = (inp[8]) ? node151 : node144;
									assign node144 = (inp[12]) ? node146 : 1'b1;
										assign node146 = (inp[1]) ? node148 : 1'b1;
											assign node148 = (inp[7]) ? 1'b1 : 1'b1;
									assign node151 = (inp[0]) ? node157 : node152;
										assign node152 = (inp[7]) ? node154 : 1'b1;
											assign node154 = (inp[5]) ? 1'b1 : 1'b1;
										assign node157 = (inp[14]) ? node161 : node158;
											assign node158 = (inp[3]) ? 1'b1 : 1'b1;
											assign node161 = (inp[5]) ? 1'b0 : 1'b1;
							assign node164 = (inp[12]) ? node186 : node165;
								assign node165 = (inp[8]) ? node173 : node166;
									assign node166 = (inp[1]) ? node168 : 1'b1;
										assign node168 = (inp[5]) ? node170 : 1'b1;
											assign node170 = (inp[14]) ? 1'b1 : 1'b1;
									assign node173 = (inp[2]) ? node179 : node174;
										assign node174 = (inp[7]) ? node176 : 1'b1;
											assign node176 = (inp[1]) ? 1'b1 : 1'b1;
										assign node179 = (inp[7]) ? node183 : node180;
											assign node180 = (inp[3]) ? 1'b1 : 1'b1;
											assign node183 = (inp[0]) ? 1'b0 : 1'b1;
								assign node186 = (inp[5]) ? node200 : node187;
									assign node187 = (inp[3]) ? node193 : node188;
										assign node188 = (inp[1]) ? node190 : 1'b1;
											assign node190 = (inp[0]) ? 1'b1 : 1'b1;
										assign node193 = (inp[0]) ? node197 : node194;
											assign node194 = (inp[7]) ? 1'b1 : 1'b1;
											assign node197 = (inp[8]) ? 1'b0 : 1'b1;
									assign node200 = (inp[0]) ? node208 : node201;
										assign node201 = (inp[7]) ? node205 : node202;
											assign node202 = (inp[2]) ? 1'b1 : 1'b1;
											assign node205 = (inp[2]) ? 1'b0 : 1'b1;
										assign node208 = (inp[1]) ? node212 : node209;
											assign node209 = (inp[3]) ? 1'b0 : 1'b1;
											assign node212 = (inp[7]) ? 1'b0 : 1'b0;
						assign node215 = (inp[14]) ? node267 : node216;
							assign node216 = (inp[8]) ? node238 : node217;
								assign node217 = (inp[5]) ? node225 : node218;
									assign node218 = (inp[11]) ? node220 : 1'b1;
										assign node220 = (inp[12]) ? node222 : 1'b1;
											assign node222 = (inp[2]) ? 1'b1 : 1'b1;
									assign node225 = (inp[3]) ? node231 : node226;
										assign node226 = (inp[11]) ? node228 : 1'b1;
											assign node228 = (inp[7]) ? 1'b1 : 1'b1;
										assign node231 = (inp[0]) ? node235 : node232;
											assign node232 = (inp[1]) ? 1'b1 : 1'b1;
											assign node235 = (inp[11]) ? 1'b0 : 1'b1;
								assign node238 = (inp[1]) ? node252 : node239;
									assign node239 = (inp[12]) ? node245 : node240;
										assign node240 = (inp[7]) ? node242 : 1'b1;
											assign node242 = (inp[5]) ? 1'b1 : 1'b1;
										assign node245 = (inp[2]) ? node249 : node246;
											assign node246 = (inp[5]) ? 1'b1 : 1'b1;
											assign node249 = (inp[7]) ? 1'b0 : 1'b1;
									assign node252 = (inp[3]) ? node260 : node253;
										assign node253 = (inp[2]) ? node257 : node254;
											assign node254 = (inp[7]) ? 1'b1 : 1'b1;
											assign node257 = (inp[5]) ? 1'b0 : 1'b1;
										assign node260 = (inp[2]) ? node264 : node261;
											assign node261 = (inp[11]) ? 1'b0 : 1'b1;
											assign node264 = (inp[5]) ? 1'b0 : 1'b0;
							assign node267 = (inp[1]) ? node297 : node268;
								assign node268 = (inp[7]) ? node282 : node269;
									assign node269 = (inp[8]) ? node275 : node270;
										assign node270 = (inp[11]) ? node272 : 1'b1;
											assign node272 = (inp[5]) ? 1'b1 : 1'b1;
										assign node275 = (inp[2]) ? node279 : node276;
											assign node276 = (inp[5]) ? 1'b1 : 1'b1;
											assign node279 = (inp[5]) ? 1'b0 : 1'b1;
									assign node282 = (inp[11]) ? node290 : node283;
										assign node283 = (inp[5]) ? node287 : node284;
											assign node284 = (inp[8]) ? 1'b1 : 1'b1;
											assign node287 = (inp[2]) ? 1'b0 : 1'b1;
										assign node290 = (inp[5]) ? node294 : node291;
											assign node291 = (inp[8]) ? 1'b0 : 1'b1;
											assign node294 = (inp[12]) ? 1'b0 : 1'b0;
								assign node297 = (inp[0]) ? node313 : node298;
									assign node298 = (inp[5]) ? node306 : node299;
										assign node299 = (inp[8]) ? node303 : node300;
											assign node300 = (inp[12]) ? 1'b1 : 1'b1;
											assign node303 = (inp[3]) ? 1'b0 : 1'b1;
										assign node306 = (inp[2]) ? node310 : node307;
											assign node307 = (inp[3]) ? 1'b0 : 1'b1;
											assign node310 = (inp[11]) ? 1'b0 : 1'b0;
									assign node313 = (inp[2]) ? node321 : node314;
										assign node314 = (inp[8]) ? node318 : node315;
											assign node315 = (inp[12]) ? 1'b0 : 1'b1;
											assign node318 = (inp[7]) ? 1'b0 : 1'b0;
										assign node321 = (inp[7]) ? 1'b0 : node322;
											assign node322 = (inp[5]) ? 1'b0 : 1'b0;
				assign node326 = (inp[7]) ? node522 : node327;
					assign node327 = (inp[12]) ? node411 : node328;
						assign node328 = (inp[0]) ? node360 : node329;
							assign node329 = (inp[8]) ? node339 : node330;
								assign node330 = (inp[10]) ? node332 : 1'b1;
									assign node332 = (inp[14]) ? node334 : 1'b1;
										assign node334 = (inp[2]) ? node336 : 1'b1;
											assign node336 = (inp[4]) ? 1'b1 : 1'b1;
								assign node339 = (inp[14]) ? node347 : node340;
									assign node340 = (inp[3]) ? node342 : 1'b1;
										assign node342 = (inp[5]) ? node344 : 1'b1;
											assign node344 = (inp[10]) ? 1'b0 : 1'b1;
									assign node347 = (inp[10]) ? node353 : node348;
										assign node348 = (inp[5]) ? node350 : 1'b1;
											assign node350 = (inp[3]) ? 1'b1 : 1'b1;
										assign node353 = (inp[11]) ? node357 : node354;
											assign node354 = (inp[5]) ? 1'b1 : 1'b1;
											assign node357 = (inp[1]) ? 1'b0 : 1'b1;
							assign node360 = (inp[4]) ? node382 : node361;
								assign node361 = (inp[10]) ? node369 : node362;
									assign node362 = (inp[2]) ? node364 : 1'b1;
										assign node364 = (inp[11]) ? node366 : 1'b1;
											assign node366 = (inp[14]) ? 1'b1 : 1'b1;
									assign node369 = (inp[3]) ? node375 : node370;
										assign node370 = (inp[11]) ? node372 : 1'b1;
											assign node372 = (inp[8]) ? 1'b1 : 1'b1;
										assign node375 = (inp[2]) ? node379 : node376;
											assign node376 = (inp[11]) ? 1'b1 : 1'b1;
											assign node379 = (inp[11]) ? 1'b0 : 1'b1;
								assign node382 = (inp[8]) ? node396 : node383;
									assign node383 = (inp[1]) ? node389 : node384;
										assign node384 = (inp[2]) ? node386 : 1'b1;
											assign node386 = (inp[3]) ? 1'b1 : 1'b1;
										assign node389 = (inp[14]) ? node393 : node390;
											assign node390 = (inp[11]) ? 1'b1 : 1'b1;
											assign node393 = (inp[2]) ? 1'b0 : 1'b1;
									assign node396 = (inp[5]) ? node404 : node397;
										assign node397 = (inp[10]) ? node401 : node398;
											assign node398 = (inp[11]) ? 1'b1 : 1'b1;
											assign node401 = (inp[14]) ? 1'b0 : 1'b1;
										assign node404 = (inp[11]) ? node408 : node405;
											assign node405 = (inp[2]) ? 1'b0 : 1'b1;
											assign node408 = (inp[14]) ? 1'b0 : 1'b0;
						assign node411 = (inp[14]) ? node463 : node412;
							assign node412 = (inp[2]) ? node434 : node413;
								assign node413 = (inp[0]) ? node421 : node414;
									assign node414 = (inp[3]) ? node416 : 1'b1;
										assign node416 = (inp[10]) ? node418 : 1'b1;
											assign node418 = (inp[11]) ? 1'b1 : 1'b1;
									assign node421 = (inp[8]) ? node427 : node422;
										assign node422 = (inp[11]) ? node424 : 1'b1;
											assign node424 = (inp[4]) ? 1'b1 : 1'b1;
										assign node427 = (inp[1]) ? node431 : node428;
											assign node428 = (inp[10]) ? 1'b1 : 1'b1;
											assign node431 = (inp[3]) ? 1'b0 : 1'b1;
								assign node434 = (inp[8]) ? node448 : node435;
									assign node435 = (inp[0]) ? node441 : node436;
										assign node436 = (inp[10]) ? node438 : 1'b1;
											assign node438 = (inp[1]) ? 1'b1 : 1'b1;
										assign node441 = (inp[4]) ? node445 : node442;
											assign node442 = (inp[5]) ? 1'b1 : 1'b1;
											assign node445 = (inp[3]) ? 1'b0 : 1'b1;
									assign node448 = (inp[1]) ? node456 : node449;
										assign node449 = (inp[11]) ? node453 : node450;
											assign node450 = (inp[10]) ? 1'b1 : 1'b1;
											assign node453 = (inp[10]) ? 1'b0 : 1'b1;
										assign node456 = (inp[4]) ? node460 : node457;
											assign node457 = (inp[10]) ? 1'b0 : 1'b1;
											assign node460 = (inp[0]) ? 1'b0 : 1'b0;
							assign node463 = (inp[11]) ? node493 : node464;
								assign node464 = (inp[8]) ? node478 : node465;
									assign node465 = (inp[3]) ? node471 : node466;
										assign node466 = (inp[5]) ? node468 : 1'b1;
											assign node468 = (inp[10]) ? 1'b1 : 1'b1;
										assign node471 = (inp[10]) ? node475 : node472;
											assign node472 = (inp[1]) ? 1'b1 : 1'b1;
											assign node475 = (inp[2]) ? 1'b0 : 1'b1;
									assign node478 = (inp[0]) ? node486 : node479;
										assign node479 = (inp[4]) ? node483 : node480;
											assign node480 = (inp[3]) ? 1'b1 : 1'b1;
											assign node483 = (inp[5]) ? 1'b0 : 1'b1;
										assign node486 = (inp[5]) ? node490 : node487;
											assign node487 = (inp[10]) ? 1'b0 : 1'b1;
											assign node490 = (inp[1]) ? 1'b0 : 1'b0;
								assign node493 = (inp[0]) ? node509 : node494;
									assign node494 = (inp[10]) ? node502 : node495;
										assign node495 = (inp[5]) ? node499 : node496;
											assign node496 = (inp[2]) ? 1'b1 : 1'b1;
											assign node499 = (inp[2]) ? 1'b0 : 1'b1;
										assign node502 = (inp[2]) ? node506 : node503;
											assign node503 = (inp[1]) ? 1'b0 : 1'b1;
											assign node506 = (inp[8]) ? 1'b0 : 1'b0;
									assign node509 = (inp[3]) ? node517 : node510;
										assign node510 = (inp[2]) ? node514 : node511;
											assign node511 = (inp[8]) ? 1'b0 : 1'b1;
											assign node514 = (inp[4]) ? 1'b0 : 1'b0;
										assign node517 = (inp[1]) ? 1'b0 : node518;
											assign node518 = (inp[8]) ? 1'b0 : 1'b0;
					assign node522 = (inp[4]) ? node634 : node523;
						assign node523 = (inp[2]) ? node575 : node524;
							assign node524 = (inp[0]) ? node546 : node525;
								assign node525 = (inp[5]) ? node533 : node526;
									assign node526 = (inp[12]) ? node528 : 1'b1;
										assign node528 = (inp[11]) ? node530 : 1'b1;
											assign node530 = (inp[14]) ? 1'b1 : 1'b1;
									assign node533 = (inp[14]) ? node539 : node534;
										assign node534 = (inp[8]) ? node536 : 1'b1;
											assign node536 = (inp[10]) ? 1'b1 : 1'b1;
										assign node539 = (inp[3]) ? node543 : node540;
											assign node540 = (inp[8]) ? 1'b1 : 1'b1;
											assign node543 = (inp[10]) ? 1'b0 : 1'b1;
								assign node546 = (inp[3]) ? node560 : node547;
									assign node547 = (inp[8]) ? node553 : node548;
										assign node548 = (inp[10]) ? node550 : 1'b1;
											assign node550 = (inp[1]) ? 1'b1 : 1'b1;
										assign node553 = (inp[1]) ? node557 : node554;
											assign node554 = (inp[14]) ? 1'b1 : 1'b1;
											assign node557 = (inp[12]) ? 1'b0 : 1'b1;
									assign node560 = (inp[11]) ? node568 : node561;
										assign node561 = (inp[10]) ? node565 : node562;
											assign node562 = (inp[12]) ? 1'b1 : 1'b1;
											assign node565 = (inp[5]) ? 1'b0 : 1'b1;
										assign node568 = (inp[14]) ? node572 : node569;
											assign node569 = (inp[12]) ? 1'b0 : 1'b1;
											assign node572 = (inp[8]) ? 1'b0 : 1'b0;
							assign node575 = (inp[1]) ? node605 : node576;
								assign node576 = (inp[10]) ? node590 : node577;
									assign node577 = (inp[8]) ? node583 : node578;
										assign node578 = (inp[12]) ? node580 : 1'b1;
											assign node580 = (inp[14]) ? 1'b1 : 1'b1;
										assign node583 = (inp[5]) ? node587 : node584;
											assign node584 = (inp[3]) ? 1'b1 : 1'b1;
											assign node587 = (inp[11]) ? 1'b0 : 1'b1;
									assign node590 = (inp[3]) ? node598 : node591;
										assign node591 = (inp[0]) ? node595 : node592;
											assign node592 = (inp[5]) ? 1'b1 : 1'b1;
											assign node595 = (inp[8]) ? 1'b0 : 1'b1;
										assign node598 = (inp[0]) ? node602 : node599;
											assign node599 = (inp[14]) ? 1'b0 : 1'b1;
											assign node602 = (inp[11]) ? 1'b0 : 1'b0;
								assign node605 = (inp[5]) ? node621 : node606;
									assign node606 = (inp[8]) ? node614 : node607;
										assign node607 = (inp[14]) ? node611 : node608;
											assign node608 = (inp[0]) ? 1'b1 : 1'b1;
											assign node611 = (inp[12]) ? 1'b0 : 1'b1;
										assign node614 = (inp[10]) ? node618 : node615;
											assign node615 = (inp[0]) ? 1'b0 : 1'b1;
											assign node618 = (inp[11]) ? 1'b0 : 1'b0;
									assign node621 = (inp[0]) ? node629 : node622;
										assign node622 = (inp[11]) ? node626 : node623;
											assign node623 = (inp[10]) ? 1'b0 : 1'b1;
											assign node626 = (inp[10]) ? 1'b0 : 1'b0;
										assign node629 = (inp[8]) ? 1'b0 : node630;
											assign node630 = (inp[14]) ? 1'b0 : 1'b0;
						assign node634 = (inp[14]) ? node694 : node635;
							assign node635 = (inp[1]) ? node665 : node636;
								assign node636 = (inp[10]) ? node650 : node637;
									assign node637 = (inp[11]) ? node643 : node638;
										assign node638 = (inp[3]) ? node640 : 1'b1;
											assign node640 = (inp[0]) ? 1'b1 : 1'b1;
										assign node643 = (inp[12]) ? node647 : node644;
											assign node644 = (inp[5]) ? 1'b1 : 1'b1;
											assign node647 = (inp[2]) ? 1'b0 : 1'b1;
									assign node650 = (inp[0]) ? node658 : node651;
										assign node651 = (inp[5]) ? node655 : node652;
											assign node652 = (inp[2]) ? 1'b1 : 1'b1;
											assign node655 = (inp[8]) ? 1'b0 : 1'b1;
										assign node658 = (inp[12]) ? node662 : node659;
											assign node659 = (inp[11]) ? 1'b0 : 1'b1;
											assign node662 = (inp[5]) ? 1'b0 : 1'b0;
								assign node665 = (inp[0]) ? node681 : node666;
									assign node666 = (inp[2]) ? node674 : node667;
										assign node667 = (inp[12]) ? node671 : node668;
											assign node668 = (inp[8]) ? 1'b1 : 1'b1;
											assign node671 = (inp[3]) ? 1'b0 : 1'b1;
										assign node674 = (inp[3]) ? node678 : node675;
											assign node675 = (inp[8]) ? 1'b0 : 1'b1;
											assign node678 = (inp[10]) ? 1'b0 : 1'b0;
									assign node681 = (inp[8]) ? node689 : node682;
										assign node682 = (inp[2]) ? node686 : node683;
											assign node683 = (inp[3]) ? 1'b0 : 1'b1;
											assign node686 = (inp[5]) ? 1'b0 : 1'b0;
										assign node689 = (inp[11]) ? 1'b0 : node690;
											assign node690 = (inp[12]) ? 1'b0 : 1'b0;
							assign node694 = (inp[5]) ? node724 : node695;
								assign node695 = (inp[3]) ? node711 : node696;
									assign node696 = (inp[12]) ? node704 : node697;
										assign node697 = (inp[2]) ? node701 : node698;
											assign node698 = (inp[10]) ? 1'b1 : 1'b1;
											assign node701 = (inp[11]) ? 1'b0 : 1'b1;
										assign node704 = (inp[8]) ? node708 : node705;
											assign node705 = (inp[11]) ? 1'b0 : 1'b1;
											assign node708 = (inp[1]) ? 1'b0 : 1'b0;
									assign node711 = (inp[8]) ? node719 : node712;
										assign node712 = (inp[12]) ? node716 : node713;
											assign node713 = (inp[10]) ? 1'b0 : 1'b1;
											assign node716 = (inp[2]) ? 1'b0 : 1'b0;
										assign node719 = (inp[1]) ? 1'b0 : node720;
											assign node720 = (inp[2]) ? 1'b0 : 1'b0;
								assign node724 = (inp[1]) ? node738 : node725;
									assign node725 = (inp[8]) ? node733 : node726;
										assign node726 = (inp[11]) ? node730 : node727;
											assign node727 = (inp[10]) ? 1'b0 : 1'b1;
											assign node730 = (inp[12]) ? 1'b0 : 1'b0;
										assign node733 = (inp[12]) ? 1'b0 : node734;
											assign node734 = (inp[3]) ? 1'b0 : 1'b0;
									assign node738 = (inp[2]) ? 1'b0 : node739;
										assign node739 = (inp[0]) ? 1'b0 : node740;
											assign node740 = (inp[11]) ? 1'b0 : 1'b0;
			assign node745 = (inp[3]) ? node1165 : node746;
				assign node746 = (inp[4]) ? node942 : node747;
					assign node747 = (inp[11]) ? node831 : node748;
						assign node748 = (inp[10]) ? node780 : node749;
							assign node749 = (inp[5]) ? node759 : node750;
								assign node750 = (inp[14]) ? node752 : 1'b1;
									assign node752 = (inp[8]) ? node754 : 1'b1;
										assign node754 = (inp[2]) ? node756 : 1'b1;
											assign node756 = (inp[7]) ? 1'b1 : 1'b1;
								assign node759 = (inp[7]) ? node767 : node760;
									assign node760 = (inp[12]) ? node762 : 1'b1;
										assign node762 = (inp[2]) ? node764 : 1'b1;
											assign node764 = (inp[6]) ? 1'b1 : 1'b1;
									assign node767 = (inp[14]) ? node773 : node768;
										assign node768 = (inp[2]) ? node770 : 1'b1;
											assign node770 = (inp[8]) ? 1'b1 : 1'b1;
										assign node773 = (inp[0]) ? node777 : node774;
											assign node774 = (inp[2]) ? 1'b1 : 1'b1;
											assign node777 = (inp[6]) ? 1'b0 : 1'b1;
							assign node780 = (inp[1]) ? node802 : node781;
								assign node781 = (inp[12]) ? node789 : node782;
									assign node782 = (inp[8]) ? node784 : 1'b1;
										assign node784 = (inp[0]) ? node786 : 1'b1;
											assign node786 = (inp[2]) ? 1'b1 : 1'b1;
									assign node789 = (inp[14]) ? node795 : node790;
										assign node790 = (inp[8]) ? node792 : 1'b1;
											assign node792 = (inp[5]) ? 1'b1 : 1'b1;
										assign node795 = (inp[7]) ? node799 : node796;
											assign node796 = (inp[8]) ? 1'b1 : 1'b1;
											assign node799 = (inp[6]) ? 1'b0 : 1'b1;
								assign node802 = (inp[7]) ? node816 : node803;
									assign node803 = (inp[5]) ? node809 : node804;
										assign node804 = (inp[8]) ? node806 : 1'b1;
											assign node806 = (inp[12]) ? 1'b1 : 1'b1;
										assign node809 = (inp[14]) ? node813 : node810;
											assign node810 = (inp[8]) ? 1'b1 : 1'b1;
											assign node813 = (inp[6]) ? 1'b0 : 1'b1;
									assign node816 = (inp[2]) ? node824 : node817;
										assign node817 = (inp[14]) ? node821 : node818;
											assign node818 = (inp[5]) ? 1'b1 : 1'b1;
											assign node821 = (inp[12]) ? 1'b0 : 1'b1;
										assign node824 = (inp[6]) ? node828 : node825;
											assign node825 = (inp[0]) ? 1'b0 : 1'b1;
											assign node828 = (inp[5]) ? 1'b0 : 1'b0;
						assign node831 = (inp[7]) ? node883 : node832;
							assign node832 = (inp[8]) ? node854 : node833;
								assign node833 = (inp[5]) ? node841 : node834;
									assign node834 = (inp[10]) ? node836 : 1'b1;
										assign node836 = (inp[12]) ? node838 : 1'b1;
											assign node838 = (inp[14]) ? 1'b0 : 1'b1;
									assign node841 = (inp[2]) ? node847 : node842;
										assign node842 = (inp[12]) ? node844 : 1'b1;
											assign node844 = (inp[6]) ? 1'b1 : 1'b1;
										assign node847 = (inp[1]) ? node851 : node848;
											assign node848 = (inp[14]) ? 1'b1 : 1'b1;
											assign node851 = (inp[12]) ? 1'b0 : 1'b1;
								assign node854 = (inp[14]) ? node868 : node855;
									assign node855 = (inp[6]) ? node861 : node856;
										assign node856 = (inp[2]) ? node858 : 1'b1;
											assign node858 = (inp[10]) ? 1'b1 : 1'b1;
										assign node861 = (inp[5]) ? node865 : node862;
											assign node862 = (inp[12]) ? 1'b1 : 1'b1;
											assign node865 = (inp[0]) ? 1'b0 : 1'b1;
									assign node868 = (inp[0]) ? node876 : node869;
										assign node869 = (inp[2]) ? node873 : node870;
											assign node870 = (inp[6]) ? 1'b1 : 1'b1;
											assign node873 = (inp[5]) ? 1'b0 : 1'b1;
										assign node876 = (inp[1]) ? node880 : node877;
											assign node877 = (inp[12]) ? 1'b0 : 1'b1;
											assign node880 = (inp[2]) ? 1'b0 : 1'b0;
							assign node883 = (inp[1]) ? node913 : node884;
								assign node884 = (inp[2]) ? node898 : node885;
									assign node885 = (inp[0]) ? node891 : node886;
										assign node886 = (inp[8]) ? node888 : 1'b1;
											assign node888 = (inp[10]) ? 1'b1 : 1'b1;
										assign node891 = (inp[8]) ? node895 : node892;
											assign node892 = (inp[14]) ? 1'b1 : 1'b1;
											assign node895 = (inp[12]) ? 1'b0 : 1'b1;
									assign node898 = (inp[5]) ? node906 : node899;
										assign node899 = (inp[10]) ? node903 : node900;
											assign node900 = (inp[8]) ? 1'b1 : 1'b1;
											assign node903 = (inp[0]) ? 1'b0 : 1'b1;
										assign node906 = (inp[12]) ? node910 : node907;
											assign node907 = (inp[0]) ? 1'b0 : 1'b1;
											assign node910 = (inp[14]) ? 1'b0 : 1'b0;
								assign node913 = (inp[5]) ? node929 : node914;
									assign node914 = (inp[0]) ? node922 : node915;
										assign node915 = (inp[10]) ? node919 : node916;
											assign node916 = (inp[2]) ? 1'b1 : 1'b1;
											assign node919 = (inp[8]) ? 1'b0 : 1'b1;
										assign node922 = (inp[8]) ? node926 : node923;
											assign node923 = (inp[14]) ? 1'b0 : 1'b1;
											assign node926 = (inp[6]) ? 1'b0 : 1'b0;
									assign node929 = (inp[2]) ? node937 : node930;
										assign node930 = (inp[12]) ? node934 : node931;
											assign node931 = (inp[8]) ? 1'b0 : 1'b1;
											assign node934 = (inp[14]) ? 1'b0 : 1'b0;
										assign node937 = (inp[6]) ? 1'b0 : node938;
											assign node938 = (inp[8]) ? 1'b0 : 1'b0;
					assign node942 = (inp[2]) ? node1054 : node943;
						assign node943 = (inp[5]) ? node995 : node944;
							assign node944 = (inp[8]) ? node966 : node945;
								assign node945 = (inp[10]) ? node953 : node946;
									assign node946 = (inp[0]) ? node948 : 1'b1;
										assign node948 = (inp[7]) ? node950 : 1'b1;
											assign node950 = (inp[6]) ? 1'b1 : 1'b1;
									assign node953 = (inp[1]) ? node959 : node954;
										assign node954 = (inp[12]) ? node956 : 1'b1;
											assign node956 = (inp[14]) ? 1'b1 : 1'b1;
										assign node959 = (inp[0]) ? node963 : node960;
											assign node960 = (inp[6]) ? 1'b1 : 1'b1;
											assign node963 = (inp[12]) ? 1'b0 : 1'b1;
								assign node966 = (inp[1]) ? node980 : node967;
									assign node967 = (inp[7]) ? node973 : node968;
										assign node968 = (inp[11]) ? node970 : 1'b1;
											assign node970 = (inp[0]) ? 1'b1 : 1'b1;
										assign node973 = (inp[12]) ? node977 : node974;
											assign node974 = (inp[11]) ? 1'b1 : 1'b1;
											assign node977 = (inp[0]) ? 1'b0 : 1'b1;
									assign node980 = (inp[14]) ? node988 : node981;
										assign node981 = (inp[10]) ? node985 : node982;
											assign node982 = (inp[0]) ? 1'b1 : 1'b1;
											assign node985 = (inp[6]) ? 1'b0 : 1'b1;
										assign node988 = (inp[0]) ? node992 : node989;
											assign node989 = (inp[12]) ? 1'b0 : 1'b1;
											assign node992 = (inp[11]) ? 1'b0 : 1'b0;
							assign node995 = (inp[6]) ? node1025 : node996;
								assign node996 = (inp[1]) ? node1010 : node997;
									assign node997 = (inp[14]) ? node1003 : node998;
										assign node998 = (inp[8]) ? node1000 : 1'b1;
											assign node1000 = (inp[12]) ? 1'b1 : 1'b1;
										assign node1003 = (inp[11]) ? node1007 : node1004;
											assign node1004 = (inp[12]) ? 1'b1 : 1'b1;
											assign node1007 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1010 = (inp[8]) ? node1018 : node1011;
										assign node1011 = (inp[10]) ? node1015 : node1012;
											assign node1012 = (inp[0]) ? 1'b1 : 1'b1;
											assign node1015 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1018 = (inp[12]) ? node1022 : node1019;
											assign node1019 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1022 = (inp[0]) ? 1'b0 : 1'b0;
								assign node1025 = (inp[0]) ? node1041 : node1026;
									assign node1026 = (inp[14]) ? node1034 : node1027;
										assign node1027 = (inp[10]) ? node1031 : node1028;
											assign node1028 = (inp[11]) ? 1'b1 : 1'b1;
											assign node1031 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1034 = (inp[12]) ? node1038 : node1035;
											assign node1035 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1038 = (inp[11]) ? 1'b0 : 1'b0;
									assign node1041 = (inp[8]) ? node1049 : node1042;
										assign node1042 = (inp[14]) ? node1046 : node1043;
											assign node1043 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1046 = (inp[10]) ? 1'b0 : 1'b0;
										assign node1049 = (inp[11]) ? 1'b0 : node1050;
											assign node1050 = (inp[7]) ? 1'b0 : 1'b0;
						assign node1054 = (inp[10]) ? node1114 : node1055;
							assign node1055 = (inp[6]) ? node1085 : node1056;
								assign node1056 = (inp[7]) ? node1070 : node1057;
									assign node1057 = (inp[12]) ? node1063 : node1058;
										assign node1058 = (inp[11]) ? node1060 : 1'b1;
											assign node1060 = (inp[14]) ? 1'b1 : 1'b1;
										assign node1063 = (inp[14]) ? node1067 : node1064;
											assign node1064 = (inp[1]) ? 1'b1 : 1'b1;
											assign node1067 = (inp[8]) ? 1'b0 : 1'b1;
									assign node1070 = (inp[0]) ? node1078 : node1071;
										assign node1071 = (inp[5]) ? node1075 : node1072;
											assign node1072 = (inp[12]) ? 1'b1 : 1'b1;
											assign node1075 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1078 = (inp[8]) ? node1082 : node1079;
											assign node1079 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1082 = (inp[14]) ? 1'b0 : 1'b0;
								assign node1085 = (inp[0]) ? node1101 : node1086;
									assign node1086 = (inp[1]) ? node1094 : node1087;
										assign node1087 = (inp[5]) ? node1091 : node1088;
											assign node1088 = (inp[8]) ? 1'b1 : 1'b1;
											assign node1091 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1094 = (inp[12]) ? node1098 : node1095;
											assign node1095 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1098 = (inp[11]) ? 1'b0 : 1'b0;
									assign node1101 = (inp[7]) ? node1109 : node1102;
										assign node1102 = (inp[8]) ? node1106 : node1103;
											assign node1103 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1106 = (inp[11]) ? 1'b0 : 1'b0;
										assign node1109 = (inp[1]) ? 1'b0 : node1110;
											assign node1110 = (inp[5]) ? 1'b0 : 1'b0;
							assign node1114 = (inp[14]) ? node1144 : node1115;
								assign node1115 = (inp[12]) ? node1131 : node1116;
									assign node1116 = (inp[1]) ? node1124 : node1117;
										assign node1117 = (inp[6]) ? node1121 : node1118;
											assign node1118 = (inp[11]) ? 1'b1 : 1'b1;
											assign node1121 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1124 = (inp[8]) ? node1128 : node1125;
											assign node1125 = (inp[0]) ? 1'b0 : 1'b1;
											assign node1128 = (inp[6]) ? 1'b0 : 1'b0;
									assign node1131 = (inp[0]) ? node1139 : node1132;
										assign node1132 = (inp[7]) ? node1136 : node1133;
											assign node1133 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1136 = (inp[8]) ? 1'b0 : 1'b0;
										assign node1139 = (inp[6]) ? 1'b0 : node1140;
											assign node1140 = (inp[8]) ? 1'b0 : 1'b0;
								assign node1144 = (inp[5]) ? node1158 : node1145;
									assign node1145 = (inp[12]) ? node1153 : node1146;
										assign node1146 = (inp[7]) ? node1150 : node1147;
											assign node1147 = (inp[0]) ? 1'b0 : 1'b1;
											assign node1150 = (inp[6]) ? 1'b0 : 1'b0;
										assign node1153 = (inp[1]) ? 1'b0 : node1154;
											assign node1154 = (inp[6]) ? 1'b0 : 1'b0;
									assign node1158 = (inp[7]) ? 1'b0 : node1159;
										assign node1159 = (inp[0]) ? 1'b0 : node1160;
											assign node1160 = (inp[6]) ? 1'b0 : 1'b0;
				assign node1165 = (inp[7]) ? node1389 : node1166;
					assign node1166 = (inp[1]) ? node1278 : node1167;
						assign node1167 = (inp[8]) ? node1219 : node1168;
							assign node1168 = (inp[14]) ? node1190 : node1169;
								assign node1169 = (inp[2]) ? node1177 : node1170;
									assign node1170 = (inp[12]) ? node1172 : 1'b1;
										assign node1172 = (inp[0]) ? node1174 : 1'b1;
											assign node1174 = (inp[4]) ? 1'b1 : 1'b1;
									assign node1177 = (inp[4]) ? node1183 : node1178;
										assign node1178 = (inp[11]) ? node1180 : 1'b1;
											assign node1180 = (inp[6]) ? 1'b1 : 1'b1;
										assign node1183 = (inp[5]) ? node1187 : node1184;
											assign node1184 = (inp[12]) ? 1'b1 : 1'b1;
											assign node1187 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1190 = (inp[11]) ? node1204 : node1191;
									assign node1191 = (inp[0]) ? node1197 : node1192;
										assign node1192 = (inp[12]) ? node1194 : 1'b1;
											assign node1194 = (inp[2]) ? 1'b1 : 1'b1;
										assign node1197 = (inp[6]) ? node1201 : node1198;
											assign node1198 = (inp[2]) ? 1'b1 : 1'b1;
											assign node1201 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1204 = (inp[5]) ? node1212 : node1205;
										assign node1205 = (inp[0]) ? node1209 : node1206;
											assign node1206 = (inp[4]) ? 1'b1 : 1'b1;
											assign node1209 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1212 = (inp[0]) ? node1216 : node1213;
											assign node1213 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1216 = (inp[10]) ? 1'b0 : 1'b0;
							assign node1219 = (inp[2]) ? node1249 : node1220;
								assign node1220 = (inp[11]) ? node1234 : node1221;
									assign node1221 = (inp[5]) ? node1227 : node1222;
										assign node1222 = (inp[4]) ? node1224 : 1'b1;
											assign node1224 = (inp[10]) ? 1'b1 : 1'b1;
										assign node1227 = (inp[0]) ? node1231 : node1228;
											assign node1228 = (inp[4]) ? 1'b1 : 1'b1;
											assign node1231 = (inp[12]) ? 1'b0 : 1'b1;
									assign node1234 = (inp[12]) ? node1242 : node1235;
										assign node1235 = (inp[6]) ? node1239 : node1236;
											assign node1236 = (inp[10]) ? 1'b1 : 1'b1;
											assign node1239 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1242 = (inp[6]) ? node1246 : node1243;
											assign node1243 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1246 = (inp[14]) ? 1'b0 : 1'b0;
								assign node1249 = (inp[5]) ? node1265 : node1250;
									assign node1250 = (inp[6]) ? node1258 : node1251;
										assign node1251 = (inp[4]) ? node1255 : node1252;
											assign node1252 = (inp[10]) ? 1'b1 : 1'b1;
											assign node1255 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1258 = (inp[0]) ? node1262 : node1259;
											assign node1259 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1262 = (inp[14]) ? 1'b0 : 1'b0;
									assign node1265 = (inp[0]) ? node1273 : node1266;
										assign node1266 = (inp[14]) ? node1270 : node1267;
											assign node1267 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1270 = (inp[10]) ? 1'b0 : 1'b0;
										assign node1273 = (inp[14]) ? 1'b0 : node1274;
											assign node1274 = (inp[10]) ? 1'b0 : 1'b0;
						assign node1278 = (inp[5]) ? node1338 : node1279;
							assign node1279 = (inp[0]) ? node1309 : node1280;
								assign node1280 = (inp[2]) ? node1294 : node1281;
									assign node1281 = (inp[4]) ? node1287 : node1282;
										assign node1282 = (inp[8]) ? node1284 : 1'b1;
											assign node1284 = (inp[10]) ? 1'b1 : 1'b1;
										assign node1287 = (inp[11]) ? node1291 : node1288;
											assign node1288 = (inp[6]) ? 1'b1 : 1'b1;
											assign node1291 = (inp[14]) ? 1'b0 : 1'b1;
									assign node1294 = (inp[12]) ? node1302 : node1295;
										assign node1295 = (inp[14]) ? node1299 : node1296;
											assign node1296 = (inp[8]) ? 1'b1 : 1'b1;
											assign node1299 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1302 = (inp[6]) ? node1306 : node1303;
											assign node1303 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1306 = (inp[4]) ? 1'b0 : 1'b0;
								assign node1309 = (inp[14]) ? node1325 : node1310;
									assign node1310 = (inp[11]) ? node1318 : node1311;
										assign node1311 = (inp[12]) ? node1315 : node1312;
											assign node1312 = (inp[8]) ? 1'b1 : 1'b1;
											assign node1315 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1318 = (inp[2]) ? node1322 : node1319;
											assign node1319 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1322 = (inp[4]) ? 1'b0 : 1'b0;
									assign node1325 = (inp[4]) ? node1333 : node1326;
										assign node1326 = (inp[12]) ? node1330 : node1327;
											assign node1327 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1330 = (inp[10]) ? 1'b0 : 1'b0;
										assign node1333 = (inp[6]) ? 1'b0 : node1334;
											assign node1334 = (inp[2]) ? 1'b0 : 1'b0;
							assign node1338 = (inp[4]) ? node1368 : node1339;
								assign node1339 = (inp[6]) ? node1355 : node1340;
									assign node1340 = (inp[11]) ? node1348 : node1341;
										assign node1341 = (inp[2]) ? node1345 : node1342;
											assign node1342 = (inp[10]) ? 1'b1 : 1'b1;
											assign node1345 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1348 = (inp[10]) ? node1352 : node1349;
											assign node1349 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1352 = (inp[8]) ? 1'b0 : 1'b0;
									assign node1355 = (inp[12]) ? node1363 : node1356;
										assign node1356 = (inp[8]) ? node1360 : node1357;
											assign node1357 = (inp[0]) ? 1'b0 : 1'b1;
											assign node1360 = (inp[0]) ? 1'b0 : 1'b0;
										assign node1363 = (inp[11]) ? 1'b0 : node1364;
											assign node1364 = (inp[0]) ? 1'b0 : 1'b0;
								assign node1368 = (inp[10]) ? node1382 : node1369;
									assign node1369 = (inp[0]) ? node1377 : node1370;
										assign node1370 = (inp[11]) ? node1374 : node1371;
											assign node1371 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1374 = (inp[6]) ? 1'b0 : 1'b0;
										assign node1377 = (inp[14]) ? 1'b0 : node1378;
											assign node1378 = (inp[6]) ? 1'b0 : 1'b0;
									assign node1382 = (inp[14]) ? 1'b0 : node1383;
										assign node1383 = (inp[0]) ? 1'b0 : node1384;
											assign node1384 = (inp[6]) ? 1'b0 : 1'b0;
					assign node1389 = (inp[0]) ? node1497 : node1390;
						assign node1390 = (inp[10]) ? node1450 : node1391;
							assign node1391 = (inp[11]) ? node1421 : node1392;
								assign node1392 = (inp[12]) ? node1406 : node1393;
									assign node1393 = (inp[6]) ? node1399 : node1394;
										assign node1394 = (inp[14]) ? node1396 : 1'b1;
											assign node1396 = (inp[5]) ? 1'b1 : 1'b1;
										assign node1399 = (inp[14]) ? node1403 : node1400;
											assign node1400 = (inp[4]) ? 1'b1 : 1'b1;
											assign node1403 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1406 = (inp[1]) ? node1414 : node1407;
										assign node1407 = (inp[2]) ? node1411 : node1408;
											assign node1408 = (inp[5]) ? 1'b1 : 1'b1;
											assign node1411 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1414 = (inp[4]) ? node1418 : node1415;
											assign node1415 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1418 = (inp[5]) ? 1'b0 : 1'b0;
								assign node1421 = (inp[6]) ? node1437 : node1422;
									assign node1422 = (inp[12]) ? node1430 : node1423;
										assign node1423 = (inp[5]) ? node1427 : node1424;
											assign node1424 = (inp[2]) ? 1'b1 : 1'b1;
											assign node1427 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1430 = (inp[8]) ? node1434 : node1431;
											assign node1431 = (inp[5]) ? 1'b0 : 1'b1;
											assign node1434 = (inp[1]) ? 1'b0 : 1'b0;
									assign node1437 = (inp[8]) ? node1445 : node1438;
										assign node1438 = (inp[4]) ? node1442 : node1439;
											assign node1439 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1442 = (inp[12]) ? 1'b0 : 1'b0;
										assign node1445 = (inp[2]) ? 1'b0 : node1446;
											assign node1446 = (inp[14]) ? 1'b0 : 1'b0;
							assign node1450 = (inp[14]) ? node1480 : node1451;
								assign node1451 = (inp[5]) ? node1467 : node1452;
									assign node1452 = (inp[12]) ? node1460 : node1453;
										assign node1453 = (inp[2]) ? node1457 : node1454;
											assign node1454 = (inp[11]) ? 1'b1 : 1'b1;
											assign node1457 = (inp[6]) ? 1'b0 : 1'b1;
										assign node1460 = (inp[4]) ? node1464 : node1461;
											assign node1461 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1464 = (inp[11]) ? 1'b0 : 1'b0;
									assign node1467 = (inp[6]) ? node1475 : node1468;
										assign node1468 = (inp[1]) ? node1472 : node1469;
											assign node1469 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1472 = (inp[4]) ? 1'b0 : 1'b0;
										assign node1475 = (inp[2]) ? 1'b0 : node1476;
											assign node1476 = (inp[12]) ? 1'b0 : 1'b0;
								assign node1480 = (inp[6]) ? node1490 : node1481;
									assign node1481 = (inp[1]) ? 1'b0 : node1482;
										assign node1482 = (inp[4]) ? node1486 : node1483;
											assign node1483 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1486 = (inp[11]) ? 1'b0 : 1'b0;
									assign node1490 = (inp[12]) ? 1'b0 : node1491;
										assign node1491 = (inp[2]) ? 1'b0 : node1492;
											assign node1492 = (inp[8]) ? 1'b0 : 1'b0;
						assign node1497 = (inp[8]) ? node1549 : node1498;
							assign node1498 = (inp[2]) ? node1528 : node1499;
								assign node1499 = (inp[5]) ? node1515 : node1500;
									assign node1500 = (inp[11]) ? node1508 : node1501;
										assign node1501 = (inp[1]) ? node1505 : node1502;
											assign node1502 = (inp[10]) ? 1'b1 : 1'b1;
											assign node1505 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1508 = (inp[6]) ? node1512 : node1509;
											assign node1509 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1512 = (inp[4]) ? 1'b0 : 1'b0;
									assign node1515 = (inp[6]) ? node1523 : node1516;
										assign node1516 = (inp[12]) ? node1520 : node1517;
											assign node1517 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1520 = (inp[14]) ? 1'b0 : 1'b0;
										assign node1523 = (inp[4]) ? 1'b0 : node1524;
											assign node1524 = (inp[1]) ? 1'b0 : 1'b0;
								assign node1528 = (inp[5]) ? node1542 : node1529;
									assign node1529 = (inp[1]) ? node1537 : node1530;
										assign node1530 = (inp[6]) ? node1534 : node1531;
											assign node1531 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1534 = (inp[11]) ? 1'b0 : 1'b0;
										assign node1537 = (inp[10]) ? 1'b0 : node1538;
											assign node1538 = (inp[12]) ? 1'b0 : 1'b0;
									assign node1542 = (inp[12]) ? 1'b0 : node1543;
										assign node1543 = (inp[6]) ? 1'b0 : node1544;
											assign node1544 = (inp[14]) ? 1'b0 : 1'b0;
							assign node1549 = (inp[11]) ? node1571 : node1550;
								assign node1550 = (inp[12]) ? node1564 : node1551;
									assign node1551 = (inp[5]) ? node1559 : node1552;
										assign node1552 = (inp[2]) ? node1556 : node1553;
											assign node1553 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1556 = (inp[6]) ? 1'b0 : 1'b0;
										assign node1559 = (inp[10]) ? 1'b0 : node1560;
											assign node1560 = (inp[4]) ? 1'b0 : 1'b0;
									assign node1564 = (inp[10]) ? 1'b0 : node1565;
										assign node1565 = (inp[1]) ? 1'b0 : node1566;
											assign node1566 = (inp[14]) ? 1'b0 : 1'b0;
								assign node1571 = (inp[4]) ? 1'b0 : node1572;
									assign node1572 = (inp[14]) ? 1'b0 : node1573;
										assign node1573 = (inp[10]) ? 1'b0 : node1574;
											assign node1574 = (inp[1]) ? 1'b0 : 1'b0;
		assign node1580 = (inp[14]) ? node2418 : node1581;
			assign node1581 = (inp[11]) ? node1999 : node1582;
				assign node1582 = (inp[2]) ? node1776 : node1583;
					assign node1583 = (inp[8]) ? node1667 : node1584;
						assign node1584 = (inp[3]) ? node1616 : node1585;
							assign node1585 = (inp[12]) ? node1595 : node1586;
								assign node1586 = (inp[9]) ? node1588 : 1'b1;
									assign node1588 = (inp[6]) ? node1590 : 1'b1;
										assign node1590 = (inp[1]) ? node1592 : 1'b1;
											assign node1592 = (inp[7]) ? 1'b1 : 1'b1;
								assign node1595 = (inp[1]) ? node1603 : node1596;
									assign node1596 = (inp[7]) ? node1598 : 1'b1;
										assign node1598 = (inp[0]) ? node1600 : 1'b1;
											assign node1600 = (inp[9]) ? 1'b1 : 1'b1;
									assign node1603 = (inp[4]) ? node1609 : node1604;
										assign node1604 = (inp[7]) ? node1606 : 1'b1;
											assign node1606 = (inp[9]) ? 1'b1 : 1'b1;
										assign node1609 = (inp[5]) ? node1613 : node1610;
											assign node1610 = (inp[0]) ? 1'b1 : 1'b1;
											assign node1613 = (inp[7]) ? 1'b0 : 1'b1;
							assign node1616 = (inp[0]) ? node1638 : node1617;
								assign node1617 = (inp[4]) ? node1625 : node1618;
									assign node1618 = (inp[12]) ? node1620 : 1'b1;
										assign node1620 = (inp[9]) ? node1622 : 1'b1;
											assign node1622 = (inp[5]) ? 1'b1 : 1'b1;
									assign node1625 = (inp[10]) ? node1631 : node1626;
										assign node1626 = (inp[1]) ? node1628 : 1'b1;
											assign node1628 = (inp[6]) ? 1'b1 : 1'b1;
										assign node1631 = (inp[7]) ? node1635 : node1632;
											assign node1632 = (inp[5]) ? 1'b1 : 1'b1;
											assign node1635 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1638 = (inp[1]) ? node1652 : node1639;
									assign node1639 = (inp[4]) ? node1645 : node1640;
										assign node1640 = (inp[5]) ? node1642 : 1'b1;
											assign node1642 = (inp[12]) ? 1'b1 : 1'b1;
										assign node1645 = (inp[7]) ? node1649 : node1646;
											assign node1646 = (inp[10]) ? 1'b1 : 1'b1;
											assign node1649 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1652 = (inp[6]) ? node1660 : node1653;
										assign node1653 = (inp[5]) ? node1657 : node1654;
											assign node1654 = (inp[10]) ? 1'b1 : 1'b1;
											assign node1657 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1660 = (inp[5]) ? node1664 : node1661;
											assign node1661 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1664 = (inp[9]) ? 1'b0 : 1'b0;
						assign node1667 = (inp[7]) ? node1717 : node1668;
							assign node1668 = (inp[1]) ? node1690 : node1669;
								assign node1669 = (inp[0]) ? node1677 : node1670;
									assign node1670 = (inp[6]) ? node1672 : 1'b1;
										assign node1672 = (inp[5]) ? node1674 : 1'b1;
											assign node1674 = (inp[3]) ? 1'b1 : 1'b1;
									assign node1677 = (inp[12]) ? node1683 : node1678;
										assign node1678 = (inp[6]) ? node1680 : 1'b1;
											assign node1680 = (inp[3]) ? 1'b1 : 1'b1;
										assign node1683 = (inp[10]) ? node1687 : node1684;
											assign node1684 = (inp[3]) ? 1'b1 : 1'b1;
											assign node1687 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1690 = (inp[12]) ? node1704 : node1691;
									assign node1691 = (inp[6]) ? node1697 : node1692;
										assign node1692 = (inp[10]) ? node1694 : 1'b1;
											assign node1694 = (inp[4]) ? 1'b1 : 1'b1;
										assign node1697 = (inp[9]) ? node1701 : node1698;
											assign node1698 = (inp[5]) ? 1'b1 : 1'b1;
											assign node1701 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1704 = (inp[5]) ? node1712 : node1705;
										assign node1705 = (inp[10]) ? node1709 : node1706;
											assign node1706 = (inp[0]) ? 1'b1 : 1'b1;
											assign node1709 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1712 = (inp[3]) ? 1'b0 : node1713;
											assign node1713 = (inp[9]) ? 1'b0 : 1'b1;
							assign node1717 = (inp[3]) ? node1747 : node1718;
								assign node1718 = (inp[5]) ? node1732 : node1719;
									assign node1719 = (inp[6]) ? node1725 : node1720;
										assign node1720 = (inp[4]) ? node1722 : 1'b1;
											assign node1722 = (inp[12]) ? 1'b1 : 1'b1;
										assign node1725 = (inp[9]) ? node1729 : node1726;
											assign node1726 = (inp[12]) ? 1'b1 : 1'b1;
											assign node1729 = (inp[0]) ? 1'b0 : 1'b1;
									assign node1732 = (inp[4]) ? node1740 : node1733;
										assign node1733 = (inp[9]) ? node1737 : node1734;
											assign node1734 = (inp[12]) ? 1'b1 : 1'b1;
											assign node1737 = (inp[1]) ? 1'b0 : 1'b1;
										assign node1740 = (inp[12]) ? node1744 : node1741;
											assign node1741 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1744 = (inp[9]) ? 1'b0 : 1'b0;
								assign node1747 = (inp[9]) ? node1763 : node1748;
									assign node1748 = (inp[1]) ? node1756 : node1749;
										assign node1749 = (inp[12]) ? node1753 : node1750;
											assign node1750 = (inp[10]) ? 1'b1 : 1'b1;
											assign node1753 = (inp[0]) ? 1'b0 : 1'b1;
										assign node1756 = (inp[4]) ? node1760 : node1757;
											assign node1757 = (inp[6]) ? 1'b0 : 1'b1;
											assign node1760 = (inp[10]) ? 1'b0 : 1'b0;
									assign node1763 = (inp[6]) ? node1771 : node1764;
										assign node1764 = (inp[12]) ? node1768 : node1765;
											assign node1765 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1768 = (inp[10]) ? 1'b0 : 1'b0;
										assign node1771 = (inp[10]) ? 1'b0 : node1772;
											assign node1772 = (inp[5]) ? 1'b0 : 1'b0;
					assign node1776 = (inp[9]) ? node1888 : node1777;
						assign node1777 = (inp[0]) ? node1829 : node1778;
							assign node1778 = (inp[10]) ? node1800 : node1779;
								assign node1779 = (inp[6]) ? node1787 : node1780;
									assign node1780 = (inp[1]) ? node1782 : 1'b1;
										assign node1782 = (inp[7]) ? node1784 : 1'b1;
											assign node1784 = (inp[12]) ? 1'b1 : 1'b1;
									assign node1787 = (inp[7]) ? node1793 : node1788;
										assign node1788 = (inp[5]) ? node1790 : 1'b1;
											assign node1790 = (inp[4]) ? 1'b1 : 1'b1;
										assign node1793 = (inp[12]) ? node1797 : node1794;
											assign node1794 = (inp[4]) ? 1'b1 : 1'b1;
											assign node1797 = (inp[8]) ? 1'b0 : 1'b1;
								assign node1800 = (inp[8]) ? node1814 : node1801;
									assign node1801 = (inp[5]) ? node1807 : node1802;
										assign node1802 = (inp[7]) ? node1804 : 1'b1;
											assign node1804 = (inp[3]) ? 1'b1 : 1'b1;
										assign node1807 = (inp[6]) ? node1811 : node1808;
											assign node1808 = (inp[12]) ? 1'b1 : 1'b1;
											assign node1811 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1814 = (inp[7]) ? node1822 : node1815;
										assign node1815 = (inp[6]) ? node1819 : node1816;
											assign node1816 = (inp[5]) ? 1'b1 : 1'b1;
											assign node1819 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1822 = (inp[6]) ? node1826 : node1823;
											assign node1823 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1826 = (inp[1]) ? 1'b0 : 1'b0;
							assign node1829 = (inp[5]) ? node1859 : node1830;
								assign node1830 = (inp[12]) ? node1844 : node1831;
									assign node1831 = (inp[3]) ? node1837 : node1832;
										assign node1832 = (inp[6]) ? node1834 : 1'b1;
											assign node1834 = (inp[10]) ? 1'b1 : 1'b1;
										assign node1837 = (inp[8]) ? node1841 : node1838;
											assign node1838 = (inp[7]) ? 1'b1 : 1'b1;
											assign node1841 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1844 = (inp[4]) ? node1852 : node1845;
										assign node1845 = (inp[1]) ? node1849 : node1846;
											assign node1846 = (inp[10]) ? 1'b1 : 1'b1;
											assign node1849 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1852 = (inp[1]) ? node1856 : node1853;
											assign node1853 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1856 = (inp[6]) ? 1'b0 : 1'b0;
								assign node1859 = (inp[1]) ? node1875 : node1860;
									assign node1860 = (inp[6]) ? node1868 : node1861;
										assign node1861 = (inp[4]) ? node1865 : node1862;
											assign node1862 = (inp[3]) ? 1'b1 : 1'b1;
											assign node1865 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1868 = (inp[3]) ? node1872 : node1869;
											assign node1869 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1872 = (inp[7]) ? 1'b0 : 1'b0;
									assign node1875 = (inp[10]) ? node1883 : node1876;
										assign node1876 = (inp[6]) ? node1880 : node1877;
											assign node1877 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1880 = (inp[4]) ? 1'b0 : 1'b0;
										assign node1883 = (inp[3]) ? 1'b0 : node1884;
											assign node1884 = (inp[12]) ? 1'b0 : 1'b0;
						assign node1888 = (inp[7]) ? node1948 : node1889;
							assign node1889 = (inp[8]) ? node1919 : node1890;
								assign node1890 = (inp[10]) ? node1904 : node1891;
									assign node1891 = (inp[3]) ? node1897 : node1892;
										assign node1892 = (inp[5]) ? node1894 : 1'b1;
											assign node1894 = (inp[1]) ? 1'b1 : 1'b1;
										assign node1897 = (inp[6]) ? node1901 : node1898;
											assign node1898 = (inp[0]) ? 1'b1 : 1'b1;
											assign node1901 = (inp[5]) ? 1'b0 : 1'b1;
									assign node1904 = (inp[6]) ? node1912 : node1905;
										assign node1905 = (inp[5]) ? node1909 : node1906;
											assign node1906 = (inp[4]) ? 1'b1 : 1'b1;
											assign node1909 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1912 = (inp[0]) ? node1916 : node1913;
											assign node1913 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1916 = (inp[1]) ? 1'b0 : 1'b0;
								assign node1919 = (inp[10]) ? node1935 : node1920;
									assign node1920 = (inp[12]) ? node1928 : node1921;
										assign node1921 = (inp[6]) ? node1925 : node1922;
											assign node1922 = (inp[1]) ? 1'b1 : 1'b1;
											assign node1925 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1928 = (inp[1]) ? node1932 : node1929;
											assign node1929 = (inp[5]) ? 1'b0 : 1'b1;
											assign node1932 = (inp[0]) ? 1'b0 : 1'b0;
									assign node1935 = (inp[1]) ? node1943 : node1936;
										assign node1936 = (inp[0]) ? node1940 : node1937;
											assign node1937 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1940 = (inp[3]) ? 1'b0 : 1'b0;
										assign node1943 = (inp[6]) ? 1'b0 : node1944;
											assign node1944 = (inp[4]) ? 1'b0 : 1'b0;
							assign node1948 = (inp[5]) ? node1978 : node1949;
								assign node1949 = (inp[3]) ? node1965 : node1950;
									assign node1950 = (inp[1]) ? node1958 : node1951;
										assign node1951 = (inp[6]) ? node1955 : node1952;
											assign node1952 = (inp[12]) ? 1'b1 : 1'b1;
											assign node1955 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1958 = (inp[6]) ? node1962 : node1959;
											assign node1959 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1962 = (inp[0]) ? 1'b0 : 1'b0;
									assign node1965 = (inp[12]) ? node1973 : node1966;
										assign node1966 = (inp[10]) ? node1970 : node1967;
											assign node1967 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1970 = (inp[4]) ? 1'b0 : 1'b0;
										assign node1973 = (inp[8]) ? 1'b0 : node1974;
											assign node1974 = (inp[6]) ? 1'b0 : 1'b0;
								assign node1978 = (inp[4]) ? node1992 : node1979;
									assign node1979 = (inp[12]) ? node1987 : node1980;
										assign node1980 = (inp[3]) ? node1984 : node1981;
											assign node1981 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1984 = (inp[10]) ? 1'b0 : 1'b0;
										assign node1987 = (inp[0]) ? 1'b0 : node1988;
											assign node1988 = (inp[10]) ? 1'b0 : 1'b0;
									assign node1992 = (inp[12]) ? 1'b0 : node1993;
										assign node1993 = (inp[1]) ? 1'b0 : node1994;
											assign node1994 = (inp[6]) ? 1'b0 : 1'b0;
				assign node1999 = (inp[12]) ? node2223 : node2000;
					assign node2000 = (inp[3]) ? node2112 : node2001;
						assign node2001 = (inp[5]) ? node2053 : node2002;
							assign node2002 = (inp[6]) ? node2024 : node2003;
								assign node2003 = (inp[2]) ? node2011 : node2004;
									assign node2004 = (inp[10]) ? node2006 : 1'b1;
										assign node2006 = (inp[8]) ? node2008 : 1'b1;
											assign node2008 = (inp[4]) ? 1'b1 : 1'b1;
									assign node2011 = (inp[8]) ? node2017 : node2012;
										assign node2012 = (inp[0]) ? node2014 : 1'b1;
											assign node2014 = (inp[1]) ? 1'b1 : 1'b1;
										assign node2017 = (inp[4]) ? node2021 : node2018;
											assign node2018 = (inp[9]) ? 1'b1 : 1'b1;
											assign node2021 = (inp[1]) ? 1'b0 : 1'b1;
								assign node2024 = (inp[4]) ? node2038 : node2025;
									assign node2025 = (inp[9]) ? node2031 : node2026;
										assign node2026 = (inp[8]) ? node2028 : 1'b1;
											assign node2028 = (inp[10]) ? 1'b1 : 1'b1;
										assign node2031 = (inp[10]) ? node2035 : node2032;
											assign node2032 = (inp[8]) ? 1'b1 : 1'b1;
											assign node2035 = (inp[8]) ? 1'b0 : 1'b1;
									assign node2038 = (inp[0]) ? node2046 : node2039;
										assign node2039 = (inp[2]) ? node2043 : node2040;
											assign node2040 = (inp[10]) ? 1'b1 : 1'b1;
											assign node2043 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2046 = (inp[7]) ? node2050 : node2047;
											assign node2047 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2050 = (inp[9]) ? 1'b0 : 1'b0;
							assign node2053 = (inp[9]) ? node2083 : node2054;
								assign node2054 = (inp[8]) ? node2068 : node2055;
									assign node2055 = (inp[0]) ? node2061 : node2056;
										assign node2056 = (inp[1]) ? node2058 : 1'b1;
											assign node2058 = (inp[6]) ? 1'b1 : 1'b1;
										assign node2061 = (inp[10]) ? node2065 : node2062;
											assign node2062 = (inp[1]) ? 1'b1 : 1'b1;
											assign node2065 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2068 = (inp[10]) ? node2076 : node2069;
										assign node2069 = (inp[1]) ? node2073 : node2070;
											assign node2070 = (inp[6]) ? 1'b1 : 1'b1;
											assign node2073 = (inp[6]) ? 1'b0 : 1'b1;
										assign node2076 = (inp[6]) ? node2080 : node2077;
											assign node2077 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2080 = (inp[0]) ? 1'b0 : 1'b0;
								assign node2083 = (inp[4]) ? node2099 : node2084;
									assign node2084 = (inp[1]) ? node2092 : node2085;
										assign node2085 = (inp[2]) ? node2089 : node2086;
											assign node2086 = (inp[6]) ? 1'b1 : 1'b1;
											assign node2089 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2092 = (inp[6]) ? node2096 : node2093;
											assign node2093 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2096 = (inp[7]) ? 1'b0 : 1'b0;
									assign node2099 = (inp[0]) ? node2107 : node2100;
										assign node2100 = (inp[7]) ? node2104 : node2101;
											assign node2101 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2104 = (inp[6]) ? 1'b0 : 1'b0;
										assign node2107 = (inp[10]) ? 1'b0 : node2108;
											assign node2108 = (inp[1]) ? 1'b0 : 1'b0;
						assign node2112 = (inp[10]) ? node2172 : node2113;
							assign node2113 = (inp[0]) ? node2143 : node2114;
								assign node2114 = (inp[6]) ? node2128 : node2115;
									assign node2115 = (inp[4]) ? node2121 : node2116;
										assign node2116 = (inp[1]) ? node2118 : 1'b1;
											assign node2118 = (inp[2]) ? 1'b1 : 1'b1;
										assign node2121 = (inp[2]) ? node2125 : node2122;
											assign node2122 = (inp[8]) ? 1'b1 : 1'b1;
											assign node2125 = (inp[1]) ? 1'b0 : 1'b1;
									assign node2128 = (inp[4]) ? node2136 : node2129;
										assign node2129 = (inp[8]) ? node2133 : node2130;
											assign node2130 = (inp[2]) ? 1'b1 : 1'b1;
											assign node2133 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2136 = (inp[8]) ? node2140 : node2137;
											assign node2137 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2140 = (inp[7]) ? 1'b0 : 1'b0;
								assign node2143 = (inp[8]) ? node2159 : node2144;
									assign node2144 = (inp[1]) ? node2152 : node2145;
										assign node2145 = (inp[5]) ? node2149 : node2146;
											assign node2146 = (inp[2]) ? 1'b1 : 1'b1;
											assign node2149 = (inp[4]) ? 1'b0 : 1'b1;
										assign node2152 = (inp[9]) ? node2156 : node2153;
											assign node2153 = (inp[6]) ? 1'b0 : 1'b1;
											assign node2156 = (inp[7]) ? 1'b0 : 1'b0;
									assign node2159 = (inp[9]) ? node2167 : node2160;
										assign node2160 = (inp[4]) ? node2164 : node2161;
											assign node2161 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2164 = (inp[2]) ? 1'b0 : 1'b0;
										assign node2167 = (inp[5]) ? 1'b0 : node2168;
											assign node2168 = (inp[6]) ? 1'b0 : 1'b0;
							assign node2172 = (inp[8]) ? node2202 : node2173;
								assign node2173 = (inp[7]) ? node2189 : node2174;
									assign node2174 = (inp[2]) ? node2182 : node2175;
										assign node2175 = (inp[5]) ? node2179 : node2176;
											assign node2176 = (inp[1]) ? 1'b1 : 1'b1;
											assign node2179 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2182 = (inp[4]) ? node2186 : node2183;
											assign node2183 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2186 = (inp[6]) ? 1'b0 : 1'b0;
									assign node2189 = (inp[9]) ? node2197 : node2190;
										assign node2190 = (inp[1]) ? node2194 : node2191;
											assign node2191 = (inp[2]) ? 1'b0 : 1'b1;
											assign node2194 = (inp[6]) ? 1'b0 : 1'b0;
										assign node2197 = (inp[4]) ? 1'b0 : node2198;
											assign node2198 = (inp[6]) ? 1'b0 : 1'b0;
								assign node2202 = (inp[1]) ? node2216 : node2203;
									assign node2203 = (inp[4]) ? node2211 : node2204;
										assign node2204 = (inp[5]) ? node2208 : node2205;
											assign node2205 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2208 = (inp[7]) ? 1'b0 : 1'b0;
										assign node2211 = (inp[0]) ? 1'b0 : node2212;
											assign node2212 = (inp[9]) ? 1'b0 : 1'b0;
									assign node2216 = (inp[5]) ? 1'b0 : node2217;
										assign node2217 = (inp[2]) ? 1'b0 : node2218;
											assign node2218 = (inp[0]) ? 1'b0 : 1'b0;
					assign node2223 = (inp[6]) ? node2335 : node2224;
						assign node2224 = (inp[2]) ? node2284 : node2225;
							assign node2225 = (inp[5]) ? node2255 : node2226;
								assign node2226 = (inp[7]) ? node2240 : node2227;
									assign node2227 = (inp[1]) ? node2233 : node2228;
										assign node2228 = (inp[4]) ? node2230 : 1'b1;
											assign node2230 = (inp[0]) ? 1'b1 : 1'b1;
										assign node2233 = (inp[3]) ? node2237 : node2234;
											assign node2234 = (inp[4]) ? 1'b1 : 1'b1;
											assign node2237 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2240 = (inp[0]) ? node2248 : node2241;
										assign node2241 = (inp[8]) ? node2245 : node2242;
											assign node2242 = (inp[4]) ? 1'b1 : 1'b1;
											assign node2245 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2248 = (inp[9]) ? node2252 : node2249;
											assign node2249 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2252 = (inp[10]) ? 1'b0 : 1'b0;
								assign node2255 = (inp[9]) ? node2271 : node2256;
									assign node2256 = (inp[0]) ? node2264 : node2257;
										assign node2257 = (inp[8]) ? node2261 : node2258;
											assign node2258 = (inp[7]) ? 1'b1 : 1'b1;
											assign node2261 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2264 = (inp[1]) ? node2268 : node2265;
											assign node2265 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2268 = (inp[4]) ? 1'b0 : 1'b0;
									assign node2271 = (inp[10]) ? node2279 : node2272;
										assign node2272 = (inp[3]) ? node2276 : node2273;
											assign node2273 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2276 = (inp[4]) ? 1'b0 : 1'b0;
										assign node2279 = (inp[8]) ? 1'b0 : node2280;
											assign node2280 = (inp[3]) ? 1'b0 : 1'b0;
							assign node2284 = (inp[3]) ? node2314 : node2285;
								assign node2285 = (inp[7]) ? node2301 : node2286;
									assign node2286 = (inp[0]) ? node2294 : node2287;
										assign node2287 = (inp[9]) ? node2291 : node2288;
											assign node2288 = (inp[5]) ? 1'b1 : 1'b1;
											assign node2291 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2294 = (inp[1]) ? node2298 : node2295;
											assign node2295 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2298 = (inp[5]) ? 1'b0 : 1'b0;
									assign node2301 = (inp[4]) ? node2309 : node2302;
										assign node2302 = (inp[10]) ? node2306 : node2303;
											assign node2303 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2306 = (inp[1]) ? 1'b0 : 1'b0;
										assign node2309 = (inp[0]) ? 1'b0 : node2310;
											assign node2310 = (inp[10]) ? 1'b0 : 1'b0;
								assign node2314 = (inp[10]) ? node2328 : node2315;
									assign node2315 = (inp[4]) ? node2323 : node2316;
										assign node2316 = (inp[8]) ? node2320 : node2317;
											assign node2317 = (inp[0]) ? 1'b0 : 1'b1;
											assign node2320 = (inp[0]) ? 1'b0 : 1'b0;
										assign node2323 = (inp[5]) ? 1'b0 : node2324;
											assign node2324 = (inp[1]) ? 1'b0 : 1'b0;
									assign node2328 = (inp[0]) ? 1'b0 : node2329;
										assign node2329 = (inp[5]) ? 1'b0 : node2330;
											assign node2330 = (inp[8]) ? 1'b0 : 1'b0;
						assign node2335 = (inp[3]) ? node2387 : node2336;
							assign node2336 = (inp[10]) ? node2366 : node2337;
								assign node2337 = (inp[2]) ? node2353 : node2338;
									assign node2338 = (inp[5]) ? node2346 : node2339;
										assign node2339 = (inp[8]) ? node2343 : node2340;
											assign node2340 = (inp[7]) ? 1'b1 : 1'b1;
											assign node2343 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2346 = (inp[9]) ? node2350 : node2347;
											assign node2347 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2350 = (inp[0]) ? 1'b0 : 1'b0;
									assign node2353 = (inp[8]) ? node2361 : node2354;
										assign node2354 = (inp[0]) ? node2358 : node2355;
											assign node2355 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2358 = (inp[4]) ? 1'b0 : 1'b0;
										assign node2361 = (inp[4]) ? 1'b0 : node2362;
											assign node2362 = (inp[0]) ? 1'b0 : 1'b0;
								assign node2366 = (inp[5]) ? node2380 : node2367;
									assign node2367 = (inp[9]) ? node2375 : node2368;
										assign node2368 = (inp[1]) ? node2372 : node2369;
											assign node2369 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2372 = (inp[0]) ? 1'b0 : 1'b0;
										assign node2375 = (inp[4]) ? 1'b0 : node2376;
											assign node2376 = (inp[8]) ? 1'b0 : 1'b0;
									assign node2380 = (inp[7]) ? 1'b0 : node2381;
										assign node2381 = (inp[4]) ? 1'b0 : node2382;
											assign node2382 = (inp[9]) ? 1'b0 : 1'b0;
							assign node2387 = (inp[4]) ? node2409 : node2388;
								assign node2388 = (inp[8]) ? node2402 : node2389;
									assign node2389 = (inp[2]) ? node2397 : node2390;
										assign node2390 = (inp[0]) ? node2394 : node2391;
											assign node2391 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2394 = (inp[10]) ? 1'b0 : 1'b0;
										assign node2397 = (inp[5]) ? 1'b0 : node2398;
											assign node2398 = (inp[1]) ? 1'b0 : 1'b0;
									assign node2402 = (inp[9]) ? 1'b0 : node2403;
										assign node2403 = (inp[7]) ? 1'b0 : node2404;
											assign node2404 = (inp[10]) ? 1'b0 : 1'b0;
								assign node2409 = (inp[5]) ? 1'b0 : node2410;
									assign node2410 = (inp[9]) ? 1'b0 : node2411;
										assign node2411 = (inp[0]) ? 1'b0 : node2412;
											assign node2412 = (inp[7]) ? 1'b0 : 1'b0;
			assign node2418 = (inp[2]) ? node2838 : node2419;
				assign node2419 = (inp[9]) ? node2643 : node2420;
					assign node2420 = (inp[3]) ? node2532 : node2421;
						assign node2421 = (inp[6]) ? node2473 : node2422;
							assign node2422 = (inp[7]) ? node2444 : node2423;
								assign node2423 = (inp[4]) ? node2431 : node2424;
									assign node2424 = (inp[12]) ? node2426 : 1'b1;
										assign node2426 = (inp[8]) ? node2428 : 1'b1;
											assign node2428 = (inp[5]) ? 1'b1 : 1'b1;
									assign node2431 = (inp[5]) ? node2437 : node2432;
										assign node2432 = (inp[12]) ? node2434 : 1'b1;
											assign node2434 = (inp[1]) ? 1'b1 : 1'b1;
										assign node2437 = (inp[12]) ? node2441 : node2438;
											assign node2438 = (inp[10]) ? 1'b1 : 1'b1;
											assign node2441 = (inp[10]) ? 1'b0 : 1'b1;
								assign node2444 = (inp[11]) ? node2458 : node2445;
									assign node2445 = (inp[5]) ? node2451 : node2446;
										assign node2446 = (inp[8]) ? node2448 : 1'b1;
											assign node2448 = (inp[12]) ? 1'b1 : 1'b1;
										assign node2451 = (inp[10]) ? node2455 : node2452;
											assign node2452 = (inp[0]) ? 1'b1 : 1'b1;
											assign node2455 = (inp[0]) ? 1'b0 : 1'b1;
									assign node2458 = (inp[8]) ? node2466 : node2459;
										assign node2459 = (inp[5]) ? node2463 : node2460;
											assign node2460 = (inp[10]) ? 1'b1 : 1'b1;
											assign node2463 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2466 = (inp[12]) ? node2470 : node2467;
											assign node2467 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2470 = (inp[1]) ? 1'b0 : 1'b0;
							assign node2473 = (inp[10]) ? node2503 : node2474;
								assign node2474 = (inp[1]) ? node2488 : node2475;
									assign node2475 = (inp[7]) ? node2481 : node2476;
										assign node2476 = (inp[4]) ? node2478 : 1'b1;
											assign node2478 = (inp[11]) ? 1'b1 : 1'b1;
										assign node2481 = (inp[11]) ? node2485 : node2482;
											assign node2482 = (inp[5]) ? 1'b1 : 1'b1;
											assign node2485 = (inp[12]) ? 1'b0 : 1'b1;
									assign node2488 = (inp[11]) ? node2496 : node2489;
										assign node2489 = (inp[4]) ? node2493 : node2490;
											assign node2490 = (inp[0]) ? 1'b1 : 1'b1;
											assign node2493 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2496 = (inp[4]) ? node2500 : node2497;
											assign node2497 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2500 = (inp[0]) ? 1'b0 : 1'b0;
								assign node2503 = (inp[12]) ? node2519 : node2504;
									assign node2504 = (inp[0]) ? node2512 : node2505;
										assign node2505 = (inp[11]) ? node2509 : node2506;
											assign node2506 = (inp[7]) ? 1'b1 : 1'b1;
											assign node2509 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2512 = (inp[11]) ? node2516 : node2513;
											assign node2513 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2516 = (inp[1]) ? 1'b0 : 1'b0;
									assign node2519 = (inp[4]) ? node2527 : node2520;
										assign node2520 = (inp[7]) ? node2524 : node2521;
											assign node2521 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2524 = (inp[0]) ? 1'b0 : 1'b0;
										assign node2527 = (inp[1]) ? 1'b0 : node2528;
											assign node2528 = (inp[11]) ? 1'b0 : 1'b0;
						assign node2532 = (inp[4]) ? node2592 : node2533;
							assign node2533 = (inp[8]) ? node2563 : node2534;
								assign node2534 = (inp[7]) ? node2548 : node2535;
									assign node2535 = (inp[6]) ? node2541 : node2536;
										assign node2536 = (inp[1]) ? node2538 : 1'b1;
											assign node2538 = (inp[12]) ? 1'b1 : 1'b1;
										assign node2541 = (inp[5]) ? node2545 : node2542;
											assign node2542 = (inp[12]) ? 1'b1 : 1'b1;
											assign node2545 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2548 = (inp[10]) ? node2556 : node2549;
										assign node2549 = (inp[6]) ? node2553 : node2550;
											assign node2550 = (inp[11]) ? 1'b1 : 1'b1;
											assign node2553 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2556 = (inp[0]) ? node2560 : node2557;
											assign node2557 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2560 = (inp[1]) ? 1'b0 : 1'b0;
								assign node2563 = (inp[0]) ? node2579 : node2564;
									assign node2564 = (inp[5]) ? node2572 : node2565;
										assign node2565 = (inp[7]) ? node2569 : node2566;
											assign node2566 = (inp[10]) ? 1'b1 : 1'b1;
											assign node2569 = (inp[1]) ? 1'b0 : 1'b1;
										assign node2572 = (inp[11]) ? node2576 : node2573;
											assign node2573 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2576 = (inp[1]) ? 1'b0 : 1'b0;
									assign node2579 = (inp[6]) ? node2587 : node2580;
										assign node2580 = (inp[7]) ? node2584 : node2581;
											assign node2581 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2584 = (inp[11]) ? 1'b0 : 1'b0;
										assign node2587 = (inp[5]) ? 1'b0 : node2588;
											assign node2588 = (inp[7]) ? 1'b0 : 1'b0;
							assign node2592 = (inp[11]) ? node2622 : node2593;
								assign node2593 = (inp[1]) ? node2609 : node2594;
									assign node2594 = (inp[10]) ? node2602 : node2595;
										assign node2595 = (inp[0]) ? node2599 : node2596;
											assign node2596 = (inp[7]) ? 1'b1 : 1'b1;
											assign node2599 = (inp[12]) ? 1'b0 : 1'b1;
										assign node2602 = (inp[7]) ? node2606 : node2603;
											assign node2603 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2606 = (inp[6]) ? 1'b0 : 1'b0;
									assign node2609 = (inp[12]) ? node2617 : node2610;
										assign node2610 = (inp[5]) ? node2614 : node2611;
											assign node2611 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2614 = (inp[6]) ? 1'b0 : 1'b0;
										assign node2617 = (inp[7]) ? 1'b0 : node2618;
											assign node2618 = (inp[8]) ? 1'b0 : 1'b0;
								assign node2622 = (inp[0]) ? node2636 : node2623;
									assign node2623 = (inp[12]) ? node2631 : node2624;
										assign node2624 = (inp[8]) ? node2628 : node2625;
											assign node2625 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2628 = (inp[5]) ? 1'b0 : 1'b0;
										assign node2631 = (inp[5]) ? 1'b0 : node2632;
											assign node2632 = (inp[7]) ? 1'b0 : 1'b0;
									assign node2636 = (inp[6]) ? 1'b0 : node2637;
										assign node2637 = (inp[7]) ? 1'b0 : node2638;
											assign node2638 = (inp[1]) ? 1'b0 : 1'b0;
					assign node2643 = (inp[6]) ? node2755 : node2644;
						assign node2644 = (inp[12]) ? node2704 : node2645;
							assign node2645 = (inp[8]) ? node2675 : node2646;
								assign node2646 = (inp[5]) ? node2660 : node2647;
									assign node2647 = (inp[10]) ? node2653 : node2648;
										assign node2648 = (inp[0]) ? node2650 : 1'b1;
											assign node2650 = (inp[11]) ? 1'b1 : 1'b1;
										assign node2653 = (inp[3]) ? node2657 : node2654;
											assign node2654 = (inp[4]) ? 1'b1 : 1'b1;
											assign node2657 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2660 = (inp[1]) ? node2668 : node2661;
										assign node2661 = (inp[4]) ? node2665 : node2662;
											assign node2662 = (inp[0]) ? 1'b1 : 1'b1;
											assign node2665 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2668 = (inp[7]) ? node2672 : node2669;
											assign node2669 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2672 = (inp[10]) ? 1'b0 : 1'b0;
								assign node2675 = (inp[1]) ? node2691 : node2676;
									assign node2676 = (inp[4]) ? node2684 : node2677;
										assign node2677 = (inp[10]) ? node2681 : node2678;
											assign node2678 = (inp[11]) ? 1'b1 : 1'b1;
											assign node2681 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2684 = (inp[7]) ? node2688 : node2685;
											assign node2685 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2688 = (inp[5]) ? 1'b0 : 1'b0;
									assign node2691 = (inp[0]) ? node2699 : node2692;
										assign node2692 = (inp[5]) ? node2696 : node2693;
											assign node2693 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2696 = (inp[11]) ? 1'b0 : 1'b0;
										assign node2699 = (inp[7]) ? 1'b0 : node2700;
											assign node2700 = (inp[4]) ? 1'b0 : 1'b0;
							assign node2704 = (inp[3]) ? node2734 : node2705;
								assign node2705 = (inp[7]) ? node2721 : node2706;
									assign node2706 = (inp[5]) ? node2714 : node2707;
										assign node2707 = (inp[10]) ? node2711 : node2708;
											assign node2708 = (inp[8]) ? 1'b1 : 1'b1;
											assign node2711 = (inp[4]) ? 1'b0 : 1'b1;
										assign node2714 = (inp[10]) ? node2718 : node2715;
											assign node2715 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2718 = (inp[8]) ? 1'b0 : 1'b0;
									assign node2721 = (inp[10]) ? node2729 : node2722;
										assign node2722 = (inp[0]) ? node2726 : node2723;
											assign node2723 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2726 = (inp[8]) ? 1'b0 : 1'b0;
										assign node2729 = (inp[5]) ? 1'b0 : node2730;
											assign node2730 = (inp[1]) ? 1'b0 : 1'b0;
								assign node2734 = (inp[7]) ? node2748 : node2735;
									assign node2735 = (inp[4]) ? node2743 : node2736;
										assign node2736 = (inp[8]) ? node2740 : node2737;
											assign node2737 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2740 = (inp[1]) ? 1'b0 : 1'b0;
										assign node2743 = (inp[1]) ? 1'b0 : node2744;
											assign node2744 = (inp[11]) ? 1'b0 : 1'b0;
									assign node2748 = (inp[4]) ? 1'b0 : node2749;
										assign node2749 = (inp[10]) ? 1'b0 : node2750;
											assign node2750 = (inp[0]) ? 1'b0 : 1'b0;
						assign node2755 = (inp[3]) ? node2807 : node2756;
							assign node2756 = (inp[1]) ? node2786 : node2757;
								assign node2757 = (inp[10]) ? node2773 : node2758;
									assign node2758 = (inp[5]) ? node2766 : node2759;
										assign node2759 = (inp[11]) ? node2763 : node2760;
											assign node2760 = (inp[0]) ? 1'b1 : 1'b1;
											assign node2763 = (inp[4]) ? 1'b0 : 1'b1;
										assign node2766 = (inp[12]) ? node2770 : node2767;
											assign node2767 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2770 = (inp[11]) ? 1'b0 : 1'b0;
									assign node2773 = (inp[8]) ? node2781 : node2774;
										assign node2774 = (inp[7]) ? node2778 : node2775;
											assign node2775 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2778 = (inp[11]) ? 1'b0 : 1'b0;
										assign node2781 = (inp[4]) ? 1'b0 : node2782;
											assign node2782 = (inp[12]) ? 1'b0 : 1'b0;
								assign node2786 = (inp[12]) ? node2800 : node2787;
									assign node2787 = (inp[0]) ? node2795 : node2788;
										assign node2788 = (inp[8]) ? node2792 : node2789;
											assign node2789 = (inp[5]) ? 1'b0 : 1'b1;
											assign node2792 = (inp[11]) ? 1'b0 : 1'b0;
										assign node2795 = (inp[11]) ? 1'b0 : node2796;
											assign node2796 = (inp[5]) ? 1'b0 : 1'b0;
									assign node2800 = (inp[5]) ? 1'b0 : node2801;
										assign node2801 = (inp[0]) ? 1'b0 : node2802;
											assign node2802 = (inp[8]) ? 1'b0 : 1'b0;
							assign node2807 = (inp[7]) ? node2829 : node2808;
								assign node2808 = (inp[4]) ? node2822 : node2809;
									assign node2809 = (inp[10]) ? node2817 : node2810;
										assign node2810 = (inp[12]) ? node2814 : node2811;
											assign node2811 = (inp[0]) ? 1'b0 : 1'b1;
											assign node2814 = (inp[8]) ? 1'b0 : 1'b0;
										assign node2817 = (inp[0]) ? 1'b0 : node2818;
											assign node2818 = (inp[11]) ? 1'b0 : 1'b0;
									assign node2822 = (inp[11]) ? 1'b0 : node2823;
										assign node2823 = (inp[5]) ? 1'b0 : node2824;
											assign node2824 = (inp[10]) ? 1'b0 : 1'b0;
								assign node2829 = (inp[5]) ? 1'b0 : node2830;
									assign node2830 = (inp[1]) ? 1'b0 : node2831;
										assign node2831 = (inp[4]) ? 1'b0 : node2832;
											assign node2832 = (inp[11]) ? 1'b0 : 1'b0;
				assign node2838 = (inp[6]) ? node3034 : node2839;
					assign node2839 = (inp[4]) ? node2951 : node2840;
						assign node2840 = (inp[8]) ? node2900 : node2841;
							assign node2841 = (inp[0]) ? node2871 : node2842;
								assign node2842 = (inp[10]) ? node2856 : node2843;
									assign node2843 = (inp[3]) ? node2849 : node2844;
										assign node2844 = (inp[1]) ? node2846 : 1'b1;
											assign node2846 = (inp[11]) ? 1'b1 : 1'b1;
										assign node2849 = (inp[1]) ? node2853 : node2850;
											assign node2850 = (inp[7]) ? 1'b1 : 1'b1;
											assign node2853 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2856 = (inp[12]) ? node2864 : node2857;
										assign node2857 = (inp[7]) ? node2861 : node2858;
											assign node2858 = (inp[9]) ? 1'b1 : 1'b1;
											assign node2861 = (inp[11]) ? 1'b0 : 1'b1;
										assign node2864 = (inp[5]) ? node2868 : node2865;
											assign node2865 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2868 = (inp[7]) ? 1'b0 : 1'b0;
								assign node2871 = (inp[1]) ? node2887 : node2872;
									assign node2872 = (inp[11]) ? node2880 : node2873;
										assign node2873 = (inp[10]) ? node2877 : node2874;
											assign node2874 = (inp[7]) ? 1'b1 : 1'b1;
											assign node2877 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2880 = (inp[10]) ? node2884 : node2881;
											assign node2881 = (inp[12]) ? 1'b0 : 1'b1;
											assign node2884 = (inp[9]) ? 1'b0 : 1'b0;
									assign node2887 = (inp[9]) ? node2895 : node2888;
										assign node2888 = (inp[11]) ? node2892 : node2889;
											assign node2889 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2892 = (inp[12]) ? 1'b0 : 1'b0;
										assign node2895 = (inp[7]) ? 1'b0 : node2896;
											assign node2896 = (inp[3]) ? 1'b0 : 1'b0;
							assign node2900 = (inp[9]) ? node2930 : node2901;
								assign node2901 = (inp[0]) ? node2917 : node2902;
									assign node2902 = (inp[7]) ? node2910 : node2903;
										assign node2903 = (inp[3]) ? node2907 : node2904;
											assign node2904 = (inp[10]) ? 1'b1 : 1'b1;
											assign node2907 = (inp[12]) ? 1'b0 : 1'b1;
										assign node2910 = (inp[3]) ? node2914 : node2911;
											assign node2911 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2914 = (inp[11]) ? 1'b0 : 1'b0;
									assign node2917 = (inp[5]) ? node2925 : node2918;
										assign node2918 = (inp[1]) ? node2922 : node2919;
											assign node2919 = (inp[7]) ? 1'b0 : 1'b1;
											assign node2922 = (inp[12]) ? 1'b0 : 1'b0;
										assign node2925 = (inp[3]) ? 1'b0 : node2926;
											assign node2926 = (inp[11]) ? 1'b0 : 1'b0;
								assign node2930 = (inp[1]) ? node2944 : node2931;
									assign node2931 = (inp[10]) ? node2939 : node2932;
										assign node2932 = (inp[5]) ? node2936 : node2933;
											assign node2933 = (inp[0]) ? 1'b0 : 1'b1;
											assign node2936 = (inp[7]) ? 1'b0 : 1'b0;
										assign node2939 = (inp[11]) ? 1'b0 : node2940;
											assign node2940 = (inp[5]) ? 1'b0 : 1'b0;
									assign node2944 = (inp[3]) ? 1'b0 : node2945;
										assign node2945 = (inp[5]) ? 1'b0 : node2946;
											assign node2946 = (inp[11]) ? 1'b0 : 1'b0;
						assign node2951 = (inp[12]) ? node3003 : node2952;
							assign node2952 = (inp[11]) ? node2982 : node2953;
								assign node2953 = (inp[9]) ? node2969 : node2954;
									assign node2954 = (inp[7]) ? node2962 : node2955;
										assign node2955 = (inp[1]) ? node2959 : node2956;
											assign node2956 = (inp[5]) ? 1'b1 : 1'b1;
											assign node2959 = (inp[0]) ? 1'b0 : 1'b1;
										assign node2962 = (inp[10]) ? node2966 : node2963;
											assign node2963 = (inp[1]) ? 1'b0 : 1'b1;
											assign node2966 = (inp[5]) ? 1'b0 : 1'b0;
									assign node2969 = (inp[8]) ? node2977 : node2970;
										assign node2970 = (inp[3]) ? node2974 : node2971;
											assign node2971 = (inp[10]) ? 1'b0 : 1'b1;
											assign node2974 = (inp[0]) ? 1'b0 : 1'b0;
										assign node2977 = (inp[0]) ? 1'b0 : node2978;
											assign node2978 = (inp[3]) ? 1'b0 : 1'b0;
								assign node2982 = (inp[8]) ? node2996 : node2983;
									assign node2983 = (inp[10]) ? node2991 : node2984;
										assign node2984 = (inp[7]) ? node2988 : node2985;
											assign node2985 = (inp[0]) ? 1'b0 : 1'b1;
											assign node2988 = (inp[1]) ? 1'b0 : 1'b0;
										assign node2991 = (inp[0]) ? 1'b0 : node2992;
											assign node2992 = (inp[9]) ? 1'b0 : 1'b0;
									assign node2996 = (inp[7]) ? 1'b0 : node2997;
										assign node2997 = (inp[0]) ? 1'b0 : node2998;
											assign node2998 = (inp[9]) ? 1'b0 : 1'b0;
							assign node3003 = (inp[1]) ? node3025 : node3004;
								assign node3004 = (inp[8]) ? node3018 : node3005;
									assign node3005 = (inp[5]) ? node3013 : node3006;
										assign node3006 = (inp[7]) ? node3010 : node3007;
											assign node3007 = (inp[11]) ? 1'b0 : 1'b1;
											assign node3010 = (inp[10]) ? 1'b0 : 1'b0;
										assign node3013 = (inp[11]) ? 1'b0 : node3014;
											assign node3014 = (inp[10]) ? 1'b0 : 1'b0;
									assign node3018 = (inp[10]) ? 1'b0 : node3019;
										assign node3019 = (inp[11]) ? 1'b0 : node3020;
											assign node3020 = (inp[3]) ? 1'b0 : 1'b0;
								assign node3025 = (inp[7]) ? 1'b0 : node3026;
									assign node3026 = (inp[10]) ? 1'b0 : node3027;
										assign node3027 = (inp[9]) ? 1'b0 : node3028;
											assign node3028 = (inp[0]) ? 1'b0 : 1'b0;
					assign node3034 = (inp[12]) ? node3118 : node3035;
						assign node3035 = (inp[9]) ? node3087 : node3036;
							assign node3036 = (inp[5]) ? node3066 : node3037;
								assign node3037 = (inp[0]) ? node3053 : node3038;
									assign node3038 = (inp[10]) ? node3046 : node3039;
										assign node3039 = (inp[1]) ? node3043 : node3040;
											assign node3040 = (inp[3]) ? 1'b1 : 1'b1;
											assign node3043 = (inp[4]) ? 1'b0 : 1'b1;
										assign node3046 = (inp[11]) ? node3050 : node3047;
											assign node3047 = (inp[7]) ? 1'b0 : 1'b1;
											assign node3050 = (inp[4]) ? 1'b0 : 1'b0;
									assign node3053 = (inp[1]) ? node3061 : node3054;
										assign node3054 = (inp[3]) ? node3058 : node3055;
											assign node3055 = (inp[8]) ? 1'b0 : 1'b1;
											assign node3058 = (inp[11]) ? 1'b0 : 1'b0;
										assign node3061 = (inp[8]) ? 1'b0 : node3062;
											assign node3062 = (inp[7]) ? 1'b0 : 1'b0;
								assign node3066 = (inp[8]) ? node3080 : node3067;
									assign node3067 = (inp[1]) ? node3075 : node3068;
										assign node3068 = (inp[0]) ? node3072 : node3069;
											assign node3069 = (inp[10]) ? 1'b0 : 1'b1;
											assign node3072 = (inp[4]) ? 1'b0 : 1'b0;
										assign node3075 = (inp[11]) ? 1'b0 : node3076;
											assign node3076 = (inp[0]) ? 1'b0 : 1'b0;
									assign node3080 = (inp[11]) ? 1'b0 : node3081;
										assign node3081 = (inp[10]) ? 1'b0 : node3082;
											assign node3082 = (inp[3]) ? 1'b0 : 1'b0;
							assign node3087 = (inp[5]) ? node3109 : node3088;
								assign node3088 = (inp[0]) ? node3102 : node3089;
									assign node3089 = (inp[10]) ? node3097 : node3090;
										assign node3090 = (inp[8]) ? node3094 : node3091;
											assign node3091 = (inp[11]) ? 1'b0 : 1'b1;
											assign node3094 = (inp[11]) ? 1'b0 : 1'b0;
										assign node3097 = (inp[7]) ? 1'b0 : node3098;
											assign node3098 = (inp[11]) ? 1'b0 : 1'b0;
									assign node3102 = (inp[1]) ? 1'b0 : node3103;
										assign node3103 = (inp[7]) ? 1'b0 : node3104;
											assign node3104 = (inp[3]) ? 1'b0 : 1'b0;
								assign node3109 = (inp[8]) ? 1'b0 : node3110;
									assign node3110 = (inp[3]) ? 1'b0 : node3111;
										assign node3111 = (inp[10]) ? 1'b0 : node3112;
											assign node3112 = (inp[1]) ? 1'b0 : 1'b0;
						assign node3118 = (inp[3]) ? node3150 : node3119;
							assign node3119 = (inp[5]) ? node3141 : node3120;
								assign node3120 = (inp[7]) ? node3134 : node3121;
									assign node3121 = (inp[10]) ? node3129 : node3122;
										assign node3122 = (inp[4]) ? node3126 : node3123;
											assign node3123 = (inp[8]) ? 1'b0 : 1'b1;
											assign node3126 = (inp[11]) ? 1'b0 : 1'b0;
										assign node3129 = (inp[0]) ? 1'b0 : node3130;
											assign node3130 = (inp[1]) ? 1'b0 : 1'b0;
									assign node3134 = (inp[1]) ? 1'b0 : node3135;
										assign node3135 = (inp[11]) ? 1'b0 : node3136;
											assign node3136 = (inp[0]) ? 1'b0 : 1'b0;
								assign node3141 = (inp[10]) ? 1'b0 : node3142;
									assign node3142 = (inp[1]) ? 1'b0 : node3143;
										assign node3143 = (inp[0]) ? 1'b0 : node3144;
											assign node3144 = (inp[8]) ? 1'b0 : 1'b0;
							assign node3150 = (inp[1]) ? 1'b0 : node3151;
								assign node3151 = (inp[0]) ? 1'b0 : node3152;
									assign node3152 = (inp[8]) ? 1'b0 : node3153;
										assign node3153 = (inp[7]) ? 1'b0 : node3154;
											assign node3154 = (inp[10]) ? 1'b0 : 1'b0;

endmodule