module dtc_split5_bm50 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node5;
	wire [2-1:0] node9;
	wire [2-1:0] node10;
	wire [2-1:0] node14;
	wire [2-1:0] node15;
	wire [2-1:0] node16;
	wire [2-1:0] node19;
	wire [2-1:0] node22;
	wire [2-1:0] node23;
	wire [2-1:0] node26;
	wire [2-1:0] node29;
	wire [2-1:0] node30;
	wire [2-1:0] node31;
	wire [2-1:0] node32;
	wire [2-1:0] node36;
	wire [2-1:0] node37;
	wire [2-1:0] node40;
	wire [2-1:0] node43;
	wire [2-1:0] node44;
	wire [2-1:0] node45;
	wire [2-1:0] node49;
	wire [2-1:0] node50;
	wire [2-1:0] node53;
	wire [2-1:0] node56;
	wire [2-1:0] node57;
	wire [2-1:0] node58;
	wire [2-1:0] node59;
	wire [2-1:0] node61;
	wire [2-1:0] node64;
	wire [2-1:0] node66;
	wire [2-1:0] node69;
	wire [2-1:0] node70;
	wire [2-1:0] node71;
	wire [2-1:0] node75;
	wire [2-1:0] node77;
	wire [2-1:0] node80;
	wire [2-1:0] node81;
	wire [2-1:0] node82;
	wire [2-1:0] node84;
	wire [2-1:0] node87;
	wire [2-1:0] node88;
	wire [2-1:0] node91;
	wire [2-1:0] node94;
	wire [2-1:0] node95;
	wire [2-1:0] node96;
	wire [2-1:0] node99;
	wire [2-1:0] node102;
	wire [2-1:0] node103;
	wire [2-1:0] node106;

	assign outp = (inp[5]) ? node56 : node1;
		assign node1 = (inp[1]) ? node29 : node2;
			assign node2 = (inp[4]) ? node14 : node3;
				assign node3 = (inp[3]) ? node9 : node4;
					assign node4 = (inp[6]) ? 2'b11 : node5;
						assign node5 = (inp[2]) ? 2'b11 : 2'b10;
					assign node9 = (inp[0]) ? 2'b01 : node10;
						assign node10 = (inp[2]) ? 2'b01 : 2'b10;
				assign node14 = (inp[7]) ? node22 : node15;
					assign node15 = (inp[0]) ? node19 : node16;
						assign node16 = (inp[2]) ? 2'b00 : 2'b01;
						assign node19 = (inp[6]) ? 2'b01 : 2'b00;
					assign node22 = (inp[0]) ? node26 : node23;
						assign node23 = (inp[2]) ? 2'b01 : 2'b00;
						assign node26 = (inp[6]) ? 2'b00 : 2'b00;
			assign node29 = (inp[3]) ? node43 : node30;
				assign node30 = (inp[4]) ? node36 : node31;
					assign node31 = (inp[6]) ? 2'b00 : node32;
						assign node32 = (inp[2]) ? 2'b00 : 2'b01;
					assign node36 = (inp[7]) ? node40 : node37;
						assign node37 = (inp[0]) ? 2'b00 : 2'b00;
						assign node40 = (inp[0]) ? 2'b10 : 2'b11;
				assign node43 = (inp[7]) ? node49 : node44;
					assign node44 = (inp[4]) ? 2'b10 : node45;
						assign node45 = (inp[2]) ? 2'b00 : 2'b01;
					assign node49 = (inp[0]) ? node53 : node50;
						assign node50 = (inp[6]) ? 2'b11 : 2'b10;
						assign node53 = (inp[2]) ? 2'b10 : 2'b10;
		assign node56 = (inp[0]) ? node80 : node57;
			assign node57 = (inp[7]) ? node69 : node58;
				assign node58 = (inp[1]) ? node64 : node59;
					assign node59 = (inp[4]) ? node61 : 2'b00;
						assign node61 = (inp[3]) ? 2'b10 : 2'b00;
					assign node64 = (inp[3]) ? node66 : 2'b10;
						assign node66 = (inp[4]) ? 2'b00 : 2'b10;
				assign node69 = (inp[2]) ? node75 : node70;
					assign node70 = (inp[6]) ? 2'b11 : node71;
						assign node71 = (inp[3]) ? 2'b10 : 2'b00;
					assign node75 = (inp[1]) ? node77 : 2'b11;
						assign node77 = (inp[3]) ? 2'b01 : 2'b11;
			assign node80 = (inp[7]) ? node94 : node81;
				assign node81 = (inp[6]) ? node87 : node82;
					assign node82 = (inp[2]) ? node84 : 2'b10;
						assign node84 = (inp[4]) ? 2'b11 : 2'b01;
					assign node87 = (inp[1]) ? node91 : node88;
						assign node88 = (inp[3]) ? 2'b11 : 2'b01;
						assign node91 = (inp[4]) ? 2'b01 : 2'b01;
				assign node94 = (inp[6]) ? node102 : node95;
					assign node95 = (inp[2]) ? node99 : node96;
						assign node96 = (inp[1]) ? 2'b01 : 2'b11;
						assign node99 = (inp[4]) ? 2'b00 : 2'b10;
					assign node102 = (inp[1]) ? node106 : node103;
						assign node103 = (inp[3]) ? 2'b10 : 2'b00;
						assign node106 = (inp[3]) ? 2'b00 : 2'b10;

endmodule