module dtc_split05_bm22 (
	input  wire [11-1:0] inp,
	output wire [11-1:0] outp
);

	wire [11-1:0] node1;
	wire [11-1:0] node2;
	wire [11-1:0] node3;
	wire [11-1:0] node4;
	wire [11-1:0] node5;
	wire [11-1:0] node6;
	wire [11-1:0] node8;
	wire [11-1:0] node11;
	wire [11-1:0] node14;
	wire [11-1:0] node15;
	wire [11-1:0] node19;
	wire [11-1:0] node21;
	wire [11-1:0] node23;
	wire [11-1:0] node26;
	wire [11-1:0] node27;
	wire [11-1:0] node28;
	wire [11-1:0] node31;
	wire [11-1:0] node34;
	wire [11-1:0] node35;
	wire [11-1:0] node36;
	wire [11-1:0] node40;
	wire [11-1:0] node42;
	wire [11-1:0] node43;
	wire [11-1:0] node47;
	wire [11-1:0] node48;
	wire [11-1:0] node49;
	wire [11-1:0] node50;
	wire [11-1:0] node54;
	wire [11-1:0] node57;
	wire [11-1:0] node58;
	wire [11-1:0] node60;
	wire [11-1:0] node63;
	wire [11-1:0] node66;
	wire [11-1:0] node67;
	wire [11-1:0] node68;
	wire [11-1:0] node69;
	wire [11-1:0] node70;
	wire [11-1:0] node71;
	wire [11-1:0] node75;
	wire [11-1:0] node78;
	wire [11-1:0] node81;
	wire [11-1:0] node82;
	wire [11-1:0] node83;
	wire [11-1:0] node86;
	wire [11-1:0] node87;
	wire [11-1:0] node91;
	wire [11-1:0] node92;
	wire [11-1:0] node93;
	wire [11-1:0] node97;
	wire [11-1:0] node99;
	wire [11-1:0] node102;
	wire [11-1:0] node103;
	wire [11-1:0] node104;
	wire [11-1:0] node107;
	wire [11-1:0] node108;
	wire [11-1:0] node111;
	wire [11-1:0] node114;
	wire [11-1:0] node115;
	wire [11-1:0] node116;
	wire [11-1:0] node117;
	wire [11-1:0] node119;
	wire [11-1:0] node123;
	wire [11-1:0] node125;
	wire [11-1:0] node128;

	assign outp = (inp[4]) ? node66 : node1;
		assign node1 = (inp[1]) ? node47 : node2;
			assign node2 = (inp[5]) ? node26 : node3;
				assign node3 = (inp[9]) ? node19 : node4;
					assign node4 = (inp[7]) ? node14 : node5;
						assign node5 = (inp[6]) ? node11 : node6;
							assign node6 = (inp[3]) ? node8 : 11'b01111111111;
								assign node8 = (inp[0]) ? 11'b00111111111 : 11'b01111111111;
							assign node11 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
						assign node14 = (inp[10]) ? 11'b00001111111 : node15;
							assign node15 = (inp[8]) ? 11'b00001111111 : 11'b00011111111;
					assign node19 = (inp[7]) ? node21 : 11'b00001111111;
						assign node21 = (inp[6]) ? node23 : 11'b00000111111;
							assign node23 = (inp[8]) ? 11'b00000111111 : 11'b00001111111;
				assign node26 = (inp[3]) ? node34 : node27;
					assign node27 = (inp[7]) ? node31 : node28;
						assign node28 = (inp[0]) ? 11'b00001111111 : 11'b00011111111;
						assign node31 = (inp[6]) ? 11'b00001111111 : 11'b00000111111;
					assign node34 = (inp[10]) ? node40 : node35;
						assign node35 = (inp[8]) ? 11'b00000111111 : node36;
							assign node36 = (inp[6]) ? 11'b00000111111 : 11'b00011111111;
						assign node40 = (inp[0]) ? node42 : 11'b00001111111;
							assign node42 = (inp[7]) ? 11'b00000011111 : node43;
								assign node43 = (inp[2]) ? 11'b00000011111 : 11'b00000111111;
			assign node47 = (inp[10]) ? node57 : node48;
				assign node48 = (inp[0]) ? node54 : node49;
					assign node49 = (inp[6]) ? 11'b00000111111 : node50;
						assign node50 = (inp[5]) ? 11'b00011111111 : 11'b00001111111;
					assign node54 = (inp[9]) ? 11'b00000001111 : 11'b00000111111;
				assign node57 = (inp[6]) ? node63 : node58;
					assign node58 = (inp[0]) ? node60 : 11'b00000111111;
						assign node60 = (inp[7]) ? 11'b00000011111 : 11'b00000001111;
					assign node63 = (inp[8]) ? 11'b00000001111 : 11'b00000000111;
		assign node66 = (inp[2]) ? node102 : node67;
			assign node67 = (inp[3]) ? node81 : node68;
				assign node68 = (inp[7]) ? node78 : node69;
					assign node69 = (inp[1]) ? node75 : node70;
						assign node70 = (inp[10]) ? 11'b00001111111 : node71;
							assign node71 = (inp[8]) ? 11'b00001111111 : 11'b00111111111;
						assign node75 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
					assign node78 = (inp[5]) ? 11'b00000001111 : 11'b00000111111;
				assign node81 = (inp[1]) ? node91 : node82;
					assign node82 = (inp[10]) ? node86 : node83;
						assign node83 = (inp[6]) ? 11'b00000011111 : 11'b00000111111;
						assign node86 = (inp[7]) ? 11'b00000000111 : node87;
							assign node87 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
					assign node91 = (inp[5]) ? node97 : node92;
						assign node92 = (inp[0]) ? 11'b00000001111 : node93;
							assign node93 = (inp[9]) ? 11'b00000011111 : 11'b00000111111;
						assign node97 = (inp[8]) ? node99 : 11'b00000001111;
							assign node99 = (inp[6]) ? 11'b00000000111 : 11'b00000000011;
			assign node102 = (inp[9]) ? node114 : node103;
				assign node103 = (inp[5]) ? node107 : node104;
					assign node104 = (inp[10]) ? 11'b00000011111 : 11'b00000111111;
					assign node107 = (inp[1]) ? node111 : node108;
						assign node108 = (inp[7]) ? 11'b00000001111 : 11'b00000011111;
						assign node111 = (inp[0]) ? 11'b00000000111 : 11'b00000001111;
				assign node114 = (inp[7]) ? node128 : node115;
					assign node115 = (inp[3]) ? node123 : node116;
						assign node116 = (inp[0]) ? 11'b00000001111 : node117;
							assign node117 = (inp[10]) ? node119 : 11'b00000011111;
								assign node119 = (inp[6]) ? 11'b00000001111 : 11'b00000011111;
						assign node123 = (inp[1]) ? node125 : 11'b00000001111;
							assign node125 = (inp[6]) ? 11'b00000000011 : 11'b00000001111;
					assign node128 = (inp[10]) ? 11'b00000000111 : 11'b00000001111;

endmodule