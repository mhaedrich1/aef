module dtc_split25_bm89 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node263;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node274;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node412;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node486;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node502;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node532;
	wire [3-1:0] node534;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node606;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node636;
	wire [3-1:0] node639;
	wire [3-1:0] node641;
	wire [3-1:0] node643;
	wire [3-1:0] node646;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;

	assign outp = (inp[6]) ? node382 : node1;
		assign node1 = (inp[3]) ? node185 : node2;
			assign node2 = (inp[7]) ? node48 : node3;
				assign node3 = (inp[9]) ? 3'b111 : node4;
					assign node4 = (inp[4]) ? node16 : node5;
						assign node5 = (inp[10]) ? 3'b111 : node6;
							assign node6 = (inp[11]) ? node10 : node7;
								assign node7 = (inp[5]) ? 3'b011 : 3'b101;
								assign node10 = (inp[5]) ? 3'b101 : node11;
									assign node11 = (inp[2]) ? 3'b011 : 3'b101;
						assign node16 = (inp[10]) ? node30 : node17;
							assign node17 = (inp[11]) ? node21 : node18;
								assign node18 = (inp[8]) ? 3'b100 : 3'b010;
								assign node21 = (inp[2]) ? node25 : node22;
									assign node22 = (inp[5]) ? 3'b110 : 3'b001;
									assign node25 = (inp[1]) ? node27 : 3'b110;
										assign node27 = (inp[8]) ? 3'b010 : 3'b110;
							assign node30 = (inp[8]) ? node38 : node31;
								assign node31 = (inp[11]) ? 3'b011 : node32;
									assign node32 = (inp[1]) ? node34 : 3'b101;
										assign node34 = (inp[2]) ? 3'b001 : 3'b101;
								assign node38 = (inp[11]) ? node44 : node39;
									assign node39 = (inp[1]) ? node41 : 3'b001;
										assign node41 = (inp[2]) ? 3'b110 : 3'b001;
									assign node44 = (inp[5]) ? 3'b001 : 3'b101;
				assign node48 = (inp[10]) ? node122 : node49;
					assign node49 = (inp[5]) ? node93 : node50;
						assign node50 = (inp[4]) ? node74 : node51;
							assign node51 = (inp[11]) ? node61 : node52;
								assign node52 = (inp[2]) ? node54 : 3'b110;
									assign node54 = (inp[8]) ? 3'b010 : node55;
										assign node55 = (inp[9]) ? 3'b110 : node56;
											assign node56 = (inp[0]) ? 3'b110 : 3'b010;
								assign node61 = (inp[9]) ? node69 : node62;
									assign node62 = (inp[2]) ? node66 : node63;
										assign node63 = (inp[8]) ? 3'b001 : 3'b011;
										assign node66 = (inp[8]) ? 3'b101 : 3'b111;
									assign node69 = (inp[8]) ? node71 : 3'b110;
										assign node71 = (inp[0]) ? 3'b110 : 3'b000;
							assign node74 = (inp[9]) ? node86 : node75;
								assign node75 = (inp[0]) ? node81 : node76;
									assign node76 = (inp[11]) ? node78 : 3'b100;
										assign node78 = (inp[1]) ? 3'b100 : 3'b000;
									assign node81 = (inp[8]) ? node83 : 3'b010;
										assign node83 = (inp[11]) ? 3'b100 : 3'b000;
								assign node86 = (inp[8]) ? node88 : 3'b101;
									assign node88 = (inp[11]) ? node90 : 3'b111;
										assign node90 = (inp[0]) ? 3'b100 : 3'b110;
						assign node93 = (inp[4]) ? node107 : node94;
							assign node94 = (inp[11]) ? node102 : node95;
								assign node95 = (inp[9]) ? 3'b000 : node96;
									assign node96 = (inp[8]) ? 3'b000 : node97;
										assign node97 = (inp[0]) ? 3'b010 : 3'b110;
								assign node102 = (inp[8]) ? 3'b110 : node103;
									assign node103 = (inp[1]) ? 3'b110 : 3'b000;
							assign node107 = (inp[9]) ? node119 : node108;
								assign node108 = (inp[8]) ? node112 : node109;
									assign node109 = (inp[1]) ? 3'b000 : 3'b010;
									assign node112 = (inp[0]) ? 3'b000 : node113;
										assign node113 = (inp[1]) ? node115 : 3'b100;
											assign node115 = (inp[2]) ? 3'b000 : 3'b100;
								assign node119 = (inp[1]) ? 3'b001 : 3'b101;
					assign node122 = (inp[4]) ? node146 : node123;
						assign node123 = (inp[9]) ? 3'b100 : node124;
							assign node124 = (inp[11]) ? node132 : node125;
								assign node125 = (inp[2]) ? node127 : 3'b101;
									assign node127 = (inp[5]) ? 3'b010 : node128;
										assign node128 = (inp[8]) ? 3'b001 : 3'b101;
								assign node132 = (inp[5]) ? node140 : node133;
									assign node133 = (inp[8]) ? node137 : node134;
										assign node134 = (inp[2]) ? 3'b011 : 3'b001;
										assign node137 = (inp[2]) ? 3'b111 : 3'b011;
									assign node140 = (inp[0]) ? node142 : 3'b011;
										assign node142 = (inp[2]) ? 3'b101 : 3'b111;
						assign node146 = (inp[9]) ? node168 : node147;
							assign node147 = (inp[11]) ? node157 : node148;
								assign node148 = (inp[8]) ? node154 : node149;
									assign node149 = (inp[0]) ? node151 : 3'b110;
										assign node151 = (inp[5]) ? 3'b010 : 3'b110;
									assign node154 = (inp[2]) ? 3'b100 : 3'b010;
								assign node157 = (inp[8]) ? node163 : node158;
									assign node158 = (inp[5]) ? node160 : 3'b001;
										assign node160 = (inp[0]) ? 3'b110 : 3'b001;
									assign node163 = (inp[1]) ? node165 : 3'b110;
										assign node165 = (inp[5]) ? 3'b110 : 3'b010;
							assign node168 = (inp[8]) ? node176 : node169;
								assign node169 = (inp[11]) ? 3'b001 : node170;
									assign node170 = (inp[5]) ? 3'b011 : node171;
										assign node171 = (inp[0]) ? 3'b111 : 3'b011;
								assign node176 = (inp[1]) ? node182 : node177;
									assign node177 = (inp[0]) ? node179 : 3'b011;
										assign node179 = (inp[5]) ? 3'b101 : 3'b011;
									assign node182 = (inp[11]) ? 3'b111 : 3'b101;
			assign node185 = (inp[9]) ? node267 : node186;
				assign node186 = (inp[7]) ? node248 : node187;
					assign node187 = (inp[4]) ? node243 : node188;
						assign node188 = (inp[10]) ? node210 : node189;
							assign node189 = (inp[11]) ? node197 : node190;
								assign node190 = (inp[8]) ? 3'b000 : node191;
									assign node191 = (inp[5]) ? node193 : 3'b100;
										assign node193 = (inp[0]) ? 3'b000 : 3'b100;
								assign node197 = (inp[8]) ? node205 : node198;
									assign node198 = (inp[1]) ? node200 : 3'b010;
										assign node200 = (inp[5]) ? node202 : 3'b010;
											assign node202 = (inp[0]) ? 3'b100 : 3'b010;
									assign node205 = (inp[5]) ? 3'b100 : node206;
										assign node206 = (inp[1]) ? 3'b010 : 3'b110;
							assign node210 = (inp[11]) ? node230 : node211;
								assign node211 = (inp[1]) ? node221 : node212;
									assign node212 = (inp[5]) ? node218 : node213;
										assign node213 = (inp[2]) ? node215 : 3'b110;
											assign node215 = (inp[8]) ? 3'b010 : 3'b110;
										assign node218 = (inp[8]) ? 3'b000 : 3'b110;
									assign node221 = (inp[2]) ? node225 : node222;
										assign node222 = (inp[0]) ? 3'b010 : 3'b110;
										assign node225 = (inp[5]) ? node227 : 3'b010;
											assign node227 = (inp[8]) ? 3'b000 : 3'b010;
								assign node230 = (inp[5]) ? node238 : node231;
									assign node231 = (inp[0]) ? node235 : node232;
										assign node232 = (inp[8]) ? 3'b101 : 3'b111;
										assign node235 = (inp[1]) ? 3'b011 : 3'b001;
									assign node238 = (inp[8]) ? 3'b110 : node239;
										assign node239 = (inp[1]) ? 3'b110 : 3'b011;
						assign node243 = (inp[11]) ? node245 : 3'b000;
							assign node245 = (inp[10]) ? 3'b100 : 3'b000;
					assign node248 = (inp[10]) ? node250 : 3'b000;
						assign node250 = (inp[4]) ? 3'b000 : node251;
							assign node251 = (inp[11]) ? node261 : node252;
								assign node252 = (inp[8]) ? node256 : node253;
									assign node253 = (inp[0]) ? 3'b000 : 3'b100;
									assign node256 = (inp[0]) ? node258 : 3'b000;
										assign node258 = (inp[2]) ? 3'b000 : 3'b100;
								assign node261 = (inp[2]) ? node263 : 3'b000;
									assign node263 = (inp[1]) ? 3'b100 : 3'b010;
				assign node267 = (inp[4]) ? node327 : node268;
					assign node268 = (inp[7]) ? node288 : node269;
						assign node269 = (inp[10]) ? 3'b111 : node270;
							assign node270 = (inp[11]) ? node278 : node271;
								assign node271 = (inp[5]) ? 3'b011 : node272;
									assign node272 = (inp[8]) ? node274 : 3'b101;
										assign node274 = (inp[0]) ? 3'b011 : 3'b101;
								assign node278 = (inp[2]) ? node282 : node279;
									assign node279 = (inp[0]) ? 3'b101 : 3'b011;
									assign node282 = (inp[0]) ? 3'b011 : node283;
										assign node283 = (inp[8]) ? 3'b011 : 3'b101;
						assign node288 = (inp[10]) ? node312 : node289;
							assign node289 = (inp[11]) ? node301 : node290;
								assign node290 = (inp[5]) ? node296 : node291;
									assign node291 = (inp[0]) ? 3'b110 : node292;
										assign node292 = (inp[8]) ? 3'b110 : 3'b010;
									assign node296 = (inp[8]) ? node298 : 3'b010;
										assign node298 = (inp[2]) ? 3'b100 : 3'b000;
								assign node301 = (inp[8]) ? node309 : node302;
									assign node302 = (inp[1]) ? node306 : node303;
										assign node303 = (inp[5]) ? 3'b001 : 3'b011;
										assign node306 = (inp[2]) ? 3'b001 : 3'b100;
									assign node309 = (inp[0]) ? 3'b110 : 3'b001;
							assign node312 = (inp[8]) ? node318 : node313;
								assign node313 = (inp[1]) ? 3'b001 : node314;
									assign node314 = (inp[2]) ? 3'b001 : 3'b101;
								assign node318 = (inp[5]) ? node324 : node319;
									assign node319 = (inp[11]) ? node321 : 3'b101;
										assign node321 = (inp[2]) ? 3'b111 : 3'b011;
									assign node324 = (inp[0]) ? 3'b110 : 3'b010;
					assign node327 = (inp[10]) ? node351 : node328;
						assign node328 = (inp[7]) ? node338 : node329;
							assign node329 = (inp[11]) ? node333 : node330;
								assign node330 = (inp[8]) ? 3'b100 : 3'b010;
								assign node333 = (inp[8]) ? node335 : 3'b110;
									assign node335 = (inp[1]) ? 3'b010 : 3'b110;
							assign node338 = (inp[0]) ? node348 : node339;
								assign node339 = (inp[8]) ? 3'b100 : node340;
									assign node340 = (inp[2]) ? node344 : node341;
										assign node341 = (inp[11]) ? 3'b100 : 3'b000;
										assign node344 = (inp[1]) ? 3'b100 : 3'b010;
								assign node348 = (inp[8]) ? 3'b000 : 3'b010;
						assign node351 = (inp[7]) ? node365 : node352;
							assign node352 = (inp[2]) ? node360 : node353;
								assign node353 = (inp[11]) ? 3'b101 : node354;
									assign node354 = (inp[0]) ? 3'b001 : node355;
										assign node355 = (inp[8]) ? 3'b001 : 3'b101;
								assign node360 = (inp[8]) ? 3'b110 : node361;
									assign node361 = (inp[0]) ? 3'b101 : 3'b011;
							assign node365 = (inp[5]) ? node373 : node366;
								assign node366 = (inp[11]) ? node368 : 3'b010;
									assign node368 = (inp[8]) ? node370 : 3'b001;
										assign node370 = (inp[2]) ? 3'b010 : 3'b001;
								assign node373 = (inp[2]) ? node375 : 3'b110;
									assign node375 = (inp[1]) ? 3'b010 : node376;
										assign node376 = (inp[11]) ? 3'b110 : node377;
											assign node377 = (inp[8]) ? 3'b010 : 3'b010;
		assign node382 = (inp[9]) ? node460 : node383;
			assign node383 = (inp[3]) ? 3'b000 : node384;
				assign node384 = (inp[10]) ? node406 : node385;
					assign node385 = (inp[7]) ? 3'b000 : node386;
						assign node386 = (inp[4]) ? 3'b000 : node387;
							assign node387 = (inp[11]) ? node393 : node388;
								assign node388 = (inp[8]) ? 3'b000 : node389;
									assign node389 = (inp[0]) ? 3'b000 : 3'b100;
								assign node393 = (inp[5]) ? node397 : node394;
									assign node394 = (inp[8]) ? 3'b010 : 3'b110;
									assign node397 = (inp[8]) ? node399 : 3'b010;
										assign node399 = (inp[0]) ? node401 : 3'b100;
											assign node401 = (inp[2]) ? 3'b000 : 3'b100;
					assign node406 = (inp[7]) ? node444 : node407;
						assign node407 = (inp[11]) ? node427 : node408;
							assign node408 = (inp[8]) ? node418 : node409;
								assign node409 = (inp[4]) ? node415 : node410;
									assign node410 = (inp[2]) ? node412 : 3'b110;
										assign node412 = (inp[0]) ? 3'b110 : 3'b010;
									assign node415 = (inp[0]) ? 3'b000 : 3'b100;
								assign node418 = (inp[1]) ? 3'b100 : node419;
									assign node419 = (inp[2]) ? node421 : 3'b000;
										assign node421 = (inp[4]) ? 3'b000 : node422;
											assign node422 = (inp[5]) ? 3'b000 : 3'b010;
							assign node427 = (inp[4]) ? node441 : node428;
								assign node428 = (inp[8]) ? node438 : node429;
									assign node429 = (inp[0]) ? node435 : node430;
										assign node430 = (inp[5]) ? node432 : 3'b111;
											assign node432 = (inp[2]) ? 3'b011 : 3'b001;
										assign node435 = (inp[1]) ? 3'b110 : 3'b001;
									assign node438 = (inp[0]) ? 3'b110 : 3'b101;
								assign node441 = (inp[0]) ? 3'b010 : 3'b110;
						assign node444 = (inp[4]) ? 3'b000 : node445;
							assign node445 = (inp[11]) ? node451 : node446;
								assign node446 = (inp[2]) ? 3'b000 : node447;
									assign node447 = (inp[0]) ? 3'b000 : 3'b100;
								assign node451 = (inp[5]) ? 3'b100 : node452;
									assign node452 = (inp[8]) ? 3'b010 : node453;
										assign node453 = (inp[2]) ? 3'b010 : 3'b110;
			assign node460 = (inp[3]) ? node576 : node461;
				assign node461 = (inp[10]) ? node519 : node462;
					assign node462 = (inp[4]) ? node498 : node463;
						assign node463 = (inp[7]) ? node479 : node464;
							assign node464 = (inp[8]) ? node474 : node465;
								assign node465 = (inp[5]) ? node469 : node466;
									assign node466 = (inp[2]) ? 3'b011 : 3'b001;
									assign node469 = (inp[2]) ? node471 : 3'b011;
										assign node471 = (inp[11]) ? 3'b001 : 3'b011;
								assign node474 = (inp[5]) ? 3'b001 : node475;
									assign node475 = (inp[11]) ? 3'b011 : 3'b001;
							assign node479 = (inp[11]) ? node489 : node480;
								assign node480 = (inp[5]) ? node482 : 3'b010;
									assign node482 = (inp[8]) ? node484 : 3'b110;
										assign node484 = (inp[2]) ? node486 : 3'b000;
											assign node486 = (inp[1]) ? 3'b100 : 3'b000;
								assign node489 = (inp[5]) ? node493 : node490;
									assign node490 = (inp[2]) ? 3'b101 : 3'b001;
									assign node493 = (inp[8]) ? 3'b110 : node494;
										assign node494 = (inp[2]) ? 3'b011 : 3'b001;
						assign node498 = (inp[8]) ? node508 : node499;
							assign node499 = (inp[11]) ? node505 : node500;
								assign node500 = (inp[7]) ? node502 : 3'b010;
									assign node502 = (inp[5]) ? 3'b000 : 3'b010;
								assign node505 = (inp[7]) ? 3'b010 : 3'b110;
							assign node508 = (inp[11]) ? node512 : node509;
								assign node509 = (inp[7]) ? 3'b000 : 3'b100;
								assign node512 = (inp[7]) ? node516 : node513;
									assign node513 = (inp[1]) ? 3'b010 : 3'b110;
									assign node516 = (inp[1]) ? 3'b100 : 3'b110;
					assign node519 = (inp[4]) ? node537 : node520;
						assign node520 = (inp[5]) ? node526 : node521;
							assign node521 = (inp[11]) ? 3'b011 : node522;
								assign node522 = (inp[7]) ? 3'b001 : 3'b011;
							assign node526 = (inp[11]) ? node532 : node527;
								assign node527 = (inp[8]) ? 3'b110 : node528;
									assign node528 = (inp[7]) ? 3'b111 : 3'b011;
								assign node532 = (inp[2]) ? node534 : 3'b101;
									assign node534 = (inp[1]) ? 3'b001 : 3'b011;
						assign node537 = (inp[7]) ? node563 : node538;
							assign node538 = (inp[1]) ? node550 : node539;
								assign node539 = (inp[8]) ? node541 : 3'b101;
									assign node541 = (inp[0]) ? node543 : 3'b001;
										assign node543 = (inp[2]) ? node547 : node544;
											assign node544 = (inp[11]) ? 3'b001 : 3'b000;
											assign node547 = (inp[5]) ? 3'b001 : 3'b001;
								assign node550 = (inp[11]) ? node556 : node551;
									assign node551 = (inp[0]) ? 3'b110 : node552;
										assign node552 = (inp[5]) ? 3'b101 : 3'b001;
									assign node556 = (inp[8]) ? node560 : node557;
										assign node557 = (inp[5]) ? 3'b101 : 3'b011;
										assign node560 = (inp[5]) ? 3'b001 : 3'b101;
							assign node563 = (inp[11]) ? node571 : node564;
								assign node564 = (inp[8]) ? node566 : 3'b110;
									assign node566 = (inp[0]) ? 3'b010 : node567;
										assign node567 = (inp[5]) ? 3'b010 : 3'b110;
								assign node571 = (inp[5]) ? node573 : 3'b001;
									assign node573 = (inp[1]) ? 3'b101 : 3'b110;
				assign node576 = (inp[7]) ? node646 : node577;
					assign node577 = (inp[10]) ? node599 : node578;
						assign node578 = (inp[4]) ? 3'b000 : node579;
							assign node579 = (inp[11]) ? node585 : node580;
								assign node580 = (inp[8]) ? 3'b000 : node581;
									assign node581 = (inp[1]) ? 3'b000 : 3'b100;
								assign node585 = (inp[8]) ? node595 : node586;
									assign node586 = (inp[2]) ? node592 : node587;
										assign node587 = (inp[0]) ? 3'b100 : node588;
											assign node588 = (inp[5]) ? 3'b010 : 3'b110;
										assign node592 = (inp[0]) ? 3'b010 : 3'b110;
									assign node595 = (inp[2]) ? 3'b100 : 3'b010;
						assign node599 = (inp[5]) ? node625 : node600;
							assign node600 = (inp[0]) ? node614 : node601;
								assign node601 = (inp[8]) ? node609 : node602;
									assign node602 = (inp[4]) ? node606 : node603;
										assign node603 = (inp[1]) ? 3'b111 : 3'b010;
										assign node606 = (inp[11]) ? 3'b110 : 3'b100;
									assign node609 = (inp[11]) ? 3'b010 : node610;
										assign node610 = (inp[2]) ? 3'b010 : 3'b110;
								assign node614 = (inp[11]) ? node618 : node615;
									assign node615 = (inp[4]) ? 3'b000 : 3'b010;
									assign node618 = (inp[4]) ? 3'b010 : node619;
										assign node619 = (inp[8]) ? 3'b001 : node620;
											assign node620 = (inp[2]) ? 3'b001 : 3'b011;
							assign node625 = (inp[4]) ? node639 : node626;
								assign node626 = (inp[2]) ? node636 : node627;
									assign node627 = (inp[11]) ? node631 : node628;
										assign node628 = (inp[0]) ? 3'b010 : 3'b110;
										assign node631 = (inp[8]) ? 3'b110 : node632;
											assign node632 = (inp[1]) ? 3'b100 : 3'b001;
									assign node636 = (inp[0]) ? 3'b100 : 3'b000;
								assign node639 = (inp[1]) ? node641 : 3'b100;
									assign node641 = (inp[11]) ? node643 : 3'b000;
										assign node643 = (inp[2]) ? 3'b000 : 3'b100;
					assign node646 = (inp[10]) ? node648 : 3'b000;
						assign node648 = (inp[4]) ? node656 : node649;
							assign node649 = (inp[11]) ? node653 : node650;
								assign node650 = (inp[5]) ? 3'b000 : 3'b100;
								assign node653 = (inp[5]) ? 3'b100 : 3'b110;
							assign node656 = (inp[5]) ? 3'b000 : node657;
								assign node657 = (inp[8]) ? 3'b000 : node658;
									assign node658 = (inp[11]) ? 3'b100 : 3'b000;

endmodule