module dtc_split5_bm48 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node6;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node13;
	wire [14-1:0] node14;
	wire [14-1:0] node20;
	wire [14-1:0] node21;
	wire [14-1:0] node22;
	wire [14-1:0] node23;
	wire [14-1:0] node26;
	wire [14-1:0] node28;
	wire [14-1:0] node29;
	wire [14-1:0] node33;
	wire [14-1:0] node35;
	wire [14-1:0] node37;
	wire [14-1:0] node40;
	wire [14-1:0] node42;
	wire [14-1:0] node44;
	wire [14-1:0] node45;
	wire [14-1:0] node49;
	wire [14-1:0] node50;
	wire [14-1:0] node51;
	wire [14-1:0] node52;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node55;
	wire [14-1:0] node57;
	wire [14-1:0] node59;
	wire [14-1:0] node62;
	wire [14-1:0] node63;
	wire [14-1:0] node67;
	wire [14-1:0] node68;
	wire [14-1:0] node69;
	wire [14-1:0] node75;
	wire [14-1:0] node77;
	wire [14-1:0] node78;
	wire [14-1:0] node80;
	wire [14-1:0] node85;
	wire [14-1:0] node86;
	wire [14-1:0] node88;
	wire [14-1:0] node89;
	wire [14-1:0] node90;
	wire [14-1:0] node91;
	wire [14-1:0] node93;
	wire [14-1:0] node96;
	wire [14-1:0] node97;
	wire [14-1:0] node101;
	wire [14-1:0] node102;
	wire [14-1:0] node103;
	wire [14-1:0] node104;
	wire [14-1:0] node111;
	wire [14-1:0] node112;
	wire [14-1:0] node114;
	wire [14-1:0] node115;
	wire [14-1:0] node116;
	wire [14-1:0] node117;
	wire [14-1:0] node123;
	wire [14-1:0] node124;
	wire [14-1:0] node128;
	wire [14-1:0] node129;
	wire [14-1:0] node131;
	wire [14-1:0] node132;
	wire [14-1:0] node133;
	wire [14-1:0] node135;
	wire [14-1:0] node136;
	wire [14-1:0] node138;
	wire [14-1:0] node139;
	wire [14-1:0] node144;
	wire [14-1:0] node146;
	wire [14-1:0] node147;
	wire [14-1:0] node148;
	wire [14-1:0] node150;
	wire [14-1:0] node152;
	wire [14-1:0] node155;
	wire [14-1:0] node156;
	wire [14-1:0] node157;
	wire [14-1:0] node159;
	wire [14-1:0] node164;
	wire [14-1:0] node166;
	wire [14-1:0] node168;
	wire [14-1:0] node171;
	wire [14-1:0] node172;
	wire [14-1:0] node173;
	wire [14-1:0] node175;
	wire [14-1:0] node176;
	wire [14-1:0] node179;
	wire [14-1:0] node180;
	wire [14-1:0] node185;
	wire [14-1:0] node186;
	wire [14-1:0] node187;
	wire [14-1:0] node188;
	wire [14-1:0] node193;
	wire [14-1:0] node195;
	wire [14-1:0] node196;
	wire [14-1:0] node200;
	wire [14-1:0] node201;
	wire [14-1:0] node202;
	wire [14-1:0] node204;
	wire [14-1:0] node206;
	wire [14-1:0] node209;
	wire [14-1:0] node210;
	wire [14-1:0] node211;
	wire [14-1:0] node214;
	wire [14-1:0] node215;
	wire [14-1:0] node216;
	wire [14-1:0] node218;
	wire [14-1:0] node223;
	wire [14-1:0] node224;
	wire [14-1:0] node225;
	wire [14-1:0] node227;
	wire [14-1:0] node228;
	wire [14-1:0] node234;
	wire [14-1:0] node235;
	wire [14-1:0] node237;
	wire [14-1:0] node239;
	wire [14-1:0] node240;
	wire [14-1:0] node241;
	wire [14-1:0] node242;
	wire [14-1:0] node248;
	wire [14-1:0] node249;
	wire [14-1:0] node250;
	wire [14-1:0] node251;
	wire [14-1:0] node253;
	wire [14-1:0] node254;
	wire [14-1:0] node259;
	wire [14-1:0] node260;
	wire [14-1:0] node261;
	wire [14-1:0] node263;
	wire [14-1:0] node265;
	wire [14-1:0] node266;
	wire [14-1:0] node272;
	wire [14-1:0] node273;
	wire [14-1:0] node275;
	wire [14-1:0] node276;
	wire [14-1:0] node280;
	wire [14-1:0] node282;
	wire [14-1:0] node284;
	wire [14-1:0] node287;
	wire [14-1:0] node288;
	wire [14-1:0] node289;
	wire [14-1:0] node291;
	wire [14-1:0] node292;
	wire [14-1:0] node293;
	wire [14-1:0] node294;
	wire [14-1:0] node296;
	wire [14-1:0] node301;
	wire [14-1:0] node302;
	wire [14-1:0] node304;
	wire [14-1:0] node306;
	wire [14-1:0] node307;
	wire [14-1:0] node308;
	wire [14-1:0] node314;
	wire [14-1:0] node315;
	wire [14-1:0] node316;
	wire [14-1:0] node317;
	wire [14-1:0] node318;
	wire [14-1:0] node321;
	wire [14-1:0] node322;
	wire [14-1:0] node323;
	wire [14-1:0] node324;
	wire [14-1:0] node330;
	wire [14-1:0] node331;
	wire [14-1:0] node332;
	wire [14-1:0] node333;
	wire [14-1:0] node335;
	wire [14-1:0] node337;
	wire [14-1:0] node339;
	wire [14-1:0] node342;
	wire [14-1:0] node344;
	wire [14-1:0] node349;
	wire [14-1:0] node351;
	wire [14-1:0] node352;
	wire [14-1:0] node353;
	wire [14-1:0] node355;
	wire [14-1:0] node356;
	wire [14-1:0] node359;
	wire [14-1:0] node364;
	wire [14-1:0] node366;
	wire [14-1:0] node368;
	wire [14-1:0] node370;
	wire [14-1:0] node371;
	wire [14-1:0] node372;
	wire [14-1:0] node374;
	wire [14-1:0] node375;
	wire [14-1:0] node379;
	wire [14-1:0] node382;
	wire [14-1:0] node384;
	wire [14-1:0] node387;
	wire [14-1:0] node388;
	wire [14-1:0] node389;
	wire [14-1:0] node391;
	wire [14-1:0] node392;
	wire [14-1:0] node393;
	wire [14-1:0] node394;
	wire [14-1:0] node395;
	wire [14-1:0] node397;
	wire [14-1:0] node400;
	wire [14-1:0] node401;
	wire [14-1:0] node405;
	wire [14-1:0] node406;
	wire [14-1:0] node408;
	wire [14-1:0] node412;
	wire [14-1:0] node413;
	wire [14-1:0] node415;
	wire [14-1:0] node419;
	wire [14-1:0] node420;
	wire [14-1:0] node422;
	wire [14-1:0] node423;
	wire [14-1:0] node425;
	wire [14-1:0] node430;
	wire [14-1:0] node431;
	wire [14-1:0] node432;
	wire [14-1:0] node433;
	wire [14-1:0] node435;
	wire [14-1:0] node437;
	wire [14-1:0] node438;
	wire [14-1:0] node439;
	wire [14-1:0] node443;
	wire [14-1:0] node444;
	wire [14-1:0] node450;
	wire [14-1:0] node451;
	wire [14-1:0] node452;
	wire [14-1:0] node453;
	wire [14-1:0] node454;
	wire [14-1:0] node455;
	wire [14-1:0] node461;
	wire [14-1:0] node464;
	wire [14-1:0] node466;
	wire [14-1:0] node467;
	wire [14-1:0] node469;
	wire [14-1:0] node473;
	wire [14-1:0] node474;
	wire [14-1:0] node475;
	wire [14-1:0] node477;
	wire [14-1:0] node478;
	wire [14-1:0] node479;
	wire [14-1:0] node480;
	wire [14-1:0] node483;
	wire [14-1:0] node488;
	wire [14-1:0] node489;
	wire [14-1:0] node490;
	wire [14-1:0] node492;
	wire [14-1:0] node493;
	wire [14-1:0] node495;
	wire [14-1:0] node496;
	wire [14-1:0] node499;
	wire [14-1:0] node501;
	wire [14-1:0] node504;
	wire [14-1:0] node508;
	wire [14-1:0] node510;
	wire [14-1:0] node512;
	wire [14-1:0] node514;
	wire [14-1:0] node518;
	wire [14-1:0] node519;
	wire [14-1:0] node520;
	wire [14-1:0] node521;
	wire [14-1:0] node522;
	wire [14-1:0] node523;
	wire [14-1:0] node528;
	wire [14-1:0] node530;
	wire [14-1:0] node532;
	wire [14-1:0] node535;
	wire [14-1:0] node536;
	wire [14-1:0] node537;
	wire [14-1:0] node538;
	wire [14-1:0] node539;
	wire [14-1:0] node544;
	wire [14-1:0] node546;
	wire [14-1:0] node548;
	wire [14-1:0] node551;
	wire [14-1:0] node552;
	wire [14-1:0] node553;
	wire [14-1:0] node554;
	wire [14-1:0] node558;
	wire [14-1:0] node560;
	wire [14-1:0] node561;
	wire [14-1:0] node562;
	wire [14-1:0] node564;
	wire [14-1:0] node565;
	wire [14-1:0] node566;
	wire [14-1:0] node573;
	wire [14-1:0] node574;
	wire [14-1:0] node575;
	wire [14-1:0] node576;
	wire [14-1:0] node577;
	wire [14-1:0] node578;
	wire [14-1:0] node579;
	wire [14-1:0] node585;
	wire [14-1:0] node588;
	wire [14-1:0] node589;
	wire [14-1:0] node593;
	wire [14-1:0] node594;
	wire [14-1:0] node595;
	wire [14-1:0] node596;
	wire [14-1:0] node597;
	wire [14-1:0] node598;
	wire [14-1:0] node599;
	wire [14-1:0] node606;
	wire [14-1:0] node609;
	wire [14-1:0] node610;
	wire [14-1:0] node613;
	wire [14-1:0] node616;
	wire [14-1:0] node617;
	wire [14-1:0] node618;
	wire [14-1:0] node619;
	wire [14-1:0] node621;
	wire [14-1:0] node622;
	wire [14-1:0] node623;
	wire [14-1:0] node624;
	wire [14-1:0] node625;
	wire [14-1:0] node626;
	wire [14-1:0] node630;
	wire [14-1:0] node632;
	wire [14-1:0] node637;
	wire [14-1:0] node639;
	wire [14-1:0] node640;
	wire [14-1:0] node642;
	wire [14-1:0] node643;
	wire [14-1:0] node647;
	wire [14-1:0] node649;
	wire [14-1:0] node650;
	wire [14-1:0] node651;
	wire [14-1:0] node654;
	wire [14-1:0] node658;
	wire [14-1:0] node659;
	wire [14-1:0] node660;
	wire [14-1:0] node661;
	wire [14-1:0] node662;
	wire [14-1:0] node664;
	wire [14-1:0] node666;
	wire [14-1:0] node667;
	wire [14-1:0] node671;
	wire [14-1:0] node672;
	wire [14-1:0] node677;
	wire [14-1:0] node678;
	wire [14-1:0] node679;
	wire [14-1:0] node680;
	wire [14-1:0] node681;
	wire [14-1:0] node684;
	wire [14-1:0] node687;
	wire [14-1:0] node688;
	wire [14-1:0] node691;
	wire [14-1:0] node694;
	wire [14-1:0] node695;
	wire [14-1:0] node696;
	wire [14-1:0] node701;
	wire [14-1:0] node702;
	wire [14-1:0] node704;
	wire [14-1:0] node708;
	wire [14-1:0] node709;
	wire [14-1:0] node711;
	wire [14-1:0] node713;
	wire [14-1:0] node715;
	wire [14-1:0] node719;
	wire [14-1:0] node720;
	wire [14-1:0] node721;
	wire [14-1:0] node722;
	wire [14-1:0] node723;
	wire [14-1:0] node724;
	wire [14-1:0] node725;
	wire [14-1:0] node727;
	wire [14-1:0] node731;
	wire [14-1:0] node733;
	wire [14-1:0] node734;
	wire [14-1:0] node738;
	wire [14-1:0] node739;
	wire [14-1:0] node741;
	wire [14-1:0] node744;
	wire [14-1:0] node746;
	wire [14-1:0] node749;
	wire [14-1:0] node751;
	wire [14-1:0] node752;
	wire [14-1:0] node754;
	wire [14-1:0] node756;
	wire [14-1:0] node757;
	wire [14-1:0] node761;
	wire [14-1:0] node762;
	wire [14-1:0] node763;
	wire [14-1:0] node767;
	wire [14-1:0] node769;
	wire [14-1:0] node772;
	wire [14-1:0] node774;
	wire [14-1:0] node776;
	wire [14-1:0] node778;
	wire [14-1:0] node780;
	wire [14-1:0] node782;
	wire [14-1:0] node783;
	wire [14-1:0] node787;
	wire [14-1:0] node788;
	wire [14-1:0] node789;
	wire [14-1:0] node790;
	wire [14-1:0] node791;
	wire [14-1:0] node792;
	wire [14-1:0] node793;
	wire [14-1:0] node794;
	wire [14-1:0] node801;
	wire [14-1:0] node803;
	wire [14-1:0] node805;
	wire [14-1:0] node807;
	wire [14-1:0] node810;
	wire [14-1:0] node811;
	wire [14-1:0] node812;
	wire [14-1:0] node813;
	wire [14-1:0] node814;
	wire [14-1:0] node822;
	wire [14-1:0] node823;
	wire [14-1:0] node824;
	wire [14-1:0] node825;
	wire [14-1:0] node826;
	wire [14-1:0] node827;
	wire [14-1:0] node829;
	wire [14-1:0] node831;
	wire [14-1:0] node835;
	wire [14-1:0] node836;
	wire [14-1:0] node838;
	wire [14-1:0] node839;
	wire [14-1:0] node842;
	wire [14-1:0] node844;
	wire [14-1:0] node845;
	wire [14-1:0] node848;
	wire [14-1:0] node851;
	wire [14-1:0] node853;
	wire [14-1:0] node854;
	wire [14-1:0] node855;
	wire [14-1:0] node860;
	wire [14-1:0] node861;
	wire [14-1:0] node862;
	wire [14-1:0] node863;
	wire [14-1:0] node865;
	wire [14-1:0] node870;
	wire [14-1:0] node872;
	wire [14-1:0] node874;
	wire [14-1:0] node876;
	wire [14-1:0] node879;
	wire [14-1:0] node880;
	wire [14-1:0] node881;
	wire [14-1:0] node882;
	wire [14-1:0] node884;
	wire [14-1:0] node885;
	wire [14-1:0] node887;
	wire [14-1:0] node891;
	wire [14-1:0] node893;
	wire [14-1:0] node895;
	wire [14-1:0] node897;
	wire [14-1:0] node898;
	wire [14-1:0] node902;
	wire [14-1:0] node903;
	wire [14-1:0] node905;
	wire [14-1:0] node906;
	wire [14-1:0] node911;
	wire [14-1:0] node912;
	wire [14-1:0] node913;
	wire [14-1:0] node914;
	wire [14-1:0] node915;
	wire [14-1:0] node921;
	wire [14-1:0] node922;
	wire [14-1:0] node923;
	wire [14-1:0] node925;
	wire [14-1:0] node926;
	wire [14-1:0] node931;
	wire [14-1:0] node932;
	wire [14-1:0] node934;
	wire [14-1:0] node936;
	wire [14-1:0] node939;
	wire [14-1:0] node940;
	wire [14-1:0] node944;
	wire [14-1:0] node945;
	wire [14-1:0] node946;
	wire [14-1:0] node948;
	wire [14-1:0] node949;
	wire [14-1:0] node950;
	wire [14-1:0] node951;
	wire [14-1:0] node954;
	wire [14-1:0] node956;
	wire [14-1:0] node958;
	wire [14-1:0] node963;
	wire [14-1:0] node964;
	wire [14-1:0] node965;
	wire [14-1:0] node966;
	wire [14-1:0] node967;
	wire [14-1:0] node968;
	wire [14-1:0] node975;
	wire [14-1:0] node977;
	wire [14-1:0] node979;
	wire [14-1:0] node981;
	wire [14-1:0] node984;
	wire [14-1:0] node985;
	wire [14-1:0] node986;
	wire [14-1:0] node987;
	wire [14-1:0] node988;
	wire [14-1:0] node989;
	wire [14-1:0] node991;
	wire [14-1:0] node995;
	wire [14-1:0] node996;
	wire [14-1:0] node1000;
	wire [14-1:0] node1001;
	wire [14-1:0] node1002;
	wire [14-1:0] node1003;
	wire [14-1:0] node1004;
	wire [14-1:0] node1011;
	wire [14-1:0] node1013;
	wire [14-1:0] node1015;
	wire [14-1:0] node1017;

	assign outp = (inp[10]) ? node518 : node1;
		assign node1 = (inp[13]) ? node287 : node2;
			assign node2 = (inp[11]) ? node128 : node3;
				assign node3 = (inp[12]) ? node49 : node4;
					assign node4 = (inp[8]) ? node6 : 14'b00000100000011;
						assign node6 = (inp[1]) ? node8 : 14'b00000000000000;
							assign node8 = (inp[3]) ? node20 : node9;
								assign node9 = (inp[2]) ? node11 : 14'b00000000000000;
									assign node11 = (inp[4]) ? 14'b00000000000000 : node12;
										assign node12 = (inp[9]) ? 14'b00000000000000 : node13;
											assign node13 = (inp[6]) ? 14'b00000000000000 : node14;
												assign node14 = (inp[0]) ? 14'b10000000011010 : 14'b00000000000000;
								assign node20 = (inp[0]) ? node40 : node21;
									assign node21 = (inp[2]) ? node33 : node22;
										assign node22 = (inp[6]) ? node26 : node23;
											assign node23 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
											assign node26 = (inp[7]) ? node28 : 14'b00000000000000;
												assign node28 = (inp[5]) ? 14'b00000000011100 : node29;
													assign node29 = (inp[9]) ? 14'b01000000010000 : 14'b00000000000000;
										assign node33 = (inp[6]) ? node35 : 14'b00000000000000;
											assign node35 = (inp[9]) ? node37 : 14'b00000000000000;
												assign node37 = (inp[5]) ? 14'b00000000011100 : 14'b01001000000100;
									assign node40 = (inp[9]) ? node42 : 14'b00000000000000;
										assign node42 = (inp[6]) ? node44 : 14'b00000000000000;
											assign node44 = (inp[2]) ? 14'b00000000000000 : node45;
												assign node45 = (inp[5]) ? 14'b00000000011100 : 14'b00000000000000;
					assign node49 = (inp[8]) ? node85 : node50;
						assign node50 = (inp[9]) ? 14'b00000000000000 : node51;
							assign node51 = (inp[5]) ? node75 : node52;
								assign node52 = (inp[7]) ? 14'b00000000000000 : node53;
									assign node53 = (inp[2]) ? node67 : node54;
										assign node54 = (inp[6]) ? node62 : node55;
											assign node55 = (inp[1]) ? node57 : 14'b00000000000000;
												assign node57 = (inp[0]) ? node59 : 14'b00000000000000;
													assign node59 = (inp[3]) ? 14'b00000000000000 : 14'b00100000000011;
											assign node62 = (inp[0]) ? 14'b00000000000000 : node63;
												assign node63 = (inp[1]) ? 14'b00000000000000 : 14'b00100000000011;
										assign node67 = (inp[6]) ? 14'b00000000000000 : node68;
											assign node68 = (inp[3]) ? 14'b00000000000000 : node69;
												assign node69 = (inp[4]) ? 14'b00000000000000 : 14'b00100000000011;
								assign node75 = (inp[6]) ? node77 : 14'b00000000000000;
									assign node77 = (inp[0]) ? 14'b00000000000000 : node78;
										assign node78 = (inp[7]) ? node80 : 14'b00000000000000;
											assign node80 = (inp[1]) ? 14'b00001000000101 : 14'b00000000000000;
						assign node85 = (inp[6]) ? node111 : node86;
							assign node86 = (inp[1]) ? node88 : 14'b00000000000000;
								assign node88 = (inp[2]) ? 14'b00000000000000 : node89;
									assign node89 = (inp[0]) ? node101 : node90;
										assign node90 = (inp[9]) ? node96 : node91;
											assign node91 = (inp[3]) ? node93 : 14'b00100000000011;
												assign node93 = (inp[4]) ? 14'b00000000000000 : 14'b00001000000000;
											assign node96 = (inp[7]) ? 14'b00000000000000 : node97;
												assign node97 = (inp[3]) ? 14'b00001000000101 : 14'b00000000000000;
										assign node101 = (inp[3]) ? 14'b00000000000000 : node102;
											assign node102 = (inp[4]) ? 14'b00000000000000 : node103;
												assign node103 = (inp[9]) ? 14'b00000000000000 : node104;
													assign node104 = (inp[5]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node111 = (inp[3]) ? node123 : node112;
								assign node112 = (inp[1]) ? node114 : 14'b00000000000000;
									assign node114 = (inp[0]) ? 14'b00000000000000 : node115;
										assign node115 = (inp[4]) ? 14'b00000000000000 : node116;
											assign node116 = (inp[9]) ? 14'b00000000000000 : node117;
												assign node117 = (inp[2]) ? 14'b00000000000000 : 14'b10100100111111;
								assign node123 = (inp[1]) ? 14'b00000000000000 : node124;
									assign node124 = (inp[9]) ? 14'b11110111110010 : 14'b00000000000000;
				assign node128 = (inp[12]) ? node200 : node129;
					assign node129 = (inp[1]) ? node131 : 14'b00000000000000;
						assign node131 = (inp[8]) ? node171 : node132;
							assign node132 = (inp[3]) ? node144 : node133;
								assign node133 = (inp[0]) ? node135 : 14'b00000000000000;
									assign node135 = (inp[4]) ? 14'b00000000000000 : node136;
										assign node136 = (inp[2]) ? node138 : 14'b00000000000000;
											assign node138 = (inp[6]) ? 14'b00000000000000 : node139;
												assign node139 = (inp[9]) ? 14'b00000000000000 : 14'b00100000000011;
								assign node144 = (inp[7]) ? node146 : 14'b00000000000000;
									assign node146 = (inp[2]) ? node164 : node147;
										assign node147 = (inp[0]) ? node155 : node148;
											assign node148 = (inp[6]) ? node150 : 14'b10010000001101;
												assign node150 = (inp[9]) ? node152 : 14'b00000000000000;
													assign node152 = (inp[4]) ? 14'b10100000101010 : 14'b10100000111010;
											assign node155 = (inp[4]) ? 14'b00000000000000 : node156;
												assign node156 = (inp[5]) ? 14'b00000000000000 : node157;
													assign node157 = (inp[9]) ? node159 : 14'b00000000000000;
														assign node159 = (inp[6]) ? 14'b01001000000100 : 14'b00000000000000;
										assign node164 = (inp[9]) ? node166 : 14'b00000000000000;
											assign node166 = (inp[6]) ? node168 : 14'b00000000000000;
												assign node168 = (inp[5]) ? 14'b00000000000000 : 14'b01001000000100;
							assign node171 = (inp[3]) ? node185 : node172;
								assign node172 = (inp[9]) ? 14'b00000000000000 : node173;
									assign node173 = (inp[6]) ? node175 : 14'b01001000000100;
										assign node175 = (inp[7]) ? node179 : node176;
											assign node176 = (inp[5]) ? 14'b00000000000000 : 14'b11000000000100;
											assign node179 = (inp[0]) ? 14'b00000000000000 : node180;
												assign node180 = (inp[4]) ? 14'b11000000000100 : 14'b00000000000000;
								assign node185 = (inp[7]) ? node193 : node186;
									assign node186 = (inp[0]) ? 14'b00000000000000 : node187;
										assign node187 = (inp[2]) ? 14'b00000000000000 : node188;
											assign node188 = (inp[6]) ? 14'b00000000000000 : 14'b00000100000001;
									assign node193 = (inp[9]) ? node195 : 14'b00000000000000;
										assign node195 = (inp[5]) ? 14'b00000000000000 : node196;
											assign node196 = (inp[6]) ? 14'b01100000001010 : 14'b00000000000000;
					assign node200 = (inp[9]) ? node234 : node201;
						assign node201 = (inp[1]) ? node209 : node202;
							assign node202 = (inp[6]) ? node204 : 14'b00000000000000;
								assign node204 = (inp[3]) ? node206 : 14'b00000000000000;
									assign node206 = (inp[8]) ? 14'b00000000000000 : 14'b01100000001010;
							assign node209 = (inp[3]) ? node223 : node210;
								assign node210 = (inp[6]) ? node214 : node211;
									assign node211 = (inp[8]) ? 14'b00100100011111 : 14'b10000100011000;
									assign node214 = (inp[8]) ? 14'b01000100000100 : node215;
										assign node215 = (inp[2]) ? 14'b00000000000000 : node216;
											assign node216 = (inp[5]) ? node218 : 14'b00000000000000;
												assign node218 = (inp[0]) ? 14'b00000000000000 : 14'b10100000001000;
								assign node223 = (inp[6]) ? 14'b00000000000000 : node224;
									assign node224 = (inp[2]) ? 14'b00000000000000 : node225;
										assign node225 = (inp[7]) ? node227 : 14'b00000000000000;
											assign node227 = (inp[0]) ? 14'b00000000000000 : node228;
												assign node228 = (inp[8]) ? 14'b00000000000000 : 14'b01001000000101;
						assign node234 = (inp[3]) ? node248 : node235;
							assign node235 = (inp[7]) ? node237 : 14'b00000000000000;
								assign node237 = (inp[1]) ? node239 : 14'b00000000000000;
									assign node239 = (inp[8]) ? 14'b00000000000000 : node240;
										assign node240 = (inp[0]) ? 14'b00000000000000 : node241;
											assign node241 = (inp[2]) ? 14'b00000000000000 : node242;
												assign node242 = (inp[6]) ? 14'b00000000000000 : 14'b01001000000100;
							assign node248 = (inp[6]) ? node272 : node249;
								assign node249 = (inp[8]) ? node259 : node250;
									assign node250 = (inp[2]) ? 14'b00000000000000 : node251;
										assign node251 = (inp[1]) ? node253 : 14'b00000000000000;
											assign node253 = (inp[0]) ? 14'b00000000000000 : node254;
												assign node254 = (inp[7]) ? 14'b01001000000100 : 14'b00000000000000;
									assign node259 = (inp[7]) ? 14'b00000000000000 : node260;
										assign node260 = (inp[2]) ? 14'b00000000000000 : node261;
											assign node261 = (inp[1]) ? node263 : 14'b00000000000000;
												assign node263 = (inp[5]) ? node265 : 14'b00000000000000;
													assign node265 = (inp[0]) ? 14'b00000000000000 : node266;
														assign node266 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
								assign node272 = (inp[8]) ? node280 : node273;
									assign node273 = (inp[5]) ? node275 : 14'b00000000000000;
										assign node275 = (inp[7]) ? 14'b00000000000000 : node276;
											assign node276 = (inp[1]) ? 14'b01001000001100 : 14'b00000000000000;
									assign node280 = (inp[1]) ? node282 : 14'b10100010001100;
										assign node282 = (inp[7]) ? node284 : 14'b00000000000000;
											assign node284 = (inp[5]) ? 14'b10000000011010 : 14'b00000000000000;
			assign node287 = (inp[12]) ? node387 : node288;
				assign node288 = (inp[1]) ? node314 : node289;
					assign node289 = (inp[3]) ? node291 : 14'b00000000000000;
						assign node291 = (inp[8]) ? node301 : node292;
							assign node292 = (inp[7]) ? 14'b00000000000000 : node293;
								assign node293 = (inp[9]) ? 14'b00000000000000 : node294;
									assign node294 = (inp[6]) ? node296 : 14'b00000000000000;
										assign node296 = (inp[11]) ? 14'b00000000000000 : 14'b11000000000100;
							assign node301 = (inp[2]) ? 14'b00000000000000 : node302;
								assign node302 = (inp[6]) ? node304 : 14'b00000000000000;
									assign node304 = (inp[11]) ? node306 : 14'b00000000000000;
										assign node306 = (inp[9]) ? 14'b00000000000000 : node307;
											assign node307 = (inp[0]) ? 14'b00000000000000 : node308;
												assign node308 = (inp[7]) ? 14'b00000000000000 : 14'b00100000000011;
					assign node314 = (inp[6]) ? node364 : node315;
						assign node315 = (inp[9]) ? node349 : node316;
							assign node316 = (inp[3]) ? node330 : node317;
								assign node317 = (inp[11]) ? node321 : node318;
									assign node318 = (inp[8]) ? 14'b00000000000000 : 14'b11000000000100;
									assign node321 = (inp[8]) ? 14'b00000000011100 : node322;
										assign node322 = (inp[4]) ? 14'b00000000000000 : node323;
											assign node323 = (inp[2]) ? 14'b10110101111111 : node324;
												assign node324 = (inp[7]) ? 14'b01001000000100 : 14'b00000000000000;
								assign node330 = (inp[2]) ? 14'b00000000000000 : node331;
									assign node331 = (inp[0]) ? 14'b00000000000000 : node332;
										assign node332 = (inp[11]) ? node342 : node333;
											assign node333 = (inp[8]) ? node335 : 14'b00000000000000;
												assign node335 = (inp[5]) ? node337 : 14'b00000000000000;
													assign node337 = (inp[7]) ? node339 : 14'b00000000000000;
														assign node339 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
											assign node342 = (inp[8]) ? node344 : 14'b10000100101010;
												assign node344 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node349 = (inp[11]) ? node351 : 14'b00000000000000;
								assign node351 = (inp[0]) ? 14'b00000000000000 : node352;
									assign node352 = (inp[2]) ? 14'b00000000000000 : node353;
										assign node353 = (inp[3]) ? node355 : 14'b00000000000000;
											assign node355 = (inp[8]) ? node359 : node356;
												assign node356 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
												assign node359 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
						assign node364 = (inp[7]) ? node366 : 14'b00000000000000;
							assign node366 = (inp[3]) ? node368 : 14'b00000000000000;
								assign node368 = (inp[9]) ? node370 : 14'b00000000000000;
									assign node370 = (inp[5]) ? node382 : node371;
										assign node371 = (inp[11]) ? node379 : node372;
											assign node372 = (inp[8]) ? node374 : 14'b01100000000110;
												assign node374 = (inp[4]) ? 14'b00000000000000 : node375;
													assign node375 = (inp[0]) ? 14'b00000000000000 : 14'b00000000011100;
											assign node379 = (inp[8]) ? 14'b10100010001100 : 14'b10000010001100;
										assign node382 = (inp[11]) ? node384 : 14'b00000000000000;
											assign node384 = (inp[8]) ? 14'b00000000000000 : 14'b01001000000101;
				assign node387 = (inp[8]) ? node473 : node388;
					assign node388 = (inp[3]) ? node430 : node389;
						assign node389 = (inp[1]) ? node391 : 14'b00000000000000;
							assign node391 = (inp[6]) ? node419 : node392;
								assign node392 = (inp[4]) ? node412 : node393;
									assign node393 = (inp[2]) ? node405 : node394;
										assign node394 = (inp[7]) ? node400 : node395;
											assign node395 = (inp[0]) ? node397 : 14'b00000000000000;
												assign node397 = (inp[9]) ? 14'b00000000000000 : 14'b01001000000101;
											assign node400 = (inp[0]) ? 14'b00000000000000 : node401;
												assign node401 = (inp[11]) ? 14'b10100010001100 : 14'b11110111110010;
										assign node405 = (inp[9]) ? 14'b00000000000000 : node406;
											assign node406 = (inp[0]) ? node408 : 14'b00000000000000;
												assign node408 = (inp[11]) ? 14'b00000000000000 : 14'b10000000101100;
									assign node412 = (inp[0]) ? 14'b00000000000000 : node413;
										assign node413 = (inp[9]) ? node415 : 14'b00000000000000;
											assign node415 = (inp[7]) ? 14'b10100010001100 : 14'b00000000000000;
								assign node419 = (inp[9]) ? 14'b00000000000000 : node420;
									assign node420 = (inp[5]) ? node422 : 14'b00000000000000;
										assign node422 = (inp[0]) ? 14'b00000000000000 : node423;
											assign node423 = (inp[7]) ? node425 : 14'b00000000000000;
												assign node425 = (inp[2]) ? 14'b00000000000000 : 14'b01001000000101;
						assign node430 = (inp[6]) ? node450 : node431;
							assign node431 = (inp[0]) ? 14'b00000000000000 : node432;
								assign node432 = (inp[2]) ? 14'b00000000000000 : node433;
									assign node433 = (inp[7]) ? node435 : 14'b00000000000000;
										assign node435 = (inp[1]) ? node437 : 14'b00000000000000;
											assign node437 = (inp[11]) ? node443 : node438;
												assign node438 = (inp[9]) ? 14'b11110111110010 : node439;
													assign node439 = (inp[5]) ? 14'b11110111110010 : 14'b00000000000000;
												assign node443 = (inp[9]) ? 14'b10100010001100 : node444;
													assign node444 = (inp[5]) ? 14'b10100010001100 : 14'b10010101111110;
							assign node450 = (inp[1]) ? node464 : node451;
								assign node451 = (inp[11]) ? node461 : node452;
									assign node452 = (inp[7]) ? 14'b00000000000000 : node453;
										assign node453 = (inp[2]) ? 14'b00000000000000 : node454;
											assign node454 = (inp[0]) ? 14'b00000000000000 : node455;
												assign node455 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
									assign node461 = (inp[9]) ? 14'b00000000000000 : 14'b00100100001101;
								assign node464 = (inp[5]) ? node466 : 14'b00000000000000;
									assign node466 = (inp[7]) ? 14'b00000000000000 : node467;
										assign node467 = (inp[9]) ? node469 : 14'b00000000000000;
											assign node469 = (inp[11]) ? 14'b00000000011100 : 14'b00000000011101;
					assign node473 = (inp[11]) ? 14'b01000000010100 : node474;
						assign node474 = (inp[6]) ? node488 : node475;
							assign node475 = (inp[1]) ? node477 : 14'b00000000000000;
								assign node477 = (inp[2]) ? 14'b00000000000000 : node478;
									assign node478 = (inp[0]) ? 14'b00000000000000 : node479;
										assign node479 = (inp[3]) ? node483 : node480;
											assign node480 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
											assign node483 = (inp[7]) ? 14'b00000000000000 : 14'b10000100101010;
							assign node488 = (inp[3]) ? node508 : node489;
								assign node489 = (inp[9]) ? 14'b00000000000000 : node490;
									assign node490 = (inp[1]) ? node492 : 14'b00000000000000;
										assign node492 = (inp[5]) ? node504 : node493;
											assign node493 = (inp[7]) ? node495 : 14'b10010100011100;
												assign node495 = (inp[2]) ? node499 : node496;
													assign node496 = (inp[0]) ? 14'b00000000000000 : 14'b10010010001100;
													assign node499 = (inp[0]) ? node501 : 14'b00000000000000;
														assign node501 = (inp[4]) ? 14'b10010010001100 : 14'b00000000000000;
											assign node504 = (inp[7]) ? 14'b11100100010100 : 14'b11100100000100;
								assign node508 = (inp[9]) ? node510 : 14'b00000000000000;
									assign node510 = (inp[1]) ? node512 : 14'b01001000000100;
										assign node512 = (inp[5]) ? node514 : 14'b00000000000000;
											assign node514 = (inp[7]) ? 14'b01001000001001 : 14'b00000000000000;
		assign node518 = (inp[1]) ? node616 : node519;
			assign node519 = (inp[3]) ? node535 : node520;
				assign node520 = (inp[11]) ? node528 : node521;
					assign node521 = (inp[12]) ? 14'b00000000000000 : node522;
						assign node522 = (inp[13]) ? 14'b00000000000000 : node523;
							assign node523 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
					assign node528 = (inp[8]) ? node530 : 14'b00000000000000;
						assign node530 = (inp[12]) ? node532 : 14'b00000000000000;
							assign node532 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
				assign node535 = (inp[6]) ? node551 : node536;
					assign node536 = (inp[12]) ? node544 : node537;
						assign node537 = (inp[13]) ? 14'b00000000000000 : node538;
							assign node538 = (inp[8]) ? 14'b00000000000000 : node539;
								assign node539 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
						assign node544 = (inp[13]) ? node546 : 14'b00000000000000;
							assign node546 = (inp[11]) ? node548 : 14'b00000000000000;
								assign node548 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node551 = (inp[12]) ? node573 : node552;
						assign node552 = (inp[11]) ? node558 : node553;
							assign node553 = (inp[13]) ? 14'b00000000000000 : node554;
								assign node554 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
							assign node558 = (inp[13]) ? node560 : 14'b00000000000000;
								assign node560 = (inp[0]) ? 14'b00000000000000 : node561;
									assign node561 = (inp[9]) ? 14'b00000000000000 : node562;
										assign node562 = (inp[8]) ? node564 : 14'b00000000000000;
											assign node564 = (inp[7]) ? 14'b00000000000000 : node565;
												assign node565 = (inp[2]) ? 14'b00000000000000 : node566;
													assign node566 = (inp[5]) ? 14'b10000100101010 : 14'b10000100111010;
						assign node573 = (inp[13]) ? node593 : node574;
							assign node574 = (inp[11]) ? node588 : node575;
								assign node575 = (inp[8]) ? node585 : node576;
									assign node576 = (inp[9]) ? 14'b00000000000000 : node577;
										assign node577 = (inp[7]) ? 14'b00000000000000 : node578;
											assign node578 = (inp[2]) ? 14'b00000000000000 : node579;
												assign node579 = (inp[0]) ? 14'b00000000000000 : 14'b10100100111000;
									assign node585 = (inp[9]) ? 14'b01100000001010 : 14'b00000000000000;
								assign node588 = (inp[8]) ? 14'b00000000000000 : node589;
									assign node589 = (inp[9]) ? 14'b00000000000000 : 14'b01001000000101;
							assign node593 = (inp[11]) ? node609 : node594;
								assign node594 = (inp[9]) ? node606 : node595;
									assign node595 = (inp[0]) ? 14'b00000000000000 : node596;
										assign node596 = (inp[7]) ? 14'b00000000000000 : node597;
											assign node597 = (inp[2]) ? 14'b00000000000000 : node598;
												assign node598 = (inp[8]) ? 14'b00000000000000 : node599;
													assign node599 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
									assign node606 = (inp[8]) ? 14'b00100100001101 : 14'b00000000000000;
								assign node609 = (inp[9]) ? node613 : node610;
									assign node610 = (inp[8]) ? 14'b10000100001000 : 14'b10010101111110;
									assign node613 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
			assign node616 = (inp[13]) ? node822 : node617;
				assign node617 = (inp[12]) ? node719 : node618;
					assign node618 = (inp[11]) ? node658 : node619;
						assign node619 = (inp[8]) ? node621 : 14'b10000100001000;
							assign node621 = (inp[3]) ? node637 : node622;
								assign node622 = (inp[9]) ? 14'b00000000000000 : node623;
									assign node623 = (inp[6]) ? 14'b00000000000000 : node624;
										assign node624 = (inp[0]) ? node630 : node625;
											assign node625 = (inp[4]) ? 14'b00100000000011 : node626;
												assign node626 = (inp[2]) ? 14'b00000000000000 : 14'b00100000000011;
											assign node630 = (inp[2]) ? node632 : 14'b00000000000000;
												assign node632 = (inp[4]) ? 14'b00000000000000 : 14'b00100000000011;
								assign node637 = (inp[7]) ? node639 : 14'b00000000000000;
									assign node639 = (inp[9]) ? node647 : node640;
										assign node640 = (inp[5]) ? node642 : 14'b00000000000000;
											assign node642 = (inp[0]) ? 14'b00000000000000 : node643;
												assign node643 = (inp[2]) ? 14'b00000000000000 : 14'b00000000011100;
										assign node647 = (inp[6]) ? node649 : 14'b00000000000000;
											assign node649 = (inp[5]) ? 14'b10100000001000 : node650;
												assign node650 = (inp[2]) ? node654 : node651;
													assign node651 = (inp[0]) ? 14'b00000000000000 : 14'b00100000001010;
													assign node654 = (inp[4]) ? 14'b00000000000000 : 14'b10010010001101;
						assign node658 = (inp[6]) ? node708 : node659;
							assign node659 = (inp[8]) ? node677 : node660;
								assign node660 = (inp[2]) ? 14'b00000000000000 : node661;
									assign node661 = (inp[3]) ? node671 : node662;
										assign node662 = (inp[0]) ? node664 : 14'b00000000000000;
											assign node664 = (inp[7]) ? node666 : 14'b00000000000000;
												assign node666 = (inp[4]) ? 14'b00000000000000 : node667;
													assign node667 = (inp[9]) ? 14'b00000000000000 : 14'b01100000001010;
										assign node671 = (inp[0]) ? 14'b00000000000000 : node672;
											assign node672 = (inp[7]) ? 14'b00000000000000 : 14'b00100000000011;
								assign node677 = (inp[9]) ? node701 : node678;
									assign node678 = (inp[3]) ? node694 : node679;
										assign node679 = (inp[0]) ? node687 : node680;
											assign node680 = (inp[2]) ? node684 : node681;
												assign node681 = (inp[4]) ? 14'b10000010001101 : 14'b10000001001101;
												assign node684 = (inp[7]) ? 14'b00000000000000 : 14'b10000100001101;
											assign node687 = (inp[4]) ? node691 : node688;
												assign node688 = (inp[2]) ? 14'b10010000001101 : 14'b00000000000000;
												assign node691 = (inp[2]) ? 14'b00000000000000 : 14'b10000000011101;
										assign node694 = (inp[2]) ? 14'b00000000000000 : node695;
											assign node695 = (inp[7]) ? 14'b00000000000000 : node696;
												assign node696 = (inp[0]) ? 14'b00000000000000 : 14'b00100000001010;
									assign node701 = (inp[2]) ? 14'b00000000000000 : node702;
										assign node702 = (inp[3]) ? node704 : 14'b00000000000000;
											assign node704 = (inp[0]) ? 14'b00000000000000 : 14'b00100000001010;
							assign node708 = (inp[5]) ? 14'b00000000000000 : node709;
								assign node709 = (inp[3]) ? node711 : 14'b00000000000000;
									assign node711 = (inp[7]) ? node713 : 14'b00000000000000;
										assign node713 = (inp[9]) ? node715 : 14'b00000000000000;
											assign node715 = (inp[8]) ? 14'b01001000000100 : 14'b00000100001111;
					assign node719 = (inp[0]) ? node787 : node720;
						assign node720 = (inp[2]) ? node772 : node721;
							assign node721 = (inp[6]) ? node749 : node722;
								assign node722 = (inp[3]) ? node738 : node723;
									assign node723 = (inp[11]) ? node731 : node724;
										assign node724 = (inp[9]) ? 14'b00000000000000 : node725;
											assign node725 = (inp[8]) ? node727 : 14'b00000000000000;
												assign node727 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
										assign node731 = (inp[9]) ? node733 : 14'b00000000000000;
											assign node733 = (inp[5]) ? 14'b00000000000000 : node734;
												assign node734 = (inp[8]) ? 14'b00000000000000 : 14'b00100100001101;
									assign node738 = (inp[7]) ? node744 : node739;
										assign node739 = (inp[8]) ? node741 : 14'b00000000000000;
											assign node741 = (inp[11]) ? 14'b00000000000000 : 14'b00000000011100;
										assign node744 = (inp[11]) ? node746 : 14'b00000000000000;
											assign node746 = (inp[8]) ? 14'b00000000000000 : 14'b00100100001101;
								assign node749 = (inp[5]) ? node751 : 14'b00000000000000;
									assign node751 = (inp[7]) ? node761 : node752;
										assign node752 = (inp[9]) ? node754 : 14'b00000000000000;
											assign node754 = (inp[3]) ? node756 : 14'b00000000000000;
												assign node756 = (inp[8]) ? 14'b00000000000000 : node757;
													assign node757 = (inp[11]) ? 14'b00000100001111 : 14'b00001000001100;
										assign node761 = (inp[11]) ? node767 : node762;
											assign node762 = (inp[8]) ? 14'b01100000000110 : node763;
												assign node763 = (inp[3]) ? 14'b00000000000000 : 14'b00000100001101;
											assign node767 = (inp[4]) ? node769 : 14'b00000000000000;
												assign node769 = (inp[9]) ? 14'b00000000000000 : 14'b01100000000010;
							assign node772 = (inp[5]) ? node774 : 14'b00000000000000;
								assign node774 = (inp[9]) ? node776 : 14'b00000000000000;
									assign node776 = (inp[6]) ? node778 : 14'b00000000000000;
										assign node778 = (inp[3]) ? node780 : 14'b00000000000000;
											assign node780 = (inp[7]) ? node782 : 14'b00000100001111;
												assign node782 = (inp[4]) ? 14'b00000000000000 : node783;
													assign node783 = (inp[8]) ? 14'b01100000000110 : 14'b00000000000000;
						assign node787 = (inp[8]) ? 14'b00000000000000 : node788;
							assign node788 = (inp[7]) ? node810 : node789;
								assign node789 = (inp[5]) ? node801 : node790;
									assign node790 = (inp[4]) ? 14'b00000000000000 : node791;
										assign node791 = (inp[3]) ? 14'b00000000000000 : node792;
											assign node792 = (inp[6]) ? 14'b00000000000000 : node793;
												assign node793 = (inp[9]) ? 14'b00000000000000 : node794;
													assign node794 = (inp[11]) ? 14'b00001000000101 : 14'b01001000000100;
									assign node801 = (inp[6]) ? node803 : 14'b00000000000000;
										assign node803 = (inp[9]) ? node805 : 14'b00000000000000;
											assign node805 = (inp[3]) ? node807 : 14'b00000000000000;
												assign node807 = (inp[4]) ? 14'b00000100001111 : 14'b00001000001100;
								assign node810 = (inp[3]) ? 14'b00000000000000 : node811;
									assign node811 = (inp[5]) ? 14'b00000000000000 : node812;
										assign node812 = (inp[9]) ? 14'b00000000000000 : node813;
											assign node813 = (inp[4]) ? 14'b00000000000000 : node814;
												assign node814 = (inp[6]) ? 14'b00000000000000 : 14'b00001000000101;
				assign node822 = (inp[8]) ? node944 : node823;
					assign node823 = (inp[12]) ? node879 : node824;
						assign node824 = (inp[2]) ? node860 : node825;
							assign node825 = (inp[7]) ? node835 : node826;
								assign node826 = (inp[0]) ? 14'b00000000000000 : node827;
									assign node827 = (inp[3]) ? node829 : 14'b00000000000000;
										assign node829 = (inp[11]) ? node831 : 14'b00000000000000;
											assign node831 = (inp[6]) ? 14'b00000000000000 : 14'b00100000000011;
								assign node835 = (inp[0]) ? node851 : node836;
									assign node836 = (inp[9]) ? node838 : 14'b00000000000000;
										assign node838 = (inp[6]) ? node842 : node839;
											assign node839 = (inp[11]) ? 14'b00000000000000 : 14'b00001000000100;
											assign node842 = (inp[3]) ? node844 : 14'b00000000000000;
												assign node844 = (inp[5]) ? node848 : node845;
													assign node845 = (inp[11]) ? 14'b00001000001001 : 14'b00000000011101;
													assign node848 = (inp[11]) ? 14'b10100101111111 : 14'b00000000000000;
									assign node851 = (inp[11]) ? node853 : 14'b00000000000000;
										assign node853 = (inp[6]) ? 14'b00000000000000 : node854;
											assign node854 = (inp[9]) ? 14'b00000000000000 : node855;
												assign node855 = (inp[4]) ? 14'b00000000000000 : 14'b10000100001101;
							assign node860 = (inp[9]) ? node870 : node861;
								assign node861 = (inp[6]) ? 14'b00000000000000 : node862;
									assign node862 = (inp[3]) ? 14'b00000000000000 : node863;
										assign node863 = (inp[0]) ? node865 : 14'b00000000000000;
											assign node865 = (inp[11]) ? 14'b00000000011100 : 14'b00000000000000;
								assign node870 = (inp[6]) ? node872 : 14'b00000000000000;
									assign node872 = (inp[3]) ? node874 : 14'b00000000000000;
										assign node874 = (inp[7]) ? node876 : 14'b00000000000000;
											assign node876 = (inp[11]) ? 14'b01000100000010 : 14'b00000000000000;
						assign node879 = (inp[9]) ? node911 : node880;
							assign node880 = (inp[3]) ? node902 : node881;
								assign node881 = (inp[6]) ? node891 : node882;
									assign node882 = (inp[11]) ? node884 : 14'b00000000011101;
										assign node884 = (inp[2]) ? 14'b00000000000000 : node885;
											assign node885 = (inp[7]) ? node887 : 14'b00000000000000;
												assign node887 = (inp[5]) ? 14'b00000000000000 : 14'b10000000001111;
									assign node891 = (inp[11]) ? node893 : 14'b00000000000000;
										assign node893 = (inp[5]) ? node895 : 14'b00000000000000;
											assign node895 = (inp[4]) ? node897 : 14'b00000000000000;
												assign node897 = (inp[0]) ? 14'b00000000000000 : node898;
													assign node898 = (inp[2]) ? 14'b00000000000000 : 14'b01001000000101;
								assign node902 = (inp[11]) ? 14'b00000000000000 : node903;
									assign node903 = (inp[7]) ? node905 : 14'b00000000000000;
										assign node905 = (inp[2]) ? 14'b00000000000000 : node906;
											assign node906 = (inp[4]) ? 14'b01100000001010 : 14'b00000000000000;
							assign node911 = (inp[3]) ? node921 : node912;
								assign node912 = (inp[0]) ? 14'b00000000000000 : node913;
									assign node913 = (inp[2]) ? 14'b00000000000000 : node914;
										assign node914 = (inp[11]) ? 14'b00000000000000 : node915;
											assign node915 = (inp[7]) ? 14'b01100000001010 : 14'b00000000000000;
								assign node921 = (inp[5]) ? node931 : node922;
									assign node922 = (inp[2]) ? 14'b00000000000000 : node923;
										assign node923 = (inp[7]) ? node925 : 14'b00000000000000;
											assign node925 = (inp[0]) ? 14'b00000000000000 : node926;
												assign node926 = (inp[11]) ? 14'b00000000000000 : 14'b01100000001010;
									assign node931 = (inp[6]) ? node939 : node932;
										assign node932 = (inp[7]) ? node934 : 14'b00000000000000;
											assign node934 = (inp[4]) ? node936 : 14'b00000000000000;
												assign node936 = (inp[11]) ? 14'b00000000000000 : 14'b01100000001010;
										assign node939 = (inp[7]) ? 14'b00000000000000 : node940;
											assign node940 = (inp[11]) ? 14'b10100100001000 : 14'b10100000001000;
					assign node944 = (inp[11]) ? node984 : node945;
						assign node945 = (inp[12]) ? node963 : node946;
							assign node946 = (inp[3]) ? node948 : 14'b00000000000000;
								assign node948 = (inp[0]) ? 14'b00000000000000 : node949;
									assign node949 = (inp[2]) ? 14'b00000000000000 : node950;
										assign node950 = (inp[6]) ? node954 : node951;
											assign node951 = (inp[7]) ? 14'b00000000000000 : 14'b00001000001001;
											assign node954 = (inp[7]) ? node956 : 14'b00000000000000;
												assign node956 = (inp[9]) ? node958 : 14'b00000000000000;
													assign node958 = (inp[4]) ? 14'b10000100101000 : 14'b10000100111000;
							assign node963 = (inp[9]) ? node975 : node964;
								assign node964 = (inp[3]) ? 14'b00000000000000 : node965;
									assign node965 = (inp[6]) ? 14'b00000100001110 : node966;
										assign node966 = (inp[0]) ? 14'b00001000000100 : node967;
											assign node967 = (inp[2]) ? 14'b00001000000100 : node968;
												assign node968 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
								assign node975 = (inp[3]) ? node977 : 14'b00000000000000;
									assign node977 = (inp[7]) ? node979 : 14'b00000000000000;
										assign node979 = (inp[5]) ? node981 : 14'b00000000000000;
											assign node981 = (inp[6]) ? 14'b00000000011100 : 14'b00000000000000;
						assign node984 = (inp[12]) ? 14'b10000100001000 : node985;
							assign node985 = (inp[6]) ? node1011 : node986;
								assign node986 = (inp[9]) ? node1000 : node987;
									assign node987 = (inp[3]) ? node995 : node988;
										assign node988 = (inp[0]) ? 14'b10100100011000 : node989;
											assign node989 = (inp[2]) ? node991 : 14'b10000000001010;
												assign node991 = (inp[4]) ? 14'b10100100011000 : 14'b00000000000000;
										assign node995 = (inp[0]) ? 14'b00000000000000 : node996;
											assign node996 = (inp[5]) ? 14'b10100100101000 : 14'b00000000000000;
									assign node1000 = (inp[7]) ? 14'b00000000000000 : node1001;
										assign node1001 = (inp[5]) ? 14'b00000000000000 : node1002;
											assign node1002 = (inp[0]) ? 14'b00000000000000 : node1003;
												assign node1003 = (inp[2]) ? 14'b00000000000000 : node1004;
													assign node1004 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
								assign node1011 = (inp[7]) ? node1013 : 14'b00000000000000;
									assign node1013 = (inp[3]) ? node1015 : 14'b00000000000000;
										assign node1015 = (inp[9]) ? node1017 : 14'b00000000000000;
											assign node1017 = (inp[5]) ? 14'b00000000000000 : 14'b00100100001101;

endmodule