module dtc_split75_bm58 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node35;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node278;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node304;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node324;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node341;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[0]) ? node214 : node3;
			assign node3 = (inp[4]) ? node89 : node4;
				assign node4 = (inp[9]) ? node40 : node5;
					assign node5 = (inp[1]) ? 3'b000 : node6;
						assign node6 = (inp[11]) ? node22 : node7;
							assign node7 = (inp[8]) ? 3'b100 : node8;
								assign node8 = (inp[3]) ? node16 : node9;
									assign node9 = (inp[10]) ? 3'b100 : node10;
										assign node10 = (inp[2]) ? 3'b100 : node11;
											assign node11 = (inp[7]) ? 3'b000 : 3'b100;
									assign node16 = (inp[10]) ? node18 : 3'b000;
										assign node18 = (inp[2]) ? 3'b100 : 3'b000;
							assign node22 = (inp[8]) ? node24 : 3'b000;
								assign node24 = (inp[10]) ? node32 : node25;
									assign node25 = (inp[3]) ? 3'b000 : node26;
										assign node26 = (inp[2]) ? 3'b100 : node27;
											assign node27 = (inp[5]) ? 3'b000 : 3'b100;
									assign node32 = (inp[2]) ? 3'b100 : node33;
										assign node33 = (inp[7]) ? node35 : 3'b100;
											assign node35 = (inp[3]) ? 3'b000 : 3'b100;
					assign node40 = (inp[1]) ? node72 : node41;
						assign node41 = (inp[11]) ? node57 : node42;
							assign node42 = (inp[8]) ? node50 : node43;
								assign node43 = (inp[3]) ? node45 : 3'b000;
									assign node45 = (inp[2]) ? 3'b000 : node46;
										assign node46 = (inp[10]) ? 3'b000 : 3'b100;
								assign node50 = (inp[10]) ? 3'b100 : node51;
									assign node51 = (inp[3]) ? 3'b000 : node52;
										assign node52 = (inp[2]) ? 3'b100 : 3'b000;
							assign node57 = (inp[8]) ? node65 : node58;
								assign node58 = (inp[10]) ? node60 : 3'b100;
									assign node60 = (inp[3]) ? node62 : 3'b000;
										assign node62 = (inp[2]) ? 3'b000 : 3'b100;
								assign node65 = (inp[10]) ? node67 : 3'b000;
									assign node67 = (inp[2]) ? 3'b100 : node68;
										assign node68 = (inp[3]) ? 3'b000 : 3'b100;
						assign node72 = (inp[8]) ? node74 : 3'b100;
							assign node74 = (inp[10]) ? node82 : node75;
								assign node75 = (inp[11]) ? 3'b100 : node76;
									assign node76 = (inp[3]) ? node78 : 3'b000;
										assign node78 = (inp[2]) ? 3'b000 : 3'b100;
								assign node82 = (inp[2]) ? 3'b000 : node83;
									assign node83 = (inp[11]) ? node85 : 3'b000;
										assign node85 = (inp[3]) ? 3'b100 : 3'b000;
				assign node89 = (inp[9]) ? node127 : node90;
					assign node90 = (inp[1]) ? node92 : 3'b100;
						assign node92 = (inp[11]) ? node110 : node93;
							assign node93 = (inp[8]) ? 3'b100 : node94;
								assign node94 = (inp[3]) ? node102 : node95;
									assign node95 = (inp[10]) ? 3'b100 : node96;
										assign node96 = (inp[7]) ? node98 : 3'b100;
											assign node98 = (inp[2]) ? 3'b100 : 3'b000;
									assign node102 = (inp[10]) ? node104 : 3'b000;
										assign node104 = (inp[7]) ? node106 : 3'b100;
											assign node106 = (inp[2]) ? 3'b100 : 3'b000;
							assign node110 = (inp[8]) ? node112 : 3'b000;
								assign node112 = (inp[10]) ? node120 : node113;
									assign node113 = (inp[3]) ? 3'b000 : node114;
										assign node114 = (inp[7]) ? node116 : 3'b100;
											assign node116 = (inp[2]) ? 3'b100 : 3'b000;
									assign node120 = (inp[7]) ? node122 : 3'b100;
										assign node122 = (inp[2]) ? 3'b100 : node123;
											assign node123 = (inp[3]) ? 3'b000 : 3'b100;
					assign node127 = (inp[11]) ? node171 : node128;
						assign node128 = (inp[10]) ? node158 : node129;
							assign node129 = (inp[1]) ? node141 : node130;
								assign node130 = (inp[3]) ? node136 : node131;
									assign node131 = (inp[2]) ? 3'b101 : node132;
										assign node132 = (inp[8]) ? 3'b000 : 3'b001;
									assign node136 = (inp[2]) ? 3'b001 : node137;
										assign node137 = (inp[8]) ? 3'b100 : 3'b001;
								assign node141 = (inp[8]) ? node149 : node142;
									assign node142 = (inp[7]) ? node144 : 3'b100;
										assign node144 = (inp[3]) ? node146 : 3'b100;
											assign node146 = (inp[5]) ? 3'b100 : 3'b000;
									assign node149 = (inp[2]) ? node155 : node150;
										assign node150 = (inp[3]) ? node152 : 3'b101;
											assign node152 = (inp[7]) ? 3'b001 : 3'b101;
										assign node155 = (inp[3]) ? 3'b000 : 3'b100;
							assign node158 = (inp[8]) ? node166 : node159;
								assign node159 = (inp[2]) ? 3'b101 : node160;
									assign node160 = (inp[3]) ? node162 : 3'b001;
										assign node162 = (inp[1]) ? 3'b001 : 3'b101;
								assign node166 = (inp[2]) ? 3'b000 : node167;
									assign node167 = (inp[7]) ? 3'b011 : 3'b111;
						assign node171 = (inp[2]) ? node197 : node172;
							assign node172 = (inp[10]) ? node186 : node173;
								assign node173 = (inp[1]) ? node181 : node174;
									assign node174 = (inp[8]) ? node176 : 3'b100;
										assign node176 = (inp[3]) ? 3'b000 : node177;
											assign node177 = (inp[7]) ? 3'b000 : 3'b100;
									assign node181 = (inp[8]) ? node183 : 3'b000;
										assign node183 = (inp[3]) ? 3'b101 : 3'b001;
								assign node186 = (inp[8]) ? node194 : node187;
									assign node187 = (inp[1]) ? 3'b100 : node188;
										assign node188 = (inp[3]) ? node190 : 3'b101;
											assign node190 = (inp[5]) ? 3'b101 : 3'b001;
									assign node194 = (inp[7]) ? 3'b010 : 3'b110;
							assign node197 = (inp[8]) ? node205 : node198;
								assign node198 = (inp[10]) ? 3'b001 : node199;
									assign node199 = (inp[1]) ? node201 : 3'b001;
										assign node201 = (inp[3]) ? 3'b000 : 3'b100;
								assign node205 = (inp[10]) ? 3'b000 : node206;
									assign node206 = (inp[1]) ? node210 : node207;
										assign node207 = (inp[3]) ? 3'b001 : 3'b101;
										assign node210 = (inp[3]) ? 3'b000 : 3'b100;
			assign node214 = (inp[9]) ? node216 : 3'b000;
				assign node216 = (inp[1]) ? node292 : node217;
					assign node217 = (inp[8]) ? node251 : node218;
						assign node218 = (inp[11]) ? node242 : node219;
							assign node219 = (inp[10]) ? node233 : node220;
								assign node220 = (inp[4]) ? node228 : node221;
									assign node221 = (inp[3]) ? 3'b000 : node222;
										assign node222 = (inp[7]) ? node224 : 3'b100;
											assign node224 = (inp[2]) ? 3'b100 : 3'b000;
									assign node228 = (inp[2]) ? 3'b000 : node229;
										assign node229 = (inp[3]) ? 3'b100 : 3'b000;
								assign node233 = (inp[2]) ? 3'b100 : node234;
									assign node234 = (inp[7]) ? 3'b000 : node235;
										assign node235 = (inp[3]) ? node237 : 3'b100;
											assign node237 = (inp[4]) ? 3'b000 : 3'b100;
							assign node242 = (inp[4]) ? node244 : 3'b000;
								assign node244 = (inp[10]) ? node246 : 3'b100;
									assign node246 = (inp[2]) ? 3'b000 : node247;
										assign node247 = (inp[3]) ? 3'b100 : 3'b000;
						assign node251 = (inp[4]) ? node269 : node252;
							assign node252 = (inp[11]) ? node254 : 3'b100;
								assign node254 = (inp[3]) ? node262 : node255;
									assign node255 = (inp[7]) ? node257 : 3'b100;
										assign node257 = (inp[5]) ? 3'b100 : node258;
											assign node258 = (inp[2]) ? 3'b100 : 3'b000;
									assign node262 = (inp[10]) ? node264 : 3'b000;
										assign node264 = (inp[2]) ? 3'b100 : node265;
											assign node265 = (inp[7]) ? 3'b000 : 3'b100;
							assign node269 = (inp[10]) ? node283 : node270;
								assign node270 = (inp[3]) ? node278 : node271;
									assign node271 = (inp[2]) ? 3'b101 : node272;
										assign node272 = (inp[11]) ? 3'b100 : node273;
											assign node273 = (inp[7]) ? 3'b001 : 3'b101;
									assign node278 = (inp[11]) ? node280 : 3'b001;
										assign node280 = (inp[2]) ? 3'b001 : 3'b000;
								assign node283 = (inp[2]) ? 3'b000 : node284;
									assign node284 = (inp[7]) ? node288 : node285;
										assign node285 = (inp[11]) ? 3'b100 : 3'b101;
										assign node288 = (inp[11]) ? 3'b000 : 3'b001;
					assign node292 = (inp[4]) ? node294 : 3'b000;
						assign node294 = (inp[11]) ? node324 : node295;
							assign node295 = (inp[8]) ? node311 : node296;
								assign node296 = (inp[3]) ? node304 : node297;
									assign node297 = (inp[10]) ? 3'b100 : node298;
										assign node298 = (inp[7]) ? node300 : 3'b100;
											assign node300 = (inp[5]) ? 3'b100 : 3'b000;
									assign node304 = (inp[10]) ? node306 : 3'b000;
										assign node306 = (inp[2]) ? 3'b100 : node307;
											assign node307 = (inp[7]) ? 3'b000 : 3'b100;
								assign node311 = (inp[2]) ? node319 : node312;
									assign node312 = (inp[10]) ? node316 : node313;
										assign node313 = (inp[3]) ? 3'b100 : 3'b000;
										assign node316 = (inp[7]) ? 3'b001 : 3'b101;
									assign node319 = (inp[3]) ? 3'b000 : node320;
										assign node320 = (inp[10]) ? 3'b000 : 3'b100;
							assign node324 = (inp[8]) ? node326 : 3'b000;
								assign node326 = (inp[7]) ? node338 : node327;
									assign node327 = (inp[2]) ? node333 : node328;
										assign node328 = (inp[10]) ? 3'b100 : node329;
											assign node329 = (inp[3]) ? 3'b000 : 3'b100;
										assign node333 = (inp[10]) ? 3'b000 : node334;
											assign node334 = (inp[3]) ? 3'b000 : 3'b100;
									assign node338 = (inp[3]) ? 3'b000 : node339;
										assign node339 = (inp[2]) ? node341 : 3'b000;
											assign node341 = (inp[10]) ? 3'b000 : 3'b100;

endmodule