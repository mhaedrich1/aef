module dtc_split125_bm57 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node282;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node351;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node396;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node414;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node446;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node471;
	wire [3-1:0] node473;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node503;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node519;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node545;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node577;

	assign outp = (inp[6]) ? node322 : node1;
		assign node1 = (inp[4]) ? node173 : node2;
			assign node2 = (inp[5]) ? node88 : node3;
				assign node3 = (inp[8]) ? node51 : node4;
					assign node4 = (inp[1]) ? node24 : node5;
						assign node5 = (inp[9]) ? node11 : node6;
							assign node6 = (inp[3]) ? node8 : 3'b011;
								assign node8 = (inp[11]) ? 3'b011 : 3'b001;
							assign node11 = (inp[11]) ? node19 : node12;
								assign node12 = (inp[3]) ? node16 : node13;
									assign node13 = (inp[0]) ? 3'b010 : 3'b011;
									assign node16 = (inp[0]) ? 3'b010 : 3'b000;
								assign node19 = (inp[0]) ? 3'b000 : node20;
									assign node20 = (inp[3]) ? 3'b000 : 3'b001;
						assign node24 = (inp[0]) ? node42 : node25;
							assign node25 = (inp[7]) ? node33 : node26;
								assign node26 = (inp[11]) ? 3'b010 : node27;
									assign node27 = (inp[9]) ? 3'b000 : node28;
										assign node28 = (inp[10]) ? 3'b010 : 3'b000;
								assign node33 = (inp[3]) ? node37 : node34;
									assign node34 = (inp[2]) ? 3'b010 : 3'b011;
									assign node37 = (inp[11]) ? 3'b011 : node38;
										assign node38 = (inp[9]) ? 3'b001 : 3'b000;
							assign node42 = (inp[9]) ? node46 : node43;
								assign node43 = (inp[2]) ? 3'b000 : 3'b001;
								assign node46 = (inp[7]) ? 3'b000 : node47;
									assign node47 = (inp[2]) ? 3'b011 : 3'b010;
					assign node51 = (inp[7]) ? node77 : node52;
						assign node52 = (inp[3]) ? node66 : node53;
							assign node53 = (inp[9]) ? 3'b100 : node54;
								assign node54 = (inp[1]) ? node60 : node55;
									assign node55 = (inp[10]) ? node57 : 3'b100;
										assign node57 = (inp[11]) ? 3'b101 : 3'b100;
									assign node60 = (inp[2]) ? node62 : 3'b101;
										assign node62 = (inp[11]) ? 3'b101 : 3'b100;
							assign node66 = (inp[2]) ? node74 : node67;
								assign node67 = (inp[10]) ? node69 : 3'b111;
									assign node69 = (inp[1]) ? 3'b110 : node70;
										assign node70 = (inp[11]) ? 3'b110 : 3'b110;
								assign node74 = (inp[1]) ? 3'b111 : 3'b110;
						assign node77 = (inp[3]) ? node83 : node78;
							assign node78 = (inp[10]) ? 3'b111 : node79;
								assign node79 = (inp[1]) ? 3'b110 : 3'b111;
							assign node83 = (inp[11]) ? node85 : 3'b101;
								assign node85 = (inp[10]) ? 3'b100 : 3'b101;
				assign node88 = (inp[3]) ? node126 : node89;
					assign node89 = (inp[7]) ? node105 : node90;
						assign node90 = (inp[8]) ? node98 : node91;
							assign node91 = (inp[0]) ? node93 : 3'b110;
								assign node93 = (inp[11]) ? node95 : 3'b110;
									assign node95 = (inp[9]) ? 3'b110 : 3'b111;
							assign node98 = (inp[2]) ? 3'b100 : node99;
								assign node99 = (inp[1]) ? node101 : 3'b101;
									assign node101 = (inp[9]) ? 3'b100 : 3'b101;
						assign node105 = (inp[11]) ? node115 : node106;
							assign node106 = (inp[2]) ? 3'b111 : node107;
								assign node107 = (inp[8]) ? 3'b110 : node108;
									assign node108 = (inp[10]) ? 3'b111 : node109;
										assign node109 = (inp[0]) ? 3'b101 : 3'b100;
							assign node115 = (inp[1]) ? node121 : node116;
								assign node116 = (inp[8]) ? 3'b110 : node117;
									assign node117 = (inp[10]) ? 3'b110 : 3'b100;
								assign node121 = (inp[0]) ? 3'b111 : node122;
									assign node122 = (inp[9]) ? 3'b111 : 3'b110;
					assign node126 = (inp[7]) ? node146 : node127;
						assign node127 = (inp[8]) ? node141 : node128;
							assign node128 = (inp[2]) ? node134 : node129;
								assign node129 = (inp[11]) ? 3'b110 : node130;
									assign node130 = (inp[10]) ? 3'b100 : 3'b110;
								assign node134 = (inp[1]) ? 3'b101 : node135;
									assign node135 = (inp[9]) ? 3'b100 : node136;
										assign node136 = (inp[10]) ? 3'b111 : 3'b110;
							assign node141 = (inp[10]) ? 3'b111 : node142;
								assign node142 = (inp[0]) ? 3'b110 : 3'b111;
						assign node146 = (inp[10]) ? node160 : node147;
							assign node147 = (inp[8]) ? node153 : node148;
								assign node148 = (inp[2]) ? 3'b111 : node149;
									assign node149 = (inp[11]) ? 3'b110 : 3'b111;
								assign node153 = (inp[2]) ? 3'b101 : node154;
									assign node154 = (inp[9]) ? node156 : 3'b100;
										assign node156 = (inp[1]) ? 3'b101 : 3'b100;
							assign node160 = (inp[1]) ? node166 : node161;
								assign node161 = (inp[9]) ? 3'b101 : node162;
									assign node162 = (inp[8]) ? 3'b100 : 3'b101;
								assign node166 = (inp[2]) ? 3'b101 : node167;
									assign node167 = (inp[8]) ? 3'b100 : node168;
										assign node168 = (inp[11]) ? 3'b100 : 3'b100;
			assign node173 = (inp[8]) ? node263 : node174;
				assign node174 = (inp[5]) ? node228 : node175;
					assign node175 = (inp[7]) ? node201 : node176;
						assign node176 = (inp[0]) ? node192 : node177;
							assign node177 = (inp[3]) ? node187 : node178;
								assign node178 = (inp[2]) ? node182 : node179;
									assign node179 = (inp[11]) ? 3'b101 : 3'b100;
									assign node182 = (inp[10]) ? 3'b111 : node183;
										assign node183 = (inp[11]) ? 3'b111 : 3'b101;
								assign node187 = (inp[11]) ? 3'b111 : node188;
									assign node188 = (inp[2]) ? 3'b111 : 3'b110;
							assign node192 = (inp[2]) ? node196 : node193;
								assign node193 = (inp[3]) ? 3'b101 : 3'b111;
								assign node196 = (inp[10]) ? node198 : 3'b110;
									assign node198 = (inp[1]) ? 3'b100 : 3'b110;
						assign node201 = (inp[9]) ? node223 : node202;
							assign node202 = (inp[3]) ? node212 : node203;
								assign node203 = (inp[11]) ? 3'b111 : node204;
									assign node204 = (inp[10]) ? node208 : node205;
										assign node205 = (inp[2]) ? 3'b100 : 3'b100;
										assign node208 = (inp[1]) ? 3'b111 : 3'b110;
								assign node212 = (inp[11]) ? node218 : node213;
									assign node213 = (inp[1]) ? node215 : 3'b100;
										assign node215 = (inp[10]) ? 3'b111 : 3'b101;
									assign node218 = (inp[0]) ? 3'b100 : node219;
										assign node219 = (inp[1]) ? 3'b100 : 3'b101;
							assign node223 = (inp[10]) ? node225 : 3'b101;
								assign node225 = (inp[2]) ? 3'b100 : 3'b101;
					assign node228 = (inp[3]) ? node246 : node229;
						assign node229 = (inp[10]) ? node235 : node230;
							assign node230 = (inp[7]) ? node232 : 3'b001;
								assign node232 = (inp[2]) ? 3'b010 : 3'b011;
							assign node235 = (inp[7]) ? node241 : node236;
								assign node236 = (inp[9]) ? node238 : 3'b010;
									assign node238 = (inp[2]) ? 3'b011 : 3'b010;
								assign node241 = (inp[9]) ? 3'b001 : node242;
									assign node242 = (inp[2]) ? 3'b001 : 3'b000;
						assign node246 = (inp[10]) ? node252 : node247;
							assign node247 = (inp[7]) ? 3'b010 : node248;
								assign node248 = (inp[0]) ? 3'b000 : 3'b001;
							assign node252 = (inp[7]) ? node256 : node253;
								assign node253 = (inp[11]) ? 3'b010 : 3'b011;
								assign node256 = (inp[2]) ? node258 : 3'b001;
									assign node258 = (inp[9]) ? 3'b001 : node259;
										assign node259 = (inp[11]) ? 3'b000 : 3'b000;
				assign node263 = (inp[7]) ? node287 : node264;
					assign node264 = (inp[10]) ? node278 : node265;
						assign node265 = (inp[11]) ? node267 : 3'b011;
							assign node267 = (inp[2]) ? 3'b011 : node268;
								assign node268 = (inp[0]) ? node274 : node269;
									assign node269 = (inp[9]) ? node271 : 3'b010;
										assign node271 = (inp[1]) ? 3'b010 : 3'b011;
									assign node274 = (inp[3]) ? 3'b010 : 3'b011;
						assign node278 = (inp[3]) ? 3'b010 : node279;
							assign node279 = (inp[11]) ? 3'b011 : node280;
								assign node280 = (inp[2]) ? node282 : 3'b000;
									assign node282 = (inp[1]) ? 3'b011 : 3'b010;
					assign node287 = (inp[11]) ? node311 : node288;
						assign node288 = (inp[5]) ? node302 : node289;
							assign node289 = (inp[10]) ? node295 : node290;
								assign node290 = (inp[2]) ? node292 : 3'b010;
									assign node292 = (inp[1]) ? 3'b010 : 3'b011;
								assign node295 = (inp[3]) ? node297 : 3'b010;
									assign node297 = (inp[2]) ? 3'b011 : node298;
										assign node298 = (inp[9]) ? 3'b010 : 3'b011;
							assign node302 = (inp[0]) ? 3'b000 : node303;
								assign node303 = (inp[9]) ? 3'b001 : node304;
									assign node304 = (inp[2]) ? 3'b000 : node305;
										assign node305 = (inp[10]) ? 3'b001 : 3'b000;
						assign node311 = (inp[1]) ? node317 : node312;
							assign node312 = (inp[5]) ? 3'b001 : node313;
								assign node313 = (inp[10]) ? 3'b000 : 3'b001;
							assign node317 = (inp[10]) ? 3'b000 : node318;
								assign node318 = (inp[2]) ? 3'b000 : 3'b001;
		assign node322 = (inp[8]) ? node464 : node323;
			assign node323 = (inp[5]) ? node389 : node324;
				assign node324 = (inp[3]) ? node356 : node325;
					assign node325 = (inp[10]) ? node341 : node326;
						assign node326 = (inp[7]) ? node334 : node327;
							assign node327 = (inp[9]) ? node331 : node328;
								assign node328 = (inp[1]) ? 3'b101 : 3'b100;
								assign node331 = (inp[2]) ? 3'b100 : 3'b110;
							assign node334 = (inp[4]) ? node338 : node335;
								assign node335 = (inp[11]) ? 3'b101 : 3'b111;
								assign node338 = (inp[11]) ? 3'b111 : 3'b101;
						assign node341 = (inp[7]) ? node351 : node342;
							assign node342 = (inp[4]) ? 3'b111 : node343;
								assign node343 = (inp[1]) ? node345 : 3'b110;
									assign node345 = (inp[0]) ? 3'b111 : node346;
										assign node346 = (inp[2]) ? 3'b110 : 3'b110;
							assign node351 = (inp[4]) ? node353 : 3'b101;
								assign node353 = (inp[11]) ? 3'b101 : 3'b110;
					assign node356 = (inp[10]) ? node372 : node357;
						assign node357 = (inp[2]) ? node363 : node358;
							assign node358 = (inp[11]) ? 3'b110 : node359;
								assign node359 = (inp[9]) ? 3'b110 : 3'b100;
							assign node363 = (inp[0]) ? 3'b110 : node364;
								assign node364 = (inp[11]) ? 3'b111 : node365;
									assign node365 = (inp[4]) ? 3'b101 : node366;
										assign node366 = (inp[9]) ? 3'b111 : 3'b110;
						assign node372 = (inp[11]) ? node384 : node373;
							assign node373 = (inp[0]) ? node379 : node374;
								assign node374 = (inp[4]) ? node376 : 3'b110;
									assign node376 = (inp[2]) ? 3'b111 : 3'b110;
								assign node379 = (inp[9]) ? node381 : 3'b111;
									assign node381 = (inp[2]) ? 3'b101 : 3'b100;
							assign node384 = (inp[2]) ? 3'b100 : node385;
								assign node385 = (inp[0]) ? 3'b101 : 3'b100;
				assign node389 = (inp[10]) ? node441 : node390;
					assign node390 = (inp[4]) ? node424 : node391;
						assign node391 = (inp[0]) ? node411 : node392;
							assign node392 = (inp[2]) ? node400 : node393;
								assign node393 = (inp[11]) ? 3'b001 : node394;
									assign node394 = (inp[9]) ? node396 : 3'b000;
										assign node396 = (inp[1]) ? 3'b010 : 3'b000;
								assign node400 = (inp[9]) ? node406 : node401;
									assign node401 = (inp[1]) ? node403 : 3'b010;
										assign node403 = (inp[7]) ? 3'b000 : 3'b000;
									assign node406 = (inp[3]) ? 3'b001 : node407;
										assign node407 = (inp[11]) ? 3'b001 : 3'b010;
							assign node411 = (inp[3]) ? node419 : node412;
								assign node412 = (inp[11]) ? 3'b001 : node413;
									assign node413 = (inp[7]) ? 3'b000 : node414;
										assign node414 = (inp[9]) ? 3'b011 : 3'b010;
								assign node419 = (inp[1]) ? 3'b010 : node420;
									assign node420 = (inp[11]) ? 3'b011 : 3'b010;
						assign node424 = (inp[1]) ? node430 : node425;
							assign node425 = (inp[11]) ? node427 : 3'b011;
								assign node427 = (inp[9]) ? 3'b010 : 3'b011;
							assign node430 = (inp[11]) ? 3'b010 : node431;
								assign node431 = (inp[9]) ? node433 : 3'b010;
									assign node433 = (inp[3]) ? node437 : node434;
										assign node434 = (inp[7]) ? 3'b011 : 3'b010;
										assign node437 = (inp[0]) ? 3'b011 : 3'b010;
					assign node441 = (inp[4]) ? node457 : node442;
						assign node442 = (inp[3]) ? node450 : node443;
							assign node443 = (inp[7]) ? 3'b011 : node444;
								assign node444 = (inp[11]) ? node446 : 3'b000;
									assign node446 = (inp[2]) ? 3'b010 : 3'b011;
							assign node450 = (inp[11]) ? node454 : node451;
								assign node451 = (inp[9]) ? 3'b011 : 3'b010;
								assign node454 = (inp[9]) ? 3'b000 : 3'b001;
						assign node457 = (inp[0]) ? node461 : node458;
							assign node458 = (inp[7]) ? 3'b001 : 3'b000;
							assign node461 = (inp[11]) ? 3'b001 : 3'b000;
			assign node464 = (inp[4]) ? node534 : node465;
				assign node465 = (inp[3]) ? node493 : node466;
					assign node466 = (inp[5]) ? node476 : node467;
						assign node467 = (inp[11]) ? node471 : node468;
							assign node468 = (inp[9]) ? 3'b000 : 3'b001;
							assign node471 = (inp[10]) ? node473 : 3'b011;
								assign node473 = (inp[2]) ? 3'b011 : 3'b010;
						assign node476 = (inp[9]) ? node482 : node477;
							assign node477 = (inp[7]) ? 3'b011 : node478;
								assign node478 = (inp[2]) ? 3'b011 : 3'b010;
							assign node482 = (inp[7]) ? node490 : node483;
								assign node483 = (inp[0]) ? node485 : 3'b011;
									assign node485 = (inp[11]) ? 3'b011 : node486;
										assign node486 = (inp[10]) ? 3'b010 : 3'b010;
								assign node490 = (inp[11]) ? 3'b010 : 3'b011;
					assign node493 = (inp[5]) ? node515 : node494;
						assign node494 = (inp[11]) ? node508 : node495;
							assign node495 = (inp[10]) ? node503 : node496;
								assign node496 = (inp[9]) ? 3'b011 : node497;
									assign node497 = (inp[1]) ? 3'b010 : node498;
										assign node498 = (inp[2]) ? 3'b010 : 3'b011;
								assign node503 = (inp[9]) ? node505 : 3'b011;
									assign node505 = (inp[7]) ? 3'b011 : 3'b010;
							assign node508 = (inp[10]) ? node510 : 3'b000;
								assign node510 = (inp[7]) ? node512 : 3'b001;
									assign node512 = (inp[2]) ? 3'b001 : 3'b000;
						assign node515 = (inp[10]) ? node529 : node516;
							assign node516 = (inp[0]) ? node522 : node517;
								assign node517 = (inp[1]) ? node519 : 3'b000;
									assign node519 = (inp[2]) ? 3'b001 : 3'b000;
								assign node522 = (inp[7]) ? node524 : 3'b001;
									assign node524 = (inp[2]) ? node526 : 3'b001;
										assign node526 = (inp[1]) ? 3'b000 : 3'b000;
							assign node529 = (inp[9]) ? node531 : 3'b001;
								assign node531 = (inp[7]) ? 3'b000 : 3'b001;
				assign node534 = (inp[5]) ? node566 : node535;
					assign node535 = (inp[11]) ? node559 : node536;
						assign node536 = (inp[3]) ? node548 : node537;
							assign node537 = (inp[9]) ? node543 : node538;
								assign node538 = (inp[10]) ? node540 : 3'b010;
									assign node540 = (inp[2]) ? 3'b010 : 3'b011;
								assign node543 = (inp[10]) ? node545 : 3'b011;
									assign node545 = (inp[2]) ? 3'b010 : 3'b011;
							assign node548 = (inp[7]) ? 3'b011 : node549;
								assign node549 = (inp[0]) ? node551 : 3'b010;
									assign node551 = (inp[9]) ? node555 : node552;
										assign node552 = (inp[1]) ? 3'b011 : 3'b010;
										assign node555 = (inp[1]) ? 3'b010 : 3'b011;
						assign node559 = (inp[2]) ? 3'b000 : node560;
							assign node560 = (inp[3]) ? 3'b001 : node561;
								assign node561 = (inp[1]) ? 3'b001 : 3'b000;
					assign node566 = (inp[3]) ? node576 : node567;
						assign node567 = (inp[11]) ? node573 : node568;
							assign node568 = (inp[10]) ? 3'b001 : node569;
								assign node569 = (inp[7]) ? 3'b001 : 3'b000;
							assign node573 = (inp[7]) ? 3'b000 : 3'b001;
						assign node576 = (inp[10]) ? 3'b000 : node577;
							assign node577 = (inp[11]) ? 3'b000 : 3'b001;

endmodule