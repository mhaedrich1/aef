module dtc_split05_bm40 (
	input  wire [16-1:0] inp,
	output wire [40-1:0] outp
);

	wire [40-1:0] node1;
	wire [40-1:0] node2;
	wire [40-1:0] node4;
	wire [40-1:0] node5;
	wire [40-1:0] node7;
	wire [40-1:0] node8;
	wire [40-1:0] node9;
	wire [40-1:0] node15;
	wire [40-1:0] node16;
	wire [40-1:0] node19;
	wire [40-1:0] node20;
	wire [40-1:0] node21;
	wire [40-1:0] node22;
	wire [40-1:0] node23;
	wire [40-1:0] node26;
	wire [40-1:0] node29;
	wire [40-1:0] node30;
	wire [40-1:0] node33;
	wire [40-1:0] node36;
	wire [40-1:0] node37;
	wire [40-1:0] node38;
	wire [40-1:0] node41;
	wire [40-1:0] node44;
	wire [40-1:0] node45;
	wire [40-1:0] node48;
	wire [40-1:0] node51;
	wire [40-1:0] node52;
	wire [40-1:0] node53;
	wire [40-1:0] node54;
	wire [40-1:0] node57;
	wire [40-1:0] node60;
	wire [40-1:0] node61;
	wire [40-1:0] node64;
	wire [40-1:0] node67;
	wire [40-1:0] node68;
	wire [40-1:0] node69;
	wire [40-1:0] node72;
	wire [40-1:0] node75;
	wire [40-1:0] node76;
	wire [40-1:0] node79;
	wire [40-1:0] node82;
	wire [40-1:0] node83;
	wire [40-1:0] node85;
	wire [40-1:0] node88;
	wire [40-1:0] node89;
	wire [40-1:0] node90;
	wire [40-1:0] node91;
	wire [40-1:0] node92;
	wire [40-1:0] node93;
	wire [40-1:0] node96;
	wire [40-1:0] node100;
	wire [40-1:0] node101;
	wire [40-1:0] node102;
	wire [40-1:0] node104;
	wire [40-1:0] node106;
	wire [40-1:0] node107;
	wire [40-1:0] node111;
	wire [40-1:0] node112;
	wire [40-1:0] node113;
	wire [40-1:0] node114;
	wire [40-1:0] node118;
	wire [40-1:0] node119;
	wire [40-1:0] node122;
	wire [40-1:0] node126;
	wire [40-1:0] node128;
	wire [40-1:0] node130;
	wire [40-1:0] node132;
	wire [40-1:0] node134;
	wire [40-1:0] node137;
	wire [40-1:0] node138;
	wire [40-1:0] node139;
	wire [40-1:0] node140;
	wire [40-1:0] node143;
	wire [40-1:0] node145;
	wire [40-1:0] node146;
	wire [40-1:0] node148;
	wire [40-1:0] node149;
	wire [40-1:0] node152;
	wire [40-1:0] node155;
	wire [40-1:0] node157;
	wire [40-1:0] node160;
	wire [40-1:0] node162;
	wire [40-1:0] node164;
	wire [40-1:0] node165;
	wire [40-1:0] node167;
	wire [40-1:0] node170;
	wire [40-1:0] node172;
	wire [40-1:0] node175;
	wire [40-1:0] node176;
	wire [40-1:0] node177;
	wire [40-1:0] node180;
	wire [40-1:0] node183;
	wire [40-1:0] node185;
	wire [40-1:0] node186;
	wire [40-1:0] node188;
	wire [40-1:0] node189;
	wire [40-1:0] node192;
	wire [40-1:0] node194;
	wire [40-1:0] node195;
	wire [40-1:0] node199;
	wire [40-1:0] node200;
	wire [40-1:0] node202;
	wire [40-1:0] node205;
	wire [40-1:0] node208;
	wire [40-1:0] node210;
	wire [40-1:0] node211;
	wire [40-1:0] node212;
	wire [40-1:0] node213;
	wire [40-1:0] node214;
	wire [40-1:0] node215;
	wire [40-1:0] node217;
	wire [40-1:0] node220;
	wire [40-1:0] node221;
	wire [40-1:0] node223;
	wire [40-1:0] node226;
	wire [40-1:0] node229;
	wire [40-1:0] node230;
	wire [40-1:0] node231;
	wire [40-1:0] node232;
	wire [40-1:0] node233;
	wire [40-1:0] node238;
	wire [40-1:0] node241;
	wire [40-1:0] node242;
	wire [40-1:0] node245;
	wire [40-1:0] node247;
	wire [40-1:0] node250;
	wire [40-1:0] node252;
	wire [40-1:0] node253;
	wire [40-1:0] node254;
	wire [40-1:0] node255;
	wire [40-1:0] node258;
	wire [40-1:0] node261;
	wire [40-1:0] node262;
	wire [40-1:0] node263;
	wire [40-1:0] node266;
	wire [40-1:0] node269;
	wire [40-1:0] node271;
	wire [40-1:0] node274;
	wire [40-1:0] node275;
	wire [40-1:0] node276;
	wire [40-1:0] node279;
	wire [40-1:0] node282;
	wire [40-1:0] node283;
	wire [40-1:0] node284;
	wire [40-1:0] node288;
	wire [40-1:0] node289;
	wire [40-1:0] node293;
	wire [40-1:0] node294;
	wire [40-1:0] node295;
	wire [40-1:0] node296;
	wire [40-1:0] node297;
	wire [40-1:0] node303;
	wire [40-1:0] node304;
	wire [40-1:0] node306;
	wire [40-1:0] node308;
	wire [40-1:0] node309;
	wire [40-1:0] node310;
	wire [40-1:0] node314;
	wire [40-1:0] node317;
	wire [40-1:0] node318;
	wire [40-1:0] node320;
	wire [40-1:0] node323;
	wire [40-1:0] node324;
	wire [40-1:0] node325;
	wire [40-1:0] node327;
	wire [40-1:0] node330;
	wire [40-1:0] node333;
	wire [40-1:0] node336;
	wire [40-1:0] node337;
	wire [40-1:0] node338;
	wire [40-1:0] node340;
	wire [40-1:0] node342;
	wire [40-1:0] node343;
	wire [40-1:0] node347;
	wire [40-1:0] node348;
	wire [40-1:0] node349;
	wire [40-1:0] node351;
	wire [40-1:0] node355;
	wire [40-1:0] node356;
	wire [40-1:0] node357;
	wire [40-1:0] node358;
	wire [40-1:0] node361;
	wire [40-1:0] node362;
	wire [40-1:0] node368;
	wire [40-1:0] node369;
	wire [40-1:0] node370;
	wire [40-1:0] node372;
	wire [40-1:0] node374;
	wire [40-1:0] node375;
	wire [40-1:0] node379;
	wire [40-1:0] node380;
	wire [40-1:0] node381;
	wire [40-1:0] node384;
	wire [40-1:0] node385;
	wire [40-1:0] node386;
	wire [40-1:0] node389;
	wire [40-1:0] node392;
	wire [40-1:0] node396;
	wire [40-1:0] node397;
	wire [40-1:0] node398;
	wire [40-1:0] node400;
	wire [40-1:0] node402;
	wire [40-1:0] node404;
	wire [40-1:0] node407;
	wire [40-1:0] node410;
	wire [40-1:0] node412;
	wire [40-1:0] node413;
	wire [40-1:0] node415;
	wire [40-1:0] node416;

	assign outp = (inp[1]) ? node82 : node1;
		assign node1 = (inp[9]) ? node15 : node2;
			assign node2 = (inp[7]) ? node4 : 40'b0000000000000000000000000000000000000000;
				assign node4 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node5;
					assign node5 = (inp[4]) ? node7 : 40'b0000000000000000000000000000000000000000;
						assign node7 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node8;
							assign node8 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : node9;
								assign node9 = (inp[8]) ? 40'b0000000000000000100000000000000000000000 : 40'b0000000000000000000000000000000000000000;
			assign node15 = (inp[8]) ? node19 : node16;
				assign node16 = (inp[4]) ? 40'b0000000001000000000000000000000000000100 : 40'b0000000000000000000000000000000000000100;
				assign node19 = (inp[7]) ? node51 : node20;
					assign node20 = (inp[11]) ? node36 : node21;
						assign node21 = (inp[14]) ? node29 : node22;
							assign node22 = (inp[3]) ? node26 : node23;
								assign node23 = (inp[4]) ? 40'b0000000001000010010100100000001001000100 : 40'b0000000000000010010100100000001001000100;
								assign node26 = (inp[4]) ? 40'b0000000001000000010100100000001011000100 : 40'b0000000000000000010100100000001011000100;
							assign node29 = (inp[3]) ? node33 : node30;
								assign node30 = (inp[4]) ? 40'b0000000001001010010000100000001001000100 : 40'b0000000000001010010000100000001001000100;
								assign node33 = (inp[4]) ? 40'b0000000001001000010000100000001011000100 : 40'b0000000000001000010000100000001011000100;
						assign node36 = (inp[3]) ? node44 : node37;
							assign node37 = (inp[14]) ? node41 : node38;
								assign node38 = (inp[4]) ? 40'b0000000001000010010100100000000001000110 : 40'b0000000000000010010100100000000001000110;
								assign node41 = (inp[4]) ? 40'b0000000001001010010000100000000001000110 : 40'b0000000000001010010000100000000001000110;
							assign node44 = (inp[14]) ? node48 : node45;
								assign node45 = (inp[4]) ? 40'b0000000001000000010100100000000011000110 : 40'b0000000000000000010100100000000011000110;
								assign node48 = (inp[4]) ? 40'b0000000001001000010000100000000011000110 : 40'b0000000000001000010000100000000011000110;
					assign node51 = (inp[14]) ? node67 : node52;
						assign node52 = (inp[11]) ? node60 : node53;
							assign node53 = (inp[3]) ? node57 : node54;
								assign node54 = (inp[4]) ? 40'b0100000001000010000000101000001100000100 : 40'b0100000000000010000000101000001100000100;
								assign node57 = (inp[4]) ? 40'b0100000001000000000000101000001110000100 : 40'b0100000000000000000000101000001110000100;
							assign node60 = (inp[3]) ? node64 : node61;
								assign node61 = (inp[4]) ? 40'b0100000001000010000000101000000100000110 : 40'b0100000000000010000000101000000100000110;
								assign node64 = (inp[4]) ? 40'b0100000001000000000000101000000110000110 : 40'b0100000000000000000000101000000110000110;
						assign node67 = (inp[11]) ? node75 : node68;
							assign node68 = (inp[3]) ? node72 : node69;
								assign node69 = (inp[4]) ? 40'b0100000001000010000000100000001100000101 : 40'b0100000000000010000000100000001100000101;
								assign node72 = (inp[4]) ? 40'b0100000001000000000000100000001110000101 : 40'b0100000000000000000000100000001110000101;
							assign node75 = (inp[3]) ? node79 : node76;
								assign node76 = (inp[4]) ? 40'b0100000001000010000000100000000100000111 : 40'b0100000000000010000000100000000100000111;
								assign node79 = (inp[4]) ? 40'b0100000001000000000000100000000110000111 : 40'b0100000000000000000000100000000110000111;
		assign node82 = (inp[4]) ? node88 : node83;
			assign node83 = (inp[9]) ? node85 : 40'b0000000001000000000000000000000000000000;
				assign node85 = (inp[8]) ? 40'b0000000001000000000000000000000000000000 : 40'b0000100001000000000000000000000000000000;
			assign node88 = (inp[9]) ? node208 : node89;
				assign node89 = (inp[14]) ? node137 : node90;
					assign node90 = (inp[8]) ? node100 : node91;
						assign node91 = (inp[7]) ? 40'b0000000000000000000000000000000000000000 : node92;
							assign node92 = (inp[3]) ? node96 : node93;
								assign node93 = (inp[11]) ? 40'b0000000000000010000001000000000000000000 : 40'b0000000000000010000000000100000000000000;
								assign node96 = (inp[11]) ? 40'b0000000000000001010000000100000000000000 : 40'b0000000000100010000000000000000000000000;
						assign node100 = (inp[7]) ? node126 : node101;
							assign node101 = (inp[10]) ? node111 : node102;
								assign node102 = (inp[6]) ? node104 : 40'b0000000000000000000000000000000000000000;
									assign node104 = (inp[12]) ? node106 : 40'b0000000000000000000000000000000000000000;
										assign node106 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node107;
											assign node107 = (inp[3]) ? 40'b0000000000000010010000100000000000000010 : 40'b0000000000000000000000000000000000000000;
								assign node111 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node112;
									assign node112 = (inp[5]) ? node118 : node113;
										assign node113 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node114;
											assign node114 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000001000000000;
										assign node118 = (inp[12]) ? node122 : node119;
											assign node119 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000001000000000;
											assign node122 = (inp[6]) ? 40'b0000000000000000000000000000001000000000 : 40'b0000000000000000010000100000001010000000;
							assign node126 = (inp[10]) ? node128 : 40'b0000000000000000000000000000000000000000;
								assign node128 = (inp[13]) ? node130 : 40'b0000000000000000000000000000000000000000;
									assign node130 = (inp[3]) ? node132 : 40'b0000000000000000000000000000000000000000;
										assign node132 = (inp[0]) ? node134 : 40'b0000000000000000000000000000000000000000;
											assign node134 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000010000000100000000;
					assign node137 = (inp[8]) ? node175 : node138;
						assign node138 = (inp[7]) ? node160 : node139;
							assign node139 = (inp[11]) ? node143 : node140;
								assign node140 = (inp[3]) ? 40'b0000000000100000000000000000000010000000 : 40'b0000000000000000000000000100000010000000;
								assign node143 = (inp[3]) ? node145 : 40'b0000000000000000000001000000000010000000;
									assign node145 = (inp[6]) ? node155 : node146;
										assign node146 = (inp[0]) ? node148 : 40'b0000000000000000000000000000000000000000;
											assign node148 = (inp[10]) ? node152 : node149;
												assign node149 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010010000010000000000000000;
												assign node152 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000010000010000000010000000;
										assign node155 = (inp[12]) ? node157 : 40'b0000000000000000000000000000000000000000;
											assign node157 = (inp[0]) ? 40'b0000000000000010010000010000000000000000 : 40'b0000000000000000000000000000000000000000;
							assign node160 = (inp[11]) ? node162 : 40'b0000000000000000000000000000000000000000;
								assign node162 = (inp[3]) ? node164 : 40'b0000000000000000000000000000000000000000;
									assign node164 = (inp[10]) ? node170 : node165;
										assign node165 = (inp[13]) ? node167 : 40'b0000000000000000000000000000000000000000;
											assign node167 = (inp[0]) ? 40'b0000000000000010000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
										assign node170 = (inp[13]) ? node172 : 40'b0000000000000000000000010000000110000000;
											assign node172 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010000000010000000110000000;
						assign node175 = (inp[3]) ? node183 : node176;
							assign node176 = (inp[7]) ? node180 : node177;
								assign node177 = (inp[11]) ? 40'b0000000000001000010000100100000001000000 : 40'b0000000000000000010100100100000001000000;
								assign node180 = (inp[11]) ? 40'b0100000000000000000000100100000100000001 : 40'b0100000000000000000000101100000100000000;
							assign node183 = (inp[0]) ? node185 : 40'b0000000000000000000000000000000000000000;
								assign node185 = (inp[7]) ? node199 : node186;
									assign node186 = (inp[6]) ? node188 : 40'b0000000000000000000000000000000000000000;
										assign node188 = (inp[15]) ? node192 : node189;
											assign node189 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000010001000000000000000000001000010;
											assign node192 = (inp[11]) ? node194 : 40'b0000000010000010010100100000000001000000;
												assign node194 = (inp[13]) ? 40'b0000000010001000000000000000000001000010 : node195;
													assign node195 = (inp[2]) ? 40'b0000000000001001010000000000000001000010 : 40'b0000000010001001010000000000000001000000;
									assign node199 = (inp[10]) ? node205 : node200;
										assign node200 = (inp[6]) ? node202 : 40'b0000000000000000000000000000000000000000;
											assign node202 = (inp[12]) ? 40'b0100000000000001000000000000000100000011 : 40'b0000000000000000000000000000000000000000;
										assign node205 = (inp[2]) ? 40'b0100000000000000000000010000000100000001 : 40'b0100000000000000000000011000000100000000;
				assign node208 = (inp[8]) ? node210 : 40'b0000100000000000000000000000000000000000;
					assign node210 = (inp[7]) ? node336 : node211;
						assign node211 = (inp[3]) ? node293 : node212;
							assign node212 = (inp[14]) ? node250 : node213;
								assign node213 = (inp[0]) ? node229 : node214;
									assign node214 = (inp[6]) ? node220 : node215;
										assign node215 = (inp[11]) ? node217 : 40'b0001000000001001010110000010001000010000;
											assign node217 = (inp[13]) ? 40'b1001000000000001010110000010001000000000 : 40'b1001000000000101010110000010101000000000;
										assign node220 = (inp[10]) ? node226 : node221;
											assign node221 = (inp[5]) ? node223 : 40'b1001000000011101010010000010001000010000;
												assign node223 = (inp[11]) ? 40'b0001000000001101010010000011001000000000 : 40'b0001000000000101010010000001001000010000;
											assign node226 = (inp[15]) ? 40'b1001000000000001010010000001001000010000 : 40'b1001000000010001010010000001001000000000;
									assign node229 = (inp[15]) ? node241 : node230;
										assign node230 = (inp[11]) ? node238 : node231;
											assign node231 = (inp[5]) ? 40'b0000000000011001010110000010001000010000 : node232;
												assign node232 = (inp[6]) ? 40'b1000000000011101010010000010001000010000 : node233;
													assign node233 = (inp[12]) ? 40'b1000000000011001010010000010001000010000 : 40'b1000000000010001010010000000001000010000;
											assign node238 = (inp[10]) ? 40'b1000000000011001010010000010101000000000 : 40'b0000000000011101010010000010101000000000;
										assign node241 = (inp[10]) ? node245 : node242;
											assign node242 = (inp[11]) ? 40'b0000000000000101010110000010001000000000 : 40'b1000000000000101010110000010101000010000;
											assign node245 = (inp[5]) ? node247 : 40'b0000000000001001010010000010001000000000;
												assign node247 = (inp[6]) ? 40'b0000000000001001010010000011101000010000 : 40'b0000000000001001010110000010101000010000;
								assign node250 = (inp[11]) ? node252 : 40'b0000000000000000000000000000000000000000;
									assign node252 = (inp[10]) ? node274 : node253;
										assign node253 = (inp[5]) ? node261 : node254;
											assign node254 = (inp[15]) ? node258 : node255;
												assign node255 = (inp[2]) ? 40'b1001010000010100000000000001000000000000 : 40'b1001010000011100000000000010000000000000;
												assign node258 = (inp[2]) ? 40'b0001010000001100000000000011000000000000 : 40'b1000010000001100000000000010000000000000;
											assign node261 = (inp[6]) ? node269 : node262;
												assign node262 = (inp[0]) ? node266 : node263;
													assign node263 = (inp[12]) ? 40'b0001010000001100000100000010000000000000 : 40'b0001010000000100000100000010000000000000;
													assign node266 = (inp[15]) ? 40'b0000010000000100000100000010000000000000 : 40'b0000010000010100000100000010000000000000;
												assign node269 = (inp[2]) ? node271 : 40'b1000010000000100000000000001100000000000;
													assign node271 = (inp[12]) ? 40'b0001010000000100000000000001000000000000 : 40'b0001010000000100000100000011100000000000;
										assign node274 = (inp[15]) ? node282 : node275;
											assign node275 = (inp[5]) ? node279 : node276;
												assign node276 = (inp[12]) ? 40'b1001010000010000000000000001000000000000 : 40'b1001010000010000000100000010000000000000;
												assign node279 = (inp[2]) ? 40'b0000010000010000000100000011000000000000 : 40'b1000010000010000000100000010000000000000;
											assign node282 = (inp[12]) ? node288 : node283;
												assign node283 = (inp[2]) ? 40'b1000010000000000000100000010000000000000 : node284;
													assign node284 = (inp[13]) ? 40'b1001010000000000000000000000000000000000 : 40'b1000010000000000000000000000100000000000;
												assign node288 = (inp[6]) ? 40'b0000010000001000000000000011000000000000 : node289;
													assign node289 = (inp[0]) ? 40'b1000010000001000000000000010100000000000 : 40'b1001010000001000000000000010100000000000;
							assign node293 = (inp[11]) ? node303 : node294;
								assign node294 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node295;
									assign node295 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node296;
										assign node296 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : node297;
											assign node297 = (inp[12]) ? 40'b1000000000010100000000000001000000100000 : 40'b1000000000010100000100000010000000100000;
								assign node303 = (inp[14]) ? node317 : node304;
									assign node304 = (inp[5]) ? node306 : 40'b0000000000000000000000000000000000000000;
										assign node306 = (inp[12]) ? node308 : 40'b0000000000000000000000000000000000000000;
											assign node308 = (inp[15]) ? node314 : node309;
												assign node309 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node310;
													assign node310 = (inp[0]) ? 40'b1000000000010100001000000000000000010000 : 40'b0000000000000000000000000000000000000000;
												assign node314 = (inp[13]) ? 40'b0001000000000000001100000010000000010000 : 40'b0001000000000000001100000010100000010000;
									assign node317 = (inp[5]) ? node323 : node318;
										assign node318 = (inp[12]) ? node320 : 40'b0011000000001000000100000010000000000000;
											assign node320 = (inp[13]) ? 40'b0011000000011100000000000011000000000000 : 40'b0011000000011100000000000010100000000000;
										assign node323 = (inp[6]) ? node333 : node324;
											assign node324 = (inp[15]) ? node330 : node325;
												assign node325 = (inp[2]) ? node327 : 40'b1010000000010000000100000010000000000000;
													assign node327 = (inp[13]) ? 40'b0010000000010000000100000011000000000000 : 40'b0011000000010000000100000011100000000000;
												assign node330 = (inp[0]) ? 40'b0010000000000100000100000010100000000000 : 40'b0011000000000100000100000011000000000000;
											assign node333 = (inp[12]) ? 40'b0010000000000000000000000001100000000000 : 40'b1011000000010000000000000001000000000000;
						assign node336 = (inp[3]) ? node368 : node337;
							assign node337 = (inp[10]) ? node347 : node338;
								assign node338 = (inp[0]) ? node340 : 40'b0000000000000000000000000000000000000000;
									assign node340 = (inp[11]) ? node342 : 40'b0000000000000000000000000000000000000000;
										assign node342 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node343;
											assign node343 = (inp[6]) ? 40'b0000001000000100000100000010100000001000 : 40'b1000001000010100000000000000100000001000;
								assign node347 = (inp[15]) ? node355 : node348;
									assign node348 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : node349;
										assign node349 = (inp[13]) ? node351 : 40'b0000000000000000000000000000000000000000;
											assign node351 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000001100011000000100000010000000000000;
									assign node355 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node356;
										assign node356 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : node357;
											assign node357 = (inp[11]) ? node361 : node358;
												assign node358 = (inp[13]) ? 40'b1001001100001000000000000010000000000000 : 40'b0000000000000000000000000000000000000000;
												assign node361 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node362;
													assign node362 = (inp[13]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000000000000100000010100000001000;
							assign node368 = (inp[6]) ? node396 : node369;
								assign node369 = (inp[11]) ? node379 : node370;
									assign node370 = (inp[14]) ? node372 : 40'b0000000000000000000000000000000000000000;
										assign node372 = (inp[5]) ? node374 : 40'b1000001000000100000000000001000000000000;
											assign node374 = (inp[13]) ? 40'b0001001000010000000100000011000000000000 : node375;
												assign node375 = (inp[15]) ? 40'b1001001000000000000100000010100000000000 : 40'b1001001000010100000100000010100000000000;
									assign node379 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node380;
										assign node380 = (inp[5]) ? node384 : node381;
											assign node381 = (inp[2]) ? 40'b1000001000000000000000000001000000001000 : 40'b1000001000001100000000000010000000001000;
											assign node384 = (inp[12]) ? node392 : node385;
												assign node385 = (inp[0]) ? node389 : node386;
													assign node386 = (inp[10]) ? 40'b0001001000000000000100000010000000001000 : 40'b1001001000000100000100000010100000001000;
													assign node389 = (inp[15]) ? 40'b1000001000000000000100000010000000001000 : 40'b1000001000010000000100000010000000001000;
												assign node392 = (inp[13]) ? 40'b0000001000001000000100000010000000001000 : 40'b0000001000011000000100000010100000001000;
								assign node396 = (inp[5]) ? node410 : node397;
									assign node397 = (inp[13]) ? node407 : node398;
										assign node398 = (inp[0]) ? node400 : 40'b0001001000001000000100000010100000001000;
											assign node400 = (inp[14]) ? node402 : 40'b0000000000000000000000000000000000000000;
												assign node402 = (inp[10]) ? node404 : 40'b1000001000001100000000000010100000000000;
													assign node404 = (inp[2]) ? 40'b0000001000001000000100000010100000000000 : 40'b0000001000001000000000000010100000000000;
										assign node407 = (inp[10]) ? 40'b0001001000001000000000000011000000001000 : 40'b0000000000000000000000000000000000000000;
									assign node410 = (inp[0]) ? node412 : 40'b0000000000000000000000000000000000000000;
										assign node412 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node413;
											assign node413 = (inp[14]) ? node415 : 40'b1000001000000100000000000001100000001000;
												assign node415 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node416;
													assign node416 = (inp[10]) ? 40'b1000001000000000000000000001100000000000 : 40'b1000001000000100000000000001100000000000;

endmodule