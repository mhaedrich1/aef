module dtc_split875_bm67 (
	input  wire [10-1:0] inp,
	output wire [77-1:0] outp
);

	wire [77-1:0] node1;
	wire [77-1:0] node2;
	wire [77-1:0] node5;
	wire [77-1:0] node8;
	wire [77-1:0] node9;
	wire [77-1:0] node12;

	assign outp = (inp[8]) ? node8 : node1;
		assign node1 = (inp[1]) ? node5 : node2;
			assign node2 = (inp[6]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000100000000000 : 77'b10100010000000000001000111000000000000000000100000010100011010000110000000000;
			assign node5 = (inp[0]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000;
		assign node8 = (inp[7]) ? node12 : node9;
			assign node9 = (inp[1]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000000000000000010000000000000000000000000000000000000010000100100000000;
			assign node12 = (inp[9]) ? 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000 : 77'b00000000000000000000000000000000000000000000000000000000000000000000000000000;

endmodule