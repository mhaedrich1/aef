module dtc_split05_bm56 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node290;
	wire [3-1:0] node291;

	assign outp = (inp[11]) ? node160 : node1;
		assign node1 = (inp[2]) ? node81 : node2;
			assign node2 = (inp[7]) ? node48 : node3;
				assign node3 = (inp[9]) ? node31 : node4;
					assign node4 = (inp[0]) ? node20 : node5;
						assign node5 = (inp[6]) ? node15 : node6;
							assign node6 = (inp[5]) ? 3'b101 : node7;
								assign node7 = (inp[1]) ? node11 : node8;
									assign node8 = (inp[10]) ? 3'b001 : 3'b101;
									assign node11 = (inp[10]) ? 3'b101 : 3'b001;
							assign node15 = (inp[8]) ? 3'b011 : node16;
								assign node16 = (inp[5]) ? 3'b111 : 3'b011;
						assign node20 = (inp[1]) ? node24 : node21;
							assign node21 = (inp[10]) ? 3'b100 : 3'b001;
							assign node24 = (inp[6]) ? node26 : 3'b110;
								assign node26 = (inp[5]) ? node28 : 3'b110;
									assign node28 = (inp[8]) ? 3'b100 : 3'b110;
					assign node31 = (inp[6]) ? node41 : node32;
						assign node32 = (inp[10]) ? node34 : 3'b100;
							assign node34 = (inp[3]) ? 3'b011 : node35;
								assign node35 = (inp[8]) ? node37 : 3'b110;
									assign node37 = (inp[5]) ? 3'b110 : 3'b100;
						assign node41 = (inp[5]) ? node43 : 3'b100;
							assign node43 = (inp[0]) ? node45 : 3'b000;
								assign node45 = (inp[3]) ? 3'b100 : 3'b000;
				assign node48 = (inp[9]) ? node62 : node49;
					assign node49 = (inp[8]) ? node55 : node50;
						assign node50 = (inp[1]) ? node52 : 3'b010;
							assign node52 = (inp[5]) ? 3'b000 : 3'b100;
						assign node55 = (inp[0]) ? node59 : node56;
							assign node56 = (inp[10]) ? 3'b110 : 3'b010;
							assign node59 = (inp[10]) ? 3'b101 : 3'b111;
					assign node62 = (inp[1]) ? node70 : node63;
						assign node63 = (inp[10]) ? 3'b001 : node64;
							assign node64 = (inp[3]) ? 3'b110 : node65;
								assign node65 = (inp[5]) ? 3'b001 : 3'b011;
						assign node70 = (inp[5]) ? node78 : node71;
							assign node71 = (inp[6]) ? node75 : node72;
								assign node72 = (inp[10]) ? 3'b111 : 3'b011;
								assign node75 = (inp[4]) ? 3'b101 : 3'b010;
							assign node78 = (inp[3]) ? 3'b010 : 3'b011;
			assign node81 = (inp[8]) ? node119 : node82;
				assign node82 = (inp[6]) ? node102 : node83;
					assign node83 = (inp[0]) ? node91 : node84;
						assign node84 = (inp[4]) ? 3'b000 : node85;
							assign node85 = (inp[3]) ? node87 : 3'b010;
								assign node87 = (inp[5]) ? 3'b000 : 3'b010;
						assign node91 = (inp[1]) ? node95 : node92;
							assign node92 = (inp[9]) ? 3'b100 : 3'b110;
							assign node95 = (inp[5]) ? node97 : 3'b010;
								assign node97 = (inp[9]) ? node99 : 3'b001;
									assign node99 = (inp[4]) ? 3'b011 : 3'b010;
					assign node102 = (inp[4]) ? node116 : node103;
						assign node103 = (inp[10]) ? node107 : node104;
							assign node104 = (inp[1]) ? 3'b100 : 3'b001;
							assign node107 = (inp[5]) ? node109 : 3'b001;
								assign node109 = (inp[9]) ? node113 : node110;
									assign node110 = (inp[7]) ? 3'b001 : 3'b000;
									assign node113 = (inp[7]) ? 3'b000 : 3'b001;
						assign node116 = (inp[9]) ? 3'b111 : 3'b011;
				assign node119 = (inp[3]) ? node143 : node120;
					assign node120 = (inp[4]) ? node134 : node121;
						assign node121 = (inp[7]) ? node127 : node122;
							assign node122 = (inp[9]) ? node124 : 3'b100;
								assign node124 = (inp[0]) ? 3'b101 : 3'b100;
							assign node127 = (inp[5]) ? 3'b001 : node128;
								assign node128 = (inp[6]) ? 3'b101 : node129;
									assign node129 = (inp[10]) ? 3'b100 : 3'b100;
						assign node134 = (inp[5]) ? node136 : 3'b010;
							assign node136 = (inp[6]) ? node138 : 3'b010;
								assign node138 = (inp[10]) ? node140 : 3'b100;
									assign node140 = (inp[7]) ? 3'b000 : 3'b001;
					assign node143 = (inp[1]) ? node157 : node144;
						assign node144 = (inp[9]) ? node152 : node145;
							assign node145 = (inp[7]) ? node149 : node146;
								assign node146 = (inp[5]) ? 3'b000 : 3'b100;
								assign node149 = (inp[5]) ? 3'b001 : 3'b011;
							assign node152 = (inp[6]) ? node154 : 3'b011;
								assign node154 = (inp[0]) ? 3'b001 : 3'b011;
						assign node157 = (inp[4]) ? 3'b101 : 3'b111;
		assign node160 = (inp[8]) ? node234 : node161;
			assign node161 = (inp[6]) ? node191 : node162;
				assign node162 = (inp[10]) ? node174 : node163;
					assign node163 = (inp[7]) ? node169 : node164;
						assign node164 = (inp[4]) ? 3'b001 : node165;
							assign node165 = (inp[5]) ? 3'b001 : 3'b011;
						assign node169 = (inp[3]) ? 3'b000 : node170;
							assign node170 = (inp[4]) ? 3'b000 : 3'b010;
					assign node174 = (inp[5]) ? node184 : node175;
						assign node175 = (inp[9]) ? 3'b100 : node176;
							assign node176 = (inp[1]) ? node178 : 3'b110;
								assign node178 = (inp[3]) ? node180 : 3'b100;
									assign node180 = (inp[4]) ? 3'b110 : 3'b100;
						assign node184 = (inp[4]) ? node188 : node185;
							assign node185 = (inp[1]) ? 3'b100 : 3'b101;
							assign node188 = (inp[0]) ? 3'b110 : 3'b111;
				assign node191 = (inp[10]) ? node205 : node192;
					assign node192 = (inp[0]) ? node200 : node193;
						assign node193 = (inp[3]) ? node197 : node194;
							assign node194 = (inp[1]) ? 3'b110 : 3'b111;
							assign node197 = (inp[4]) ? 3'b110 : 3'b100;
						assign node200 = (inp[7]) ? node202 : 3'b100;
							assign node202 = (inp[3]) ? 3'b100 : 3'b110;
					assign node205 = (inp[4]) ? node215 : node206;
						assign node206 = (inp[5]) ? node210 : node207;
							assign node207 = (inp[3]) ? 3'b001 : 3'b011;
							assign node210 = (inp[2]) ? 3'b001 : node211;
								assign node211 = (inp[9]) ? 3'b000 : 3'b001;
						assign node215 = (inp[5]) ? node227 : node216;
							assign node216 = (inp[3]) ? node222 : node217;
								assign node217 = (inp[7]) ? node219 : 3'b000;
									assign node219 = (inp[9]) ? 3'b001 : 3'b000;
								assign node222 = (inp[7]) ? 3'b011 : node223;
									assign node223 = (inp[9]) ? 3'b011 : 3'b010;
							assign node227 = (inp[7]) ? node231 : node228;
								assign node228 = (inp[1]) ? 3'b011 : 3'b010;
								assign node231 = (inp[9]) ? 3'b010 : 3'b011;
			assign node234 = (inp[3]) ? node260 : node235;
				assign node235 = (inp[7]) ? node241 : node236;
					assign node236 = (inp[9]) ? node238 : 3'b110;
						assign node238 = (inp[2]) ? 3'b011 : 3'b001;
					assign node241 = (inp[10]) ? node251 : node242;
						assign node242 = (inp[0]) ? node244 : 3'b111;
							assign node244 = (inp[9]) ? node246 : 3'b111;
								assign node246 = (inp[5]) ? node248 : 3'b110;
									assign node248 = (inp[1]) ? 3'b110 : 3'b100;
						assign node251 = (inp[5]) ? node253 : 3'b100;
							assign node253 = (inp[6]) ? node257 : node254;
								assign node254 = (inp[4]) ? 3'b101 : 3'b111;
								assign node257 = (inp[4]) ? 3'b001 : 3'b011;
				assign node260 = (inp[4]) ? node276 : node261;
					assign node261 = (inp[10]) ? node269 : node262;
						assign node262 = (inp[6]) ? node266 : node263;
							assign node263 = (inp[7]) ? 3'b000 : 3'b001;
							assign node266 = (inp[9]) ? 3'b110 : 3'b111;
						assign node269 = (inp[6]) ? node271 : 3'b111;
							assign node271 = (inp[5]) ? node273 : 3'b011;
								assign node273 = (inp[9]) ? 3'b011 : 3'b010;
					assign node276 = (inp[6]) ? node290 : node277;
						assign node277 = (inp[10]) ? 3'b101 : node278;
							assign node278 = (inp[5]) ? node286 : node279;
								assign node279 = (inp[1]) ? node283 : node280;
									assign node280 = (inp[9]) ? 3'b010 : 3'b010;
									assign node283 = (inp[7]) ? 3'b011 : 3'b010;
								assign node286 = (inp[0]) ? 3'b001 : 3'b000;
						assign node290 = (inp[10]) ? 3'b000 : node291;
							assign node291 = (inp[9]) ? 3'b101 : 3'b100;

endmodule