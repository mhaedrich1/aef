module dtc_split33_bm40 (
	input  wire [16-1:0] inp,
	output wire [40-1:0] outp
);

	wire [40-1:0] node1;
	wire [40-1:0] node2;
	wire [40-1:0] node3;
	wire [40-1:0] node5;
	wire [40-1:0] node7;
	wire [40-1:0] node8;
	wire [40-1:0] node9;
	wire [40-1:0] node15;
	wire [40-1:0] node17;
	wire [40-1:0] node18;
	wire [40-1:0] node19;
	wire [40-1:0] node20;
	wire [40-1:0] node21;
	wire [40-1:0] node24;
	wire [40-1:0] node27;
	wire [40-1:0] node28;
	wire [40-1:0] node31;
	wire [40-1:0] node33;
	wire [40-1:0] node34;
	wire [40-1:0] node36;
	wire [40-1:0] node39;
	wire [40-1:0] node40;
	wire [40-1:0] node43;
	wire [40-1:0] node46;
	wire [40-1:0] node47;
	wire [40-1:0] node49;
	wire [40-1:0] node51;
	wire [40-1:0] node52;
	wire [40-1:0] node54;
	wire [40-1:0] node56;
	wire [40-1:0] node58;
	wire [40-1:0] node59;
	wire [40-1:0] node62;
	wire [40-1:0] node64;
	wire [40-1:0] node67;
	wire [40-1:0] node68;
	wire [40-1:0] node70;
	wire [40-1:0] node72;
	wire [40-1:0] node74;
	wire [40-1:0] node77;
	wire [40-1:0] node80;
	wire [40-1:0] node81;
	wire [40-1:0] node84;
	wire [40-1:0] node85;
	wire [40-1:0] node87;
	wire [40-1:0] node89;
	wire [40-1:0] node91;
	wire [40-1:0] node93;
	wire [40-1:0] node96;
	wire [40-1:0] node97;
	wire [40-1:0] node99;
	wire [40-1:0] node101;
	wire [40-1:0] node103;
	wire [40-1:0] node104;
	wire [40-1:0] node105;
	wire [40-1:0] node108;
	wire [40-1:0] node112;
	wire [40-1:0] node113;
	wire [40-1:0] node115;
	wire [40-1:0] node116;
	wire [40-1:0] node117;
	wire [40-1:0] node121;
	wire [40-1:0] node122;
	wire [40-1:0] node126;
	wire [40-1:0] node129;
	wire [40-1:0] node130;
	wire [40-1:0] node131;
	wire [40-1:0] node133;
	wire [40-1:0] node135;
	wire [40-1:0] node136;
	wire [40-1:0] node138;
	wire [40-1:0] node140;
	wire [40-1:0] node141;
	wire [40-1:0] node143;
	wire [40-1:0] node144;
	wire [40-1:0] node148;
	wire [40-1:0] node150;
	wire [40-1:0] node152;
	wire [40-1:0] node155;
	wire [40-1:0] node156;
	wire [40-1:0] node157;
	wire [40-1:0] node159;
	wire [40-1:0] node161;
	wire [40-1:0] node165;
	wire [40-1:0] node169;
	wire [40-1:0] node170;
	wire [40-1:0] node172;
	wire [40-1:0] node174;
	wire [40-1:0] node175;
	wire [40-1:0] node177;
	wire [40-1:0] node180;
	wire [40-1:0] node181;
	wire [40-1:0] node184;
	wire [40-1:0] node187;
	wire [40-1:0] node188;
	wire [40-1:0] node191;
	wire [40-1:0] node192;
	wire [40-1:0] node194;
	wire [40-1:0] node196;
	wire [40-1:0] node198;
	wire [40-1:0] node200;
	wire [40-1:0] node202;
	wire [40-1:0] node204;
	wire [40-1:0] node207;
	wire [40-1:0] node208;
	wire [40-1:0] node210;
	wire [40-1:0] node212;
	wire [40-1:0] node213;
	wire [40-1:0] node214;
	wire [40-1:0] node217;
	wire [40-1:0] node220;
	wire [40-1:0] node221;
	wire [40-1:0] node223;
	wire [40-1:0] node226;
	wire [40-1:0] node227;
	wire [40-1:0] node229;
	wire [40-1:0] node232;
	wire [40-1:0] node235;
	wire [40-1:0] node236;
	wire [40-1:0] node238;
	wire [40-1:0] node240;
	wire [40-1:0] node242;
	wire [40-1:0] node244;
	wire [40-1:0] node247;
	wire [40-1:0] node250;
	wire [40-1:0] node251;
	wire [40-1:0] node252;
	wire [40-1:0] node255;
	wire [40-1:0] node256;
	wire [40-1:0] node257;
	wire [40-1:0] node258;
	wire [40-1:0] node259;
	wire [40-1:0] node262;
	wire [40-1:0] node265;
	wire [40-1:0] node266;
	wire [40-1:0] node269;
	wire [40-1:0] node272;
	wire [40-1:0] node273;
	wire [40-1:0] node274;
	wire [40-1:0] node277;
	wire [40-1:0] node280;
	wire [40-1:0] node281;
	wire [40-1:0] node284;
	wire [40-1:0] node287;
	wire [40-1:0] node288;
	wire [40-1:0] node289;
	wire [40-1:0] node290;
	wire [40-1:0] node293;
	wire [40-1:0] node296;
	wire [40-1:0] node297;
	wire [40-1:0] node300;
	wire [40-1:0] node303;
	wire [40-1:0] node304;
	wire [40-1:0] node305;
	wire [40-1:0] node308;
	wire [40-1:0] node311;
	wire [40-1:0] node312;
	wire [40-1:0] node315;
	wire [40-1:0] node318;
	wire [40-1:0] node319;
	wire [40-1:0] node322;
	wire [40-1:0] node324;
	wire [40-1:0] node325;
	wire [40-1:0] node326;
	wire [40-1:0] node327;
	wire [40-1:0] node328;
	wire [40-1:0] node329;
	wire [40-1:0] node330;
	wire [40-1:0] node331;
	wire [40-1:0] node332;
	wire [40-1:0] node333;
	wire [40-1:0] node334;
	wire [40-1:0] node336;
	wire [40-1:0] node339;
	wire [40-1:0] node340;
	wire [40-1:0] node344;
	wire [40-1:0] node345;
	wire [40-1:0] node348;
	wire [40-1:0] node351;
	wire [40-1:0] node352;
	wire [40-1:0] node355;
	wire [40-1:0] node356;
	wire [40-1:0] node360;
	wire [40-1:0] node361;
	wire [40-1:0] node362;
	wire [40-1:0] node365;
	wire [40-1:0] node367;
	wire [40-1:0] node370;
	wire [40-1:0] node371;
	wire [40-1:0] node373;
	wire [40-1:0] node376;
	wire [40-1:0] node378;
	wire [40-1:0] node381;
	wire [40-1:0] node382;
	wire [40-1:0] node383;
	wire [40-1:0] node384;
	wire [40-1:0] node385;
	wire [40-1:0] node388;
	wire [40-1:0] node389;
	wire [40-1:0] node392;
	wire [40-1:0] node395;
	wire [40-1:0] node398;
	wire [40-1:0] node399;
	wire [40-1:0] node402;
	wire [40-1:0] node403;
	wire [40-1:0] node404;
	wire [40-1:0] node407;
	wire [40-1:0] node410;
	wire [40-1:0] node413;
	wire [40-1:0] node414;
	wire [40-1:0] node415;
	wire [40-1:0] node416;
	wire [40-1:0] node419;
	wire [40-1:0] node420;
	wire [40-1:0] node424;
	wire [40-1:0] node426;
	wire [40-1:0] node429;
	wire [40-1:0] node431;
	wire [40-1:0] node434;
	wire [40-1:0] node435;
	wire [40-1:0] node436;
	wire [40-1:0] node437;
	wire [40-1:0] node438;
	wire [40-1:0] node440;
	wire [40-1:0] node441;
	wire [40-1:0] node444;
	wire [40-1:0] node447;
	wire [40-1:0] node448;
	wire [40-1:0] node452;
	wire [40-1:0] node453;
	wire [40-1:0] node455;
	wire [40-1:0] node458;
	wire [40-1:0] node461;
	wire [40-1:0] node462;
	wire [40-1:0] node463;
	wire [40-1:0] node466;
	wire [40-1:0] node467;
	wire [40-1:0] node470;
	wire [40-1:0] node472;
	wire [40-1:0] node475;
	wire [40-1:0] node477;
	wire [40-1:0] node480;
	wire [40-1:0] node481;
	wire [40-1:0] node482;
	wire [40-1:0] node483;
	wire [40-1:0] node486;
	wire [40-1:0] node487;
	wire [40-1:0] node491;
	wire [40-1:0] node492;
	wire [40-1:0] node495;
	wire [40-1:0] node498;
	wire [40-1:0] node499;
	wire [40-1:0] node501;
	wire [40-1:0] node502;
	wire [40-1:0] node505;
	wire [40-1:0] node508;
	wire [40-1:0] node509;
	wire [40-1:0] node510;
	wire [40-1:0] node513;
	wire [40-1:0] node516;
	wire [40-1:0] node519;
	wire [40-1:0] node520;
	wire [40-1:0] node521;
	wire [40-1:0] node522;
	wire [40-1:0] node523;
	wire [40-1:0] node524;
	wire [40-1:0] node528;
	wire [40-1:0] node529;
	wire [40-1:0] node530;
	wire [40-1:0] node534;
	wire [40-1:0] node535;
	wire [40-1:0] node538;
	wire [40-1:0] node540;
	wire [40-1:0] node543;
	wire [40-1:0] node544;
	wire [40-1:0] node545;
	wire [40-1:0] node546;
	wire [40-1:0] node550;
	wire [40-1:0] node551;
	wire [40-1:0] node554;
	wire [40-1:0] node557;
	wire [40-1:0] node558;
	wire [40-1:0] node561;
	wire [40-1:0] node564;
	wire [40-1:0] node565;
	wire [40-1:0] node566;
	wire [40-1:0] node567;
	wire [40-1:0] node569;
	wire [40-1:0] node572;
	wire [40-1:0] node575;
	wire [40-1:0] node576;
	wire [40-1:0] node580;
	wire [40-1:0] node581;
	wire [40-1:0] node582;
	wire [40-1:0] node584;
	wire [40-1:0] node587;
	wire [40-1:0] node590;
	wire [40-1:0] node592;
	wire [40-1:0] node595;
	wire [40-1:0] node596;
	wire [40-1:0] node597;
	wire [40-1:0] node598;
	wire [40-1:0] node599;
	wire [40-1:0] node600;
	wire [40-1:0] node605;
	wire [40-1:0] node606;
	wire [40-1:0] node607;
	wire [40-1:0] node612;
	wire [40-1:0] node613;
	wire [40-1:0] node614;
	wire [40-1:0] node615;
	wire [40-1:0] node617;
	wire [40-1:0] node620;
	wire [40-1:0] node624;
	wire [40-1:0] node625;
	wire [40-1:0] node626;
	wire [40-1:0] node630;
	wire [40-1:0] node633;
	wire [40-1:0] node634;
	wire [40-1:0] node635;
	wire [40-1:0] node636;
	wire [40-1:0] node639;
	wire [40-1:0] node640;
	wire [40-1:0] node644;
	wire [40-1:0] node645;
	wire [40-1:0] node648;
	wire [40-1:0] node649;
	wire [40-1:0] node653;
	wire [40-1:0] node654;
	wire [40-1:0] node656;
	wire [40-1:0] node659;
	wire [40-1:0] node660;
	wire [40-1:0] node662;
	wire [40-1:0] node663;
	wire [40-1:0] node667;
	wire [40-1:0] node668;
	wire [40-1:0] node672;
	wire [40-1:0] node673;
	wire [40-1:0] node675;
	wire [40-1:0] node676;
	wire [40-1:0] node678;
	wire [40-1:0] node679;
	wire [40-1:0] node680;
	wire [40-1:0] node686;
	wire [40-1:0] node687;
	wire [40-1:0] node688;
	wire [40-1:0] node689;
	wire [40-1:0] node690;
	wire [40-1:0] node691;
	wire [40-1:0] node692;
	wire [40-1:0] node694;
	wire [40-1:0] node697;
	wire [40-1:0] node699;
	wire [40-1:0] node702;
	wire [40-1:0] node705;
	wire [40-1:0] node706;
	wire [40-1:0] node708;
	wire [40-1:0] node712;
	wire [40-1:0] node713;
	wire [40-1:0] node714;
	wire [40-1:0] node716;
	wire [40-1:0] node719;
	wire [40-1:0] node720;
	wire [40-1:0] node724;
	wire [40-1:0] node725;
	wire [40-1:0] node728;
	wire [40-1:0] node729;
	wire [40-1:0] node733;
	wire [40-1:0] node734;
	wire [40-1:0] node735;
	wire [40-1:0] node736;
	wire [40-1:0] node739;
	wire [40-1:0] node742;
	wire [40-1:0] node744;
	wire [40-1:0] node745;
	wire [40-1:0] node749;
	wire [40-1:0] node750;
	wire [40-1:0] node751;
	wire [40-1:0] node752;
	wire [40-1:0] node755;
	wire [40-1:0] node758;
	wire [40-1:0] node759;
	wire [40-1:0] node762;
	wire [40-1:0] node765;
	wire [40-1:0] node767;
	wire [40-1:0] node770;
	wire [40-1:0] node771;
	wire [40-1:0] node772;
	wire [40-1:0] node773;
	wire [40-1:0] node775;
	wire [40-1:0] node778;
	wire [40-1:0] node779;
	wire [40-1:0] node781;
	wire [40-1:0] node785;
	wire [40-1:0] node786;
	wire [40-1:0] node787;
	wire [40-1:0] node788;
	wire [40-1:0] node789;
	wire [40-1:0] node794;
	wire [40-1:0] node796;
	wire [40-1:0] node799;
	wire [40-1:0] node800;
	wire [40-1:0] node801;
	wire [40-1:0] node805;
	wire [40-1:0] node806;
	wire [40-1:0] node810;
	wire [40-1:0] node811;
	wire [40-1:0] node812;
	wire [40-1:0] node813;
	wire [40-1:0] node817;
	wire [40-1:0] node818;
	wire [40-1:0] node819;
	wire [40-1:0] node823;
	wire [40-1:0] node826;
	wire [40-1:0] node827;
	wire [40-1:0] node828;
	wire [40-1:0] node831;
	wire [40-1:0] node832;
	wire [40-1:0] node834;
	wire [40-1:0] node837;
	wire [40-1:0] node838;
	wire [40-1:0] node842;
	wire [40-1:0] node843;
	wire [40-1:0] node846;
	wire [40-1:0] node849;
	wire [40-1:0] node850;
	wire [40-1:0] node851;
	wire [40-1:0] node852;
	wire [40-1:0] node853;
	wire [40-1:0] node854;
	wire [40-1:0] node855;
	wire [40-1:0] node857;
	wire [40-1:0] node863;
	wire [40-1:0] node864;
	wire [40-1:0] node865;
	wire [40-1:0] node866;
	wire [40-1:0] node867;
	wire [40-1:0] node869;
	wire [40-1:0] node872;
	wire [40-1:0] node873;
	wire [40-1:0] node875;
	wire [40-1:0] node880;
	wire [40-1:0] node881;
	wire [40-1:0] node883;
	wire [40-1:0] node887;
	wire [40-1:0] node889;
	wire [40-1:0] node891;
	wire [40-1:0] node893;
	wire [40-1:0] node894;
	wire [40-1:0] node897;
	wire [40-1:0] node898;
	wire [40-1:0] node902;
	wire [40-1:0] node903;
	wire [40-1:0] node904;
	wire [40-1:0] node906;
	wire [40-1:0] node907;
	wire [40-1:0] node913;
	wire [40-1:0] node915;
	wire [40-1:0] node916;
	wire [40-1:0] node917;
	wire [40-1:0] node918;
	wire [40-1:0] node919;
	wire [40-1:0] node920;
	wire [40-1:0] node921;
	wire [40-1:0] node924;
	wire [40-1:0] node927;
	wire [40-1:0] node928;
	wire [40-1:0] node932;
	wire [40-1:0] node934;
	wire [40-1:0] node937;
	wire [40-1:0] node938;
	wire [40-1:0] node940;
	wire [40-1:0] node943;
	wire [40-1:0] node944;
	wire [40-1:0] node947;
	wire [40-1:0] node950;
	wire [40-1:0] node951;
	wire [40-1:0] node952;
	wire [40-1:0] node954;
	wire [40-1:0] node955;
	wire [40-1:0] node958;
	wire [40-1:0] node961;
	wire [40-1:0] node964;
	wire [40-1:0] node965;
	wire [40-1:0] node966;
	wire [40-1:0] node967;
	wire [40-1:0] node970;
	wire [40-1:0] node972;
	wire [40-1:0] node975;
	wire [40-1:0] node978;
	wire [40-1:0] node979;
	wire [40-1:0] node980;
	wire [40-1:0] node983;
	wire [40-1:0] node986;
	wire [40-1:0] node987;
	wire [40-1:0] node988;
	wire [40-1:0] node992;
	wire [40-1:0] node995;
	wire [40-1:0] node996;
	wire [40-1:0] node997;
	wire [40-1:0] node998;
	wire [40-1:0] node999;
	wire [40-1:0] node1000;
	wire [40-1:0] node1003;
	wire [40-1:0] node1007;
	wire [40-1:0] node1008;
	wire [40-1:0] node1011;
	wire [40-1:0] node1012;
	wire [40-1:0] node1015;
	wire [40-1:0] node1018;
	wire [40-1:0] node1019;
	wire [40-1:0] node1020;
	wire [40-1:0] node1021;
	wire [40-1:0] node1024;
	wire [40-1:0] node1027;
	wire [40-1:0] node1030;
	wire [40-1:0] node1031;
	wire [40-1:0] node1034;
	wire [40-1:0] node1036;
	wire [40-1:0] node1038;
	wire [40-1:0] node1041;
	wire [40-1:0] node1042;
	wire [40-1:0] node1043;
	wire [40-1:0] node1044;
	wire [40-1:0] node1045;
	wire [40-1:0] node1046;
	wire [40-1:0] node1051;
	wire [40-1:0] node1054;
	wire [40-1:0] node1055;
	wire [40-1:0] node1057;
	wire [40-1:0] node1060;
	wire [40-1:0] node1063;
	wire [40-1:0] node1064;
	wire [40-1:0] node1065;
	wire [40-1:0] node1068;
	wire [40-1:0] node1071;
	wire [40-1:0] node1072;
	wire [40-1:0] node1075;
	wire [40-1:0] node1078;
	wire [40-1:0] node1079;
	wire [40-1:0] node1080;
	wire [40-1:0] node1082;
	wire [40-1:0] node1083;
	wire [40-1:0] node1084;
	wire [40-1:0] node1086;
	wire [40-1:0] node1089;
	wire [40-1:0] node1090;
	wire [40-1:0] node1094;
	wire [40-1:0] node1095;
	wire [40-1:0] node1097;
	wire [40-1:0] node1100;
	wire [40-1:0] node1101;
	wire [40-1:0] node1105;
	wire [40-1:0] node1106;
	wire [40-1:0] node1107;
	wire [40-1:0] node1109;
	wire [40-1:0] node1111;
	wire [40-1:0] node1113;
	wire [40-1:0] node1114;
	wire [40-1:0] node1117;
	wire [40-1:0] node1120;
	wire [40-1:0] node1121;
	wire [40-1:0] node1122;
	wire [40-1:0] node1124;
	wire [40-1:0] node1126;
	wire [40-1:0] node1127;
	wire [40-1:0] node1128;
	wire [40-1:0] node1133;
	wire [40-1:0] node1134;
	wire [40-1:0] node1136;
	wire [40-1:0] node1138;
	wire [40-1:0] node1141;
	wire [40-1:0] node1142;
	wire [40-1:0] node1145;
	wire [40-1:0] node1148;
	wire [40-1:0] node1149;
	wire [40-1:0] node1150;
	wire [40-1:0] node1153;
	wire [40-1:0] node1154;
	wire [40-1:0] node1157;
	wire [40-1:0] node1160;
	wire [40-1:0] node1161;
	wire [40-1:0] node1163;
	wire [40-1:0] node1165;
	wire [40-1:0] node1167;
	wire [40-1:0] node1170;
	wire [40-1:0] node1171;
	wire [40-1:0] node1173;
	wire [40-1:0] node1174;
	wire [40-1:0] node1178;
	wire [40-1:0] node1182;
	wire [40-1:0] node1183;
	wire [40-1:0] node1185;
	wire [40-1:0] node1186;
	wire [40-1:0] node1187;
	wire [40-1:0] node1188;
	wire [40-1:0] node1189;
	wire [40-1:0] node1190;
	wire [40-1:0] node1191;
	wire [40-1:0] node1192;
	wire [40-1:0] node1196;
	wire [40-1:0] node1200;
	wire [40-1:0] node1203;
	wire [40-1:0] node1204;
	wire [40-1:0] node1205;
	wire [40-1:0] node1206;
	wire [40-1:0] node1208;
	wire [40-1:0] node1212;
	wire [40-1:0] node1215;
	wire [40-1:0] node1216;
	wire [40-1:0] node1219;
	wire [40-1:0] node1221;
	wire [40-1:0] node1224;
	wire [40-1:0] node1225;
	wire [40-1:0] node1226;
	wire [40-1:0] node1227;
	wire [40-1:0] node1228;
	wire [40-1:0] node1232;
	wire [40-1:0] node1234;
	wire [40-1:0] node1237;
	wire [40-1:0] node1238;
	wire [40-1:0] node1241;
	wire [40-1:0] node1243;
	wire [40-1:0] node1246;
	wire [40-1:0] node1247;
	wire [40-1:0] node1249;
	wire [40-1:0] node1252;
	wire [40-1:0] node1254;
	wire [40-1:0] node1255;
	wire [40-1:0] node1258;
	wire [40-1:0] node1261;
	wire [40-1:0] node1262;
	wire [40-1:0] node1263;
	wire [40-1:0] node1264;
	wire [40-1:0] node1265;
	wire [40-1:0] node1267;
	wire [40-1:0] node1271;
	wire [40-1:0] node1272;
	wire [40-1:0] node1276;
	wire [40-1:0] node1277;
	wire [40-1:0] node1278;
	wire [40-1:0] node1282;
	wire [40-1:0] node1285;
	wire [40-1:0] node1286;
	wire [40-1:0] node1287;
	wire [40-1:0] node1288;
	wire [40-1:0] node1289;
	wire [40-1:0] node1292;
	wire [40-1:0] node1294;
	wire [40-1:0] node1297;
	wire [40-1:0] node1299;
	wire [40-1:0] node1301;
	wire [40-1:0] node1304;
	wire [40-1:0] node1305;
	wire [40-1:0] node1307;
	wire [40-1:0] node1310;
	wire [40-1:0] node1311;
	wire [40-1:0] node1313;
	wire [40-1:0] node1317;
	wire [40-1:0] node1318;
	wire [40-1:0] node1319;
	wire [40-1:0] node1322;
	wire [40-1:0] node1323;
	wire [40-1:0] node1327;
	wire [40-1:0] node1328;
	wire [40-1:0] node1330;
	wire [40-1:0] node1332;
	wire [40-1:0] node1335;
	wire [40-1:0] node1336;
	wire [40-1:0] node1339;
	wire [40-1:0] node1342;
	wire [40-1:0] node1343;
	wire [40-1:0] node1344;
	wire [40-1:0] node1345;
	wire [40-1:0] node1346;
	wire [40-1:0] node1347;
	wire [40-1:0] node1350;
	wire [40-1:0] node1351;
	wire [40-1:0] node1352;
	wire [40-1:0] node1355;
	wire [40-1:0] node1359;
	wire [40-1:0] node1360;
	wire [40-1:0] node1361;
	wire [40-1:0] node1362;
	wire [40-1:0] node1363;
	wire [40-1:0] node1368;
	wire [40-1:0] node1371;
	wire [40-1:0] node1372;
	wire [40-1:0] node1373;
	wire [40-1:0] node1374;
	wire [40-1:0] node1378;
	wire [40-1:0] node1381;
	wire [40-1:0] node1382;
	wire [40-1:0] node1383;
	wire [40-1:0] node1387;
	wire [40-1:0] node1388;
	wire [40-1:0] node1392;
	wire [40-1:0] node1393;
	wire [40-1:0] node1394;
	wire [40-1:0] node1395;
	wire [40-1:0] node1398;
	wire [40-1:0] node1401;
	wire [40-1:0] node1402;
	wire [40-1:0] node1406;
	wire [40-1:0] node1407;
	wire [40-1:0] node1409;
	wire [40-1:0] node1412;
	wire [40-1:0] node1413;
	wire [40-1:0] node1416;
	wire [40-1:0] node1418;
	wire [40-1:0] node1420;
	wire [40-1:0] node1423;
	wire [40-1:0] node1424;
	wire [40-1:0] node1425;
	wire [40-1:0] node1426;
	wire [40-1:0] node1427;
	wire [40-1:0] node1428;
	wire [40-1:0] node1432;
	wire [40-1:0] node1435;
	wire [40-1:0] node1436;
	wire [40-1:0] node1437;
	wire [40-1:0] node1441;
	wire [40-1:0] node1444;
	wire [40-1:0] node1445;
	wire [40-1:0] node1446;
	wire [40-1:0] node1449;
	wire [40-1:0] node1451;
	wire [40-1:0] node1454;
	wire [40-1:0] node1455;
	wire [40-1:0] node1457;
	wire [40-1:0] node1459;
	wire [40-1:0] node1462;
	wire [40-1:0] node1465;
	wire [40-1:0] node1466;
	wire [40-1:0] node1467;
	wire [40-1:0] node1468;
	wire [40-1:0] node1469;
	wire [40-1:0] node1471;
	wire [40-1:0] node1474;
	wire [40-1:0] node1477;
	wire [40-1:0] node1478;
	wire [40-1:0] node1481;
	wire [40-1:0] node1483;
	wire [40-1:0] node1486;
	wire [40-1:0] node1488;
	wire [40-1:0] node1490;
	wire [40-1:0] node1491;
	wire [40-1:0] node1495;
	wire [40-1:0] node1496;
	wire [40-1:0] node1498;
	wire [40-1:0] node1499;
	wire [40-1:0] node1502;
	wire [40-1:0] node1505;
	wire [40-1:0] node1506;
	wire [40-1:0] node1509;
	wire [40-1:0] node1510;

	assign outp = (inp[9]) ? node250 : node1;
		assign node1 = (inp[1]) ? node15 : node2;
			assign node2 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node3;
				assign node3 = (inp[4]) ? node5 : 40'b0000000000000000000000000000000000000000;
					assign node5 = (inp[8]) ? node7 : 40'b0000000000000000000000000000000000000000;
						assign node7 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node8;
							assign node8 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : node9;
								assign node9 = (inp[7]) ? 40'b0000000000000000100000000000000000000000 : 40'b0000000000000000000000000000000000000000;
			assign node15 = (inp[4]) ? node17 : 40'b0000000001000000000000000000000000000000;
				assign node17 = (inp[7]) ? node129 : node18;
					assign node18 = (inp[8]) ? node46 : node19;
						assign node19 = (inp[14]) ? node27 : node20;
							assign node20 = (inp[3]) ? node24 : node21;
								assign node21 = (inp[11]) ? 40'b0000000000000010000001000000000000000000 : 40'b0000000000000010000000000100000000000000;
								assign node24 = (inp[11]) ? 40'b0000000000000001010000000100000000000000 : 40'b0000000000100010000000000000000000000000;
							assign node27 = (inp[3]) ? node31 : node28;
								assign node28 = (inp[11]) ? 40'b0000000000000000000001000000000010000000 : 40'b0000000000000000000000000100000010000000;
								assign node31 = (inp[11]) ? node33 : 40'b0000000000100000000000000000000010000000;
									assign node33 = (inp[0]) ? node39 : node34;
										assign node34 = (inp[10]) ? node36 : 40'b0000000000000000000000000000000000000000;
											assign node36 = (inp[13]) ? 40'b0000000000000010010000010000000010000000 : 40'b0000000000000000000000000000000000000000;
										assign node39 = (inp[13]) ? node43 : node40;
											assign node40 = (inp[10]) ? 40'b0000000000000000010000010000000010000000 : 40'b0000000000000000000000000000000000000000;
											assign node43 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010010000010000000000000000;
						assign node46 = (inp[14]) ? node80 : node47;
							assign node47 = (inp[3]) ? node49 : 40'b0000000000000000000000000000000000000000;
								assign node49 = (inp[0]) ? node51 : 40'b0000000000000000000000000000000000000000;
									assign node51 = (inp[13]) ? node67 : node52;
										assign node52 = (inp[6]) ? node54 : 40'b0000000000000000000000000000000000000000;
											assign node54 = (inp[12]) ? node56 : 40'b0000000000000000000000000000000000000000;
												assign node56 = (inp[15]) ? node58 : 40'b0000000000000000000000000000000000000000;
													assign node58 = (inp[10]) ? node62 : node59;
														assign node59 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000001010000000000010000000010;
														assign node62 = (inp[5]) ? node64 : 40'b0000000000000000000000000000000000000000;
															assign node64 = (inp[11]) ? 40'b0000000010000000010000100000010010000000 : 40'b0000000010000000010000100000000010000000;
										assign node67 = (inp[10]) ? node77 : node68;
											assign node68 = (inp[6]) ? node70 : 40'b0000000000000000000000000000000000000000;
												assign node70 = (inp[12]) ? node72 : 40'b0000000000000000000000000000000000000000;
													assign node72 = (inp[5]) ? node74 : 40'b0000000000000000000000000000000000000000;
														assign node74 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000010000010010000100000000000000000;
											assign node77 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000001000000000;
							assign node80 = (inp[3]) ? node84 : node81;
								assign node81 = (inp[11]) ? 40'b0000000000001000010000100100000001000000 : 40'b0000000000000000010100100100000001000000;
								assign node84 = (inp[0]) ? node96 : node85;
									assign node85 = (inp[12]) ? node87 : 40'b0000000000000000000000000000000000000000;
										assign node87 = (inp[10]) ? node89 : 40'b0000000000000000000000000000000000000000;
											assign node89 = (inp[2]) ? node91 : 40'b0000000000000000000000000000000000000000;
												assign node91 = (inp[15]) ? node93 : 40'b0000000000000000000000000000000000000000;
													assign node93 = (inp[6]) ? 40'b0000000000001000000000000000000001000000 : 40'b0000000000000000000000000000000000000000;
									assign node96 = (inp[13]) ? node112 : node97;
										assign node97 = (inp[12]) ? node99 : 40'b0000000000000000000000000000000000000000;
											assign node99 = (inp[15]) ? node101 : 40'b0000000000000000000000000000000000000000;
												assign node101 = (inp[5]) ? node103 : 40'b0000000000000000000000000000000000000000;
													assign node103 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node104;
														assign node104 = (inp[10]) ? node108 : node105;
															assign node105 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000001010100000000001001000000;
															assign node108 = (inp[2]) ? 40'b0000000000000000010100100000001011000000 : 40'b0000000010000000010100100000000011000000;
										assign node112 = (inp[10]) ? node126 : node113;
											assign node113 = (inp[6]) ? node115 : 40'b0000000000000000000000000000000000000000;
												assign node115 = (inp[5]) ? node121 : node116;
													assign node116 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node117;
														assign node117 = (inp[2]) ? 40'b0000000000000010010100100000000001000010 : 40'b0000000000000000000000000000000000000000;
													assign node121 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : node122;
														assign node122 = (inp[11]) ? 40'b0000000010001010010000100000000001000000 : 40'b0000000010000010010100100000000001000000;
											assign node126 = (inp[11]) ? 40'b0000000010001000000000000000000001000010 : 40'b0000000000000000000100000000001001000010;
					assign node129 = (inp[14]) ? node169 : node130;
						assign node130 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node131;
							assign node131 = (inp[0]) ? node133 : 40'b0000000000000000000000000000000000000000;
								assign node133 = (inp[8]) ? node135 : 40'b0000000000000000000000000000000000000000;
									assign node135 = (inp[13]) ? node155 : node136;
										assign node136 = (inp[12]) ? node138 : 40'b0000000000000000000000000000000000000000;
											assign node138 = (inp[15]) ? node140 : 40'b0000000000000000000000000000000000000000;
												assign node140 = (inp[10]) ? node148 : node141;
													assign node141 = (inp[3]) ? node143 : 40'b0000000000000000000000000000000000000000;
														assign node143 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : node144;
															assign node144 = (inp[5]) ? 40'b0000000010000001000000000000000100000000 : 40'b0000000000000000000000000000000000000000;
													assign node148 = (inp[2]) ? node150 : 40'b0000000010000000000000100000000110000000;
														assign node150 = (inp[6]) ? node152 : 40'b0000000000000000000000000000000000000000;
															assign node152 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000100000000110000010;
										assign node155 = (inp[3]) ? node165 : node156;
											assign node156 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node157;
												assign node157 = (inp[5]) ? node159 : 40'b0000000000000000000000000000000000000000;
													assign node159 = (inp[15]) ? node161 : 40'b0000000000000000000000000000000000000000;
														assign node161 = (inp[2]) ? 40'b0000000000000010000000100000001100000000 : 40'b0000000010000010000000100000000100000000;
											assign node165 = (inp[10]) ? 40'b0000000000000000000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
						assign node169 = (inp[8]) ? node187 : node170;
							assign node170 = (inp[3]) ? node172 : 40'b0000000000000000000000000000000000000000;
								assign node172 = (inp[11]) ? node174 : 40'b0000000000000000000000000000000000000000;
									assign node174 = (inp[10]) ? node180 : node175;
										assign node175 = (inp[13]) ? node177 : 40'b0000000000000000000000000000000000000000;
											assign node177 = (inp[0]) ? 40'b0000000000000010000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
										assign node180 = (inp[13]) ? node184 : node181;
											assign node181 = (inp[0]) ? 40'b0000000000000000000000010000000110000000 : 40'b0000000000000000000000000000000000000000;
											assign node184 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010000000010000000110000000;
							assign node187 = (inp[3]) ? node191 : node188;
								assign node188 = (inp[11]) ? 40'b0100000000000000000000100100000100000001 : 40'b0100000000000000000000101100000100000000;
								assign node191 = (inp[0]) ? node207 : node192;
									assign node192 = (inp[2]) ? node194 : 40'b0000000000000000000000000000000000000000;
										assign node194 = (inp[10]) ? node196 : 40'b0000000000000000000000000000000000000000;
											assign node196 = (inp[6]) ? node198 : 40'b0000000000000000000000000000000000000000;
												assign node198 = (inp[15]) ? node200 : 40'b0000000000000000000000000000000000000000;
													assign node200 = (inp[5]) ? node202 : 40'b0000000000000000000000000000000000000000;
														assign node202 = (inp[11]) ? node204 : 40'b0100000000000000000000001000010000000000;
															assign node204 = (inp[13]) ? 40'b0100000000000000000000000000010000000001 : 40'b0100000000000000000000000000000000000001;
									assign node207 = (inp[13]) ? node235 : node208;
										assign node208 = (inp[15]) ? node210 : 40'b0000000000000000000000000000000000000000;
											assign node210 = (inp[12]) ? node212 : 40'b0000000000000000000000000000000000000000;
												assign node212 = (inp[10]) ? node220 : node213;
													assign node213 = (inp[6]) ? node217 : node214;
														assign node214 = (inp[11]) ? 40'b0100000000000001000000000000001100000001 : 40'b0100000000000001000000001000001100000000;
														assign node217 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0100000000000001000000001000000100000010;
													assign node220 = (inp[6]) ? node226 : node221;
														assign node221 = (inp[5]) ? node223 : 40'b0000000000000000000000000000000000000000;
															assign node223 = (inp[11]) ? 40'b0100000000000000000000100000001110000001 : 40'b0000000000000000000000000000000000000000;
														assign node226 = (inp[5]) ? node232 : node227;
															assign node227 = (inp[2]) ? node229 : 40'b0000000000000000000000000000000000000000;
																assign node229 = (inp[11]) ? 40'b0100000000000000000000100000000110000011 : 40'b0100000000000000000000101000000110000010;
															assign node232 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0100000010000000000000100000000110000001;
										assign node235 = (inp[10]) ? node247 : node236;
											assign node236 = (inp[12]) ? node238 : 40'b0000000000000000000000000000000000000000;
												assign node238 = (inp[5]) ? node240 : 40'b0000000000000000000000000000000000000000;
													assign node240 = (inp[15]) ? node242 : 40'b0000000000000000000000000000000000000000;
														assign node242 = (inp[2]) ? node244 : 40'b0100000010000010000000100000000100000001;
															assign node244 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0100000000000010000000101000001100000000;
											assign node247 = (inp[11]) ? 40'b0100000000000000000000010000000100000001 : 40'b0100000000000000000000011000000100000000;
		assign node250 = (inp[1]) ? node318 : node251;
			assign node251 = (inp[8]) ? node255 : node252;
				assign node252 = (inp[4]) ? 40'b0000000001000000000000000000000000000100 : 40'b0000000000000000000000000000000000000100;
				assign node255 = (inp[7]) ? node287 : node256;
					assign node256 = (inp[3]) ? node272 : node257;
						assign node257 = (inp[11]) ? node265 : node258;
							assign node258 = (inp[14]) ? node262 : node259;
								assign node259 = (inp[4]) ? 40'b0000000001000010010100100000001001000100 : 40'b0000000000000010010100100000001001000100;
								assign node262 = (inp[4]) ? 40'b0000000001001010010000100000001001000100 : 40'b0000000000001010010000100000001001000100;
							assign node265 = (inp[14]) ? node269 : node266;
								assign node266 = (inp[4]) ? 40'b0000000001000010010100100000000001000110 : 40'b0000000000000010010100100000000001000110;
								assign node269 = (inp[4]) ? 40'b0000000001001010010000100000000001000110 : 40'b0000000000001010010000100000000001000110;
						assign node272 = (inp[11]) ? node280 : node273;
							assign node273 = (inp[14]) ? node277 : node274;
								assign node274 = (inp[4]) ? 40'b0000000001000000010100100000001011000100 : 40'b0000000000000000010100100000001011000100;
								assign node277 = (inp[4]) ? 40'b0000000001001000010000100000001011000100 : 40'b0000000000001000010000100000001011000100;
							assign node280 = (inp[14]) ? node284 : node281;
								assign node281 = (inp[4]) ? 40'b0000000001000000010100100000000011000110 : 40'b0000000000000000010100100000000011000110;
								assign node284 = (inp[4]) ? 40'b0000000001001000010000100000000011000110 : 40'b0000000000001000010000100000000011000110;
					assign node287 = (inp[3]) ? node303 : node288;
						assign node288 = (inp[14]) ? node296 : node289;
							assign node289 = (inp[11]) ? node293 : node290;
								assign node290 = (inp[4]) ? 40'b0100000001000010000000101000001100000100 : 40'b0100000000000010000000101000001100000100;
								assign node293 = (inp[4]) ? 40'b0100000001000010000000101000000100000110 : 40'b0100000000000010000000101000000100000110;
							assign node296 = (inp[11]) ? node300 : node297;
								assign node297 = (inp[4]) ? 40'b0100000001000010000000100000001100000101 : 40'b0100000000000010000000100000001100000101;
								assign node300 = (inp[4]) ? 40'b0100000001000010000000100000000100000111 : 40'b0100000000000010000000100000000100000111;
						assign node303 = (inp[11]) ? node311 : node304;
							assign node304 = (inp[14]) ? node308 : node305;
								assign node305 = (inp[4]) ? 40'b0100000001000000000000101000001110000100 : 40'b0100000000000000000000101000001110000100;
								assign node308 = (inp[4]) ? 40'b0100000001000000000000100000001110000101 : 40'b0100000000000000000000100000001110000101;
							assign node311 = (inp[14]) ? node315 : node312;
								assign node312 = (inp[4]) ? 40'b0100000001000000000000101000000110000110 : 40'b0100000000000000000000101000000110000110;
								assign node315 = (inp[4]) ? 40'b0100000001000000000000100000000110000111 : 40'b0100000000000000000000100000000110000111;
			assign node318 = (inp[4]) ? node322 : node319;
				assign node319 = (inp[8]) ? 40'b0000000001000000000000000000000000000000 : 40'b0000100001000000000000000000000000000000;
				assign node322 = (inp[8]) ? node324 : 40'b0000100000000000000000000000000000000000;
					assign node324 = (inp[7]) ? node1078 : node325;
						assign node325 = (inp[3]) ? node849 : node326;
							assign node326 = (inp[14]) ? node672 : node327;
								assign node327 = (inp[10]) ? node519 : node328;
									assign node328 = (inp[11]) ? node434 : node329;
										assign node329 = (inp[15]) ? node381 : node330;
											assign node330 = (inp[0]) ? node360 : node331;
												assign node331 = (inp[13]) ? node351 : node332;
													assign node332 = (inp[12]) ? node344 : node333;
														assign node333 = (inp[5]) ? node339 : node334;
															assign node334 = (inp[6]) ? node336 : 40'b1001000000010101010110000010101000010000;
																assign node336 = (inp[2]) ? 40'b0001000000011101010110000010101000010000 : 40'b1001000000011101010010000010101000010000;
															assign node339 = (inp[2]) ? 40'b0001000000010101010110000011101000010000 : node340;
																assign node340 = (inp[6]) ? 40'b1001000000010101010010000001101000010000 : 40'b1001000000010101010110000010101000010000;
														assign node344 = (inp[6]) ? node348 : node345;
															assign node345 = (inp[5]) ? 40'b0001000000011101010110000010101000010000 : 40'b1001000000011101010010000010101000010000;
															assign node348 = (inp[5]) ? 40'b0001000000011101010010000011101000010000 : 40'b0001000000011101010010000010101000010000;
													assign node351 = (inp[2]) ? node355 : node352;
														assign node352 = (inp[6]) ? 40'b0001000000011101010010000010001000010000 : 40'b1001000000011101010010000010001000010000;
														assign node355 = (inp[6]) ? 40'b0001000000011101010010000011001000010000 : node356;
															assign node356 = (inp[5]) ? 40'b0001000000010101010110000011001000010000 : 40'b1001000000010101010010000001001000010000;
												assign node360 = (inp[13]) ? node370 : node361;
													assign node361 = (inp[12]) ? node365 : node362;
														assign node362 = (inp[6]) ? 40'b1000000000010101010010000001101000010000 : 40'b1000000000010101010010000000101000010000;
														assign node365 = (inp[6]) ? node367 : 40'b0000000000010101010110000011101000010000;
															assign node367 = (inp[5]) ? 40'b0000000000011101010010000011101000010000 : 40'b0000000000011101010010000010101000010000;
													assign node370 = (inp[2]) ? node376 : node371;
														assign node371 = (inp[12]) ? node373 : 40'b1000000000011101010010000010001000010000;
															assign node373 = (inp[6]) ? 40'b0000000000011101010010000010001000010000 : 40'b0000000000011101010110000010001000010000;
														assign node376 = (inp[12]) ? node378 : 40'b0000000000010101010110000011001000010000;
															assign node378 = (inp[5]) ? 40'b0000000000010101010010000001001000010000 : 40'b0000000000011101010010000011001000010000;
											assign node381 = (inp[0]) ? node413 : node382;
												assign node382 = (inp[12]) ? node398 : node383;
													assign node383 = (inp[2]) ? node395 : node384;
														assign node384 = (inp[13]) ? node388 : node385;
															assign node385 = (inp[6]) ? 40'b1001000000001101010010000010101000010000 : 40'b1001000000000101010010000000101000010000;
															assign node388 = (inp[6]) ? node392 : node389;
																assign node389 = (inp[5]) ? 40'b1001000000000101010110000010001000010000 : 40'b1001000000000101010010000000001000010000;
																assign node392 = (inp[5]) ? 40'b1001000000000101010010000001001000010000 : 40'b1001000000001101010010000010001000010000;
														assign node395 = (inp[5]) ? 40'b0001000000000101010110000010101000010000 : 40'b1001000000000101010110000010101000010000;
													assign node398 = (inp[6]) ? node402 : node399;
														assign node399 = (inp[13]) ? 40'b0001000000000101010110000011001000010000 : 40'b0001000000000101010110000011101000010000;
														assign node402 = (inp[13]) ? node410 : node403;
															assign node403 = (inp[2]) ? node407 : node404;
																assign node404 = (inp[5]) ? 40'b0001000000001101010010000011101000010000 : 40'b0001000000001101010010000010101000010000;
																assign node407 = (inp[5]) ? 40'b0001000000000101010010000001101000010000 : 40'b0001000000001101010010000011101000010000;
															assign node410 = (inp[5]) ? 40'b0001000000000101010010000001001000010000 : 40'b0001000000001101010010000011001000010000;
												assign node413 = (inp[13]) ? node429 : node414;
													assign node414 = (inp[5]) ? node424 : node415;
														assign node415 = (inp[6]) ? node419 : node416;
															assign node416 = (inp[2]) ? 40'b1000000000000101010110000010101000010000 : 40'b1000000000000101010010000000101000010000;
															assign node419 = (inp[2]) ? 40'b0000000000001101010110000010101000010000 : node420;
																assign node420 = (inp[12]) ? 40'b0000000000001101010010000010101000010000 : 40'b1000000000001101010010000010101000010000;
														assign node424 = (inp[2]) ? node426 : 40'b0000000000001101010110000010101000010000;
															assign node426 = (inp[6]) ? 40'b0000000000000101010010000001101000010000 : 40'b0000000000000101010110000011101000010000;
													assign node429 = (inp[6]) ? node431 : 40'b1000000000001101010010000010001000010000;
														assign node431 = (inp[12]) ? 40'b0000000000001101010010000010001000010000 : 40'b1000000000001101010010000010001000010000;
										assign node434 = (inp[13]) ? node480 : node435;
											assign node435 = (inp[6]) ? node461 : node436;
												assign node436 = (inp[5]) ? node452 : node437;
													assign node437 = (inp[15]) ? node447 : node438;
														assign node438 = (inp[0]) ? node440 : 40'b1001000000010101010110000010101000000000;
															assign node440 = (inp[12]) ? node444 : node441;
																assign node441 = (inp[2]) ? 40'b1000000000010101010110000010101000000000 : 40'b1000000000010101010010000000101000000000;
																assign node444 = (inp[2]) ? 40'b1000000000010101010010000001101000000000 : 40'b1000000000011101010010000010101000000000;
														assign node447 = (inp[12]) ? 40'b1001000000000101010010000001101000000000 : node448;
															assign node448 = (inp[2]) ? 40'b1000000000000101010110000010101000000000 : 40'b1000000000000101010010000000101000000000;
													assign node452 = (inp[15]) ? node458 : node453;
														assign node453 = (inp[2]) ? node455 : 40'b0001000000011101010110000010101000000000;
															assign node455 = (inp[0]) ? 40'b0000000000010101010110000010101000000000 : 40'b0001000000010101010110000010101000000000;
														assign node458 = (inp[12]) ? 40'b0001000000000101010110000011101000000000 : 40'b1001000000000101010110000010101000000000;
												assign node461 = (inp[5]) ? node475 : node462;
													assign node462 = (inp[12]) ? node466 : node463;
														assign node463 = (inp[15]) ? 40'b0001000000001101010110000010101000000000 : 40'b0000000000011101010110000010101000000000;
														assign node466 = (inp[0]) ? node470 : node467;
															assign node467 = (inp[2]) ? 40'b0001000000011101010010000011101000000000 : 40'b0001000000011101010010000010101000000000;
															assign node470 = (inp[15]) ? node472 : 40'b0000000000011101010010000011101000000000;
																assign node472 = (inp[2]) ? 40'b0000000000001101010010000011101000000000 : 40'b0000000000001101010010000010101000000000;
													assign node475 = (inp[2]) ? node477 : 40'b0000000000011101010010000011101000000000;
														assign node477 = (inp[12]) ? 40'b0000000000010101010010000001101000000000 : 40'b0000000000010101010110000011101000000000;
											assign node480 = (inp[0]) ? node498 : node481;
												assign node481 = (inp[5]) ? node491 : node482;
													assign node482 = (inp[6]) ? node486 : node483;
														assign node483 = (inp[12]) ? 40'b1001000000010101010010000001001000000000 : 40'b1001000000010101010010000000001000000000;
														assign node486 = (inp[15]) ? 40'b1001000000001101010010000010001000000000 : node487;
															assign node487 = (inp[12]) ? 40'b0001000000011101010010000010001000000000 : 40'b1001000000011101010010000010001000000000;
													assign node491 = (inp[15]) ? node495 : node492;
														assign node492 = (inp[12]) ? 40'b0001000000010101010010000001001000000000 : 40'b0001000000010101010110000011001000000000;
														assign node495 = (inp[2]) ? 40'b0001000000000101010010000001001000000000 : 40'b1001000000000101010010000001001000000000;
												assign node498 = (inp[2]) ? node508 : node499;
													assign node499 = (inp[12]) ? node501 : 40'b1000000000010101010010000001001000000000;
														assign node501 = (inp[6]) ? node505 : node502;
															assign node502 = (inp[15]) ? 40'b1000000000001101010010000010001000000000 : 40'b1000000000011101010010000010001000000000;
															assign node505 = (inp[5]) ? 40'b0000000000011101010010000011001000000000 : 40'b0000000000011101010010000010001000000000;
													assign node508 = (inp[15]) ? node516 : node509;
														assign node509 = (inp[5]) ? node513 : node510;
															assign node510 = (inp[12]) ? 40'b1000000000010101010010000001001000000000 : 40'b1000000000010101010110000010001000000000;
															assign node513 = (inp[12]) ? 40'b0000000000010101010110000011001000000000 : 40'b0000000000010101010110000010001000000000;
														assign node516 = (inp[5]) ? 40'b0000000000000101010110000011001000000000 : 40'b0000000000001101010010000011001000000000;
									assign node519 = (inp[0]) ? node595 : node520;
										assign node520 = (inp[13]) ? node564 : node521;
											assign node521 = (inp[11]) ? node543 : node522;
												assign node522 = (inp[12]) ? node528 : node523;
													assign node523 = (inp[6]) ? 40'b0001000000010001010110000011101000010000 : node524;
														assign node524 = (inp[5]) ? 40'b1001000000010001010110000010101000010000 : 40'b1001000000000001010110000010101000010000;
													assign node528 = (inp[15]) ? node534 : node529;
														assign node529 = (inp[5]) ? 40'b0001000000010001010110000011101000010000 : node530;
															assign node530 = (inp[2]) ? 40'b0001000000011001010010000011101000010000 : 40'b0001000000011001010010000010101000010000;
														assign node534 = (inp[2]) ? node538 : node535;
															assign node535 = (inp[6]) ? 40'b0001000000001001010010000011101000010000 : 40'b0001000000001001010110000010101000010000;
															assign node538 = (inp[6]) ? node540 : 40'b1001000000000001010010000001101000010000;
																assign node540 = (inp[5]) ? 40'b0001000000000001010010000001101000010000 : 40'b0001000000001001010010000011101000010000;
												assign node543 = (inp[5]) ? node557 : node544;
													assign node544 = (inp[6]) ? node550 : node545;
														assign node545 = (inp[12]) ? 40'b1001000000000001010010000001101000000000 : node546;
															assign node546 = (inp[15]) ? 40'b1001000000000001010110000010101000000000 : 40'b1001000000010001010110000010101000000000;
														assign node550 = (inp[15]) ? node554 : node551;
															assign node551 = (inp[2]) ? 40'b0001000000011001010110000010101000000000 : 40'b1001000000011001010010000010101000000000;
															assign node554 = (inp[12]) ? 40'b0001000000001001010010000010101000000000 : 40'b0001000000001001010110000010101000000000;
													assign node557 = (inp[6]) ? node561 : node558;
														assign node558 = (inp[12]) ? 40'b0001000000010001010110000011101000000000 : 40'b0001000000010001010110000010101000000000;
														assign node561 = (inp[12]) ? 40'b0001000000010001010010000001101000000000 : 40'b1001000000010001010010000001101000000000;
											assign node564 = (inp[15]) ? node580 : node565;
												assign node565 = (inp[11]) ? node575 : node566;
													assign node566 = (inp[2]) ? node572 : node567;
														assign node567 = (inp[6]) ? node569 : 40'b0001000000011001010110000010001000010000;
															assign node569 = (inp[5]) ? 40'b0001000000011001010010000011001000010000 : 40'b1001000000011001010010000010001000010000;
														assign node572 = (inp[6]) ? 40'b0001000000011001010110000010001000010000 : 40'b0001000000010001010110000010001000010000;
													assign node575 = (inp[6]) ? 40'b0001000000011001010010000011001000000000 : node576;
														assign node576 = (inp[2]) ? 40'b0001000000010001010110000011001000000000 : 40'b1001000000010001010110000010001000000000;
												assign node580 = (inp[11]) ? node590 : node581;
													assign node581 = (inp[6]) ? node587 : node582;
														assign node582 = (inp[5]) ? node584 : 40'b1001000000000001010010000000001000010000;
															assign node584 = (inp[12]) ? 40'b0001000000000001010110000011001000010000 : 40'b0001000000000001010110000010001000010000;
														assign node587 = (inp[12]) ? 40'b0001000000001001010010000011001000010000 : 40'b0001000000001001010110000010001000010000;
													assign node590 = (inp[6]) ? node592 : 40'b0001000000001001010110000010001000000000;
														assign node592 = (inp[5]) ? 40'b0001000000000001010110000011001000000000 : 40'b0001000000001001010110000010001000000000;
										assign node595 = (inp[15]) ? node633 : node596;
											assign node596 = (inp[13]) ? node612 : node597;
												assign node597 = (inp[6]) ? node605 : node598;
													assign node598 = (inp[12]) ? 40'b1000000000010001010010000001101000000000 : node599;
														assign node599 = (inp[11]) ? 40'b1000000000010001010110000010101000000000 : node600;
															assign node600 = (inp[2]) ? 40'b1000000000010001010110000010101000010000 : 40'b1000000000010001010010000000101000010000;
													assign node605 = (inp[5]) ? 40'b0000000000010001010110000011101000010000 : node606;
														assign node606 = (inp[2]) ? 40'b0000000000011001010110000010101000000000 : node607;
															assign node607 = (inp[12]) ? 40'b0000000000011001010010000010101000000000 : 40'b1000000000011001010010000010101000000000;
												assign node612 = (inp[6]) ? node624 : node613;
													assign node613 = (inp[12]) ? 40'b1000000000011001010010000010001000010000 : node614;
														assign node614 = (inp[11]) ? node620 : node615;
															assign node615 = (inp[5]) ? node617 : 40'b1000000000010001010110000010001000010000;
																assign node617 = (inp[2]) ? 40'b0000000000010001010110000010001000010000 : 40'b1000000000010001010110000010001000010000;
															assign node620 = (inp[2]) ? 40'b0000000000010001010110000010001000000000 : 40'b1000000000010001010110000010001000000000;
													assign node624 = (inp[5]) ? node630 : node625;
														assign node625 = (inp[11]) ? 40'b0000000000011001010010000010001000000000 : node626;
															assign node626 = (inp[12]) ? 40'b0000000000011001010010000010001000010000 : 40'b1000000000011001010010000010001000010000;
														assign node630 = (inp[11]) ? 40'b1000000000010001010010000001001000000000 : 40'b0000000000010001010010000001001000010000;
											assign node633 = (inp[11]) ? node653 : node634;
												assign node634 = (inp[13]) ? node644 : node635;
													assign node635 = (inp[5]) ? node639 : node636;
														assign node636 = (inp[2]) ? 40'b1000000000000001010010000001101000010000 : 40'b1000000000001001010010000010101000010000;
														assign node639 = (inp[2]) ? 40'b0000000000000001010110000011101000010000 : node640;
															assign node640 = (inp[12]) ? 40'b0000000000001001010010000011101000010000 : 40'b1000000000000001010010000001101000010000;
													assign node644 = (inp[6]) ? node648 : node645;
														assign node645 = (inp[12]) ? 40'b1000000000001001010010000010001000010000 : 40'b1000000000000001010110000010001000010000;
														assign node648 = (inp[12]) ? 40'b0000000000001001010010000011001000010000 : node649;
															assign node649 = (inp[2]) ? 40'b0000000000001001010110000010001000010000 : 40'b1000000000001001010010000010001000010000;
												assign node653 = (inp[13]) ? node659 : node654;
													assign node654 = (inp[5]) ? node656 : 40'b1000000000001001010010000010101000000000;
														assign node656 = (inp[2]) ? 40'b0000000000000001010110000011101000000000 : 40'b1000000000000001010110000010101000000000;
													assign node659 = (inp[12]) ? node667 : node660;
														assign node660 = (inp[2]) ? node662 : 40'b1000000000000001010010000001001000000000;
															assign node662 = (inp[5]) ? 40'b0000000000000001010110000011001000000000 : node663;
																assign node663 = (inp[6]) ? 40'b0000000000001001010110000010001000000000 : 40'b1000000000000001010110000010001000000000;
														assign node667 = (inp[5]) ? 40'b0000000000001001010110000010001000000000 : node668;
															assign node668 = (inp[6]) ? 40'b0000000000001001010010000011001000000000 : 40'b1000000000000001010010000001001000000000;
								assign node672 = (inp[11]) ? node686 : node673;
									assign node673 = (inp[0]) ? node675 : 40'b0000000000000000000000000000000000000000;
										assign node675 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node676;
											assign node676 = (inp[2]) ? node678 : 40'b0000000000000000000000000000000000000000;
												assign node678 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node679;
													assign node679 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node680;
														assign node680 = (inp[13]) ? 40'b1000000000010100001000000000000000000000 : 40'b1000000000010100001000000000100000000000;
									assign node686 = (inp[13]) ? node770 : node687;
										assign node687 = (inp[15]) ? node733 : node688;
											assign node688 = (inp[0]) ? node712 : node689;
												assign node689 = (inp[12]) ? node705 : node690;
													assign node690 = (inp[2]) ? node702 : node691;
														assign node691 = (inp[6]) ? node697 : node692;
															assign node692 = (inp[5]) ? node694 : 40'b1001010000010100000000000000100000000000;
																assign node694 = (inp[10]) ? 40'b1001010000010000000100000010100000000000 : 40'b1001010000010100000100000010100000000000;
															assign node697 = (inp[5]) ? node699 : 40'b1001010000011100000000000010100000000000;
																assign node699 = (inp[10]) ? 40'b1001010000010000000000000001100000000000 : 40'b1001010000010100000000000001100000000000;
														assign node702 = (inp[10]) ? 40'b0001010000010000000100000011100000000000 : 40'b0001010000010100000100000011100000000000;
													assign node705 = (inp[10]) ? 40'b0001010000011000000000000010100000000000 : node706;
														assign node706 = (inp[6]) ? node708 : 40'b0001010000011100000100000010100000000000;
															assign node708 = (inp[5]) ? 40'b0001010000011100000000000011100000000000 : 40'b0001010000011100000000000010100000000000;
												assign node712 = (inp[10]) ? node724 : node713;
													assign node713 = (inp[6]) ? node719 : node714;
														assign node714 = (inp[12]) ? node716 : 40'b1000010000010100000100000010100000000000;
															assign node716 = (inp[5]) ? 40'b0000010000011100000100000010100000000000 : 40'b1000010000011100000000000010100000000000;
														assign node719 = (inp[5]) ? 40'b0000010000010100000000000001100000000000 : node720;
															assign node720 = (inp[2]) ? 40'b0000010000011100000100000010100000000000 : 40'b1000010000011100000000000010100000000000;
													assign node724 = (inp[2]) ? node728 : node725;
														assign node725 = (inp[5]) ? 40'b0000010000011000000000000011100000000000 : 40'b1000010000011000000000000010100000000000;
														assign node728 = (inp[6]) ? 40'b0000010000011000000100000010100000000000 : node729;
															assign node729 = (inp[5]) ? 40'b0000010000010000000100000011100000000000 : 40'b1000010000010000000000000001100000000000;
											assign node733 = (inp[0]) ? node749 : node734;
												assign node734 = (inp[12]) ? node742 : node735;
													assign node735 = (inp[10]) ? node739 : node736;
														assign node736 = (inp[6]) ? 40'b1001010000001100000000000010100000000000 : 40'b1001010000000100000000000000100000000000;
														assign node739 = (inp[2]) ? 40'b1001010000000000000100000010100000000000 : 40'b1001010000001000000000000010100000000000;
													assign node742 = (inp[6]) ? node744 : 40'b0001010000000100000100000011100000000000;
														assign node744 = (inp[5]) ? 40'b0001010000001100000000000011100000000000 : node745;
															assign node745 = (inp[2]) ? 40'b0001010000001100000000000011100000000000 : 40'b0001010000001100000000000010100000000000;
												assign node749 = (inp[10]) ? node765 : node750;
													assign node750 = (inp[6]) ? node758 : node751;
														assign node751 = (inp[12]) ? node755 : node752;
															assign node752 = (inp[2]) ? 40'b1000010000000100000100000010100000000000 : 40'b1000010000000100000000000000100000000000;
															assign node755 = (inp[5]) ? 40'b0000010000001100000100000010100000000000 : 40'b1000010000001100000000000010100000000000;
														assign node758 = (inp[12]) ? node762 : node759;
															assign node759 = (inp[2]) ? 40'b0000010000001100000100000010100000000000 : 40'b1000010000001100000000000010100000000000;
															assign node762 = (inp[2]) ? 40'b0000010000001100000000000011100000000000 : 40'b0000010000001100000000000010100000000000;
													assign node765 = (inp[6]) ? node767 : 40'b0000010000000000000100000011100000000000;
														assign node767 = (inp[12]) ? 40'b0000010000001000000000000010100000000000 : 40'b1000010000001000000000000010100000000000;
										assign node770 = (inp[0]) ? node810 : node771;
											assign node771 = (inp[15]) ? node785 : node772;
												assign node772 = (inp[10]) ? node778 : node773;
													assign node773 = (inp[12]) ? node775 : 40'b1001010000010100000000000001000000000000;
														assign node775 = (inp[2]) ? 40'b0001010000010100000000000001000000000000 : 40'b0001010000011100000000000011000000000000;
													assign node778 = (inp[12]) ? 40'b0001010000011000000000000011000000000000 : node779;
														assign node779 = (inp[2]) ? node781 : 40'b1001010000010000000000000000000000000000;
															assign node781 = (inp[5]) ? 40'b0001010000010000000100000010000000000000 : 40'b0001010000011000000100000010000000000000;
												assign node785 = (inp[10]) ? node799 : node786;
													assign node786 = (inp[12]) ? node794 : node787;
														assign node787 = (inp[6]) ? 40'b0001010000001100000100000010000000000000 : node788;
															assign node788 = (inp[5]) ? 40'b1001010000000100000100000010000000000000 : node789;
																assign node789 = (inp[2]) ? 40'b1001010000000100000100000010000000000000 : 40'b1001010000000100000000000000000000000000;
														assign node794 = (inp[5]) ? node796 : 40'b0001010000001100000000000011000000000000;
															assign node796 = (inp[2]) ? 40'b0001010000000100000100000011000000000000 : 40'b0001010000001100000100000010000000000000;
													assign node799 = (inp[2]) ? node805 : node800;
														assign node800 = (inp[12]) ? 40'b0001010000001000000100000010000000000000 : node801;
															assign node801 = (inp[5]) ? 40'b1001010000000000000000000001000000000000 : 40'b1001010000000000000000000000000000000000;
														assign node805 = (inp[5]) ? 40'b0001010000000000000100000011000000000000 : node806;
															assign node806 = (inp[6]) ? 40'b0001010000001000000100000010000000000000 : 40'b1001010000000000000100000010000000000000;
											assign node810 = (inp[15]) ? node826 : node811;
												assign node811 = (inp[6]) ? node817 : node812;
													assign node812 = (inp[10]) ? 40'b1000010000010000000100000010000000000000 : node813;
														assign node813 = (inp[5]) ? 40'b0000010000010100000100000010000000000000 : 40'b1000010000010100000100000010000000000000;
													assign node817 = (inp[2]) ? node823 : node818;
														assign node818 = (inp[12]) ? 40'b0000010000011000000000000010000000000000 : node819;
															assign node819 = (inp[10]) ? 40'b1000010000011000000000000010000000000000 : 40'b1000010000011100000000000010000000000000;
														assign node823 = (inp[5]) ? 40'b0000010000010000000100000011000000000000 : 40'b0000010000011000000100000010000000000000;
												assign node826 = (inp[10]) ? node842 : node827;
													assign node827 = (inp[2]) ? node831 : node828;
														assign node828 = (inp[5]) ? 40'b1000010000000100000000000001000000000000 : 40'b1000010000001100000000000010000000000000;
														assign node831 = (inp[12]) ? node837 : node832;
															assign node832 = (inp[5]) ? node834 : 40'b1000010000000100000100000010000000000000;
																assign node834 = (inp[6]) ? 40'b0000010000000100000100000011000000000000 : 40'b0000010000000100000100000010000000000000;
															assign node837 = (inp[5]) ? 40'b0000010000000100000100000011000000000000 : node838;
																assign node838 = (inp[6]) ? 40'b0000010000001100000000000011000000000000 : 40'b1000010000000100000000000001000000000000;
													assign node842 = (inp[12]) ? node846 : node843;
														assign node843 = (inp[5]) ? 40'b1000010000000000000000000001000000000000 : 40'b1000010000001000000000000010000000000000;
														assign node846 = (inp[6]) ? 40'b0000010000000000000000000001000000000000 : 40'b1000010000000000000000000001000000000000;
							assign node849 = (inp[14]) ? node913 : node850;
								assign node850 = (inp[6]) ? node902 : node851;
									assign node851 = (inp[5]) ? node863 : node852;
										assign node852 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node853;
											assign node853 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : node854;
												assign node854 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : node855;
													assign node855 = (inp[13]) ? node857 : 40'b0000000000000000000000000000000000000000;
														assign node857 = (inp[0]) ? 40'b1000000000010000000000000000000000100000 : 40'b1001000000010100000000000000000000100000;
										assign node863 = (inp[11]) ? node887 : node864;
											assign node864 = (inp[2]) ? node880 : node865;
												assign node865 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node866;
													assign node866 = (inp[13]) ? node872 : node867;
														assign node867 = (inp[15]) ? node869 : 40'b0000000000000000000000000000000000000000;
															assign node869 = (inp[10]) ? 40'b1001000000000000000100000010100000100000 : 40'b0000000000000000000000000000000000000000;
														assign node872 = (inp[15]) ? 40'b0000000000000000000000000000000000000000 : node873;
															assign node873 = (inp[0]) ? node875 : 40'b1001000000010000000100000010000000100000;
																assign node875 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000010100000100000010000000100000;
												assign node880 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : node881;
													assign node881 = (inp[15]) ? node883 : 40'b0000000000000000000000000000000000000000;
														assign node883 = (inp[10]) ? 40'b0001000000000000000100000011100000100000 : 40'b0000000000000000000000000000000000000000;
											assign node887 = (inp[2]) ? node889 : 40'b0000000000000000000000000000000000000000;
												assign node889 = (inp[12]) ? node891 : 40'b0000000000000000000000000000000000000000;
													assign node891 = (inp[15]) ? node893 : 40'b0000000000000000000000000000000000000000;
														assign node893 = (inp[0]) ? node897 : node894;
															assign node894 = (inp[10]) ? 40'b0001000000000000001100000010100000010000 : 40'b0000000000000000000000000000000000000000;
															assign node897 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node898;
																assign node898 = (inp[13]) ? 40'b0000000000000100001100000010000000010000 : 40'b0000000000000100001100000010100000010000;
									assign node902 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node903;
										assign node903 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node904;
											assign node904 = (inp[15]) ? node906 : 40'b0000000000000000000000000000000000000000;
												assign node906 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node907;
													assign node907 = (inp[0]) ? 40'b0000000000001100000100000010100000100000 : 40'b0000000000000000000000000000000000000000;
								assign node913 = (inp[11]) ? node915 : 40'b0000000000000000000000000000000000000000;
									assign node915 = (inp[15]) ? node995 : node916;
										assign node916 = (inp[10]) ? node950 : node917;
											assign node917 = (inp[0]) ? node937 : node918;
												assign node918 = (inp[5]) ? node932 : node919;
													assign node919 = (inp[6]) ? node927 : node920;
														assign node920 = (inp[2]) ? node924 : node921;
															assign node921 = (inp[13]) ? 40'b1011000000011100000000000010000000000000 : 40'b1011000000011100000000000010100000000000;
															assign node924 = (inp[13]) ? 40'b1011000000010100000000000001000000000000 : 40'b1011000000010100000000000001100000000000;
														assign node927 = (inp[2]) ? 40'b0011000000011100000100000010000000000000 : node928;
															assign node928 = (inp[12]) ? 40'b0011000000011100000000000010000000000000 : 40'b1011000000011100000000000010000000000000;
													assign node932 = (inp[2]) ? node934 : 40'b1011000000010100000000000001100000000000;
														assign node934 = (inp[13]) ? 40'b0011000000010100000100000011000000000000 : 40'b0011000000010100000100000011100000000000;
												assign node937 = (inp[13]) ? node943 : node938;
													assign node938 = (inp[12]) ? node940 : 40'b1010000000011100000000000010100000000000;
														assign node940 = (inp[6]) ? 40'b0010000000011100000000000011100000000000 : 40'b0010000000011100000100000010100000000000;
													assign node943 = (inp[12]) ? node947 : node944;
														assign node944 = (inp[6]) ? 40'b0010000000010100000100000011000000000000 : 40'b0010000000010100000100000010000000000000;
														assign node947 = (inp[6]) ? 40'b0010000000011100000000000011000000000000 : 40'b1010000000010100000000000001000000000000;
											assign node950 = (inp[13]) ? node964 : node951;
												assign node951 = (inp[6]) ? node961 : node952;
													assign node952 = (inp[0]) ? node954 : 40'b0011000000010000000100000010100000000000;
														assign node954 = (inp[2]) ? node958 : node955;
															assign node955 = (inp[5]) ? 40'b1010000000010000000100000010100000000000 : 40'b1010000000010000000000000000100000000000;
															assign node958 = (inp[5]) ? 40'b0010000000010000000100000010100000000000 : 40'b1010000000010000000100000010100000000000;
													assign node961 = (inp[2]) ? 40'b0011000000011000000100000010100000000000 : 40'b0010000000011000000000000011100000000000;
												assign node964 = (inp[0]) ? node978 : node965;
													assign node965 = (inp[12]) ? node975 : node966;
														assign node966 = (inp[2]) ? node970 : node967;
															assign node967 = (inp[6]) ? 40'b1011000000010000000000000001000000000000 : 40'b1011000000010000000000000000000000000000;
															assign node970 = (inp[6]) ? node972 : 40'b1011000000010000000100000010000000000000;
																assign node972 = (inp[5]) ? 40'b0011000000010000000100000011000000000000 : 40'b0011000000011000000100000010000000000000;
														assign node975 = (inp[5]) ? 40'b0011000000010000000000000001000000000000 : 40'b1011000000010000000000000001000000000000;
													assign node978 = (inp[5]) ? node986 : node979;
														assign node979 = (inp[6]) ? node983 : node980;
															assign node980 = (inp[12]) ? 40'b1010000000010000000000000001000000000000 : 40'b1010000000010000000000000000000000000000;
															assign node983 = (inp[12]) ? 40'b0010000000011000000000000011000000000000 : 40'b1010000000011000000000000010000000000000;
														assign node986 = (inp[6]) ? node992 : node987;
															assign node987 = (inp[12]) ? 40'b0010000000010000000100000011000000000000 : node988;
																assign node988 = (inp[2]) ? 40'b0010000000010000000100000010000000000000 : 40'b1010000000010000000100000010000000000000;
															assign node992 = (inp[2]) ? 40'b0010000000010000000100000011000000000000 : 40'b0010000000011000000000000011000000000000;
										assign node995 = (inp[13]) ? node1041 : node996;
											assign node996 = (inp[10]) ? node1018 : node997;
												assign node997 = (inp[2]) ? node1007 : node998;
													assign node998 = (inp[6]) ? 40'b1011000000000100000000000001100000000000 : node999;
														assign node999 = (inp[5]) ? node1003 : node1000;
															assign node1000 = (inp[0]) ? 40'b1010000000000100000000000000100000000000 : 40'b1011000000000100000000000000100000000000;
															assign node1003 = (inp[0]) ? 40'b1010000000000100000100000010100000000000 : 40'b1011000000000100000100000010100000000000;
													assign node1007 = (inp[0]) ? node1011 : node1008;
														assign node1008 = (inp[12]) ? 40'b0011000000001100000000000011100000000000 : 40'b0011000000000100000100000011100000000000;
														assign node1011 = (inp[5]) ? node1015 : node1012;
															assign node1012 = (inp[6]) ? 40'b0010000000001100000100000010100000000000 : 40'b1010000000000100000100000010100000000000;
															assign node1015 = (inp[6]) ? 40'b0010000000000100000000000001100000000000 : 40'b0010000000000100000100000011100000000000;
												assign node1018 = (inp[0]) ? node1030 : node1019;
													assign node1019 = (inp[12]) ? node1027 : node1020;
														assign node1020 = (inp[2]) ? node1024 : node1021;
															assign node1021 = (inp[6]) ? 40'b1011000000000000000000000001100000000000 : 40'b1011000000000000000000000000100000000000;
															assign node1024 = (inp[6]) ? 40'b0011000000001000000100000010100000000000 : 40'b1011000000000000000100000010100000000000;
														assign node1027 = (inp[2]) ? 40'b0011000000000000000100000011100000000000 : 40'b0011000000001000000100000010100000000000;
													assign node1030 = (inp[6]) ? node1034 : node1031;
														assign node1031 = (inp[12]) ? 40'b1010000000001000000000000010100000000000 : 40'b1010000000000000000100000010100000000000;
														assign node1034 = (inp[12]) ? node1036 : 40'b1010000000001000000000000010100000000000;
															assign node1036 = (inp[5]) ? node1038 : 40'b0010000000001000000000000011100000000000;
																assign node1038 = (inp[2]) ? 40'b0010000000000000000000000001100000000000 : 40'b0010000000001000000000000011100000000000;
											assign node1041 = (inp[6]) ? node1063 : node1042;
												assign node1042 = (inp[10]) ? node1054 : node1043;
													assign node1043 = (inp[12]) ? node1051 : node1044;
														assign node1044 = (inp[0]) ? 40'b1010000000000100000000000000000000000000 : node1045;
															assign node1045 = (inp[5]) ? 40'b1011000000000100000100000010000000000000 : node1046;
																assign node1046 = (inp[2]) ? 40'b1011000000000100000100000010000000000000 : 40'b1011000000000100000000000000000000000000;
														assign node1051 = (inp[2]) ? 40'b0011000000000100000100000011000000000000 : 40'b0011000000001100000100000010000000000000;
													assign node1054 = (inp[12]) ? node1060 : node1055;
														assign node1055 = (inp[0]) ? node1057 : 40'b1011000000000000000100000010000000000000;
															assign node1057 = (inp[2]) ? 40'b0010000000000000000100000010000000000000 : 40'b1010000000000000000100000010000000000000;
														assign node1060 = (inp[0]) ? 40'b1010000000001000000000000010000000000000 : 40'b1011000000001000000000000010000000000000;
												assign node1063 = (inp[0]) ? node1071 : node1064;
													assign node1064 = (inp[12]) ? node1068 : node1065;
														assign node1065 = (inp[2]) ? 40'b0011000000001000000100000010000000000000 : 40'b1011000000001000000000000010000000000000;
														assign node1068 = (inp[10]) ? 40'b0011000000001000000000000011000000000000 : 40'b0011000000001100000000000011000000000000;
													assign node1071 = (inp[12]) ? node1075 : node1072;
														assign node1072 = (inp[10]) ? 40'b1010000000001000000000000010000000000000 : 40'b1010000000001100000000000010000000000000;
														assign node1075 = (inp[10]) ? 40'b0010000000001000000000000010000000000000 : 40'b0010000000001100000000000010000000000000;
						assign node1078 = (inp[3]) ? node1182 : node1079;
							assign node1079 = (inp[14]) ? node1105 : node1080;
								assign node1080 = (inp[11]) ? node1082 : 40'b0000000000000000000000000000000000000000;
									assign node1082 = (inp[15]) ? node1094 : node1083;
										assign node1083 = (inp[10]) ? node1089 : node1084;
											assign node1084 = (inp[0]) ? node1086 : 40'b0000000000000000000000000000000000000000;
												assign node1086 = (inp[13]) ? 40'b1000001000010100000000000000000000001000 : 40'b1000001000010100000000000000100000001000;
											assign node1089 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : node1090;
												assign node1090 = (inp[13]) ? 40'b1001001000010000000000000000000000001000 : 40'b1001001000010000000000000000100000001000;
										assign node1094 = (inp[0]) ? node1100 : node1095;
											assign node1095 = (inp[10]) ? node1097 : 40'b0000000000000000000000000000000000000000;
												assign node1097 = (inp[13]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000000000000100000010100000001000;
											assign node1100 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node1101;
												assign node1101 = (inp[13]) ? 40'b0000001000000100000100000010000000001000 : 40'b0000001000000100000100000010100000001000;
								assign node1105 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node1106;
									assign node1106 = (inp[15]) ? node1120 : node1107;
										assign node1107 = (inp[10]) ? node1109 : 40'b0000000000000000000000000000000000000000;
											assign node1109 = (inp[0]) ? node1111 : 40'b0000000000000000000000000000000000000000;
												assign node1111 = (inp[13]) ? node1113 : 40'b0000000000000000000000000000000000000000;
													assign node1113 = (inp[6]) ? node1117 : node1114;
														assign node1114 = (inp[12]) ? 40'b1000001100011000000000000010000000000000 : 40'b1000001100010000000100000010000000000000;
														assign node1117 = (inp[12]) ? 40'b0000001100011000000000000011000000000000 : 40'b0000001100011000000100000010000000000000;
										assign node1120 = (inp[6]) ? node1148 : node1121;
											assign node1121 = (inp[2]) ? node1133 : node1122;
												assign node1122 = (inp[13]) ? node1124 : 40'b0000000000000000000000000000000000000000;
													assign node1124 = (inp[12]) ? node1126 : 40'b0000000000000000000000000000000000000000;
														assign node1126 = (inp[5]) ? 40'b0001001100001000000100000010000000000000 : node1127;
															assign node1127 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node1128;
																assign node1128 = (inp[0]) ? 40'b1000001100001100000000000010000000000000 : 40'b0000000000000000000000000000000000000000;
												assign node1133 = (inp[13]) ? node1141 : node1134;
													assign node1134 = (inp[5]) ? node1136 : 40'b0000000000000000000000000000000000000000;
														assign node1136 = (inp[0]) ? node1138 : 40'b0000000000000000000000000000000000000000;
															assign node1138 = (inp[12]) ? 40'b0000001100000000000100000011100000000000 : 40'b0000001100000000000100000010100000000000;
													assign node1141 = (inp[10]) ? node1145 : node1142;
														assign node1142 = (inp[5]) ? 40'b0000001100000100000100000010000000000000 : 40'b1000001100000100000100000010000000000000;
														assign node1145 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : 40'b1001001100000000000100000010000000000000;
											assign node1148 = (inp[5]) ? node1160 : node1149;
												assign node1149 = (inp[0]) ? node1153 : node1150;
													assign node1150 = (inp[2]) ? 40'b0001001100001000000000000011000000000000 : 40'b1001001100001000000000000010000000000000;
													assign node1153 = (inp[10]) ? node1157 : node1154;
														assign node1154 = (inp[13]) ? 40'b0000001100001100000000000010000000000000 : 40'b0000000000000000000000000000000000000000;
														assign node1157 = (inp[12]) ? 40'b0000001100001000000000000010100000000000 : 40'b0000001100001000000100000010100000000000;
												assign node1160 = (inp[13]) ? node1170 : node1161;
													assign node1161 = (inp[0]) ? node1163 : 40'b0000000000000000000000000000000000000000;
														assign node1163 = (inp[10]) ? node1165 : 40'b0000000000000000000000000000000000000000;
															assign node1165 = (inp[12]) ? node1167 : 40'b1000001100000000000000000001100000000000;
																assign node1167 = (inp[2]) ? 40'b0000001100000000000000000001100000000000 : 40'b0000001100001000000000000011100000000000;
													assign node1170 = (inp[10]) ? node1178 : node1171;
														assign node1171 = (inp[0]) ? node1173 : 40'b0000000000000000000000000000000000000000;
															assign node1173 = (inp[12]) ? 40'b0000001100001100000000000011000000000000 : node1174;
																assign node1174 = (inp[2]) ? 40'b0000001100000100000100000011000000000000 : 40'b1000001100000100000000000001000000000000;
														assign node1178 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : 40'b0001001100001000000000000011000000000000;
							assign node1182 = (inp[11]) ? node1342 : node1183;
								assign node1183 = (inp[14]) ? node1185 : 40'b0000000000000000000000000000000000000000;
									assign node1185 = (inp[10]) ? node1261 : node1186;
										assign node1186 = (inp[0]) ? node1224 : node1187;
											assign node1187 = (inp[15]) ? node1203 : node1188;
												assign node1188 = (inp[2]) ? node1200 : node1189;
													assign node1189 = (inp[12]) ? 40'b0001001000011100000100000010000000000000 : node1190;
														assign node1190 = (inp[5]) ? node1196 : node1191;
															assign node1191 = (inp[6]) ? 40'b1001001000011100000000000010100000000000 : node1192;
																assign node1192 = (inp[13]) ? 40'b1001001000010100000000000000000000000000 : 40'b1001001000010100000000000000100000000000;
															assign node1196 = (inp[13]) ? 40'b1001001000010100000000000001000000000000 : 40'b1001001000010100000000000001100000000000;
													assign node1200 = (inp[6]) ? 40'b0001001000010100000100000011100000000000 : 40'b0001001000010100000100000011000000000000;
												assign node1203 = (inp[13]) ? node1215 : node1204;
													assign node1204 = (inp[12]) ? node1212 : node1205;
														assign node1205 = (inp[6]) ? 40'b0001001000001100000100000010100000000000 : node1206;
															assign node1206 = (inp[5]) ? node1208 : 40'b1001001000000100000100000010100000000000;
																assign node1208 = (inp[2]) ? 40'b0001001000000100000100000010100000000000 : 40'b1001001000000100000100000010100000000000;
														assign node1212 = (inp[5]) ? 40'b0001001000001100000100000010100000000000 : 40'b1001001000001100000000000010100000000000;
													assign node1215 = (inp[5]) ? node1219 : node1216;
														assign node1216 = (inp[2]) ? 40'b1001001000000100000100000010000000000000 : 40'b1001001000000100000000000000000000000000;
														assign node1219 = (inp[2]) ? node1221 : 40'b0001001000001100000100000010000000000000;
															assign node1221 = (inp[12]) ? 40'b0001001000000100000100000011000000000000 : 40'b0001001000000100000100000010000000000000;
											assign node1224 = (inp[15]) ? node1246 : node1225;
												assign node1225 = (inp[6]) ? node1237 : node1226;
													assign node1226 = (inp[13]) ? node1232 : node1227;
														assign node1227 = (inp[12]) ? 40'b1000001000011100000000000010100000000000 : node1228;
															assign node1228 = (inp[5]) ? 40'b0000001000010100000100000010100000000000 : 40'b1000001000010100000100000010100000000000;
														assign node1232 = (inp[12]) ? node1234 : 40'b1000001000010100000100000010000000000000;
															assign node1234 = (inp[2]) ? 40'b0000001000010100000100000011000000000000 : 40'b0000001000011100000100000010000000000000;
													assign node1237 = (inp[13]) ? node1241 : node1238;
														assign node1238 = (inp[12]) ? 40'b0000001000010100000000000001100000000000 : 40'b0000001000010100000100000011100000000000;
														assign node1241 = (inp[5]) ? node1243 : 40'b0000001000011100000000000011000000000000;
															assign node1243 = (inp[2]) ? 40'b0000001000010100000000000001000000000000 : 40'b1000001000010100000000000001000000000000;
												assign node1246 = (inp[2]) ? node1252 : node1247;
													assign node1247 = (inp[12]) ? node1249 : 40'b1000001000000100000000000001100000000000;
														assign node1249 = (inp[5]) ? 40'b0000001000001100000100000010100000000000 : 40'b1000001000001100000000000010100000000000;
													assign node1252 = (inp[12]) ? node1254 : 40'b0000001000000100000100000010000000000000;
														assign node1254 = (inp[5]) ? node1258 : node1255;
															assign node1255 = (inp[13]) ? 40'b1000001000000100000000000001000000000000 : 40'b1000001000000100000000000001100000000000;
															assign node1258 = (inp[13]) ? 40'b0000001000000100000000000001000000000000 : 40'b0000001000000100000000000001100000000000;
										assign node1261 = (inp[12]) ? node1285 : node1262;
											assign node1262 = (inp[6]) ? node1276 : node1263;
												assign node1263 = (inp[15]) ? node1271 : node1264;
													assign node1264 = (inp[5]) ? 40'b0001001000010000000100000010100000000000 : node1265;
														assign node1265 = (inp[13]) ? node1267 : 40'b1000001000010000000100000010100000000000;
															assign node1267 = (inp[0]) ? 40'b1000001000010000000100000010000000000000 : 40'b1001001000010000000100000010000000000000;
													assign node1271 = (inp[13]) ? 40'b1001001000000000000100000010000000000000 : node1272;
														assign node1272 = (inp[2]) ? 40'b1001001000000000000100000010100000000000 : 40'b1000001000000000000100000010100000000000;
												assign node1276 = (inp[2]) ? node1282 : node1277;
													assign node1277 = (inp[0]) ? 40'b1000001000001000000000000010100000000000 : node1278;
														assign node1278 = (inp[15]) ? 40'b1001001000000000000000000001000000000000 : 40'b1001001000010000000000000001000000000000;
													assign node1282 = (inp[15]) ? 40'b0000001000000000000100000011000000000000 : 40'b0000001000010000000100000011000000000000;
											assign node1285 = (inp[2]) ? node1317 : node1286;
												assign node1286 = (inp[15]) ? node1304 : node1287;
													assign node1287 = (inp[13]) ? node1297 : node1288;
														assign node1288 = (inp[0]) ? node1292 : node1289;
															assign node1289 = (inp[5]) ? 40'b0001001000011000000000000011100000000000 : 40'b0001001000011000000000000010100000000000;
															assign node1292 = (inp[6]) ? node1294 : 40'b0000001000011000000100000010100000000000;
																assign node1294 = (inp[5]) ? 40'b0000001000011000000000000011100000000000 : 40'b0000001000011000000000000010100000000000;
														assign node1297 = (inp[0]) ? node1299 : 40'b0001001000011000000000000010000000000000;
															assign node1299 = (inp[6]) ? node1301 : 40'b0000001000011000000100000010000000000000;
																assign node1301 = (inp[5]) ? 40'b0000001000011000000000000011000000000000 : 40'b0000001000011000000000000010000000000000;
													assign node1304 = (inp[0]) ? node1310 : node1305;
														assign node1305 = (inp[6]) ? node1307 : 40'b1001001000001000000000000010100000000000;
															assign node1307 = (inp[5]) ? 40'b0001001000001000000000000011100000000000 : 40'b0001001000001000000000000010100000000000;
														assign node1310 = (inp[13]) ? 40'b1000001000001000000000000010000000000000 : node1311;
															assign node1311 = (inp[6]) ? node1313 : 40'b0000001000001000000100000010100000000000;
																assign node1313 = (inp[5]) ? 40'b0000001000001000000000000011100000000000 : 40'b0000001000001000000000000010100000000000;
												assign node1317 = (inp[15]) ? node1327 : node1318;
													assign node1318 = (inp[6]) ? node1322 : node1319;
														assign node1319 = (inp[0]) ? 40'b1000001000010000000000000001100000000000 : 40'b1001001000010000000000000001100000000000;
														assign node1322 = (inp[5]) ? 40'b0000001000010000000000000001100000000000 : node1323;
															assign node1323 = (inp[0]) ? 40'b0000001000011000000000000011100000000000 : 40'b0001001000011000000000000011100000000000;
													assign node1327 = (inp[0]) ? node1335 : node1328;
														assign node1328 = (inp[5]) ? node1330 : 40'b0001001000001000000000000011100000000000;
															assign node1330 = (inp[6]) ? node1332 : 40'b0001001000000000000100000011100000000000;
																assign node1332 = (inp[13]) ? 40'b0001001000000000000000000001000000000000 : 40'b0001001000000000000000000001100000000000;
														assign node1335 = (inp[6]) ? node1339 : node1336;
															assign node1336 = (inp[5]) ? 40'b0000001000000000000100000011000000000000 : 40'b1000001000000000000000000001000000000000;
															assign node1339 = (inp[13]) ? 40'b0000001000001000000000000011000000000000 : 40'b0000001000001000000000000011100000000000;
								assign node1342 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node1343;
									assign node1343 = (inp[15]) ? node1423 : node1344;
										assign node1344 = (inp[0]) ? node1392 : node1345;
											assign node1345 = (inp[13]) ? node1359 : node1346;
												assign node1346 = (inp[10]) ? node1350 : node1347;
													assign node1347 = (inp[5]) ? 40'b0001001000010100000100000011100000001000 : 40'b1001001000010100000100000010100000001000;
													assign node1350 = (inp[12]) ? 40'b0001001000011000000000000011100000001000 : node1351;
														assign node1351 = (inp[2]) ? node1355 : node1352;
															assign node1352 = (inp[5]) ? 40'b1001001000010000000000000001100000001000 : 40'b1001001000011000000000000010100000001000;
															assign node1355 = (inp[6]) ? 40'b0001001000010000000100000011100000001000 : 40'b0001001000010000000100000010100000001000;
												assign node1359 = (inp[10]) ? node1371 : node1360;
													assign node1360 = (inp[5]) ? node1368 : node1361;
														assign node1361 = (inp[2]) ? 40'b1001001000010100000100000010000000001000 : node1362;
															assign node1362 = (inp[12]) ? 40'b1001001000011100000000000010000000001000 : node1363;
																assign node1363 = (inp[6]) ? 40'b1001001000011100000000000010000000001000 : 40'b1001001000010100000000000000000000001000;
														assign node1368 = (inp[6]) ? 40'b0001001000010100000000000001000000001000 : 40'b0001001000010100000100000011000000001000;
													assign node1371 = (inp[5]) ? node1381 : node1372;
														assign node1372 = (inp[6]) ? node1378 : node1373;
															assign node1373 = (inp[12]) ? 40'b1001001000010000000000000001000000001000 : node1374;
																assign node1374 = (inp[2]) ? 40'b1001001000010000000100000010000000001000 : 40'b1001001000010000000000000000000000001000;
															assign node1378 = (inp[2]) ? 40'b0001001000011000000100000010000000001000 : 40'b1001001000011000000000000010000000001000;
														assign node1381 = (inp[6]) ? node1387 : node1382;
															assign node1382 = (inp[2]) ? 40'b0001001000010000000100000011000000001000 : node1383;
																assign node1383 = (inp[12]) ? 40'b0001001000011000000100000010000000001000 : 40'b1001001000010000000100000010000000001000;
															assign node1387 = (inp[12]) ? 40'b0001001000011000000000000011000000001000 : node1388;
																assign node1388 = (inp[2]) ? 40'b0001001000010000000100000011000000001000 : 40'b1001001000010000000000000001000000001000;
											assign node1392 = (inp[13]) ? node1406 : node1393;
												assign node1393 = (inp[12]) ? node1401 : node1394;
													assign node1394 = (inp[5]) ? node1398 : node1395;
														assign node1395 = (inp[10]) ? 40'b1000001000011000000000000010100000001000 : 40'b1000001000011100000000000010100000001000;
														assign node1398 = (inp[10]) ? 40'b1000001000010000000000000001100000001000 : 40'b1000001000010100000000000001100000001000;
													assign node1401 = (inp[6]) ? 40'b0000001000011000000000000011100000001000 : node1402;
														assign node1402 = (inp[2]) ? 40'b0000001000010000000100000011100000001000 : 40'b0000001000011000000100000010100000001000;
												assign node1406 = (inp[10]) ? node1412 : node1407;
													assign node1407 = (inp[12]) ? node1409 : 40'b0000001000011100000100000010000000001000;
														assign node1409 = (inp[2]) ? 40'b0000001000011100000000000011000000001000 : 40'b0000001000011100000000000010000000001000;
													assign node1412 = (inp[12]) ? node1416 : node1413;
														assign node1413 = (inp[6]) ? 40'b0000001000011000000100000010000000001000 : 40'b1000001000010000000100000010000000001000;
														assign node1416 = (inp[2]) ? node1418 : 40'b0000001000011000000100000010000000001000;
															assign node1418 = (inp[6]) ? node1420 : 40'b1000001000010000000000000001000000001000;
																assign node1420 = (inp[5]) ? 40'b0000001000010000000000000001000000001000 : 40'b0000001000011000000000000011000000001000;
										assign node1423 = (inp[13]) ? node1465 : node1424;
											assign node1424 = (inp[0]) ? node1444 : node1425;
												assign node1425 = (inp[2]) ? node1435 : node1426;
													assign node1426 = (inp[12]) ? node1432 : node1427;
														assign node1427 = (inp[10]) ? 40'b1001001000000000000000000001100000001000 : node1428;
															assign node1428 = (inp[5]) ? 40'b1001001000000100000000000001100000001000 : 40'b1001001000000100000000000000100000001000;
														assign node1432 = (inp[6]) ? 40'b0001001000001000000000000011100000001000 : 40'b0001001000001000000100000010100000001000;
													assign node1435 = (inp[5]) ? node1441 : node1436;
														assign node1436 = (inp[6]) ? 40'b0001001000001100000100000010100000001000 : node1437;
															assign node1437 = (inp[10]) ? 40'b1001001000000000000100000010100000001000 : 40'b1001001000000100000100000010100000001000;
														assign node1441 = (inp[10]) ? 40'b0001001000000000000100000011100000001000 : 40'b0001001000000100000100000011100000001000;
												assign node1444 = (inp[2]) ? node1454 : node1445;
													assign node1445 = (inp[6]) ? node1449 : node1446;
														assign node1446 = (inp[5]) ? 40'b1000001000000100000100000010100000001000 : 40'b1000001000000100000000000000100000001000;
														assign node1449 = (inp[12]) ? node1451 : 40'b1000001000001000000000000010100000001000;
															assign node1451 = (inp[10]) ? 40'b0000001000001000000000000011100000001000 : 40'b0000001000001100000000000010100000001000;
													assign node1454 = (inp[6]) ? node1462 : node1455;
														assign node1455 = (inp[5]) ? node1457 : 40'b1000001000000000000000000001100000001000;
															assign node1457 = (inp[10]) ? node1459 : 40'b0000001000000100000100000011100000001000;
																assign node1459 = (inp[12]) ? 40'b0000001000000000000100000011100000001000 : 40'b0000001000000000000100000010100000001000;
														assign node1462 = (inp[10]) ? 40'b0000001000000000000000000001100000001000 : 40'b0000001000000100000000000001100000001000;
											assign node1465 = (inp[0]) ? node1495 : node1466;
												assign node1466 = (inp[10]) ? node1486 : node1467;
													assign node1467 = (inp[12]) ? node1477 : node1468;
														assign node1468 = (inp[5]) ? node1474 : node1469;
															assign node1469 = (inp[2]) ? node1471 : 40'b1001001000001100000000000010000000001000;
																assign node1471 = (inp[6]) ? 40'b0001001000001100000100000010000000001000 : 40'b1001001000000100000100000010000000001000;
															assign node1474 = (inp[2]) ? 40'b0001001000000100000100000011000000001000 : 40'b1001001000000100000000000001000000001000;
														assign node1477 = (inp[6]) ? node1481 : node1478;
															assign node1478 = (inp[5]) ? 40'b0001001000000100000100000011000000001000 : 40'b1001001000000100000000000001000000001000;
															assign node1481 = (inp[2]) ? node1483 : 40'b0001001000001100000000000011000000001000;
																assign node1483 = (inp[5]) ? 40'b0001001000000100000000000001000000001000 : 40'b0001001000001100000000000011000000001000;
													assign node1486 = (inp[6]) ? node1488 : 40'b1001001000000000000000000001000000001000;
														assign node1488 = (inp[12]) ? node1490 : 40'b1001001000000000000000000001000000001000;
															assign node1490 = (inp[2]) ? 40'b0001001000001000000000000011000000001000 : node1491;
																assign node1491 = (inp[5]) ? 40'b0001001000001000000000000011000000001000 : 40'b0001001000001000000000000010000000001000;
												assign node1495 = (inp[12]) ? node1505 : node1496;
													assign node1496 = (inp[10]) ? node1498 : 40'b1000001000000100000000000000000000001000;
														assign node1498 = (inp[5]) ? node1502 : node1499;
															assign node1499 = (inp[6]) ? 40'b1000001000001000000000000010000000001000 : 40'b1000001000000000000000000000000000001000;
															assign node1502 = (inp[6]) ? 40'b1000001000000000000000000001000000001000 : 40'b1000001000000000000100000010000000001000;
													assign node1505 = (inp[6]) ? node1509 : node1506;
														assign node1506 = (inp[10]) ? 40'b0000001000001000000100000010000000001000 : 40'b0000001000001100000100000010000000001000;
														assign node1509 = (inp[2]) ? 40'b0000001000001000000000000011000000001000 : node1510;
															assign node1510 = (inp[5]) ? 40'b0000001000001100000000000011000000001000 : 40'b0000001000001100000000000010000000001000;

endmodule