module dtc_split33_bm75 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node234;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node351;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node387;
	wire [3-1:0] node390;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node460;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node473;
	wire [3-1:0] node476;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node481;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node493;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node521;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node538;
	wire [3-1:0] node541;
	wire [3-1:0] node544;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node570;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node609;
	wire [3-1:0] node612;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node633;
	wire [3-1:0] node635;
	wire [3-1:0] node638;
	wire [3-1:0] node640;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node690;
	wire [3-1:0] node692;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node734;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node741;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node787;
	wire [3-1:0] node791;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node797;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node806;
	wire [3-1:0] node808;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node824;
	wire [3-1:0] node828;
	wire [3-1:0] node830;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node887;
	wire [3-1:0] node888;
	wire [3-1:0] node890;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node902;
	wire [3-1:0] node905;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node914;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node923;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node935;
	wire [3-1:0] node938;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node959;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node968;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node975;
	wire [3-1:0] node978;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node986;
	wire [3-1:0] node988;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node997;
	wire [3-1:0] node998;
	wire [3-1:0] node1003;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1018;
	wire [3-1:0] node1020;
	wire [3-1:0] node1022;
	wire [3-1:0] node1026;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1032;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1043;
	wire [3-1:0] node1046;
	wire [3-1:0] node1049;
	wire [3-1:0] node1050;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1055;
	wire [3-1:0] node1059;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1065;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1070;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1096;
	wire [3-1:0] node1098;
	wire [3-1:0] node1100;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1108;
	wire [3-1:0] node1111;
	wire [3-1:0] node1115;
	wire [3-1:0] node1116;
	wire [3-1:0] node1119;
	wire [3-1:0] node1120;
	wire [3-1:0] node1124;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1131;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1138;
	wire [3-1:0] node1140;
	wire [3-1:0] node1142;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1148;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1159;
	wire [3-1:0] node1160;
	wire [3-1:0] node1164;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1175;
	wire [3-1:0] node1176;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1181;
	wire [3-1:0] node1183;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1205;
	wire [3-1:0] node1207;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1213;
	wire [3-1:0] node1214;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1223;
	wire [3-1:0] node1224;
	wire [3-1:0] node1226;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1234;
	wire [3-1:0] node1235;
	wire [3-1:0] node1239;
	wire [3-1:0] node1241;
	wire [3-1:0] node1244;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1258;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1268;
	wire [3-1:0] node1269;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1280;
	wire [3-1:0] node1282;
	wire [3-1:0] node1283;
	wire [3-1:0] node1285;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1290;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1296;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1305;
	wire [3-1:0] node1307;
	wire [3-1:0] node1308;
	wire [3-1:0] node1311;
	wire [3-1:0] node1314;
	wire [3-1:0] node1315;
	wire [3-1:0] node1317;
	wire [3-1:0] node1319;
	wire [3-1:0] node1321;
	wire [3-1:0] node1323;

	assign outp = (inp[3]) ? node746 : node1;
		assign node1 = (inp[9]) ? node323 : node2;
			assign node2 = (inp[4]) ? node134 : node3;
				assign node3 = (inp[6]) ? node97 : node4;
					assign node4 = (inp[0]) ? node64 : node5;
						assign node5 = (inp[5]) ? node27 : node6;
							assign node6 = (inp[8]) ? node18 : node7;
								assign node7 = (inp[10]) ? node13 : node8;
									assign node8 = (inp[11]) ? 3'b011 : node9;
										assign node9 = (inp[7]) ? 3'b111 : 3'b011;
									assign node13 = (inp[2]) ? node15 : 3'b101;
										assign node15 = (inp[7]) ? 3'b111 : 3'b011;
								assign node18 = (inp[10]) ? 3'b011 : node19;
									assign node19 = (inp[7]) ? node21 : 3'b011;
										assign node21 = (inp[11]) ? node23 : 3'b111;
											assign node23 = (inp[2]) ? 3'b111 : 3'b011;
							assign node27 = (inp[8]) ? node55 : node28;
								assign node28 = (inp[2]) ? node44 : node29;
									assign node29 = (inp[1]) ? node35 : node30;
										assign node30 = (inp[10]) ? 3'b001 : node31;
											assign node31 = (inp[7]) ? 3'b101 : 3'b001;
										assign node35 = (inp[11]) ? node41 : node36;
											assign node36 = (inp[7]) ? 3'b101 : node37;
												assign node37 = (inp[10]) ? 3'b001 : 3'b101;
											assign node41 = (inp[10]) ? 3'b101 : 3'b011;
									assign node44 = (inp[10]) ? node50 : node45;
										assign node45 = (inp[1]) ? 3'b011 : node46;
											assign node46 = (inp[11]) ? 3'b001 : 3'b101;
										assign node50 = (inp[11]) ? node52 : 3'b001;
											assign node52 = (inp[7]) ? 3'b101 : 3'b110;
								assign node55 = (inp[11]) ? 3'b101 : node56;
									assign node56 = (inp[7]) ? 3'b011 : node57;
										assign node57 = (inp[10]) ? node59 : 3'b101;
											assign node59 = (inp[1]) ? 3'b101 : 3'b001;
						assign node64 = (inp[10]) ? node74 : node65;
							assign node65 = (inp[11]) ? node67 : 3'b111;
								assign node67 = (inp[2]) ? 3'b111 : node68;
									assign node68 = (inp[8]) ? node70 : 3'b111;
										assign node70 = (inp[1]) ? 3'b111 : 3'b011;
							assign node74 = (inp[7]) ? node92 : node75;
								assign node75 = (inp[5]) ? node83 : node76;
									assign node76 = (inp[11]) ? node78 : 3'b111;
										assign node78 = (inp[1]) ? node80 : 3'b011;
											assign node80 = (inp[8]) ? 3'b111 : 3'b011;
									assign node83 = (inp[8]) ? 3'b011 : node84;
										assign node84 = (inp[11]) ? node86 : 3'b101;
											assign node86 = (inp[1]) ? 3'b101 : node87;
												assign node87 = (inp[2]) ? 3'b101 : 3'b001;
								assign node92 = (inp[1]) ? 3'b111 : node93;
									assign node93 = (inp[5]) ? 3'b011 : 3'b111;
					assign node97 = (inp[10]) ? node107 : node98;
						assign node98 = (inp[5]) ? node100 : 3'b111;
							assign node100 = (inp[8]) ? 3'b111 : node101;
								assign node101 = (inp[1]) ? 3'b111 : node102;
									assign node102 = (inp[2]) ? 3'b111 : 3'b011;
						assign node107 = (inp[1]) ? node127 : node108;
							assign node108 = (inp[5]) ? node116 : node109;
								assign node109 = (inp[11]) ? node111 : 3'b111;
									assign node111 = (inp[7]) ? 3'b111 : node112;
										assign node112 = (inp[0]) ? 3'b111 : 3'b011;
								assign node116 = (inp[8]) ? node120 : node117;
									assign node117 = (inp[0]) ? 3'b011 : 3'b101;
									assign node120 = (inp[0]) ? 3'b111 : node121;
										assign node121 = (inp[11]) ? 3'b011 : node122;
											assign node122 = (inp[7]) ? 3'b111 : 3'b011;
							assign node127 = (inp[0]) ? 3'b111 : node128;
								assign node128 = (inp[5]) ? node130 : 3'b111;
									assign node130 = (inp[11]) ? 3'b101 : 3'b111;
				assign node134 = (inp[0]) ? node252 : node135;
					assign node135 = (inp[6]) ? node197 : node136;
						assign node136 = (inp[5]) ? node166 : node137;
							assign node137 = (inp[10]) ? node151 : node138;
								assign node138 = (inp[11]) ? node146 : node139;
									assign node139 = (inp[7]) ? node143 : node140;
										assign node140 = (inp[1]) ? 3'b101 : 3'b001;
										assign node143 = (inp[1]) ? 3'b011 : 3'b101;
									assign node146 = (inp[2]) ? 3'b101 : node147;
										assign node147 = (inp[1]) ? 3'b001 : 3'b110;
								assign node151 = (inp[8]) ? node161 : node152;
									assign node152 = (inp[1]) ? node156 : node153;
										assign node153 = (inp[7]) ? 3'b110 : 3'b010;
										assign node156 = (inp[7]) ? 3'b001 : node157;
											assign node157 = (inp[2]) ? 3'b001 : 3'b110;
									assign node161 = (inp[11]) ? node163 : 3'b001;
										assign node163 = (inp[7]) ? 3'b001 : 3'b110;
							assign node166 = (inp[10]) ? node184 : node167;
								assign node167 = (inp[1]) ? node179 : node168;
									assign node168 = (inp[7]) ? node172 : node169;
										assign node169 = (inp[11]) ? 3'b010 : 3'b110;
										assign node172 = (inp[11]) ? 3'b110 : node173;
											assign node173 = (inp[8]) ? 3'b001 : node174;
												assign node174 = (inp[2]) ? 3'b001 : 3'b110;
									assign node179 = (inp[7]) ? 3'b001 : node180;
										assign node180 = (inp[11]) ? 3'b110 : 3'b001;
								assign node184 = (inp[11]) ? node192 : node185;
									assign node185 = (inp[8]) ? node187 : 3'b100;
										assign node187 = (inp[1]) ? 3'b110 : node188;
											assign node188 = (inp[2]) ? 3'b110 : 3'b010;
									assign node192 = (inp[1]) ? node194 : 3'b010;
										assign node194 = (inp[8]) ? 3'b110 : 3'b010;
						assign node197 = (inp[1]) ? node223 : node198;
							assign node198 = (inp[10]) ? node204 : node199;
								assign node199 = (inp[5]) ? node201 : 3'b101;
									assign node201 = (inp[7]) ? 3'b101 : 3'b001;
								assign node204 = (inp[5]) ? node212 : node205;
									assign node205 = (inp[7]) ? node209 : node206;
										assign node206 = (inp[11]) ? 3'b001 : 3'b101;
										assign node209 = (inp[11]) ? 3'b101 : 3'b011;
									assign node212 = (inp[7]) ? node218 : node213;
										assign node213 = (inp[2]) ? 3'b110 : node214;
											assign node214 = (inp[11]) ? 3'b110 : 3'b001;
										assign node218 = (inp[11]) ? node220 : 3'b001;
											assign node220 = (inp[2]) ? 3'b001 : 3'b110;
							assign node223 = (inp[10]) ? node239 : node224;
								assign node224 = (inp[11]) ? node234 : node225;
									assign node225 = (inp[7]) ? node231 : node226;
										assign node226 = (inp[5]) ? node228 : 3'b011;
											assign node228 = (inp[8]) ? 3'b011 : 3'b101;
										assign node231 = (inp[5]) ? 3'b011 : 3'b111;
									assign node234 = (inp[2]) ? node236 : 3'b101;
										assign node236 = (inp[5]) ? 3'b011 : 3'b111;
								assign node239 = (inp[7]) ? node249 : node240;
									assign node240 = (inp[2]) ? 3'b101 : node241;
										assign node241 = (inp[5]) ? 3'b001 : node242;
											assign node242 = (inp[8]) ? 3'b101 : node243;
												assign node243 = (inp[11]) ? 3'b001 : 3'b101;
									assign node249 = (inp[5]) ? 3'b101 : 3'b011;
					assign node252 = (inp[6]) ? node292 : node253;
						assign node253 = (inp[7]) ? node271 : node254;
							assign node254 = (inp[5]) ? node262 : node255;
								assign node255 = (inp[11]) ? node257 : 3'b101;
									assign node257 = (inp[1]) ? 3'b101 : node258;
										assign node258 = (inp[10]) ? 3'b001 : 3'b101;
								assign node262 = (inp[10]) ? node266 : node263;
									assign node263 = (inp[1]) ? 3'b101 : 3'b001;
									assign node266 = (inp[1]) ? 3'b001 : node267;
										assign node267 = (inp[2]) ? 3'b110 : 3'b010;
							assign node271 = (inp[1]) ? node283 : node272;
								assign node272 = (inp[5]) ? 3'b101 : node273;
									assign node273 = (inp[2]) ? node275 : 3'b101;
										assign node275 = (inp[10]) ? node277 : 3'b011;
											assign node277 = (inp[8]) ? node279 : 3'b101;
												assign node279 = (inp[11]) ? 3'b101 : 3'b011;
								assign node283 = (inp[10]) ? node289 : node284;
									assign node284 = (inp[11]) ? 3'b011 : node285;
										assign node285 = (inp[5]) ? 3'b011 : 3'b111;
									assign node289 = (inp[5]) ? 3'b101 : 3'b011;
						assign node292 = (inp[5]) ? node304 : node293;
							assign node293 = (inp[10]) ? node295 : 3'b111;
								assign node295 = (inp[7]) ? 3'b111 : node296;
									assign node296 = (inp[1]) ? node300 : node297;
										assign node297 = (inp[8]) ? 3'b011 : 3'b101;
										assign node300 = (inp[11]) ? 3'b011 : 3'b111;
							assign node304 = (inp[10]) ? node312 : node305;
								assign node305 = (inp[7]) ? 3'b111 : node306;
									assign node306 = (inp[11]) ? 3'b011 : node307;
										assign node307 = (inp[2]) ? 3'b111 : 3'b011;
								assign node312 = (inp[7]) ? node318 : node313;
									assign node313 = (inp[11]) ? node315 : 3'b101;
										assign node315 = (inp[1]) ? 3'b101 : 3'b001;
									assign node318 = (inp[11]) ? 3'b101 : node319;
										assign node319 = (inp[2]) ? 3'b111 : 3'b011;
			assign node323 = (inp[4]) ? node497 : node324;
				assign node324 = (inp[0]) ? node426 : node325;
					assign node325 = (inp[5]) ? node355 : node326;
						assign node326 = (inp[6]) ? node336 : node327;
							assign node327 = (inp[10]) ? node331 : node328;
								assign node328 = (inp[11]) ? 3'b001 : 3'b101;
								assign node331 = (inp[11]) ? node333 : 3'b001;
									assign node333 = (inp[7]) ? 3'b001 : 3'b110;
							assign node336 = (inp[11]) ? node342 : node337;
								assign node337 = (inp[10]) ? 3'b011 : node338;
									assign node338 = (inp[2]) ? 3'b111 : 3'b011;
								assign node342 = (inp[10]) ? node348 : node343;
									assign node343 = (inp[2]) ? 3'b011 : node344;
										assign node344 = (inp[7]) ? 3'b111 : 3'b011;
									assign node348 = (inp[2]) ? 3'b101 : node349;
										assign node349 = (inp[7]) ? node351 : 3'b001;
											assign node351 = (inp[8]) ? 3'b101 : 3'b001;
						assign node355 = (inp[6]) ? node397 : node356;
							assign node356 = (inp[10]) ? node380 : node357;
								assign node357 = (inp[8]) ? node367 : node358;
									assign node358 = (inp[11]) ? 3'b110 : node359;
										assign node359 = (inp[2]) ? 3'b001 : node360;
											assign node360 = (inp[1]) ? 3'b110 : node361;
												assign node361 = (inp[7]) ? 3'b110 : 3'b010;
									assign node367 = (inp[11]) ? node375 : node368;
										assign node368 = (inp[1]) ? node370 : 3'b001;
											assign node370 = (inp[7]) ? node372 : 3'b001;
												assign node372 = (inp[2]) ? 3'b101 : 3'b001;
										assign node375 = (inp[1]) ? 3'b001 : node376;
											assign node376 = (inp[7]) ? 3'b110 : 3'b010;
								assign node380 = (inp[2]) ? node390 : node381;
									assign node381 = (inp[11]) ? node385 : node382;
										assign node382 = (inp[7]) ? 3'b110 : 3'b100;
										assign node385 = (inp[8]) ? node387 : 3'b010;
											assign node387 = (inp[7]) ? 3'b110 : 3'b010;
									assign node390 = (inp[8]) ? node392 : 3'b010;
										assign node392 = (inp[11]) ? 3'b010 : node393;
											assign node393 = (inp[1]) ? 3'b110 : 3'b010;
							assign node397 = (inp[7]) ? node409 : node398;
								assign node398 = (inp[11]) ? node406 : node399;
									assign node399 = (inp[2]) ? node403 : node400;
										assign node400 = (inp[8]) ? 3'b101 : 3'b001;
										assign node403 = (inp[1]) ? 3'b001 : 3'b110;
									assign node406 = (inp[10]) ? 3'b110 : 3'b101;
								assign node409 = (inp[2]) ? node417 : node410;
									assign node410 = (inp[1]) ? node414 : node411;
										assign node411 = (inp[11]) ? 3'b110 : 3'b001;
										assign node414 = (inp[10]) ? 3'b001 : 3'b101;
									assign node417 = (inp[10]) ? node421 : node418;
										assign node418 = (inp[11]) ? 3'b101 : 3'b011;
										assign node421 = (inp[11]) ? node423 : 3'b101;
											assign node423 = (inp[1]) ? 3'b101 : 3'b001;
					assign node426 = (inp[6]) ? node476 : node427;
						assign node427 = (inp[10]) ? node457 : node428;
							assign node428 = (inp[1]) ? node442 : node429;
								assign node429 = (inp[11]) ? 3'b101 : node430;
									assign node430 = (inp[2]) ? node434 : node431;
										assign node431 = (inp[7]) ? 3'b101 : 3'b001;
										assign node434 = (inp[8]) ? 3'b011 : node435;
											assign node435 = (inp[5]) ? 3'b101 : node436;
												assign node436 = (inp[7]) ? 3'b011 : 3'b101;
								assign node442 = (inp[5]) ? node450 : node443;
									assign node443 = (inp[7]) ? node445 : 3'b011;
										assign node445 = (inp[11]) ? node447 : 3'b111;
											assign node447 = (inp[8]) ? 3'b111 : 3'b011;
									assign node450 = (inp[7]) ? node452 : 3'b101;
										assign node452 = (inp[2]) ? 3'b011 : node453;
											assign node453 = (inp[11]) ? 3'b101 : 3'b011;
							assign node457 = (inp[5]) ? node463 : node458;
								assign node458 = (inp[7]) ? node460 : 3'b101;
									assign node460 = (inp[2]) ? 3'b011 : 3'b101;
								assign node463 = (inp[11]) ? node469 : node464;
									assign node464 = (inp[2]) ? 3'b001 : node465;
										assign node465 = (inp[1]) ? 3'b001 : 3'b110;
									assign node469 = (inp[7]) ? node471 : 3'b110;
										assign node471 = (inp[8]) ? node473 : 3'b110;
											assign node473 = (inp[1]) ? 3'b101 : 3'b001;
						assign node476 = (inp[5]) ? node478 : 3'b111;
							assign node478 = (inp[1]) ? node488 : node479;
								assign node479 = (inp[7]) ? node481 : 3'b101;
									assign node481 = (inp[10]) ? node483 : 3'b011;
										assign node483 = (inp[8]) ? node485 : 3'b101;
											assign node485 = (inp[11]) ? 3'b101 : 3'b011;
								assign node488 = (inp[7]) ? 3'b011 : node489;
									assign node489 = (inp[11]) ? node493 : node490;
										assign node490 = (inp[10]) ? 3'b011 : 3'b111;
										assign node493 = (inp[10]) ? 3'b101 : 3'b111;
				assign node497 = (inp[0]) ? node623 : node498;
					assign node498 = (inp[6]) ? node566 : node499;
						assign node499 = (inp[10]) ? node525 : node500;
							assign node500 = (inp[1]) ? node514 : node501;
								assign node501 = (inp[7]) ? node507 : node502;
									assign node502 = (inp[11]) ? node504 : 3'b100;
										assign node504 = (inp[8]) ? 3'b010 : 3'b100;
									assign node507 = (inp[11]) ? node511 : node508;
										assign node508 = (inp[5]) ? 3'b010 : 3'b110;
										assign node511 = (inp[5]) ? 3'b100 : 3'b010;
								assign node514 = (inp[5]) ? 3'b010 : node515;
									assign node515 = (inp[7]) ? node521 : node516;
										assign node516 = (inp[11]) ? 3'b010 : node517;
											assign node517 = (inp[2]) ? 3'b010 : 3'b110;
										assign node521 = (inp[11]) ? 3'b110 : 3'b001;
							assign node525 = (inp[8]) ? node551 : node526;
								assign node526 = (inp[2]) ? node544 : node527;
									assign node527 = (inp[7]) ? node535 : node528;
										assign node528 = (inp[1]) ? node530 : 3'b000;
											assign node530 = (inp[5]) ? 3'b000 : node531;
												assign node531 = (inp[11]) ? 3'b000 : 3'b100;
										assign node535 = (inp[11]) ? node541 : node536;
											assign node536 = (inp[1]) ? node538 : 3'b100;
												assign node538 = (inp[5]) ? 3'b100 : 3'b010;
											assign node541 = (inp[1]) ? 3'b100 : 3'b000;
									assign node544 = (inp[11]) ? node546 : 3'b100;
										assign node546 = (inp[7]) ? 3'b100 : node547;
											assign node547 = (inp[1]) ? 3'b100 : 3'b000;
								assign node551 = (inp[5]) ? node557 : node552;
									assign node552 = (inp[11]) ? node554 : 3'b010;
										assign node554 = (inp[1]) ? 3'b010 : 3'b100;
									assign node557 = (inp[1]) ? node563 : node558;
										assign node558 = (inp[2]) ? node560 : 3'b000;
											assign node560 = (inp[11]) ? 3'b000 : 3'b100;
										assign node563 = (inp[2]) ? 3'b010 : 3'b100;
						assign node566 = (inp[11]) ? node586 : node567;
							assign node567 = (inp[7]) ? node573 : node568;
								assign node568 = (inp[8]) ? node570 : 3'b110;
									assign node570 = (inp[2]) ? 3'b101 : 3'b110;
								assign node573 = (inp[1]) ? 3'b001 : node574;
									assign node574 = (inp[5]) ? node582 : node575;
										assign node575 = (inp[10]) ? node577 : 3'b001;
											assign node577 = (inp[8]) ? node579 : 3'b110;
												assign node579 = (inp[2]) ? 3'b001 : 3'b110;
										assign node582 = (inp[10]) ? 3'b010 : 3'b110;
							assign node586 = (inp[7]) ? node612 : node587;
								assign node587 = (inp[5]) ? node599 : node588;
									assign node588 = (inp[1]) ? node592 : node589;
										assign node589 = (inp[10]) ? 3'b010 : 3'b110;
										assign node592 = (inp[10]) ? node596 : node593;
											assign node593 = (inp[8]) ? 3'b001 : 3'b110;
											assign node596 = (inp[8]) ? 3'b110 : 3'b010;
									assign node599 = (inp[10]) ? node603 : node600;
										assign node600 = (inp[1]) ? 3'b110 : 3'b010;
										assign node603 = (inp[1]) ? node609 : node604;
											assign node604 = (inp[8]) ? 3'b100 : node605;
												assign node605 = (inp[2]) ? 3'b100 : 3'b000;
											assign node609 = (inp[2]) ? 3'b010 : 3'b100;
								assign node612 = (inp[2]) ? 3'b110 : node613;
									assign node613 = (inp[8]) ? node617 : node614;
										assign node614 = (inp[10]) ? 3'b010 : 3'b110;
										assign node617 = (inp[1]) ? 3'b110 : node618;
											assign node618 = (inp[5]) ? 3'b110 : 3'b001;
					assign node623 = (inp[6]) ? node677 : node624;
						assign node624 = (inp[5]) ? node660 : node625;
							assign node625 = (inp[10]) ? node643 : node626;
								assign node626 = (inp[1]) ? node638 : node627;
									assign node627 = (inp[7]) ? node633 : node628;
										assign node628 = (inp[11]) ? 3'b110 : node629;
											assign node629 = (inp[8]) ? 3'b001 : 3'b110;
										assign node633 = (inp[11]) ? node635 : 3'b001;
											assign node635 = (inp[2]) ? 3'b001 : 3'b110;
									assign node638 = (inp[7]) ? node640 : 3'b001;
										assign node640 = (inp[8]) ? 3'b101 : 3'b001;
								assign node643 = (inp[11]) ? node651 : node644;
									assign node644 = (inp[2]) ? node646 : 3'b110;
										assign node646 = (inp[8]) ? 3'b110 : node647;
											assign node647 = (inp[7]) ? 3'b001 : 3'b110;
									assign node651 = (inp[1]) ? node657 : node652;
										assign node652 = (inp[7]) ? node654 : 3'b010;
											assign node654 = (inp[8]) ? 3'b110 : 3'b010;
										assign node657 = (inp[7]) ? 3'b001 : 3'b010;
							assign node660 = (inp[10]) ? node672 : node661;
								assign node661 = (inp[2]) ? node667 : node662;
									assign node662 = (inp[7]) ? 3'b110 : node663;
										assign node663 = (inp[1]) ? 3'b110 : 3'b010;
									assign node667 = (inp[8]) ? 3'b110 : node668;
										assign node668 = (inp[11]) ? 3'b010 : 3'b001;
								assign node672 = (inp[7]) ? 3'b010 : node673;
									assign node673 = (inp[8]) ? 3'b010 : 3'b100;
						assign node677 = (inp[11]) ? node709 : node678;
							assign node678 = (inp[2]) ? node688 : node679;
								assign node679 = (inp[5]) ? node683 : node680;
									assign node680 = (inp[7]) ? 3'b101 : 3'b001;
									assign node683 = (inp[10]) ? 3'b001 : node684;
										assign node684 = (inp[7]) ? 3'b011 : 3'b001;
								assign node688 = (inp[10]) ? node700 : node689;
									assign node689 = (inp[7]) ? node697 : node690;
										assign node690 = (inp[8]) ? node692 : 3'b101;
											assign node692 = (inp[5]) ? node694 : 3'b011;
												assign node694 = (inp[1]) ? 3'b101 : 3'b001;
										assign node697 = (inp[1]) ? 3'b111 : 3'b011;
									assign node700 = (inp[5]) ? node706 : node701;
										assign node701 = (inp[1]) ? 3'b101 : node702;
											assign node702 = (inp[7]) ? 3'b101 : 3'b001;
										assign node706 = (inp[7]) ? 3'b001 : 3'b110;
							assign node709 = (inp[10]) ? node727 : node710;
								assign node710 = (inp[8]) ? node716 : node711;
									assign node711 = (inp[7]) ? 3'b101 : node712;
										assign node712 = (inp[5]) ? 3'b110 : 3'b001;
									assign node716 = (inp[5]) ? node720 : node717;
										assign node717 = (inp[7]) ? 3'b011 : 3'b101;
										assign node720 = (inp[7]) ? node722 : 3'b001;
											assign node722 = (inp[2]) ? 3'b101 : node723;
												assign node723 = (inp[1]) ? 3'b101 : 3'b001;
								assign node727 = (inp[5]) ? node737 : node728;
									assign node728 = (inp[1]) ? node734 : node729;
										assign node729 = (inp[2]) ? 3'b001 : node730;
											assign node730 = (inp[7]) ? 3'b001 : 3'b110;
										assign node734 = (inp[7]) ? 3'b101 : 3'b001;
									assign node737 = (inp[7]) ? node741 : node738;
										assign node738 = (inp[2]) ? 3'b010 : 3'b110;
										assign node741 = (inp[8]) ? node743 : 3'b110;
											assign node743 = (inp[2]) ? 3'b110 : 3'b001;
		assign node746 = (inp[9]) ? node1124 : node747;
			assign node747 = (inp[4]) ? node981 : node748;
				assign node748 = (inp[6]) ? node870 : node749;
					assign node749 = (inp[0]) ? node801 : node750;
						assign node750 = (inp[10]) ? node774 : node751;
							assign node751 = (inp[5]) ? node763 : node752;
								assign node752 = (inp[1]) ? node758 : node753;
									assign node753 = (inp[7]) ? node755 : 3'b010;
										assign node755 = (inp[11]) ? 3'b010 : 3'b110;
									assign node758 = (inp[11]) ? 3'b110 : node759;
										assign node759 = (inp[2]) ? 3'b001 : 3'b110;
								assign node763 = (inp[7]) ? node769 : node764;
									assign node764 = (inp[1]) ? 3'b100 : node765;
										assign node765 = (inp[2]) ? 3'b100 : 3'b000;
									assign node769 = (inp[2]) ? 3'b010 : node770;
										assign node770 = (inp[8]) ? 3'b010 : 3'b100;
							assign node774 = (inp[5]) ? node794 : node775;
								assign node775 = (inp[11]) ? node783 : node776;
									assign node776 = (inp[7]) ? 3'b010 : node777;
										assign node777 = (inp[8]) ? 3'b010 : node778;
											assign node778 = (inp[1]) ? 3'b100 : 3'b000;
									assign node783 = (inp[1]) ? node791 : node784;
										assign node784 = (inp[7]) ? 3'b100 : node785;
											assign node785 = (inp[2]) ? node787 : 3'b000;
												assign node787 = (inp[8]) ? 3'b100 : 3'b000;
										assign node791 = (inp[8]) ? 3'b010 : 3'b100;
								assign node794 = (inp[11]) ? 3'b000 : node795;
									assign node795 = (inp[7]) ? node797 : 3'b000;
										assign node797 = (inp[2]) ? 3'b000 : 3'b100;
						assign node801 = (inp[5]) ? node833 : node802;
							assign node802 = (inp[7]) ? node822 : node803;
								assign node803 = (inp[1]) ? node811 : node804;
									assign node804 = (inp[10]) ? node806 : 3'b110;
										assign node806 = (inp[8]) ? node808 : 3'b100;
											assign node808 = (inp[2]) ? 3'b110 : 3'b010;
									assign node811 = (inp[10]) ? node819 : node812;
										assign node812 = (inp[2]) ? node816 : node813;
											assign node813 = (inp[11]) ? 3'b110 : 3'b001;
											assign node816 = (inp[8]) ? 3'b101 : 3'b001;
										assign node819 = (inp[11]) ? 3'b010 : 3'b110;
								assign node822 = (inp[10]) ? node828 : node823;
									assign node823 = (inp[11]) ? 3'b001 : node824;
										assign node824 = (inp[1]) ? 3'b101 : 3'b001;
									assign node828 = (inp[1]) ? node830 : 3'b110;
										assign node830 = (inp[11]) ? 3'b110 : 3'b001;
							assign node833 = (inp[10]) ? node851 : node834;
								assign node834 = (inp[11]) ? node846 : node835;
									assign node835 = (inp[7]) ? node841 : node836;
										assign node836 = (inp[2]) ? 3'b110 : node837;
											assign node837 = (inp[8]) ? 3'b110 : 3'b010;
										assign node841 = (inp[8]) ? 3'b001 : node842;
											assign node842 = (inp[1]) ? 3'b001 : 3'b110;
									assign node846 = (inp[7]) ? 3'b110 : node847;
										assign node847 = (inp[8]) ? 3'b110 : 3'b010;
								assign node851 = (inp[8]) ? node857 : node852;
									assign node852 = (inp[2]) ? 3'b100 : node853;
										assign node853 = (inp[11]) ? 3'b000 : 3'b100;
									assign node857 = (inp[11]) ? node863 : node858;
										assign node858 = (inp[1]) ? node860 : 3'b010;
											assign node860 = (inp[7]) ? 3'b110 : 3'b010;
										assign node863 = (inp[7]) ? node865 : 3'b100;
											assign node865 = (inp[1]) ? 3'b010 : node866;
												assign node866 = (inp[2]) ? 3'b010 : 3'b100;
					assign node870 = (inp[0]) ? node930 : node871;
						assign node871 = (inp[5]) ? node909 : node872;
							assign node872 = (inp[2]) ? node894 : node873;
								assign node873 = (inp[10]) ? node887 : node874;
									assign node874 = (inp[11]) ? node876 : 3'b001;
										assign node876 = (inp[8]) ? node882 : node877;
											assign node877 = (inp[7]) ? node879 : 3'b110;
												assign node879 = (inp[1]) ? 3'b001 : 3'b110;
											assign node882 = (inp[7]) ? 3'b001 : node883;
												assign node883 = (inp[1]) ? 3'b001 : 3'b110;
									assign node887 = (inp[7]) ? 3'b110 : node888;
										assign node888 = (inp[1]) ? node890 : 3'b010;
											assign node890 = (inp[8]) ? 3'b110 : 3'b010;
								assign node894 = (inp[1]) ? node900 : node895;
									assign node895 = (inp[8]) ? node897 : 3'b110;
										assign node897 = (inp[10]) ? 3'b001 : 3'b101;
									assign node900 = (inp[10]) ? 3'b001 : node901;
										assign node901 = (inp[11]) ? node905 : node902;
											assign node902 = (inp[7]) ? 3'b011 : 3'b101;
											assign node905 = (inp[7]) ? 3'b101 : 3'b001;
							assign node909 = (inp[1]) ? node919 : node910;
								assign node910 = (inp[11]) ? 3'b010 : node911;
									assign node911 = (inp[2]) ? 3'b110 : node912;
										assign node912 = (inp[7]) ? node914 : 3'b010;
											assign node914 = (inp[10]) ? 3'b010 : 3'b110;
								assign node919 = (inp[11]) ? node923 : node920;
									assign node920 = (inp[10]) ? 3'b110 : 3'b001;
									assign node923 = (inp[10]) ? node925 : 3'b110;
										assign node925 = (inp[7]) ? 3'b010 : node926;
											assign node926 = (inp[2]) ? 3'b010 : 3'b100;
						assign node930 = (inp[11]) ? node956 : node931;
							assign node931 = (inp[7]) ? node945 : node932;
								assign node932 = (inp[5]) ? node938 : node933;
									assign node933 = (inp[1]) ? node935 : 3'b001;
										assign node935 = (inp[2]) ? 3'b101 : 3'b001;
									assign node938 = (inp[10]) ? node940 : 3'b001;
										assign node940 = (inp[2]) ? 3'b110 : node941;
											assign node941 = (inp[8]) ? 3'b110 : 3'b010;
								assign node945 = (inp[5]) ? node951 : node946;
									assign node946 = (inp[10]) ? 3'b011 : node947;
										assign node947 = (inp[1]) ? 3'b111 : 3'b011;
									assign node951 = (inp[10]) ? 3'b001 : node952;
										assign node952 = (inp[8]) ? 3'b011 : 3'b101;
							assign node956 = (inp[1]) ? node962 : node957;
								assign node957 = (inp[8]) ? node959 : 3'b110;
									assign node959 = (inp[5]) ? 3'b110 : 3'b101;
								assign node962 = (inp[2]) ? node972 : node963;
									assign node963 = (inp[10]) ? node965 : 3'b101;
										assign node965 = (inp[8]) ? 3'b001 : node966;
											assign node966 = (inp[5]) ? node968 : 3'b001;
												assign node968 = (inp[7]) ? 3'b001 : 3'b110;
									assign node972 = (inp[10]) ? node978 : node973;
										assign node973 = (inp[5]) ? node975 : 3'b011;
											assign node975 = (inp[8]) ? 3'b101 : 3'b001;
										assign node978 = (inp[8]) ? 3'b101 : 3'b110;
				assign node981 = (inp[6]) ? node1035 : node982;
					assign node982 = (inp[0]) ? node992 : node983;
						assign node983 = (inp[10]) ? 3'b000 : node984;
							assign node984 = (inp[1]) ? node986 : 3'b000;
								assign node986 = (inp[2]) ? node988 : 3'b000;
									assign node988 = (inp[5]) ? 3'b000 : 3'b100;
						assign node992 = (inp[5]) ? node1012 : node993;
							assign node993 = (inp[10]) ? node1003 : node994;
								assign node994 = (inp[1]) ? 3'b010 : node995;
									assign node995 = (inp[7]) ? node997 : 3'b100;
										assign node997 = (inp[2]) ? 3'b010 : node998;
											assign node998 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1003 = (inp[11]) ? node1005 : 3'b100;
									assign node1005 = (inp[2]) ? node1009 : node1006;
										assign node1006 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1009 = (inp[1]) ? 3'b010 : 3'b000;
							assign node1012 = (inp[11]) ? node1026 : node1013;
								assign node1013 = (inp[8]) ? 3'b100 : node1014;
									assign node1014 = (inp[10]) ? node1018 : node1015;
										assign node1015 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1018 = (inp[1]) ? node1020 : 3'b000;
											assign node1020 = (inp[2]) ? node1022 : 3'b000;
												assign node1022 = (inp[7]) ? 3'b100 : 3'b000;
								assign node1026 = (inp[7]) ? node1028 : 3'b000;
									assign node1028 = (inp[2]) ? node1032 : node1029;
										assign node1029 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1032 = (inp[10]) ? 3'b000 : 3'b010;
					assign node1035 = (inp[0]) ? node1087 : node1036;
						assign node1036 = (inp[10]) ? node1062 : node1037;
							assign node1037 = (inp[5]) ? node1049 : node1038;
								assign node1038 = (inp[11]) ? node1046 : node1039;
									assign node1039 = (inp[7]) ? node1043 : node1040;
										assign node1040 = (inp[8]) ? 3'b110 : 3'b100;
										assign node1043 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1046 = (inp[7]) ? 3'b110 : 3'b010;
								assign node1049 = (inp[7]) ? node1053 : node1050;
									assign node1050 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1053 = (inp[2]) ? node1059 : node1054;
										assign node1054 = (inp[8]) ? 3'b100 : node1055;
											assign node1055 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1059 = (inp[8]) ? 3'b010 : 3'b100;
							assign node1062 = (inp[1]) ? node1074 : node1063;
								assign node1063 = (inp[8]) ? node1065 : 3'b000;
									assign node1065 = (inp[5]) ? 3'b000 : node1066;
										assign node1066 = (inp[11]) ? node1070 : node1067;
											assign node1067 = (inp[7]) ? 3'b010 : 3'b100;
											assign node1070 = (inp[7]) ? 3'b100 : 3'b000;
								assign node1074 = (inp[8]) ? node1080 : node1075;
									assign node1075 = (inp[7]) ? 3'b100 : node1076;
										assign node1076 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1080 = (inp[7]) ? node1084 : node1081;
										assign node1081 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1084 = (inp[5]) ? 3'b100 : 3'b010;
						assign node1087 = (inp[5]) ? node1103 : node1088;
							assign node1088 = (inp[11]) ? node1096 : node1089;
								assign node1089 = (inp[1]) ? node1091 : 3'b110;
									assign node1091 = (inp[10]) ? 3'b110 : node1092;
										assign node1092 = (inp[7]) ? 3'b101 : 3'b001;
								assign node1096 = (inp[10]) ? node1098 : 3'b110;
									assign node1098 = (inp[7]) ? node1100 : 3'b010;
										assign node1100 = (inp[1]) ? 3'b110 : 3'b010;
							assign node1103 = (inp[10]) ? node1115 : node1104;
								assign node1104 = (inp[1]) ? 3'b010 : node1105;
									assign node1105 = (inp[11]) ? node1111 : node1106;
										assign node1106 = (inp[2]) ? node1108 : 3'b010;
											assign node1108 = (inp[7]) ? 3'b110 : 3'b010;
										assign node1111 = (inp[7]) ? 3'b110 : 3'b100;
								assign node1115 = (inp[11]) ? node1119 : node1116;
									assign node1116 = (inp[7]) ? 3'b010 : 3'b100;
									assign node1119 = (inp[1]) ? 3'b100 : node1120;
										assign node1120 = (inp[7]) ? 3'b100 : 3'b000;
			assign node1124 = (inp[4]) ? node1280 : node1125;
				assign node1125 = (inp[6]) ? node1175 : node1126;
					assign node1126 = (inp[0]) ? node1136 : node1127;
						assign node1127 = (inp[10]) ? 3'b000 : node1128;
							assign node1128 = (inp[5]) ? 3'b000 : node1129;
								assign node1129 = (inp[1]) ? node1131 : 3'b000;
									assign node1131 = (inp[7]) ? 3'b100 : 3'b000;
						assign node1136 = (inp[5]) ? node1156 : node1137;
							assign node1137 = (inp[1]) ? node1145 : node1138;
								assign node1138 = (inp[2]) ? node1140 : 3'b100;
									assign node1140 = (inp[10]) ? node1142 : 3'b010;
										assign node1142 = (inp[8]) ? 3'b100 : 3'b000;
								assign node1145 = (inp[10]) ? node1151 : node1146;
									assign node1146 = (inp[7]) ? node1148 : 3'b010;
										assign node1148 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1151 = (inp[8]) ? 3'b100 : node1152;
										assign node1152 = (inp[11]) ? 3'b000 : 3'b010;
							assign node1156 = (inp[7]) ? node1164 : node1157;
								assign node1157 = (inp[8]) ? node1159 : 3'b000;
									assign node1159 = (inp[10]) ? 3'b000 : node1160;
										assign node1160 = (inp[1]) ? 3'b100 : 3'b000;
								assign node1164 = (inp[10]) ? node1170 : node1165;
									assign node1165 = (inp[11]) ? 3'b100 : node1166;
										assign node1166 = (inp[1]) ? 3'b010 : 3'b100;
									assign node1170 = (inp[11]) ? 3'b000 : node1171;
										assign node1171 = (inp[8]) ? 3'b100 : 3'b000;
					assign node1175 = (inp[10]) ? node1231 : node1176;
						assign node1176 = (inp[5]) ? node1210 : node1177;
							assign node1177 = (inp[2]) ? node1195 : node1178;
								assign node1178 = (inp[0]) ? node1186 : node1179;
									assign node1179 = (inp[1]) ? node1181 : 3'b000;
										assign node1181 = (inp[7]) ? node1183 : 3'b010;
											assign node1183 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1186 = (inp[7]) ? 3'b110 : node1187;
										assign node1187 = (inp[11]) ? 3'b010 : node1188;
											assign node1188 = (inp[8]) ? 3'b110 : node1189;
												assign node1189 = (inp[1]) ? 3'b110 : 3'b010;
								assign node1195 = (inp[8]) ? node1199 : node1196;
									assign node1196 = (inp[0]) ? 3'b001 : 3'b010;
									assign node1199 = (inp[7]) ? node1205 : node1200;
										assign node1200 = (inp[0]) ? 3'b110 : node1201;
											assign node1201 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1205 = (inp[0]) ? node1207 : 3'b110;
											assign node1207 = (inp[1]) ? 3'b101 : 3'b001;
							assign node1210 = (inp[0]) ? node1218 : node1211;
								assign node1211 = (inp[11]) ? node1213 : 3'b100;
									assign node1213 = (inp[2]) ? 3'b010 : node1214;
										assign node1214 = (inp[7]) ? 3'b100 : 3'b000;
								assign node1218 = (inp[7]) ? 3'b110 : node1219;
									assign node1219 = (inp[2]) ? node1223 : node1220;
										assign node1220 = (inp[11]) ? 3'b100 : 3'b110;
										assign node1223 = (inp[8]) ? 3'b010 : node1224;
											assign node1224 = (inp[11]) ? node1226 : 3'b010;
												assign node1226 = (inp[1]) ? 3'b010 : 3'b100;
						assign node1231 = (inp[0]) ? node1251 : node1232;
							assign node1232 = (inp[5]) ? node1244 : node1233;
								assign node1233 = (inp[8]) ? node1239 : node1234;
									assign node1234 = (inp[7]) ? 3'b010 : node1235;
										assign node1235 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1239 = (inp[11]) ? node1241 : 3'b100;
										assign node1241 = (inp[1]) ? 3'b100 : 3'b000;
								assign node1244 = (inp[2]) ? node1246 : 3'b000;
									assign node1246 = (inp[8]) ? 3'b000 : node1247;
										assign node1247 = (inp[11]) ? 3'b000 : 3'b100;
							assign node1251 = (inp[5]) ? node1265 : node1252;
								assign node1252 = (inp[7]) ? node1258 : node1253;
									assign node1253 = (inp[8]) ? 3'b010 : node1254;
										assign node1254 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1258 = (inp[11]) ? 3'b010 : node1259;
										assign node1259 = (inp[8]) ? 3'b110 : node1260;
											assign node1260 = (inp[2]) ? 3'b110 : 3'b010;
								assign node1265 = (inp[2]) ? node1273 : node1266;
									assign node1266 = (inp[1]) ? node1268 : 3'b000;
										assign node1268 = (inp[8]) ? 3'b010 : node1269;
											assign node1269 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1273 = (inp[8]) ? 3'b100 : node1274;
										assign node1274 = (inp[1]) ? 3'b100 : node1275;
											assign node1275 = (inp[7]) ? 3'b100 : 3'b000;
				assign node1280 = (inp[6]) ? node1282 : 3'b000;
					assign node1282 = (inp[0]) ? node1294 : node1283;
						assign node1283 = (inp[8]) ? node1285 : 3'b000;
							assign node1285 = (inp[1]) ? node1287 : 3'b000;
								assign node1287 = (inp[5]) ? 3'b000 : node1288;
									assign node1288 = (inp[2]) ? node1290 : 3'b000;
										assign node1290 = (inp[7]) ? 3'b100 : 3'b000;
						assign node1294 = (inp[10]) ? node1314 : node1295;
							assign node1295 = (inp[7]) ? node1299 : node1296;
								assign node1296 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1299 = (inp[5]) ? node1305 : node1300;
									assign node1300 = (inp[2]) ? 3'b010 : node1301;
										assign node1301 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1305 = (inp[2]) ? node1307 : 3'b100;
										assign node1307 = (inp[8]) ? node1311 : node1308;
											assign node1308 = (inp[1]) ? 3'b100 : 3'b000;
											assign node1311 = (inp[1]) ? 3'b010 : 3'b100;
							assign node1314 = (inp[11]) ? 3'b000 : node1315;
								assign node1315 = (inp[1]) ? node1317 : 3'b000;
									assign node1317 = (inp[7]) ? node1319 : 3'b000;
										assign node1319 = (inp[5]) ? node1321 : 3'b100;
											assign node1321 = (inp[8]) ? node1323 : 3'b000;
												assign node1323 = (inp[2]) ? 3'b100 : 3'b000;

endmodule