module dtc_split75_bm50 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node5;
	wire [2-1:0] node6;
	wire [2-1:0] node9;
	wire [2-1:0] node12;
	wire [2-1:0] node13;
	wire [2-1:0] node16;
	wire [2-1:0] node19;
	wire [2-1:0] node20;
	wire [2-1:0] node21;
	wire [2-1:0] node22;
	wire [2-1:0] node25;
	wire [2-1:0] node28;
	wire [2-1:0] node30;
	wire [2-1:0] node33;
	wire [2-1:0] node35;
	wire [2-1:0] node36;
	wire [2-1:0] node39;
	wire [2-1:0] node42;
	wire [2-1:0] node43;
	wire [2-1:0] node44;
	wire [2-1:0] node46;
	wire [2-1:0] node47;
	wire [2-1:0] node50;
	wire [2-1:0] node53;
	wire [2-1:0] node54;
	wire [2-1:0] node55;
	wire [2-1:0] node58;
	wire [2-1:0] node61;
	wire [2-1:0] node62;
	wire [2-1:0] node65;
	wire [2-1:0] node68;
	wire [2-1:0] node69;
	wire [2-1:0] node70;
	wire [2-1:0] node72;
	wire [2-1:0] node75;
	wire [2-1:0] node78;
	wire [2-1:0] node79;
	wire [2-1:0] node80;
	wire [2-1:0] node83;
	wire [2-1:0] node87;
	wire [2-1:0] node88;
	wire [2-1:0] node89;
	wire [2-1:0] node90;
	wire [2-1:0] node92;
	wire [2-1:0] node93;
	wire [2-1:0] node97;
	wire [2-1:0] node98;
	wire [2-1:0] node101;
	wire [2-1:0] node102;
	wire [2-1:0] node105;
	wire [2-1:0] node108;
	wire [2-1:0] node109;
	wire [2-1:0] node110;
	wire [2-1:0] node115;
	wire [2-1:0] node116;
	wire [2-1:0] node117;
	wire [2-1:0] node118;
	wire [2-1:0] node121;
	wire [2-1:0] node124;
	wire [2-1:0] node125;
	wire [2-1:0] node128;
	wire [2-1:0] node131;
	wire [2-1:0] node132;
	wire [2-1:0] node133;
	wire [2-1:0] node136;
	wire [2-1:0] node139;
	wire [2-1:0] node140;
	wire [2-1:0] node141;
	wire [2-1:0] node145;
	wire [2-1:0] node146;
	wire [2-1:0] node149;
	wire [2-1:0] node152;
	wire [2-1:0] node153;
	wire [2-1:0] node154;
	wire [2-1:0] node155;
	wire [2-1:0] node156;
	wire [2-1:0] node157;
	wire [2-1:0] node159;
	wire [2-1:0] node162;
	wire [2-1:0] node163;
	wire [2-1:0] node166;
	wire [2-1:0] node169;
	wire [2-1:0] node170;
	wire [2-1:0] node173;
	wire [2-1:0] node176;
	wire [2-1:0] node177;
	wire [2-1:0] node178;
	wire [2-1:0] node182;
	wire [2-1:0] node185;
	wire [2-1:0] node186;
	wire [2-1:0] node187;
	wire [2-1:0] node188;
	wire [2-1:0] node191;
	wire [2-1:0] node194;
	wire [2-1:0] node195;
	wire [2-1:0] node198;
	wire [2-1:0] node201;
	wire [2-1:0] node202;
	wire [2-1:0] node204;
	wire [2-1:0] node207;
	wire [2-1:0] node208;
	wire [2-1:0] node209;
	wire [2-1:0] node213;
	wire [2-1:0] node216;
	wire [2-1:0] node217;
	wire [2-1:0] node218;
	wire [2-1:0] node219;
	wire [2-1:0] node220;
	wire [2-1:0] node224;
	wire [2-1:0] node225;
	wire [2-1:0] node229;
	wire [2-1:0] node230;
	wire [2-1:0] node231;
	wire [2-1:0] node232;
	wire [2-1:0] node236;
	wire [2-1:0] node239;
	wire [2-1:0] node241;
	wire [2-1:0] node243;
	wire [2-1:0] node246;
	wire [2-1:0] node247;
	wire [2-1:0] node248;
	wire [2-1:0] node249;
	wire [2-1:0] node252;
	wire [2-1:0] node255;
	wire [2-1:0] node256;
	wire [2-1:0] node259;
	wire [2-1:0] node262;
	wire [2-1:0] node263;
	wire [2-1:0] node264;
	wire [2-1:0] node267;

	assign outp = (inp[2]) ? node152 : node1;
		assign node1 = (inp[7]) ? node87 : node2;
			assign node2 = (inp[4]) ? node42 : node3;
				assign node3 = (inp[6]) ? node19 : node4;
					assign node4 = (inp[0]) ? node12 : node5;
						assign node5 = (inp[1]) ? node9 : node6;
							assign node6 = (inp[5]) ? 2'b01 : 2'b11;
							assign node9 = (inp[5]) ? 2'b11 : 2'b01;
						assign node12 = (inp[5]) ? node16 : node13;
							assign node13 = (inp[1]) ? 2'b00 : 2'b10;
							assign node16 = (inp[1]) ? 2'b10 : 2'b00;
					assign node19 = (inp[0]) ? node33 : node20;
						assign node20 = (inp[3]) ? node28 : node21;
							assign node21 = (inp[1]) ? node25 : node22;
								assign node22 = (inp[5]) ? 2'b00 : 2'b10;
								assign node25 = (inp[5]) ? 2'b10 : 2'b00;
							assign node28 = (inp[1]) ? node30 : 2'b10;
								assign node30 = (inp[5]) ? 2'b10 : 2'b00;
						assign node33 = (inp[5]) ? node35 : 2'b11;
							assign node35 = (inp[1]) ? node39 : node36;
								assign node36 = (inp[3]) ? 2'b11 : 2'b01;
								assign node39 = (inp[3]) ? 2'b01 : 2'b11;
				assign node42 = (inp[5]) ? node68 : node43;
					assign node43 = (inp[1]) ? node53 : node44;
						assign node44 = (inp[3]) ? node46 : 2'b10;
							assign node46 = (inp[6]) ? node50 : node47;
								assign node47 = (inp[0]) ? 2'b00 : 2'b01;
								assign node50 = (inp[0]) ? 2'b01 : 2'b00;
						assign node53 = (inp[3]) ? node61 : node54;
							assign node54 = (inp[6]) ? node58 : node55;
								assign node55 = (inp[0]) ? 2'b00 : 2'b01;
								assign node58 = (inp[0]) ? 2'b11 : 2'b00;
							assign node61 = (inp[0]) ? node65 : node62;
								assign node62 = (inp[6]) ? 2'b10 : 2'b11;
								assign node65 = (inp[6]) ? 2'b11 : 2'b10;
					assign node68 = (inp[1]) ? node78 : node69;
						assign node69 = (inp[0]) ? node75 : node70;
							assign node70 = (inp[6]) ? node72 : 2'b11;
								assign node72 = (inp[3]) ? 2'b10 : 2'b00;
							assign node75 = (inp[6]) ? 2'b11 : 2'b10;
						assign node78 = (inp[3]) ? 2'b00 : node79;
							assign node79 = (inp[6]) ? node83 : node80;
								assign node80 = (inp[0]) ? 2'b10 : 2'b11;
								assign node83 = (inp[0]) ? 2'b01 : 2'b10;
			assign node87 = (inp[4]) ? node115 : node88;
				assign node88 = (inp[1]) ? node108 : node89;
					assign node89 = (inp[6]) ? node97 : node90;
						assign node90 = (inp[0]) ? node92 : 2'b00;
							assign node92 = (inp[5]) ? 2'b11 : node93;
								assign node93 = (inp[3]) ? 2'b01 : 2'b11;
						assign node97 = (inp[0]) ? node101 : node98;
							assign node98 = (inp[5]) ? 2'b01 : 2'b11;
							assign node101 = (inp[5]) ? node105 : node102;
								assign node102 = (inp[3]) ? 2'b00 : 2'b10;
								assign node105 = (inp[3]) ? 2'b10 : 2'b00;
					assign node108 = (inp[6]) ? 2'b00 : node109;
						assign node109 = (inp[0]) ? 2'b11 : node110;
							assign node110 = (inp[5]) ? 2'b10 : 2'b00;
				assign node115 = (inp[0]) ? node131 : node116;
					assign node116 = (inp[6]) ? node124 : node117;
						assign node117 = (inp[5]) ? node121 : node118;
							assign node118 = (inp[3]) ? 2'b00 : 2'b10;
							assign node121 = (inp[3]) ? 2'b10 : 2'b00;
						assign node124 = (inp[5]) ? node128 : node125;
							assign node125 = (inp[1]) ? 2'b11 : 2'b01;
							assign node128 = (inp[1]) ? 2'b01 : 2'b11;
					assign node131 = (inp[6]) ? node139 : node132;
						assign node132 = (inp[1]) ? node136 : node133;
							assign node133 = (inp[5]) ? 2'b11 : 2'b01;
							assign node136 = (inp[3]) ? 2'b11 : 2'b01;
						assign node139 = (inp[3]) ? node145 : node140;
							assign node140 = (inp[1]) ? 2'b00 : node141;
								assign node141 = (inp[5]) ? 2'b10 : 2'b00;
							assign node145 = (inp[1]) ? node149 : node146;
								assign node146 = (inp[5]) ? 2'b10 : 2'b00;
								assign node149 = (inp[5]) ? 2'b00 : 2'b10;
		assign node152 = (inp[5]) ? node216 : node153;
			assign node153 = (inp[1]) ? node185 : node154;
				assign node154 = (inp[4]) ? node176 : node155;
					assign node155 = (inp[3]) ? node169 : node156;
						assign node156 = (inp[6]) ? node162 : node157;
							assign node157 = (inp[7]) ? node159 : 2'b11;
								assign node159 = (inp[0]) ? 2'b10 : 2'b11;
							assign node162 = (inp[7]) ? node166 : node163;
								assign node163 = (inp[0]) ? 2'b11 : 2'b10;
								assign node166 = (inp[0]) ? 2'b10 : 2'b11;
						assign node169 = (inp[7]) ? node173 : node170;
							assign node170 = (inp[0]) ? 2'b01 : 2'b10;
							assign node173 = (inp[0]) ? 2'b00 : 2'b01;
					assign node176 = (inp[7]) ? node182 : node177;
						assign node177 = (inp[0]) ? 2'b01 : node178;
							assign node178 = (inp[3]) ? 2'b00 : 2'b10;
						assign node182 = (inp[0]) ? 2'b00 : 2'b01;
				assign node185 = (inp[3]) ? node201 : node186;
					assign node186 = (inp[4]) ? node194 : node187;
						assign node187 = (inp[7]) ? node191 : node188;
							assign node188 = (inp[0]) ? 2'b01 : 2'b00;
							assign node191 = (inp[0]) ? 2'b00 : 2'b01;
						assign node194 = (inp[0]) ? node198 : node195;
							assign node195 = (inp[7]) ? 2'b11 : 2'b00;
							assign node198 = (inp[7]) ? 2'b10 : 2'b11;
					assign node201 = (inp[6]) ? node207 : node202;
						assign node202 = (inp[7]) ? node204 : 2'b11;
							assign node204 = (inp[0]) ? 2'b10 : 2'b11;
						assign node207 = (inp[0]) ? node213 : node208;
							assign node208 = (inp[7]) ? 2'b11 : node209;
								assign node209 = (inp[4]) ? 2'b10 : 2'b00;
							assign node213 = (inp[7]) ? 2'b10 : 2'b11;
			assign node216 = (inp[1]) ? node246 : node217;
				assign node217 = (inp[4]) ? node229 : node218;
					assign node218 = (inp[3]) ? node224 : node219;
						assign node219 = (inp[0]) ? 2'b00 : node220;
							assign node220 = (inp[7]) ? 2'b01 : 2'b00;
						assign node224 = (inp[0]) ? 2'b11 : node225;
							assign node225 = (inp[7]) ? 2'b11 : 2'b00;
					assign node229 = (inp[6]) ? node239 : node230;
						assign node230 = (inp[7]) ? node236 : node231;
							assign node231 = (inp[0]) ? 2'b11 : node232;
								assign node232 = (inp[3]) ? 2'b10 : 2'b00;
							assign node236 = (inp[0]) ? 2'b10 : 2'b11;
						assign node239 = (inp[3]) ? node241 : 2'b11;
							assign node241 = (inp[0]) ? node243 : 2'b11;
								assign node243 = (inp[7]) ? 2'b10 : 2'b11;
				assign node246 = (inp[4]) ? node262 : node247;
					assign node247 = (inp[3]) ? node255 : node248;
						assign node248 = (inp[7]) ? node252 : node249;
							assign node249 = (inp[0]) ? 2'b11 : 2'b10;
							assign node252 = (inp[0]) ? 2'b10 : 2'b11;
						assign node255 = (inp[0]) ? node259 : node256;
							assign node256 = (inp[7]) ? 2'b01 : 2'b10;
							assign node259 = (inp[7]) ? 2'b00 : 2'b01;
					assign node262 = (inp[3]) ? 2'b01 : node263;
						assign node263 = (inp[0]) ? node267 : node264;
							assign node264 = (inp[7]) ? 2'b01 : 2'b10;
							assign node267 = (inp[7]) ? 2'b00 : 2'b01;

endmodule