module dtc_split875_bm79 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node215;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node334;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node377;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node415;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node449;
	wire [3-1:0] node451;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node461;
	wire [3-1:0] node463;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node492;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node509;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node521;
	wire [3-1:0] node523;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node534;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node544;
	wire [3-1:0] node548;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node584;
	wire [3-1:0] node586;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node614;
	wire [3-1:0] node616;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node674;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node682;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node689;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node697;
	wire [3-1:0] node699;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node724;
	wire [3-1:0] node728;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node747;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node759;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node780;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node785;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node812;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node822;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node835;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node849;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node856;
	wire [3-1:0] node857;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node864;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node882;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node895;
	wire [3-1:0] node897;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node903;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node912;
	wire [3-1:0] node916;
	wire [3-1:0] node918;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node930;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node943;
	wire [3-1:0] node947;
	wire [3-1:0] node949;
	wire [3-1:0] node952;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node961;
	wire [3-1:0] node964;
	wire [3-1:0] node966;
	wire [3-1:0] node968;
	wire [3-1:0] node971;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node978;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node985;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1001;
	wire [3-1:0] node1005;
	wire [3-1:0] node1007;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1021;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1034;
	wire [3-1:0] node1036;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1045;
	wire [3-1:0] node1047;
	wire [3-1:0] node1050;
	wire [3-1:0] node1051;
	wire [3-1:0] node1055;
	wire [3-1:0] node1057;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1064;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1080;
	wire [3-1:0] node1082;
	wire [3-1:0] node1086;
	wire [3-1:0] node1089;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1092;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1107;
	wire [3-1:0] node1108;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1117;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1124;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1138;
	wire [3-1:0] node1139;
	wire [3-1:0] node1141;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1155;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1162;
	wire [3-1:0] node1163;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1168;
	wire [3-1:0] node1172;
	wire [3-1:0] node1174;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1180;
	wire [3-1:0] node1182;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1189;
	wire [3-1:0] node1193;
	wire [3-1:0] node1194;
	wire [3-1:0] node1195;
	wire [3-1:0] node1197;
	wire [3-1:0] node1201;
	wire [3-1:0] node1202;
	wire [3-1:0] node1204;
	wire [3-1:0] node1206;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1214;
	wire [3-1:0] node1215;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1224;
	wire [3-1:0] node1226;
	wire [3-1:0] node1227;
	wire [3-1:0] node1231;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1242;
	wire [3-1:0] node1243;
	wire [3-1:0] node1244;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1250;
	wire [3-1:0] node1252;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1259;
	wire [3-1:0] node1263;
	wire [3-1:0] node1265;
	wire [3-1:0] node1267;
	wire [3-1:0] node1270;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1276;
	wire [3-1:0] node1279;
	wire [3-1:0] node1281;
	wire [3-1:0] node1283;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1292;
	wire [3-1:0] node1294;
	wire [3-1:0] node1295;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1306;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1314;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1329;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1333;
	wire [3-1:0] node1334;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;

	assign outp = (inp[6]) ? node394 : node1;
		assign node1 = (inp[9]) ? node351 : node2;
			assign node2 = (inp[0]) ? node262 : node3;
				assign node3 = (inp[7]) ? node103 : node4;
					assign node4 = (inp[10]) ? node78 : node5;
						assign node5 = (inp[1]) ? node53 : node6;
							assign node6 = (inp[11]) ? node32 : node7;
								assign node7 = (inp[2]) ? node17 : node8;
									assign node8 = (inp[4]) ? 3'b110 : node9;
										assign node9 = (inp[5]) ? 3'b110 : node10;
											assign node10 = (inp[8]) ? node12 : 3'b100;
												assign node12 = (inp[3]) ? 3'b110 : 3'b010;
									assign node17 = (inp[3]) ? node25 : node18;
										assign node18 = (inp[8]) ? 3'b110 : node19;
											assign node19 = (inp[5]) ? node21 : 3'b110;
												assign node21 = (inp[4]) ? 3'b010 : 3'b110;
										assign node25 = (inp[5]) ? 3'b000 : node26;
											assign node26 = (inp[8]) ? node28 : 3'b010;
												assign node28 = (inp[4]) ? 3'b010 : 3'b110;
								assign node32 = (inp[8]) ? node46 : node33;
									assign node33 = (inp[2]) ? node39 : node34;
										assign node34 = (inp[3]) ? 3'b100 : node35;
											assign node35 = (inp[4]) ? 3'b100 : 3'b110;
										assign node39 = (inp[3]) ? 3'b000 : node40;
											assign node40 = (inp[4]) ? node42 : 3'b100;
												assign node42 = (inp[5]) ? 3'b000 : 3'b100;
									assign node46 = (inp[3]) ? 3'b010 : node47;
										assign node47 = (inp[4]) ? 3'b010 : node48;
											assign node48 = (inp[2]) ? 3'b010 : 3'b110;
							assign node53 = (inp[8]) ? node63 : node54;
								assign node54 = (inp[11]) ? 3'b000 : node55;
									assign node55 = (inp[2]) ? node57 : 3'b100;
										assign node57 = (inp[3]) ? 3'b000 : node58;
											assign node58 = (inp[4]) ? 3'b000 : 3'b100;
								assign node63 = (inp[11]) ? node73 : node64;
									assign node64 = (inp[2]) ? node66 : 3'b010;
										assign node66 = (inp[3]) ? 3'b100 : node67;
											assign node67 = (inp[4]) ? node69 : 3'b010;
												assign node69 = (inp[5]) ? 3'b100 : 3'b010;
									assign node73 = (inp[2]) ? node75 : 3'b100;
										assign node75 = (inp[3]) ? 3'b000 : 3'b100;
						assign node78 = (inp[8]) ? node80 : 3'b000;
							assign node80 = (inp[1]) ? 3'b000 : node81;
								assign node81 = (inp[11]) ? node93 : node82;
									assign node82 = (inp[2]) ? node88 : node83;
										assign node83 = (inp[3]) ? 3'b100 : node84;
											assign node84 = (inp[4]) ? 3'b100 : 3'b000;
										assign node88 = (inp[4]) ? node90 : 3'b100;
											assign node90 = (inp[3]) ? 3'b000 : 3'b100;
									assign node93 = (inp[2]) ? 3'b000 : node94;
										assign node94 = (inp[3]) ? 3'b000 : node95;
											assign node95 = (inp[4]) ? node97 : 3'b100;
												assign node97 = (inp[5]) ? 3'b000 : 3'b100;
					assign node103 = (inp[10]) ? node193 : node104;
						assign node104 = (inp[1]) ? node150 : node105;
							assign node105 = (inp[8]) ? node131 : node106;
								assign node106 = (inp[11]) ? node118 : node107;
									assign node107 = (inp[2]) ? node113 : node108;
										assign node108 = (inp[3]) ? 3'b001 : node109;
											assign node109 = (inp[4]) ? 3'b001 : 3'b101;
										assign node113 = (inp[4]) ? node115 : 3'b001;
											assign node115 = (inp[3]) ? 3'b110 : 3'b001;
									assign node118 = (inp[2]) ? node126 : node119;
										assign node119 = (inp[3]) ? 3'b110 : node120;
											assign node120 = (inp[4]) ? node122 : 3'b001;
												assign node122 = (inp[5]) ? 3'b110 : 3'b001;
										assign node126 = (inp[3]) ? node128 : 3'b110;
											assign node128 = (inp[4]) ? 3'b010 : 3'b110;
								assign node131 = (inp[11]) ? node139 : node132;
									assign node132 = (inp[2]) ? node134 : 3'b101;
										assign node134 = (inp[5]) ? node136 : 3'b101;
											assign node136 = (inp[3]) ? 3'b001 : 3'b101;
									assign node139 = (inp[3]) ? node143 : node140;
										assign node140 = (inp[2]) ? 3'b001 : 3'b101;
										assign node143 = (inp[2]) ? node145 : 3'b001;
											assign node145 = (inp[4]) ? node147 : 3'b001;
												assign node147 = (inp[5]) ? 3'b110 : 3'b001;
							assign node150 = (inp[8]) ? node166 : node151;
								assign node151 = (inp[11]) ? node161 : node152;
									assign node152 = (inp[2]) ? node154 : 3'b110;
										assign node154 = (inp[3]) ? 3'b010 : node155;
											assign node155 = (inp[4]) ? node157 : 3'b110;
												assign node157 = (inp[5]) ? 3'b010 : 3'b110;
									assign node161 = (inp[3]) ? node163 : 3'b010;
										assign node163 = (inp[2]) ? 3'b100 : 3'b010;
								assign node166 = (inp[11]) ? node178 : node167;
									assign node167 = (inp[2]) ? node175 : node168;
										assign node168 = (inp[3]) ? 3'b001 : node169;
											assign node169 = (inp[4]) ? 3'b001 : node170;
												assign node170 = (inp[5]) ? 3'b001 : 3'b101;
										assign node175 = (inp[3]) ? 3'b110 : 3'b001;
									assign node178 = (inp[3]) ? node186 : node179;
										assign node179 = (inp[4]) ? 3'b110 : node180;
											assign node180 = (inp[2]) ? 3'b110 : node181;
												assign node181 = (inp[5]) ? 3'b110 : 3'b001;
										assign node186 = (inp[2]) ? node188 : 3'b110;
											assign node188 = (inp[4]) ? 3'b010 : node189;
												assign node189 = (inp[5]) ? 3'b010 : 3'b110;
						assign node193 = (inp[1]) ? node231 : node194;
							assign node194 = (inp[8]) ? node220 : node195;
								assign node195 = (inp[11]) ? node211 : node196;
									assign node196 = (inp[2]) ? node204 : node197;
										assign node197 = (inp[3]) ? 3'b010 : node198;
											assign node198 = (inp[5]) ? node200 : 3'b110;
												assign node200 = (inp[4]) ? 3'b010 : 3'b110;
										assign node204 = (inp[5]) ? node206 : 3'b010;
											assign node206 = (inp[4]) ? node208 : 3'b010;
												assign node208 = (inp[3]) ? 3'b100 : 3'b010;
									assign node211 = (inp[3]) ? node215 : node212;
										assign node212 = (inp[2]) ? 3'b100 : 3'b010;
										assign node215 = (inp[2]) ? node217 : 3'b100;
											assign node217 = (inp[5]) ? 3'b000 : 3'b100;
								assign node220 = (inp[11]) ? node226 : node221;
									assign node221 = (inp[3]) ? 3'b110 : node222;
										assign node222 = (inp[2]) ? 3'b110 : 3'b001;
									assign node226 = (inp[3]) ? 3'b010 : node227;
										assign node227 = (inp[2]) ? 3'b010 : 3'b110;
							assign node231 = (inp[8]) ? node239 : node232;
								assign node232 = (inp[11]) ? 3'b000 : node233;
									assign node233 = (inp[3]) ? node235 : 3'b100;
										assign node235 = (inp[2]) ? 3'b000 : 3'b100;
								assign node239 = (inp[11]) ? node249 : node240;
									assign node240 = (inp[2]) ? node246 : node241;
										assign node241 = (inp[4]) ? 3'b010 : node242;
											assign node242 = (inp[3]) ? 3'b010 : 3'b110;
										assign node246 = (inp[3]) ? 3'b100 : 3'b010;
									assign node249 = (inp[3]) ? node255 : node250;
										assign node250 = (inp[2]) ? 3'b100 : node251;
											assign node251 = (inp[4]) ? 3'b100 : 3'b010;
										assign node255 = (inp[2]) ? node257 : 3'b100;
											assign node257 = (inp[4]) ? 3'b000 : node258;
												assign node258 = (inp[5]) ? 3'b000 : 3'b100;
				assign node262 = (inp[7]) ? node278 : node263;
					assign node263 = (inp[10]) ? 3'b000 : node264;
						assign node264 = (inp[8]) ? node266 : 3'b000;
							assign node266 = (inp[1]) ? 3'b000 : node267;
								assign node267 = (inp[2]) ? 3'b000 : node268;
									assign node268 = (inp[11]) ? 3'b000 : node269;
										assign node269 = (inp[4]) ? node271 : 3'b100;
											assign node271 = (inp[3]) ? 3'b000 : 3'b100;
					assign node278 = (inp[10]) ? node338 : node279;
						assign node279 = (inp[1]) ? node313 : node280;
							assign node280 = (inp[8]) ? node298 : node281;
								assign node281 = (inp[11]) ? node289 : node282;
									assign node282 = (inp[2]) ? 3'b100 : node283;
										assign node283 = (inp[5]) ? node285 : 3'b010;
											assign node285 = (inp[3]) ? 3'b100 : 3'b010;
									assign node289 = (inp[2]) ? node291 : 3'b100;
										assign node291 = (inp[5]) ? 3'b000 : node292;
											assign node292 = (inp[4]) ? 3'b000 : node293;
												assign node293 = (inp[3]) ? 3'b000 : 3'b100;
								assign node298 = (inp[11]) ? node306 : node299;
									assign node299 = (inp[2]) ? node301 : 3'b110;
										assign node301 = (inp[3]) ? 3'b010 : node302;
											assign node302 = (inp[4]) ? 3'b010 : 3'b110;
									assign node306 = (inp[2]) ? node308 : 3'b010;
										assign node308 = (inp[4]) ? 3'b100 : node309;
											assign node309 = (inp[3]) ? 3'b100 : 3'b010;
							assign node313 = (inp[8]) ? node321 : node314;
								assign node314 = (inp[2]) ? 3'b000 : node315;
									assign node315 = (inp[3]) ? 3'b000 : node316;
										assign node316 = (inp[11]) ? 3'b000 : 3'b100;
								assign node321 = (inp[11]) ? node331 : node322;
									assign node322 = (inp[2]) ? 3'b100 : node323;
										assign node323 = (inp[3]) ? node325 : 3'b010;
											assign node325 = (inp[5]) ? 3'b100 : node326;
												assign node326 = (inp[4]) ? 3'b100 : 3'b010;
									assign node331 = (inp[2]) ? 3'b000 : node332;
										assign node332 = (inp[4]) ? node334 : 3'b100;
											assign node334 = (inp[3]) ? 3'b000 : 3'b100;
						assign node338 = (inp[11]) ? 3'b000 : node339;
							assign node339 = (inp[8]) ? node341 : 3'b000;
								assign node341 = (inp[1]) ? 3'b000 : node342;
									assign node342 = (inp[2]) ? node344 : 3'b100;
										assign node344 = (inp[3]) ? 3'b000 : node345;
											assign node345 = (inp[4]) ? 3'b000 : 3'b100;
			assign node351 = (inp[0]) ? 3'b000 : node352;
				assign node352 = (inp[7]) ? node354 : 3'b000;
					assign node354 = (inp[10]) ? 3'b000 : node355;
						assign node355 = (inp[1]) ? node381 : node356;
							assign node356 = (inp[8]) ? node364 : node357;
								assign node357 = (inp[11]) ? 3'b000 : node358;
									assign node358 = (inp[2]) ? 3'b000 : node359;
										assign node359 = (inp[3]) ? 3'b000 : 3'b100;
								assign node364 = (inp[11]) ? node374 : node365;
									assign node365 = (inp[2]) ? 3'b100 : node366;
										assign node366 = (inp[3]) ? node368 : 3'b010;
											assign node368 = (inp[4]) ? 3'b100 : node369;
												assign node369 = (inp[5]) ? 3'b100 : 3'b010;
									assign node374 = (inp[2]) ? 3'b000 : node375;
										assign node375 = (inp[3]) ? node377 : 3'b100;
											assign node377 = (inp[4]) ? 3'b000 : 3'b100;
							assign node381 = (inp[3]) ? 3'b000 : node382;
								assign node382 = (inp[11]) ? 3'b000 : node383;
									assign node383 = (inp[8]) ? node385 : 3'b000;
										assign node385 = (inp[2]) ? 3'b000 : node386;
											assign node386 = (inp[4]) ? 3'b000 : 3'b100;
		assign node394 = (inp[9]) ? node952 : node395;
			assign node395 = (inp[0]) ? node647 : node396;
				assign node396 = (inp[7]) ? node564 : node397;
					assign node397 = (inp[10]) ? node479 : node398;
						assign node398 = (inp[1]) ? node426 : node399;
							assign node399 = (inp[8]) ? node415 : node400;
								assign node400 = (inp[11]) ? node406 : node401;
									assign node401 = (inp[2]) ? 3'b011 : node402;
										assign node402 = (inp[3]) ? 3'b011 : 3'b111;
									assign node406 = (inp[2]) ? 3'b101 : node407;
										assign node407 = (inp[3]) ? node409 : 3'b011;
											assign node409 = (inp[4]) ? 3'b101 : node410;
												assign node410 = (inp[5]) ? 3'b101 : 3'b011;
								assign node415 = (inp[11]) ? node417 : 3'b111;
									assign node417 = (inp[2]) ? 3'b011 : node418;
										assign node418 = (inp[3]) ? node420 : 3'b111;
											assign node420 = (inp[5]) ? 3'b011 : node421;
												assign node421 = (inp[4]) ? 3'b011 : 3'b111;
							assign node426 = (inp[8]) ? node454 : node427;
								assign node427 = (inp[11]) ? node443 : node428;
									assign node428 = (inp[4]) ? node438 : node429;
										assign node429 = (inp[3]) ? node433 : node430;
											assign node430 = (inp[5]) ? 3'b101 : 3'b011;
											assign node433 = (inp[5]) ? node435 : 3'b101;
												assign node435 = (inp[2]) ? 3'b001 : 3'b101;
										assign node438 = (inp[3]) ? node440 : 3'b101;
											assign node440 = (inp[2]) ? 3'b001 : 3'b101;
									assign node443 = (inp[4]) ? node449 : node444;
										assign node444 = (inp[3]) ? 3'b001 : node445;
											assign node445 = (inp[2]) ? 3'b001 : 3'b101;
										assign node449 = (inp[2]) ? node451 : 3'b001;
											assign node451 = (inp[3]) ? 3'b110 : 3'b001;
								assign node454 = (inp[11]) ? node466 : node455;
									assign node455 = (inp[4]) ? node461 : node456;
										assign node456 = (inp[2]) ? 3'b011 : node457;
											assign node457 = (inp[3]) ? 3'b011 : 3'b111;
										assign node461 = (inp[2]) ? node463 : 3'b011;
											assign node463 = (inp[3]) ? 3'b101 : 3'b011;
									assign node466 = (inp[3]) ? node474 : node467;
										assign node467 = (inp[2]) ? 3'b101 : node468;
											assign node468 = (inp[4]) ? node470 : 3'b011;
												assign node470 = (inp[5]) ? 3'b101 : 3'b011;
										assign node474 = (inp[2]) ? node476 : 3'b101;
											assign node476 = (inp[4]) ? 3'b001 : 3'b101;
						assign node479 = (inp[1]) ? node513 : node480;
							assign node480 = (inp[11]) ? node496 : node481;
								assign node481 = (inp[8]) ? node489 : node482;
									assign node482 = (inp[2]) ? 3'b001 : node483;
										assign node483 = (inp[3]) ? node485 : 3'b101;
											assign node485 = (inp[5]) ? 3'b001 : 3'b101;
									assign node489 = (inp[2]) ? 3'b101 : node490;
										assign node490 = (inp[4]) ? node492 : 3'b011;
											assign node492 = (inp[3]) ? 3'b101 : 3'b011;
								assign node496 = (inp[8]) ? node506 : node497;
									assign node497 = (inp[2]) ? 3'b110 : node498;
										assign node498 = (inp[3]) ? node500 : 3'b001;
											assign node500 = (inp[4]) ? 3'b110 : node501;
												assign node501 = (inp[5]) ? 3'b110 : 3'b001;
									assign node506 = (inp[2]) ? 3'b001 : node507;
										assign node507 = (inp[4]) ? node509 : 3'b101;
											assign node509 = (inp[3]) ? 3'b001 : 3'b101;
							assign node513 = (inp[8]) ? node539 : node514;
								assign node514 = (inp[11]) ? node526 : node515;
									assign node515 = (inp[4]) ? node521 : node516;
										assign node516 = (inp[2]) ? 3'b110 : node517;
											assign node517 = (inp[3]) ? 3'b110 : 3'b001;
										assign node521 = (inp[2]) ? node523 : 3'b110;
											assign node523 = (inp[3]) ? 3'b010 : 3'b110;
									assign node526 = (inp[3]) ? node534 : node527;
										assign node527 = (inp[2]) ? 3'b010 : node528;
											assign node528 = (inp[4]) ? node530 : 3'b110;
												assign node530 = (inp[5]) ? 3'b010 : 3'b110;
										assign node534 = (inp[2]) ? node536 : 3'b010;
											assign node536 = (inp[4]) ? 3'b100 : 3'b010;
								assign node539 = (inp[11]) ? node555 : node540;
									assign node540 = (inp[3]) ? node548 : node541;
										assign node541 = (inp[2]) ? 3'b001 : node542;
											assign node542 = (inp[5]) ? node544 : 3'b101;
												assign node544 = (inp[4]) ? 3'b001 : 3'b101;
										assign node548 = (inp[4]) ? node550 : 3'b001;
											assign node550 = (inp[2]) ? node552 : 3'b001;
												assign node552 = (inp[5]) ? 3'b110 : 3'b001;
									assign node555 = (inp[3]) ? node559 : node556;
										assign node556 = (inp[2]) ? 3'b110 : 3'b001;
										assign node559 = (inp[5]) ? node561 : 3'b110;
											assign node561 = (inp[4]) ? 3'b010 : 3'b110;
					assign node564 = (inp[10]) ? node590 : node565;
						assign node565 = (inp[8]) ? 3'b111 : node566;
							assign node566 = (inp[1]) ? node568 : 3'b111;
								assign node568 = (inp[11]) ? node578 : node569;
									assign node569 = (inp[5]) ? node571 : 3'b111;
										assign node571 = (inp[3]) ? node573 : 3'b111;
											assign node573 = (inp[2]) ? node575 : 3'b111;
												assign node575 = (inp[4]) ? 3'b011 : 3'b111;
									assign node578 = (inp[2]) ? node582 : node579;
										assign node579 = (inp[3]) ? 3'b011 : 3'b111;
										assign node582 = (inp[4]) ? node584 : 3'b011;
											assign node584 = (inp[3]) ? node586 : 3'b011;
												assign node586 = (inp[5]) ? 3'b101 : 3'b011;
						assign node590 = (inp[1]) ? node620 : node591;
							assign node591 = (inp[8]) ? node609 : node592;
								assign node592 = (inp[11]) ? node596 : node593;
									assign node593 = (inp[2]) ? 3'b011 : 3'b111;
									assign node596 = (inp[2]) ? node602 : node597;
										assign node597 = (inp[5]) ? node599 : 3'b011;
											assign node599 = (inp[3]) ? 3'b101 : 3'b011;
										assign node602 = (inp[3]) ? 3'b101 : node603;
											assign node603 = (inp[5]) ? 3'b101 : node604;
												assign node604 = (inp[4]) ? 3'b101 : 3'b011;
								assign node609 = (inp[11]) ? node611 : 3'b111;
									assign node611 = (inp[2]) ? node613 : 3'b111;
										assign node613 = (inp[3]) ? 3'b011 : node614;
											assign node614 = (inp[4]) ? node616 : 3'b111;
												assign node616 = (inp[5]) ? 3'b011 : 3'b111;
							assign node620 = (inp[8]) ? node632 : node621;
								assign node621 = (inp[11]) ? node627 : node622;
									assign node622 = (inp[2]) ? 3'b101 : node623;
										assign node623 = (inp[3]) ? 3'b101 : 3'b011;
									assign node627 = (inp[2]) ? 3'b001 : node628;
										assign node628 = (inp[3]) ? 3'b001 : 3'b101;
								assign node632 = (inp[11]) ? node638 : node633;
									assign node633 = (inp[2]) ? 3'b011 : node634;
										assign node634 = (inp[3]) ? 3'b011 : 3'b111;
									assign node638 = (inp[2]) ? 3'b101 : node639;
										assign node639 = (inp[3]) ? node641 : 3'b011;
											assign node641 = (inp[5]) ? 3'b101 : node642;
												assign node642 = (inp[4]) ? 3'b101 : 3'b011;
				assign node647 = (inp[7]) ? node789 : node648;
					assign node648 = (inp[10]) ? node716 : node649;
						assign node649 = (inp[1]) ? node677 : node650;
							assign node650 = (inp[8]) ? node666 : node651;
								assign node651 = (inp[11]) ? node659 : node652;
									assign node652 = (inp[2]) ? node654 : 3'b001;
										assign node654 = (inp[3]) ? 3'b110 : node655;
											assign node655 = (inp[4]) ? 3'b110 : 3'b001;
									assign node659 = (inp[2]) ? node661 : 3'b110;
										assign node661 = (inp[3]) ? 3'b010 : node662;
											assign node662 = (inp[4]) ? 3'b010 : 3'b110;
								assign node666 = (inp[11]) ? node672 : node667;
									assign node667 = (inp[2]) ? node669 : 3'b101;
										assign node669 = (inp[3]) ? 3'b001 : 3'b101;
									assign node672 = (inp[2]) ? node674 : 3'b001;
										assign node674 = (inp[3]) ? 3'b110 : 3'b001;
							assign node677 = (inp[11]) ? node693 : node678;
								assign node678 = (inp[8]) ? node686 : node679;
									assign node679 = (inp[2]) ? 3'b010 : node680;
										assign node680 = (inp[3]) ? node682 : 3'b110;
											assign node682 = (inp[4]) ? 3'b010 : 3'b110;
									assign node686 = (inp[2]) ? 3'b110 : node687;
										assign node687 = (inp[5]) ? node689 : 3'b001;
											assign node689 = (inp[4]) ? 3'b110 : 3'b001;
								assign node693 = (inp[8]) ? node703 : node694;
									assign node694 = (inp[2]) ? 3'b100 : node695;
										assign node695 = (inp[3]) ? node697 : 3'b010;
											assign node697 = (inp[5]) ? node699 : 3'b010;
												assign node699 = (inp[4]) ? 3'b100 : 3'b010;
									assign node703 = (inp[2]) ? node709 : node704;
										assign node704 = (inp[4]) ? node706 : 3'b110;
											assign node706 = (inp[5]) ? 3'b010 : 3'b110;
										assign node709 = (inp[5]) ? 3'b010 : node710;
											assign node710 = (inp[4]) ? 3'b010 : node711;
												assign node711 = (inp[3]) ? 3'b010 : 3'b110;
						assign node716 = (inp[1]) ? node754 : node717;
							assign node717 = (inp[8]) ? node733 : node718;
								assign node718 = (inp[11]) ? node728 : node719;
									assign node719 = (inp[2]) ? node721 : 3'b010;
										assign node721 = (inp[3]) ? 3'b100 : node722;
											assign node722 = (inp[4]) ? node724 : 3'b010;
												assign node724 = (inp[5]) ? 3'b100 : 3'b010;
									assign node728 = (inp[2]) ? node730 : 3'b100;
										assign node730 = (inp[3]) ? 3'b000 : 3'b100;
								assign node733 = (inp[11]) ? node739 : node734;
									assign node734 = (inp[3]) ? node736 : 3'b110;
										assign node736 = (inp[2]) ? 3'b010 : 3'b110;
									assign node739 = (inp[3]) ? node747 : node740;
										assign node740 = (inp[4]) ? 3'b010 : node741;
											assign node741 = (inp[5]) ? 3'b010 : node742;
												assign node742 = (inp[2]) ? 3'b010 : 3'b110;
										assign node747 = (inp[2]) ? node749 : 3'b010;
											assign node749 = (inp[5]) ? 3'b100 : node750;
												assign node750 = (inp[4]) ? 3'b100 : 3'b010;
							assign node754 = (inp[8]) ? node772 : node755;
								assign node755 = (inp[11]) ? 3'b000 : node756;
									assign node756 = (inp[2]) ? node764 : node757;
										assign node757 = (inp[3]) ? node759 : 3'b100;
											assign node759 = (inp[4]) ? node761 : 3'b100;
												assign node761 = (inp[5]) ? 3'b000 : 3'b100;
										assign node764 = (inp[3]) ? 3'b000 : node765;
											assign node765 = (inp[5]) ? 3'b000 : node766;
												assign node766 = (inp[4]) ? 3'b000 : 3'b100;
								assign node772 = (inp[11]) ? node780 : node773;
									assign node773 = (inp[2]) ? node775 : 3'b010;
										assign node775 = (inp[5]) ? 3'b100 : node776;
											assign node776 = (inp[4]) ? 3'b100 : 3'b010;
									assign node780 = (inp[2]) ? node782 : 3'b100;
										assign node782 = (inp[3]) ? 3'b000 : node783;
											assign node783 = (inp[5]) ? node785 : 3'b100;
												assign node785 = (inp[4]) ? 3'b000 : 3'b100;
					assign node789 = (inp[10]) ? node871 : node790;
						assign node790 = (inp[1]) ? node840 : node791;
							assign node791 = (inp[8]) ? node819 : node792;
								assign node792 = (inp[11]) ? node804 : node793;
									assign node793 = (inp[2]) ? node801 : node794;
										assign node794 = (inp[4]) ? 3'b011 : node795;
											assign node795 = (inp[5]) ? 3'b011 : node796;
												assign node796 = (inp[3]) ? 3'b011 : 3'b111;
										assign node801 = (inp[3]) ? 3'b101 : 3'b011;
									assign node804 = (inp[2]) ? node812 : node805;
										assign node805 = (inp[3]) ? 3'b101 : node806;
											assign node806 = (inp[5]) ? 3'b101 : node807;
												assign node807 = (inp[4]) ? 3'b101 : 3'b011;
										assign node812 = (inp[3]) ? node814 : 3'b101;
											assign node814 = (inp[5]) ? 3'b001 : node815;
												assign node815 = (inp[4]) ? 3'b001 : 3'b101;
								assign node819 = (inp[11]) ? node829 : node820;
									assign node820 = (inp[3]) ? node822 : 3'b111;
										assign node822 = (inp[2]) ? node824 : 3'b111;
											assign node824 = (inp[5]) ? 3'b011 : node825;
												assign node825 = (inp[4]) ? 3'b011 : 3'b111;
									assign node829 = (inp[3]) ? node835 : node830;
										assign node830 = (inp[4]) ? 3'b011 : node831;
											assign node831 = (inp[2]) ? 3'b011 : 3'b111;
										assign node835 = (inp[4]) ? node837 : 3'b011;
											assign node837 = (inp[2]) ? 3'b101 : 3'b011;
							assign node840 = (inp[8]) ? node856 : node841;
								assign node841 = (inp[11]) ? node849 : node842;
									assign node842 = (inp[2]) ? node844 : 3'b101;
										assign node844 = (inp[3]) ? 3'b001 : node845;
											assign node845 = (inp[4]) ? 3'b001 : 3'b101;
									assign node849 = (inp[2]) ? node851 : 3'b001;
										assign node851 = (inp[4]) ? 3'b110 : node852;
											assign node852 = (inp[3]) ? 3'b110 : 3'b001;
								assign node856 = (inp[11]) ? node864 : node857;
									assign node857 = (inp[2]) ? node859 : 3'b011;
										assign node859 = (inp[4]) ? 3'b101 : node860;
											assign node860 = (inp[3]) ? 3'b101 : 3'b011;
									assign node864 = (inp[2]) ? node866 : 3'b101;
										assign node866 = (inp[5]) ? 3'b001 : node867;
											assign node867 = (inp[3]) ? 3'b001 : 3'b101;
						assign node871 = (inp[1]) ? node921 : node872;
							assign node872 = (inp[11]) ? node900 : node873;
								assign node873 = (inp[8]) ? node889 : node874;
									assign node874 = (inp[3]) ? node882 : node875;
										assign node875 = (inp[2]) ? 3'b001 : node876;
											assign node876 = (inp[4]) ? 3'b001 : node877;
												assign node877 = (inp[5]) ? 3'b001 : 3'b101;
										assign node882 = (inp[2]) ? node884 : 3'b001;
											assign node884 = (inp[4]) ? 3'b110 : node885;
												assign node885 = (inp[5]) ? 3'b110 : 3'b001;
									assign node889 = (inp[2]) ? node895 : node890;
										assign node890 = (inp[3]) ? 3'b101 : node891;
											assign node891 = (inp[4]) ? 3'b101 : 3'b011;
										assign node895 = (inp[3]) ? node897 : 3'b101;
											assign node897 = (inp[4]) ? 3'b001 : 3'b101;
								assign node900 = (inp[8]) ? node908 : node901;
									assign node901 = (inp[2]) ? node903 : 3'b110;
										assign node903 = (inp[3]) ? node905 : 3'b110;
											assign node905 = (inp[4]) ? 3'b010 : 3'b110;
									assign node908 = (inp[2]) ? node916 : node909;
										assign node909 = (inp[3]) ? 3'b001 : node910;
											assign node910 = (inp[5]) ? node912 : 3'b101;
												assign node912 = (inp[4]) ? 3'b001 : 3'b101;
										assign node916 = (inp[4]) ? node918 : 3'b001;
											assign node918 = (inp[3]) ? 3'b110 : 3'b011;
							assign node921 = (inp[11]) ? node937 : node922;
								assign node922 = (inp[8]) ? node930 : node923;
									assign node923 = (inp[2]) ? node925 : 3'b110;
										assign node925 = (inp[3]) ? 3'b010 : node926;
											assign node926 = (inp[4]) ? 3'b010 : 3'b110;
									assign node930 = (inp[2]) ? node932 : 3'b001;
										assign node932 = (inp[3]) ? 3'b110 : node933;
											assign node933 = (inp[4]) ? 3'b110 : 3'b001;
								assign node937 = (inp[8]) ? node947 : node938;
									assign node938 = (inp[2]) ? node940 : 3'b010;
										assign node940 = (inp[3]) ? 3'b100 : node941;
											assign node941 = (inp[4]) ? node943 : 3'b010;
												assign node943 = (inp[5]) ? 3'b100 : 3'b010;
									assign node947 = (inp[2]) ? node949 : 3'b110;
										assign node949 = (inp[3]) ? 3'b010 : 3'b110;
			assign node952 = (inp[0]) ? node1210 : node953;
				assign node953 = (inp[7]) ? node1073 : node954;
					assign node954 = (inp[10]) ? node1030 : node955;
						assign node955 = (inp[1]) ? node995 : node956;
							assign node956 = (inp[11]) ? node974 : node957;
								assign node957 = (inp[2]) ? node971 : node958;
									assign node958 = (inp[8]) ? node964 : node959;
										assign node959 = (inp[4]) ? node961 : 3'b110;
											assign node961 = (inp[3]) ? 3'b010 : 3'b110;
										assign node964 = (inp[3]) ? node966 : 3'b001;
											assign node966 = (inp[5]) ? node968 : 3'b001;
												assign node968 = (inp[4]) ? 3'b110 : 3'b001;
									assign node971 = (inp[8]) ? 3'b110 : 3'b010;
								assign node974 = (inp[8]) ? node982 : node975;
									assign node975 = (inp[2]) ? 3'b100 : node976;
										assign node976 = (inp[4]) ? node978 : 3'b010;
											assign node978 = (inp[3]) ? 3'b100 : 3'b010;
									assign node982 = (inp[2]) ? node990 : node983;
										assign node983 = (inp[4]) ? node985 : 3'b110;
											assign node985 = (inp[3]) ? node987 : 3'b110;
												assign node987 = (inp[5]) ? 3'b010 : 3'b110;
										assign node990 = (inp[3]) ? 3'b010 : node991;
											assign node991 = (inp[5]) ? 3'b010 : 3'b110;
							assign node995 = (inp[8]) ? node1019 : node996;
								assign node996 = (inp[11]) ? node1012 : node997;
									assign node997 = (inp[3]) ? node1005 : node998;
										assign node998 = (inp[2]) ? 3'b100 : node999;
											assign node999 = (inp[4]) ? node1001 : 3'b010;
												assign node1001 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1005 = (inp[4]) ? node1007 : 3'b100;
											assign node1007 = (inp[2]) ? node1009 : 3'b100;
												assign node1009 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1012 = (inp[3]) ? 3'b000 : node1013;
										assign node1013 = (inp[2]) ? 3'b000 : node1014;
											assign node1014 = (inp[4]) ? 3'b000 : 3'b100;
								assign node1019 = (inp[11]) ? node1025 : node1020;
									assign node1020 = (inp[2]) ? 3'b010 : node1021;
										assign node1021 = (inp[3]) ? 3'b010 : 3'b110;
									assign node1025 = (inp[2]) ? 3'b100 : node1026;
										assign node1026 = (inp[3]) ? 3'b100 : 3'b010;
						assign node1030 = (inp[1]) ? node1064 : node1031;
							assign node1031 = (inp[8]) ? node1041 : node1032;
								assign node1032 = (inp[11]) ? 3'b000 : node1033;
									assign node1033 = (inp[2]) ? 3'b000 : node1034;
										assign node1034 = (inp[4]) ? node1036 : 3'b100;
											assign node1036 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1041 = (inp[11]) ? node1055 : node1042;
									assign node1042 = (inp[2]) ? node1050 : node1043;
										assign node1043 = (inp[5]) ? node1045 : 3'b010;
											assign node1045 = (inp[3]) ? node1047 : 3'b010;
												assign node1047 = (inp[4]) ? 3'b100 : 3'b010;
										assign node1050 = (inp[4]) ? 3'b100 : node1051;
											assign node1051 = (inp[3]) ? 3'b100 : 3'b010;
									assign node1055 = (inp[2]) ? node1057 : 3'b100;
										assign node1057 = (inp[5]) ? 3'b000 : node1058;
											assign node1058 = (inp[3]) ? 3'b000 : node1059;
												assign node1059 = (inp[4]) ? 3'b000 : 3'b100;
							assign node1064 = (inp[8]) ? node1066 : 3'b000;
								assign node1066 = (inp[11]) ? 3'b000 : node1067;
									assign node1067 = (inp[2]) ? 3'b000 : node1068;
										assign node1068 = (inp[3]) ? 3'b000 : 3'b100;
					assign node1073 = (inp[10]) ? node1145 : node1074;
						assign node1074 = (inp[1]) ? node1112 : node1075;
							assign node1075 = (inp[2]) ? node1089 : node1076;
								assign node1076 = (inp[8]) ? node1086 : node1077;
									assign node1077 = (inp[11]) ? 3'b001 : node1078;
										assign node1078 = (inp[3]) ? node1080 : 3'b101;
											assign node1080 = (inp[5]) ? node1082 : 3'b101;
												assign node1082 = (inp[4]) ? 3'b001 : 3'b101;
									assign node1086 = (inp[11]) ? 3'b101 : 3'b011;
								assign node1089 = (inp[8]) ? node1101 : node1090;
									assign node1090 = (inp[11]) ? node1096 : node1091;
										assign node1091 = (inp[4]) ? 3'b001 : node1092;
											assign node1092 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1096 = (inp[5]) ? 3'b110 : node1097;
											assign node1097 = (inp[3]) ? 3'b110 : 3'b001;
									assign node1101 = (inp[11]) ? node1107 : node1102;
										assign node1102 = (inp[3]) ? 3'b101 : node1103;
											assign node1103 = (inp[4]) ? 3'b101 : 3'b011;
										assign node1107 = (inp[3]) ? 3'b001 : node1108;
											assign node1108 = (inp[4]) ? 3'b001 : 3'b101;
							assign node1112 = (inp[11]) ? node1128 : node1113;
								assign node1113 = (inp[8]) ? node1121 : node1114;
									assign node1114 = (inp[2]) ? 3'b110 : node1115;
										assign node1115 = (inp[3]) ? node1117 : 3'b001;
											assign node1117 = (inp[4]) ? 3'b110 : 3'b001;
									assign node1121 = (inp[2]) ? 3'b001 : node1122;
										assign node1122 = (inp[3]) ? node1124 : 3'b101;
											assign node1124 = (inp[4]) ? 3'b001 : 3'b101;
								assign node1128 = (inp[8]) ? node1138 : node1129;
									assign node1129 = (inp[2]) ? 3'b010 : node1130;
										assign node1130 = (inp[3]) ? node1132 : 3'b110;
											assign node1132 = (inp[5]) ? 3'b010 : node1133;
												assign node1133 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1138 = (inp[2]) ? 3'b110 : node1139;
										assign node1139 = (inp[3]) ? node1141 : 3'b001;
											assign node1141 = (inp[4]) ? 3'b110 : 3'b001;
						assign node1145 = (inp[1]) ? node1177 : node1146;
							assign node1146 = (inp[11]) ? node1162 : node1147;
								assign node1147 = (inp[8]) ? node1155 : node1148;
									assign node1148 = (inp[2]) ? node1150 : 3'b110;
										assign node1150 = (inp[4]) ? 3'b010 : node1151;
											assign node1151 = (inp[3]) ? 3'b010 : 3'b110;
									assign node1155 = (inp[2]) ? node1157 : 3'b001;
										assign node1157 = (inp[3]) ? 3'b110 : node1158;
											assign node1158 = (inp[5]) ? 3'b110 : 3'b001;
								assign node1162 = (inp[8]) ? node1172 : node1163;
									assign node1163 = (inp[2]) ? node1165 : 3'b010;
										assign node1165 = (inp[3]) ? 3'b100 : node1166;
											assign node1166 = (inp[4]) ? node1168 : 3'b010;
												assign node1168 = (inp[5]) ? 3'b100 : 3'b010;
									assign node1172 = (inp[2]) ? node1174 : 3'b110;
										assign node1174 = (inp[3]) ? 3'b010 : 3'b110;
							assign node1177 = (inp[8]) ? node1193 : node1178;
								assign node1178 = (inp[11]) ? node1186 : node1179;
									assign node1179 = (inp[2]) ? 3'b100 : node1180;
										assign node1180 = (inp[3]) ? node1182 : 3'b010;
											assign node1182 = (inp[4]) ? 3'b100 : 3'b010;
									assign node1186 = (inp[2]) ? 3'b000 : node1187;
										assign node1187 = (inp[3]) ? node1189 : 3'b100;
											assign node1189 = (inp[4]) ? 3'b000 : 3'b100;
								assign node1193 = (inp[11]) ? node1201 : node1194;
									assign node1194 = (inp[2]) ? 3'b010 : node1195;
										assign node1195 = (inp[3]) ? node1197 : 3'b110;
											assign node1197 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1201 = (inp[2]) ? 3'b100 : node1202;
										assign node1202 = (inp[4]) ? node1204 : 3'b010;
											assign node1204 = (inp[5]) ? node1206 : 3'b010;
												assign node1206 = (inp[3]) ? 3'b100 : 3'b010;
				assign node1210 = (inp[7]) ? node1240 : node1211;
					assign node1211 = (inp[1]) ? 3'b000 : node1212;
						assign node1212 = (inp[8]) ? node1214 : 3'b000;
							assign node1214 = (inp[10]) ? 3'b000 : node1215;
								assign node1215 = (inp[11]) ? node1231 : node1216;
									assign node1216 = (inp[3]) ? node1224 : node1217;
										assign node1217 = (inp[4]) ? 3'b100 : node1218;
											assign node1218 = (inp[2]) ? 3'b100 : node1219;
												assign node1219 = (inp[5]) ? 3'b100 : 3'b010;
										assign node1224 = (inp[2]) ? node1226 : 3'b100;
											assign node1226 = (inp[4]) ? 3'b000 : node1227;
												assign node1227 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1231 = (inp[4]) ? 3'b000 : node1232;
										assign node1232 = (inp[3]) ? 3'b000 : node1233;
											assign node1233 = (inp[2]) ? 3'b000 : 3'b100;
					assign node1240 = (inp[10]) ? node1328 : node1241;
						assign node1241 = (inp[1]) ? node1299 : node1242;
							assign node1242 = (inp[11]) ? node1270 : node1243;
								assign node1243 = (inp[8]) ? node1255 : node1244;
									assign node1244 = (inp[4]) ? node1250 : node1245;
										assign node1245 = (inp[2]) ? 3'b010 : node1246;
											assign node1246 = (inp[3]) ? 3'b010 : 3'b110;
										assign node1250 = (inp[3]) ? node1252 : 3'b010;
											assign node1252 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1255 = (inp[2]) ? node1263 : node1256;
										assign node1256 = (inp[3]) ? 3'b110 : node1257;
											assign node1257 = (inp[4]) ? node1259 : 3'b001;
												assign node1259 = (inp[5]) ? 3'b110 : 3'b001;
										assign node1263 = (inp[5]) ? node1265 : 3'b110;
											assign node1265 = (inp[3]) ? node1267 : 3'b110;
												assign node1267 = (inp[4]) ? 3'b010 : 3'b110;
								assign node1270 = (inp[8]) ? node1286 : node1271;
									assign node1271 = (inp[5]) ? node1279 : node1272;
										assign node1272 = (inp[2]) ? node1276 : node1273;
											assign node1273 = (inp[3]) ? 3'b100 : 3'b010;
											assign node1276 = (inp[3]) ? 3'b000 : 3'b100;
										assign node1279 = (inp[4]) ? node1281 : 3'b100;
											assign node1281 = (inp[2]) ? node1283 : 3'b100;
												assign node1283 = (inp[3]) ? 3'b000 : 3'b100;
									assign node1286 = (inp[3]) ? node1292 : node1287;
										assign node1287 = (inp[2]) ? 3'b010 : node1288;
											assign node1288 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1292 = (inp[2]) ? node1294 : 3'b010;
											assign node1294 = (inp[4]) ? 3'b100 : node1295;
												assign node1295 = (inp[5]) ? 3'b000 : 3'b010;
							assign node1299 = (inp[8]) ? node1311 : node1300;
								assign node1300 = (inp[11]) ? 3'b000 : node1301;
									assign node1301 = (inp[2]) ? node1303 : 3'b100;
										assign node1303 = (inp[3]) ? 3'b000 : node1304;
											assign node1304 = (inp[5]) ? node1306 : 3'b100;
												assign node1306 = (inp[4]) ? 3'b000 : 3'b100;
								assign node1311 = (inp[11]) ? node1317 : node1312;
									assign node1312 = (inp[2]) ? node1314 : 3'b010;
										assign node1314 = (inp[3]) ? 3'b100 : 3'b010;
									assign node1317 = (inp[3]) ? node1325 : node1318;
										assign node1318 = (inp[2]) ? 3'b100 : node1319;
											assign node1319 = (inp[4]) ? 3'b000 : node1320;
												assign node1320 = (inp[5]) ? 3'b000 : 3'b010;
										assign node1325 = (inp[2]) ? 3'b000 : 3'b100;
						assign node1328 = (inp[1]) ? 3'b000 : node1329;
							assign node1329 = (inp[8]) ? node1331 : 3'b000;
								assign node1331 = (inp[11]) ? node1339 : node1332;
									assign node1332 = (inp[2]) ? 3'b100 : node1333;
										assign node1333 = (inp[3]) ? 3'b100 : node1334;
											assign node1334 = (inp[5]) ? 3'b010 : 3'b011;
									assign node1339 = (inp[2]) ? 3'b000 : node1340;
										assign node1340 = (inp[3]) ? 3'b000 : 3'b100;

endmodule