module dtc_split25_bm47 (
	input  wire [16-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node15;
	wire [1-1:0] node16;
	wire [1-1:0] node20;
	wire [1-1:0] node21;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node31;
	wire [1-1:0] node34;
	wire [1-1:0] node35;
	wire [1-1:0] node39;
	wire [1-1:0] node40;
	wire [1-1:0] node44;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node53;
	wire [1-1:0] node55;
	wire [1-1:0] node58;
	wire [1-1:0] node60;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node66;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node70;
	wire [1-1:0] node73;
	wire [1-1:0] node74;
	wire [1-1:0] node78;
	wire [1-1:0] node80;
	wire [1-1:0] node84;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node90;
	wire [1-1:0] node92;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node96;
	wire [1-1:0] node97;
	wire [1-1:0] node101;
	wire [1-1:0] node105;
	wire [1-1:0] node106;
	wire [1-1:0] node108;
	wire [1-1:0] node110;
	wire [1-1:0] node112;
	wire [1-1:0] node115;
	wire [1-1:0] node117;
	wire [1-1:0] node119;
	wire [1-1:0] node121;
	wire [1-1:0] node124;
	wire [1-1:0] node126;
	wire [1-1:0] node128;
	wire [1-1:0] node129;
	wire [1-1:0] node130;
	wire [1-1:0] node135;
	wire [1-1:0] node136;
	wire [1-1:0] node138;
	wire [1-1:0] node139;
	wire [1-1:0] node143;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node146;
	wire [1-1:0] node147;
	wire [1-1:0] node151;
	wire [1-1:0] node154;
	wire [1-1:0] node156;
	wire [1-1:0] node157;
	wire [1-1:0] node160;
	wire [1-1:0] node163;
	wire [1-1:0] node164;
	wire [1-1:0] node165;
	wire [1-1:0] node167;
	wire [1-1:0] node168;
	wire [1-1:0] node172;
	wire [1-1:0] node174;
	wire [1-1:0] node175;
	wire [1-1:0] node179;
	wire [1-1:0] node180;
	wire [1-1:0] node182;
	wire [1-1:0] node183;
	wire [1-1:0] node184;
	wire [1-1:0] node190;
	wire [1-1:0] node191;
	wire [1-1:0] node192;
	wire [1-1:0] node194;
	wire [1-1:0] node195;
	wire [1-1:0] node196;
	wire [1-1:0] node197;
	wire [1-1:0] node201;
	wire [1-1:0] node202;
	wire [1-1:0] node206;
	wire [1-1:0] node208;
	wire [1-1:0] node212;
	wire [1-1:0] node213;
	wire [1-1:0] node214;
	wire [1-1:0] node215;
	wire [1-1:0] node216;
	wire [1-1:0] node219;
	wire [1-1:0] node221;
	wire [1-1:0] node223;
	wire [1-1:0] node227;
	wire [1-1:0] node228;
	wire [1-1:0] node229;
	wire [1-1:0] node232;
	wire [1-1:0] node235;
	wire [1-1:0] node236;
	wire [1-1:0] node240;
	wire [1-1:0] node242;
	wire [1-1:0] node243;
	wire [1-1:0] node244;
	wire [1-1:0] node245;
	wire [1-1:0] node247;
	wire [1-1:0] node250;
	wire [1-1:0] node251;
	wire [1-1:0] node257;
	wire [1-1:0] node258;
	wire [1-1:0] node259;
	wire [1-1:0] node260;
	wire [1-1:0] node262;
	wire [1-1:0] node263;
	wire [1-1:0] node264;
	wire [1-1:0] node265;
	wire [1-1:0] node266;
	wire [1-1:0] node269;
	wire [1-1:0] node273;
	wire [1-1:0] node275;
	wire [1-1:0] node279;
	wire [1-1:0] node280;
	wire [1-1:0] node281;
	wire [1-1:0] node282;
	wire [1-1:0] node283;
	wire [1-1:0] node284;
	wire [1-1:0] node288;
	wire [1-1:0] node290;
	wire [1-1:0] node294;
	wire [1-1:0] node296;
	wire [1-1:0] node297;
	wire [1-1:0] node298;
	wire [1-1:0] node299;
	wire [1-1:0] node305;
	wire [1-1:0] node306;
	wire [1-1:0] node308;
	wire [1-1:0] node311;
	wire [1-1:0] node312;
	wire [1-1:0] node313;
	wire [1-1:0] node318;
	wire [1-1:0] node319;
	wire [1-1:0] node320;
	wire [1-1:0] node322;
	wire [1-1:0] node323;
	wire [1-1:0] node324;
	wire [1-1:0] node326;
	wire [1-1:0] node329;
	wire [1-1:0] node333;
	wire [1-1:0] node334;
	wire [1-1:0] node335;
	wire [1-1:0] node336;
	wire [1-1:0] node340;
	wire [1-1:0] node341;
	wire [1-1:0] node343;
	wire [1-1:0] node346;
	wire [1-1:0] node347;
	wire [1-1:0] node349;
	wire [1-1:0] node352;
	wire [1-1:0] node355;
	wire [1-1:0] node357;
	wire [1-1:0] node358;
	wire [1-1:0] node359;
	wire [1-1:0] node364;
	wire [1-1:0] node366;
	wire [1-1:0] node367;
	wire [1-1:0] node368;
	wire [1-1:0] node370;
	wire [1-1:0] node372;
	wire [1-1:0] node375;
	wire [1-1:0] node377;
	wire [1-1:0] node381;
	wire [1-1:0] node382;
	wire [1-1:0] node383;
	wire [1-1:0] node384;
	wire [1-1:0] node386;
	wire [1-1:0] node387;
	wire [1-1:0] node388;
	wire [1-1:0] node392;
	wire [1-1:0] node393;
	wire [1-1:0] node398;
	wire [1-1:0] node399;
	wire [1-1:0] node400;
	wire [1-1:0] node401;
	wire [1-1:0] node403;
	wire [1-1:0] node406;
	wire [1-1:0] node408;
	wire [1-1:0] node410;
	wire [1-1:0] node411;
	wire [1-1:0] node415;
	wire [1-1:0] node416;
	wire [1-1:0] node420;
	wire [1-1:0] node422;
	wire [1-1:0] node423;
	wire [1-1:0] node426;
	wire [1-1:0] node428;
	wire [1-1:0] node431;
	wire [1-1:0] node432;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node438;
	wire [1-1:0] node439;
	wire [1-1:0] node440;
	wire [1-1:0] node445;
	wire [1-1:0] node446;
	wire [1-1:0] node448;
	wire [1-1:0] node452;
	wire [1-1:0] node454;
	wire [1-1:0] node458;
	wire [1-1:0] node459;
	wire [1-1:0] node460;
	wire [1-1:0] node462;
	wire [1-1:0] node463;
	wire [1-1:0] node464;
	wire [1-1:0] node465;
	wire [1-1:0] node466;
	wire [1-1:0] node470;
	wire [1-1:0] node472;
	wire [1-1:0] node475;
	wire [1-1:0] node477;
	wire [1-1:0] node481;
	wire [1-1:0] node482;
	wire [1-1:0] node483;
	wire [1-1:0] node484;
	wire [1-1:0] node485;
	wire [1-1:0] node487;
	wire [1-1:0] node491;
	wire [1-1:0] node492;
	wire [1-1:0] node496;
	wire [1-1:0] node497;
	wire [1-1:0] node498;
	wire [1-1:0] node499;
	wire [1-1:0] node501;
	wire [1-1:0] node502;
	wire [1-1:0] node506;
	wire [1-1:0] node507;
	wire [1-1:0] node509;
	wire [1-1:0] node512;
	wire [1-1:0] node513;
	wire [1-1:0] node514;
	wire [1-1:0] node517;
	wire [1-1:0] node522;
	wire [1-1:0] node523;
	wire [1-1:0] node524;
	wire [1-1:0] node528;
	wire [1-1:0] node530;
	wire [1-1:0] node533;
	wire [1-1:0] node535;
	wire [1-1:0] node536;
	wire [1-1:0] node537;
	wire [1-1:0] node539;
	wire [1-1:0] node540;
	wire [1-1:0] node543;
	wire [1-1:0] node546;
	wire [1-1:0] node547;
	wire [1-1:0] node552;
	wire [1-1:0] node553;
	wire [1-1:0] node554;
	wire [1-1:0] node556;
	wire [1-1:0] node557;
	wire [1-1:0] node558;
	wire [1-1:0] node559;
	wire [1-1:0] node563;
	wire [1-1:0] node564;
	wire [1-1:0] node566;
	wire [1-1:0] node569;
	wire [1-1:0] node571;
	wire [1-1:0] node575;
	wire [1-1:0] node576;
	wire [1-1:0] node577;
	wire [1-1:0] node578;
	wire [1-1:0] node579;
	wire [1-1:0] node582;
	wire [1-1:0] node584;
	wire [1-1:0] node587;
	wire [1-1:0] node588;
	wire [1-1:0] node592;
	wire [1-1:0] node594;
	wire [1-1:0] node595;
	wire [1-1:0] node597;
	wire [1-1:0] node600;
	wire [1-1:0] node601;
	wire [1-1:0] node605;
	wire [1-1:0] node606;
	wire [1-1:0] node608;
	wire [1-1:0] node610;
	wire [1-1:0] node611;
	wire [1-1:0] node612;
	wire [1-1:0] node616;
	wire [1-1:0] node617;
	wire [1-1:0] node622;
	wire [1-1:0] node623;
	wire [1-1:0] node624;
	wire [1-1:0] node626;
	wire [1-1:0] node627;
	wire [1-1:0] node628;
	wire [1-1:0] node630;
	wire [1-1:0] node633;
	wire [1-1:0] node634;
	wire [1-1:0] node638;
	wire [1-1:0] node640;
	wire [1-1:0] node642;
	wire [1-1:0] node646;
	wire [1-1:0] node647;
	wire [1-1:0] node648;
	wire [1-1:0] node649;
	wire [1-1:0] node651;
	wire [1-1:0] node654;
	wire [1-1:0] node655;
	wire [1-1:0] node657;
	wire [1-1:0] node660;
	wire [1-1:0] node662;
	wire [1-1:0] node665;
	wire [1-1:0] node667;
	wire [1-1:0] node668;
	wire [1-1:0] node669;
	wire [1-1:0] node670;
	wire [1-1:0] node674;
	wire [1-1:0] node676;
	wire [1-1:0] node679;
	wire [1-1:0] node681;
	wire [1-1:0] node684;
	wire [1-1:0] node685;
	wire [1-1:0] node687;
	wire [1-1:0] node689;
	wire [1-1:0] node690;
	wire [1-1:0] node692;
	wire [1-1:0] node695;
	wire [1-1:0] node696;
	wire [1-1:0] node697;
	wire [1-1:0] node701;
	wire [1-1:0] node705;
	wire [1-1:0] node706;
	wire [1-1:0] node708;
	wire [1-1:0] node709;
	wire [1-1:0] node710;
	wire [1-1:0] node711;
	wire [1-1:0] node712;
	wire [1-1:0] node716;
	wire [1-1:0] node718;
	wire [1-1:0] node721;
	wire [1-1:0] node723;
	wire [1-1:0] node727;
	wire [1-1:0] node728;
	wire [1-1:0] node729;
	wire [1-1:0] node730;
	wire [1-1:0] node731;
	wire [1-1:0] node732;
	wire [1-1:0] node736;
	wire [1-1:0] node737;
	wire [1-1:0] node741;
	wire [1-1:0] node742;
	wire [1-1:0] node746;
	wire [1-1:0] node748;
	wire [1-1:0] node749;
	wire [1-1:0] node750;
	wire [1-1:0] node751;
	wire [1-1:0] node755;
	wire [1-1:0] node757;
	wire [1-1:0] node760;
	wire [1-1:0] node762;
	wire [1-1:0] node765;
	wire [1-1:0] node766;
	wire [1-1:0] node768;
	wire [1-1:0] node769;
	wire [1-1:0] node770;
	wire [1-1:0] node772;
	wire [1-1:0] node775;
	wire [1-1:0] node776;
	wire [1-1:0] node780;
	wire [1-1:0] node782;
	wire [1-1:0] node786;
	wire [1-1:0] node787;
	wire [1-1:0] node788;
	wire [1-1:0] node789;
	wire [1-1:0] node790;
	wire [1-1:0] node791;
	wire [1-1:0] node792;
	wire [1-1:0] node794;
	wire [1-1:0] node795;
	wire [1-1:0] node796;
	wire [1-1:0] node797;
	wire [1-1:0] node801;
	wire [1-1:0] node802;
	wire [1-1:0] node804;
	wire [1-1:0] node809;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node812;
	wire [1-1:0] node813;
	wire [1-1:0] node815;
	wire [1-1:0] node819;
	wire [1-1:0] node821;
	wire [1-1:0] node823;
	wire [1-1:0] node826;
	wire [1-1:0] node828;
	wire [1-1:0] node829;
	wire [1-1:0] node831;
	wire [1-1:0] node835;
	wire [1-1:0] node836;
	wire [1-1:0] node838;
	wire [1-1:0] node839;
	wire [1-1:0] node840;
	wire [1-1:0] node845;
	wire [1-1:0] node846;
	wire [1-1:0] node847;
	wire [1-1:0] node849;
	wire [1-1:0] node851;
	wire [1-1:0] node854;
	wire [1-1:0] node856;
	wire [1-1:0] node857;
	wire [1-1:0] node860;
	wire [1-1:0] node863;
	wire [1-1:0] node865;
	wire [1-1:0] node866;
	wire [1-1:0] node867;
	wire [1-1:0] node871;
	wire [1-1:0] node872;
	wire [1-1:0] node876;
	wire [1-1:0] node877;
	wire [1-1:0] node878;
	wire [1-1:0] node879;
	wire [1-1:0] node880;
	wire [1-1:0] node882;
	wire [1-1:0] node883;
	wire [1-1:0] node884;
	wire [1-1:0] node890;
	wire [1-1:0] node891;
	wire [1-1:0] node893;
	wire [1-1:0] node896;
	wire [1-1:0] node897;
	wire [1-1:0] node898;
	wire [1-1:0] node901;
	wire [1-1:0] node904;
	wire [1-1:0] node906;
	wire [1-1:0] node909;
	wire [1-1:0] node910;
	wire [1-1:0] node911;
	wire [1-1:0] node913;
	wire [1-1:0] node916;
	wire [1-1:0] node917;
	wire [1-1:0] node919;
	wire [1-1:0] node920;
	wire [1-1:0] node924;
	wire [1-1:0] node926;
	wire [1-1:0] node927;
	wire [1-1:0] node931;
	wire [1-1:0] node932;
	wire [1-1:0] node934;
	wire [1-1:0] node936;
	wire [1-1:0] node940;
	wire [1-1:0] node941;
	wire [1-1:0] node942;
	wire [1-1:0] node943;
	wire [1-1:0] node945;
	wire [1-1:0] node946;
	wire [1-1:0] node948;
	wire [1-1:0] node951;
	wire [1-1:0] node955;
	wire [1-1:0] node956;
	wire [1-1:0] node957;
	wire [1-1:0] node959;
	wire [1-1:0] node962;
	wire [1-1:0] node963;
	wire [1-1:0] node966;
	wire [1-1:0] node969;
	wire [1-1:0] node971;
	wire [1-1:0] node972;
	wire [1-1:0] node976;
	wire [1-1:0] node977;
	wire [1-1:0] node979;
	wire [1-1:0] node980;
	wire [1-1:0] node981;
	wire [1-1:0] node984;
	wire [1-1:0] node986;
	wire [1-1:0] node989;
	wire [1-1:0] node990;
	wire [1-1:0] node995;
	wire [1-1:0] node996;
	wire [1-1:0] node997;
	wire [1-1:0] node998;
	wire [1-1:0] node1000;
	wire [1-1:0] node1001;
	wire [1-1:0] node1002;
	wire [1-1:0] node1004;
	wire [1-1:0] node1007;
	wire [1-1:0] node1009;
	wire [1-1:0] node1011;
	wire [1-1:0] node1015;
	wire [1-1:0] node1016;
	wire [1-1:0] node1017;
	wire [1-1:0] node1018;
	wire [1-1:0] node1019;
	wire [1-1:0] node1021;
	wire [1-1:0] node1022;
	wire [1-1:0] node1025;
	wire [1-1:0] node1030;
	wire [1-1:0] node1031;
	wire [1-1:0] node1033;
	wire [1-1:0] node1036;
	wire [1-1:0] node1037;
	wire [1-1:0] node1040;
	wire [1-1:0] node1043;
	wire [1-1:0] node1045;
	wire [1-1:0] node1046;
	wire [1-1:0] node1047;
	wire [1-1:0] node1050;
	wire [1-1:0] node1054;
	wire [1-1:0] node1055;
	wire [1-1:0] node1056;
	wire [1-1:0] node1058;
	wire [1-1:0] node1059;
	wire [1-1:0] node1062;
	wire [1-1:0] node1064;
	wire [1-1:0] node1068;
	wire [1-1:0] node1069;
	wire [1-1:0] node1070;
	wire [1-1:0] node1071;
	wire [1-1:0] node1072;
	wire [1-1:0] node1077;
	wire [1-1:0] node1079;
	wire [1-1:0] node1082;
	wire [1-1:0] node1084;
	wire [1-1:0] node1085;
	wire [1-1:0] node1088;
	wire [1-1:0] node1090;
	wire [1-1:0] node1091;
	wire [1-1:0] node1094;
	wire [1-1:0] node1096;
	wire [1-1:0] node1099;
	wire [1-1:0] node1100;
	wire [1-1:0] node1101;
	wire [1-1:0] node1102;
	wire [1-1:0] node1104;
	wire [1-1:0] node1105;
	wire [1-1:0] node1106;
	wire [1-1:0] node1110;
	wire [1-1:0] node1112;
	wire [1-1:0] node1116;
	wire [1-1:0] node1117;
	wire [1-1:0] node1118;
	wire [1-1:0] node1119;
	wire [1-1:0] node1121;
	wire [1-1:0] node1124;
	wire [1-1:0] node1125;
	wire [1-1:0] node1130;
	wire [1-1:0] node1131;
	wire [1-1:0] node1132;
	wire [1-1:0] node1133;
	wire [1-1:0] node1135;
	wire [1-1:0] node1137;
	wire [1-1:0] node1141;
	wire [1-1:0] node1143;
	wire [1-1:0] node1144;
	wire [1-1:0] node1147;
	wire [1-1:0] node1150;
	wire [1-1:0] node1152;
	wire [1-1:0] node1155;
	wire [1-1:0] node1156;
	wire [1-1:0] node1158;
	wire [1-1:0] node1159;
	wire [1-1:0] node1161;
	wire [1-1:0] node1164;
	wire [1-1:0] node1165;
	wire [1-1:0] node1166;
	wire [1-1:0] node1170;
	wire [1-1:0] node1174;
	wire [1-1:0] node1175;
	wire [1-1:0] node1176;
	wire [1-1:0] node1177;
	wire [1-1:0] node1178;
	wire [1-1:0] node1180;
	wire [1-1:0] node1181;
	wire [1-1:0] node1182;
	wire [1-1:0] node1183;
	wire [1-1:0] node1187;
	wire [1-1:0] node1189;
	wire [1-1:0] node1192;
	wire [1-1:0] node1193;
	wire [1-1:0] node1195;
	wire [1-1:0] node1200;
	wire [1-1:0] node1201;
	wire [1-1:0] node1202;
	wire [1-1:0] node1203;
	wire [1-1:0] node1204;
	wire [1-1:0] node1206;
	wire [1-1:0] node1210;
	wire [1-1:0] node1212;
	wire [1-1:0] node1216;
	wire [1-1:0] node1217;
	wire [1-1:0] node1219;
	wire [1-1:0] node1222;
	wire [1-1:0] node1223;
	wire [1-1:0] node1226;
	wire [1-1:0] node1227;
	wire [1-1:0] node1230;
	wire [1-1:0] node1233;
	wire [1-1:0] node1234;
	wire [1-1:0] node1236;
	wire [1-1:0] node1237;
	wire [1-1:0] node1238;
	wire [1-1:0] node1242;
	wire [1-1:0] node1243;
	wire [1-1:0] node1244;
	wire [1-1:0] node1248;
	wire [1-1:0] node1250;
	wire [1-1:0] node1254;
	wire [1-1:0] node1255;
	wire [1-1:0] node1256;
	wire [1-1:0] node1257;
	wire [1-1:0] node1259;
	wire [1-1:0] node1260;
	wire [1-1:0] node1261;
	wire [1-1:0] node1264;
	wire [1-1:0] node1266;
	wire [1-1:0] node1269;
	wire [1-1:0] node1271;
	wire [1-1:0] node1275;
	wire [1-1:0] node1276;
	wire [1-1:0] node1277;
	wire [1-1:0] node1278;
	wire [1-1:0] node1280;
	wire [1-1:0] node1283;
	wire [1-1:0] node1284;
	wire [1-1:0] node1285;
	wire [1-1:0] node1287;
	wire [1-1:0] node1290;
	wire [1-1:0] node1291;
	wire [1-1:0] node1295;
	wire [1-1:0] node1298;
	wire [1-1:0] node1300;
	wire [1-1:0] node1301;
	wire [1-1:0] node1302;
	wire [1-1:0] node1305;
	wire [1-1:0] node1308;
	wire [1-1:0] node1309;
	wire [1-1:0] node1313;
	wire [1-1:0] node1315;
	wire [1-1:0] node1316;
	wire [1-1:0] node1317;
	wire [1-1:0] node1318;
	wire [1-1:0] node1320;
	wire [1-1:0] node1321;
	wire [1-1:0] node1325;
	wire [1-1:0] node1326;
	wire [1-1:0] node1328;
	wire [1-1:0] node1331;
	wire [1-1:0] node1334;
	wire [1-1:0] node1336;
	wire [1-1:0] node1340;
	wire [1-1:0] node1341;
	wire [1-1:0] node1343;
	wire [1-1:0] node1344;
	wire [1-1:0] node1345;
	wire [1-1:0] node1346;
	wire [1-1:0] node1349;
	wire [1-1:0] node1350;
	wire [1-1:0] node1354;
	wire [1-1:0] node1355;
	wire [1-1:0] node1360;
	wire [1-1:0] node1361;
	wire [1-1:0] node1362;
	wire [1-1:0] node1363;
	wire [1-1:0] node1364;
	wire [1-1:0] node1365;
	wire [1-1:0] node1368;
	wire [1-1:0] node1372;
	wire [1-1:0] node1373;
	wire [1-1:0] node1377;
	wire [1-1:0] node1378;
	wire [1-1:0] node1379;
	wire [1-1:0] node1381;
	wire [1-1:0] node1385;
	wire [1-1:0] node1387;
	wire [1-1:0] node1390;
	wire [1-1:0] node1391;
	wire [1-1:0] node1393;
	wire [1-1:0] node1395;
	wire [1-1:0] node1396;
	wire [1-1:0] node1397;
	wire [1-1:0] node1401;
	wire [1-1:0] node1405;
	wire [1-1:0] node1406;
	wire [1-1:0] node1407;
	wire [1-1:0] node1408;
	wire [1-1:0] node1410;
	wire [1-1:0] node1411;
	wire [1-1:0] node1412;
	wire [1-1:0] node1413;
	wire [1-1:0] node1417;
	wire [1-1:0] node1419;
	wire [1-1:0] node1422;
	wire [1-1:0] node1423;
	wire [1-1:0] node1428;
	wire [1-1:0] node1429;
	wire [1-1:0] node1430;
	wire [1-1:0] node1431;
	wire [1-1:0] node1432;
	wire [1-1:0] node1433;
	wire [1-1:0] node1436;
	wire [1-1:0] node1437;
	wire [1-1:0] node1441;
	wire [1-1:0] node1442;
	wire [1-1:0] node1447;
	wire [1-1:0] node1448;
	wire [1-1:0] node1450;
	wire [1-1:0] node1453;
	wire [1-1:0] node1454;
	wire [1-1:0] node1456;
	wire [1-1:0] node1459;
	wire [1-1:0] node1461;
	wire [1-1:0] node1464;
	wire [1-1:0] node1466;
	wire [1-1:0] node1467;
	wire [1-1:0] node1468;
	wire [1-1:0] node1469;
	wire [1-1:0] node1470;
	wire [1-1:0] node1474;
	wire [1-1:0] node1475;
	wire [1-1:0] node1479;
	wire [1-1:0] node1480;
	wire [1-1:0] node1485;
	wire [1-1:0] node1486;
	wire [1-1:0] node1487;
	wire [1-1:0] node1488;
	wire [1-1:0] node1489;
	wire [1-1:0] node1490;
	wire [1-1:0] node1492;
	wire [1-1:0] node1493;
	wire [1-1:0] node1497;
	wire [1-1:0] node1498;
	wire [1-1:0] node1499;
	wire [1-1:0] node1500;
	wire [1-1:0] node1504;
	wire [1-1:0] node1507;
	wire [1-1:0] node1508;
	wire [1-1:0] node1509;
	wire [1-1:0] node1510;
	wire [1-1:0] node1514;
	wire [1-1:0] node1517;
	wire [1-1:0] node1520;
	wire [1-1:0] node1521;
	wire [1-1:0] node1522;
	wire [1-1:0] node1523;
	wire [1-1:0] node1524;
	wire [1-1:0] node1525;
	wire [1-1:0] node1529;
	wire [1-1:0] node1531;
	wire [1-1:0] node1534;
	wire [1-1:0] node1535;
	wire [1-1:0] node1539;
	wire [1-1:0] node1541;
	wire [1-1:0] node1544;
	wire [1-1:0] node1545;
	wire [1-1:0] node1546;
	wire [1-1:0] node1548;
	wire [1-1:0] node1550;
	wire [1-1:0] node1551;
	wire [1-1:0] node1555;
	wire [1-1:0] node1557;
	wire [1-1:0] node1560;
	wire [1-1:0] node1562;
	wire [1-1:0] node1564;
	wire [1-1:0] node1566;
	wire [1-1:0] node1567;
	wire [1-1:0] node1571;
	wire [1-1:0] node1572;
	wire [1-1:0] node1574;
	wire [1-1:0] node1575;
	wire [1-1:0] node1576;
	wire [1-1:0] node1577;
	wire [1-1:0] node1583;
	wire [1-1:0] node1584;
	wire [1-1:0] node1585;
	wire [1-1:0] node1587;
	wire [1-1:0] node1589;
	wire [1-1:0] node1592;
	wire [1-1:0] node1594;
	wire [1-1:0] node1597;
	wire [1-1:0] node1598;
	wire [1-1:0] node1599;
	wire [1-1:0] node1601;
	wire [1-1:0] node1604;
	wire [1-1:0] node1605;
	wire [1-1:0] node1608;
	wire [1-1:0] node1611;
	wire [1-1:0] node1613;
	wire [1-1:0] node1614;
	wire [1-1:0] node1616;
	wire [1-1:0] node1620;
	wire [1-1:0] node1621;
	wire [1-1:0] node1622;
	wire [1-1:0] node1623;
	wire [1-1:0] node1625;
	wire [1-1:0] node1626;
	wire [1-1:0] node1630;
	wire [1-1:0] node1631;
	wire [1-1:0] node1632;
	wire [1-1:0] node1635;
	wire [1-1:0] node1637;
	wire [1-1:0] node1640;
	wire [1-1:0] node1642;
	wire [1-1:0] node1644;
	wire [1-1:0] node1647;
	wire [1-1:0] node1648;
	wire [1-1:0] node1649;
	wire [1-1:0] node1653;
	wire [1-1:0] node1654;
	wire [1-1:0] node1655;
	wire [1-1:0] node1657;
	wire [1-1:0] node1660;
	wire [1-1:0] node1662;
	wire [1-1:0] node1663;
	wire [1-1:0] node1664;
	wire [1-1:0] node1669;
	wire [1-1:0] node1670;
	wire [1-1:0] node1672;
	wire [1-1:0] node1673;
	wire [1-1:0] node1678;
	wire [1-1:0] node1679;
	wire [1-1:0] node1681;
	wire [1-1:0] node1682;
	wire [1-1:0] node1683;
	wire [1-1:0] node1685;
	wire [1-1:0] node1688;
	wire [1-1:0] node1689;
	wire [1-1:0] node1691;
	wire [1-1:0] node1693;
	wire [1-1:0] node1696;
	wire [1-1:0] node1698;
	wire [1-1:0] node1702;
	wire [1-1:0] node1703;
	wire [1-1:0] node1704;
	wire [1-1:0] node1706;
	wire [1-1:0] node1707;
	wire [1-1:0] node1708;
	wire [1-1:0] node1711;
	wire [1-1:0] node1715;
	wire [1-1:0] node1716;
	wire [1-1:0] node1718;
	wire [1-1:0] node1720;
	wire [1-1:0] node1723;
	wire [1-1:0] node1725;
	wire [1-1:0] node1728;
	wire [1-1:0] node1729;
	wire [1-1:0] node1730;
	wire [1-1:0] node1731;
	wire [1-1:0] node1733;
	wire [1-1:0] node1737;
	wire [1-1:0] node1738;
	wire [1-1:0] node1742;
	wire [1-1:0] node1744;
	wire [1-1:0] node1747;
	wire [1-1:0] node1748;
	wire [1-1:0] node1749;
	wire [1-1:0] node1750;
	wire [1-1:0] node1751;
	wire [1-1:0] node1752;
	wire [1-1:0] node1753;
	wire [1-1:0] node1755;
	wire [1-1:0] node1758;
	wire [1-1:0] node1760;
	wire [1-1:0] node1763;
	wire [1-1:0] node1765;
	wire [1-1:0] node1768;
	wire [1-1:0] node1770;
	wire [1-1:0] node1771;
	wire [1-1:0] node1772;
	wire [1-1:0] node1777;
	wire [1-1:0] node1779;
	wire [1-1:0] node1780;
	wire [1-1:0] node1781;
	wire [1-1:0] node1782;
	wire [1-1:0] node1784;
	wire [1-1:0] node1789;
	wire [1-1:0] node1790;
	wire [1-1:0] node1791;
	wire [1-1:0] node1795;
	wire [1-1:0] node1796;
	wire [1-1:0] node1798;
	wire [1-1:0] node1801;
	wire [1-1:0] node1803;
	wire [1-1:0] node1806;
	wire [1-1:0] node1807;
	wire [1-1:0] node1809;
	wire [1-1:0] node1810;
	wire [1-1:0] node1811;
	wire [1-1:0] node1812;
	wire [1-1:0] node1813;
	wire [1-1:0] node1818;
	wire [1-1:0] node1819;
	wire [1-1:0] node1824;
	wire [1-1:0] node1825;
	wire [1-1:0] node1826;
	wire [1-1:0] node1827;
	wire [1-1:0] node1829;
	wire [1-1:0] node1833;
	wire [1-1:0] node1835;
	wire [1-1:0] node1836;
	wire [1-1:0] node1837;
	wire [1-1:0] node1841;
	wire [1-1:0] node1844;
	wire [1-1:0] node1845;
	wire [1-1:0] node1847;
	wire [1-1:0] node1848;
	wire [1-1:0] node1850;
	wire [1-1:0] node1851;
	wire [1-1:0] node1857;
	wire [1-1:0] node1858;
	wire [1-1:0] node1860;
	wire [1-1:0] node1861;
	wire [1-1:0] node1862;
	wire [1-1:0] node1864;
	wire [1-1:0] node1867;
	wire [1-1:0] node1868;
	wire [1-1:0] node1870;
	wire [1-1:0] node1875;
	wire [1-1:0] node1876;
	wire [1-1:0] node1877;
	wire [1-1:0] node1878;
	wire [1-1:0] node1880;
	wire [1-1:0] node1883;
	wire [1-1:0] node1884;
	wire [1-1:0] node1885;
	wire [1-1:0] node1890;
	wire [1-1:0] node1892;
	wire [1-1:0] node1894;
	wire [1-1:0] node1895;
	wire [1-1:0] node1897;
	wire [1-1:0] node1900;
	wire [1-1:0] node1903;
	wire [1-1:0] node1904;
	wire [1-1:0] node1906;
	wire [1-1:0] node1907;
	wire [1-1:0] node1909;
	wire [1-1:0] node1912;
	wire [1-1:0] node1913;
	wire [1-1:0] node1914;
	wire [1-1:0] node1915;
	wire [1-1:0] node1919;
	wire [1-1:0] node1920;
	wire [1-1:0] node1926;
	wire [1-1:0] node1927;
	wire [1-1:0] node1928;
	wire [1-1:0] node1929;
	wire [1-1:0] node1930;
	wire [1-1:0] node1932;
	wire [1-1:0] node1933;
	wire [1-1:0] node1935;
	wire [1-1:0] node1938;
	wire [1-1:0] node1939;
	wire [1-1:0] node1940;
	wire [1-1:0] node1944;
	wire [1-1:0] node1946;
	wire [1-1:0] node1950;
	wire [1-1:0] node1951;
	wire [1-1:0] node1952;
	wire [1-1:0] node1953;
	wire [1-1:0] node1954;
	wire [1-1:0] node1958;
	wire [1-1:0] node1959;
	wire [1-1:0] node1963;
	wire [1-1:0] node1965;
	wire [1-1:0] node1968;
	wire [1-1:0] node1970;
	wire [1-1:0] node1971;
	wire [1-1:0] node1972;
	wire [1-1:0] node1976;
	wire [1-1:0] node1977;
	wire [1-1:0] node1979;
	wire [1-1:0] node1982;
	wire [1-1:0] node1983;
	wire [1-1:0] node1987;
	wire [1-1:0] node1989;
	wire [1-1:0] node1990;
	wire [1-1:0] node1991;
	wire [1-1:0] node1992;
	wire [1-1:0] node1994;
	wire [1-1:0] node1997;
	wire [1-1:0] node1998;
	wire [1-1:0] node2002;
	wire [1-1:0] node2003;
	wire [1-1:0] node2008;
	wire [1-1:0] node2009;
	wire [1-1:0] node2010;
	wire [1-1:0] node2011;
	wire [1-1:0] node2012;
	wire [1-1:0] node2013;
	wire [1-1:0] node2014;
	wire [1-1:0] node2016;
	wire [1-1:0] node2017;
	wire [1-1:0] node2019;
	wire [1-1:0] node2023;
	wire [1-1:0] node2024;
	wire [1-1:0] node2025;
	wire [1-1:0] node2026;
	wire [1-1:0] node2027;
	wire [1-1:0] node2029;
	wire [1-1:0] node2034;
	wire [1-1:0] node2035;
	wire [1-1:0] node2038;
	wire [1-1:0] node2039;
	wire [1-1:0] node2040;
	wire [1-1:0] node2044;
	wire [1-1:0] node2046;
	wire [1-1:0] node2049;
	wire [1-1:0] node2051;
	wire [1-1:0] node2052;
	wire [1-1:0] node2053;
	wire [1-1:0] node2058;
	wire [1-1:0] node2059;
	wire [1-1:0] node2061;
	wire [1-1:0] node2062;
	wire [1-1:0] node2064;
	wire [1-1:0] node2066;
	wire [1-1:0] node2069;
	wire [1-1:0] node2070;
	wire [1-1:0] node2074;
	wire [1-1:0] node2075;
	wire [1-1:0] node2076;
	wire [1-1:0] node2078;
	wire [1-1:0] node2082;
	wire [1-1:0] node2083;
	wire [1-1:0] node2085;
	wire [1-1:0] node2088;
	wire [1-1:0] node2089;
	wire [1-1:0] node2090;
	wire [1-1:0] node2093;
	wire [1-1:0] node2095;
	wire [1-1:0] node2099;
	wire [1-1:0] node2100;
	wire [1-1:0] node2101;
	wire [1-1:0] node2103;
	wire [1-1:0] node2104;
	wire [1-1:0] node2106;
	wire [1-1:0] node2111;
	wire [1-1:0] node2112;
	wire [1-1:0] node2113;
	wire [1-1:0] node2115;
	wire [1-1:0] node2117;
	wire [1-1:0] node2118;
	wire [1-1:0] node2121;
	wire [1-1:0] node2124;
	wire [1-1:0] node2126;
	wire [1-1:0] node2128;
	wire [1-1:0] node2131;
	wire [1-1:0] node2132;
	wire [1-1:0] node2134;
	wire [1-1:0] node2138;
	wire [1-1:0] node2139;
	wire [1-1:0] node2140;
	wire [1-1:0] node2141;
	wire [1-1:0] node2142;
	wire [1-1:0] node2144;
	wire [1-1:0] node2146;
	wire [1-1:0] node2150;
	wire [1-1:0] node2151;
	wire [1-1:0] node2152;
	wire [1-1:0] node2153;
	wire [1-1:0] node2157;
	wire [1-1:0] node2159;
	wire [1-1:0] node2162;
	wire [1-1:0] node2164;
	wire [1-1:0] node2166;
	wire [1-1:0] node2169;
	wire [1-1:0] node2171;
	wire [1-1:0] node2172;
	wire [1-1:0] node2174;
	wire [1-1:0] node2176;
	wire [1-1:0] node2180;
	wire [1-1:0] node2181;
	wire [1-1:0] node2182;
	wire [1-1:0] node2183;
	wire [1-1:0] node2185;
	wire [1-1:0] node2187;
	wire [1-1:0] node2191;
	wire [1-1:0] node2192;
	wire [1-1:0] node2194;
	wire [1-1:0] node2197;
	wire [1-1:0] node2198;
	wire [1-1:0] node2199;
	wire [1-1:0] node2203;
	wire [1-1:0] node2204;
	wire [1-1:0] node2208;
	wire [1-1:0] node2209;
	wire [1-1:0] node2211;
	wire [1-1:0] node2212;
	wire [1-1:0] node2214;
	wire [1-1:0] node2215;
	wire [1-1:0] node2220;
	wire [1-1:0] node2221;
	wire [1-1:0] node2222;
	wire [1-1:0] node2223;
	wire [1-1:0] node2224;
	wire [1-1:0] node2230;
	wire [1-1:0] node2231;
	wire [1-1:0] node2233;
	wire [1-1:0] node2236;
	wire [1-1:0] node2237;
	wire [1-1:0] node2241;
	wire [1-1:0] node2242;
	wire [1-1:0] node2243;
	wire [1-1:0] node2244;
	wire [1-1:0] node2246;
	wire [1-1:0] node2247;
	wire [1-1:0] node2248;
	wire [1-1:0] node2249;
	wire [1-1:0] node2253;
	wire [1-1:0] node2254;
	wire [1-1:0] node2259;
	wire [1-1:0] node2260;
	wire [1-1:0] node2261;
	wire [1-1:0] node2262;
	wire [1-1:0] node2263;
	wire [1-1:0] node2266;
	wire [1-1:0] node2268;
	wire [1-1:0] node2270;
	wire [1-1:0] node2273;
	wire [1-1:0] node2275;
	wire [1-1:0] node2279;
	wire [1-1:0] node2280;
	wire [1-1:0] node2282;
	wire [1-1:0] node2285;
	wire [1-1:0] node2286;
	wire [1-1:0] node2288;
	wire [1-1:0] node2289;
	wire [1-1:0] node2291;
	wire [1-1:0] node2295;
	wire [1-1:0] node2296;
	wire [1-1:0] node2300;
	wire [1-1:0] node2301;
	wire [1-1:0] node2303;
	wire [1-1:0] node2304;
	wire [1-1:0] node2305;
	wire [1-1:0] node2306;
	wire [1-1:0] node2311;
	wire [1-1:0] node2312;
	wire [1-1:0] node2313;
	wire [1-1:0] node2317;
	wire [1-1:0] node2319;
	wire [1-1:0] node2320;
	wire [1-1:0] node2321;
	wire [1-1:0] node2327;
	wire [1-1:0] node2328;
	wire [1-1:0] node2329;
	wire [1-1:0] node2330;
	wire [1-1:0] node2331;
	wire [1-1:0] node2333;
	wire [1-1:0] node2334;
	wire [1-1:0] node2336;
	wire [1-1:0] node2337;
	wire [1-1:0] node2343;
	wire [1-1:0] node2344;
	wire [1-1:0] node2345;
	wire [1-1:0] node2346;
	wire [1-1:0] node2348;
	wire [1-1:0] node2351;
	wire [1-1:0] node2354;
	wire [1-1:0] node2355;
	wire [1-1:0] node2359;
	wire [1-1:0] node2362;
	wire [1-1:0] node2364;
	wire [1-1:0] node2365;
	wire [1-1:0] node2366;
	wire [1-1:0] node2367;
	wire [1-1:0] node2371;
	wire [1-1:0] node2373;
	wire [1-1:0] node2377;
	wire [1-1:0] node2378;
	wire [1-1:0] node2379;
	wire [1-1:0] node2380;
	wire [1-1:0] node2382;
	wire [1-1:0] node2383;
	wire [1-1:0] node2384;
	wire [1-1:0] node2390;
	wire [1-1:0] node2391;
	wire [1-1:0] node2393;
	wire [1-1:0] node2394;
	wire [1-1:0] node2398;
	wire [1-1:0] node2399;
	wire [1-1:0] node2401;
	wire [1-1:0] node2405;
	wire [1-1:0] node2406;
	wire [1-1:0] node2407;
	wire [1-1:0] node2409;
	wire [1-1:0] node2411;
	wire [1-1:0] node2415;
	wire [1-1:0] node2416;
	wire [1-1:0] node2418;
	wire [1-1:0] node2420;
	wire [1-1:0] node2422;
	wire [1-1:0] node2425;
	wire [1-1:0] node2426;
	wire [1-1:0] node2430;
	wire [1-1:0] node2431;
	wire [1-1:0] node2432;
	wire [1-1:0] node2434;
	wire [1-1:0] node2435;
	wire [1-1:0] node2437;
	wire [1-1:0] node2440;
	wire [1-1:0] node2441;
	wire [1-1:0] node2443;
	wire [1-1:0] node2446;
	wire [1-1:0] node2447;
	wire [1-1:0] node2452;
	wire [1-1:0] node2453;
	wire [1-1:0] node2454;
	wire [1-1:0] node2455;
	wire [1-1:0] node2456;
	wire [1-1:0] node2457;
	wire [1-1:0] node2458;
	wire [1-1:0] node2462;
	wire [1-1:0] node2463;
	wire [1-1:0] node2467;
	wire [1-1:0] node2468;
	wire [1-1:0] node2473;
	wire [1-1:0] node2474;
	wire [1-1:0] node2475;
	wire [1-1:0] node2479;
	wire [1-1:0] node2480;
	wire [1-1:0] node2481;
	wire [1-1:0] node2485;
	wire [1-1:0] node2486;
	wire [1-1:0] node2490;
	wire [1-1:0] node2491;
	wire [1-1:0] node2493;
	wire [1-1:0] node2494;
	wire [1-1:0] node2495;
	wire [1-1:0] node2496;
	wire [1-1:0] node2500;
	wire [1-1:0] node2501;
	wire [1-1:0] node2505;
	wire [1-1:0] node2506;

	assign outp = (inp[6]) ? node786 : node1;
		assign node1 = (inp[15]) ? node705 : node2;
			assign node2 = (inp[12]) ? node84 : node3;
				assign node3 = (inp[4]) ? node63 : node4;
					assign node4 = (inp[0]) ? node26 : node5;
						assign node5 = (inp[1]) ? node7 : 1'b1;
							assign node7 = (inp[8]) ? 1'b1 : node8;
								assign node8 = (inp[2]) ? node20 : node9;
									assign node9 = (inp[14]) ? node15 : node10;
										assign node10 = (inp[13]) ? node12 : 1'b0;
											assign node12 = (inp[11]) ? 1'b0 : 1'b1;
										assign node15 = (inp[11]) ? 1'b1 : node16;
											assign node16 = (inp[13]) ? 1'b0 : 1'b1;
									assign node20 = (inp[11]) ? 1'b0 : node21;
										assign node21 = (inp[13]) ? 1'b1 : 1'b0;
						assign node26 = (inp[1]) ? node44 : node27;
							assign node27 = (inp[11]) ? node39 : node28;
								assign node28 = (inp[13]) ? node34 : node29;
									assign node29 = (inp[14]) ? node31 : 1'b0;
										assign node31 = (inp[2]) ? 1'b0 : 1'b1;
									assign node34 = (inp[2]) ? 1'b1 : node35;
										assign node35 = (inp[14]) ? 1'b0 : 1'b1;
								assign node39 = (inp[2]) ? 1'b0 : node40;
									assign node40 = (inp[14]) ? 1'b1 : 1'b0;
							assign node44 = (inp[8]) ? node46 : 1'b1;
								assign node46 = (inp[11]) ? node58 : node47;
									assign node47 = (inp[13]) ? node53 : node48;
										assign node48 = (inp[2]) ? 1'b0 : node49;
											assign node49 = (inp[14]) ? 1'b1 : 1'b0;
										assign node53 = (inp[14]) ? node55 : 1'b1;
											assign node55 = (inp[2]) ? 1'b1 : 1'b0;
									assign node58 = (inp[14]) ? node60 : 1'b0;
										assign node60 = (inp[2]) ? 1'b0 : 1'b1;
					assign node63 = (inp[1]) ? node65 : 1'b1;
						assign node65 = (inp[8]) ? 1'b1 : node66;
							assign node66 = (inp[11]) ? node78 : node67;
								assign node67 = (inp[13]) ? node73 : node68;
									assign node68 = (inp[14]) ? node70 : 1'b0;
										assign node70 = (inp[2]) ? 1'b0 : 1'b1;
									assign node73 = (inp[2]) ? 1'b1 : node74;
										assign node74 = (inp[14]) ? 1'b0 : 1'b1;
								assign node78 = (inp[14]) ? node80 : 1'b0;
									assign node80 = (inp[2]) ? 1'b0 : 1'b1;
				assign node84 = (inp[10]) ? node458 : node85;
					assign node85 = (inp[9]) ? node257 : node86;
						assign node86 = (inp[7]) ? node190 : node87;
							assign node87 = (inp[3]) ? node135 : node88;
								assign node88 = (inp[4]) ? node124 : node89;
									assign node89 = (inp[0]) ? node105 : node90;
										assign node90 = (inp[1]) ? node92 : 1'b0;
											assign node92 = (inp[8]) ? 1'b0 : node93;
												assign node93 = (inp[14]) ? node101 : node94;
													assign node94 = (inp[2]) ? node96 : 1'b1;
														assign node96 = (inp[11]) ? 1'b1 : node97;
															assign node97 = (inp[13]) ? 1'b0 : 1'b1;
													assign node101 = (inp[13]) ? 1'b1 : 1'b0;
										assign node105 = (inp[14]) ? node115 : node106;
											assign node106 = (inp[13]) ? node108 : 1'b1;
												assign node108 = (inp[11]) ? node110 : 1'b0;
													assign node110 = (inp[1]) ? node112 : 1'b1;
														assign node112 = (inp[8]) ? 1'b1 : 1'b0;
											assign node115 = (inp[11]) ? node117 : 1'b0;
												assign node117 = (inp[2]) ? node119 : 1'b0;
													assign node119 = (inp[1]) ? node121 : 1'b1;
														assign node121 = (inp[13]) ? 1'b1 : 1'b0;
									assign node124 = (inp[11]) ? node126 : 1'b0;
										assign node126 = (inp[1]) ? node128 : 1'b0;
											assign node128 = (inp[8]) ? 1'b0 : node129;
												assign node129 = (inp[2]) ? 1'b1 : node130;
													assign node130 = (inp[14]) ? 1'b0 : 1'b1;
								assign node135 = (inp[1]) ? node143 : node136;
									assign node136 = (inp[0]) ? node138 : 1'b1;
										assign node138 = (inp[4]) ? 1'b1 : node139;
											assign node139 = (inp[11]) ? 1'b0 : 1'b1;
									assign node143 = (inp[13]) ? node163 : node144;
										assign node144 = (inp[14]) ? node154 : node145;
											assign node145 = (inp[8]) ? node151 : node146;
												assign node146 = (inp[4]) ? 1'b0 : node147;
													assign node147 = (inp[0]) ? 1'b1 : 1'b0;
												assign node151 = (inp[4]) ? 1'b1 : 1'b0;
											assign node154 = (inp[2]) ? node156 : 1'b1;
												assign node156 = (inp[8]) ? node160 : node157;
													assign node157 = (inp[0]) ? 1'b1 : 1'b0;
													assign node160 = (inp[0]) ? 1'b0 : 1'b1;
										assign node163 = (inp[4]) ? node179 : node164;
											assign node164 = (inp[2]) ? node172 : node165;
												assign node165 = (inp[14]) ? node167 : 1'b1;
													assign node167 = (inp[0]) ? 1'b1 : node168;
														assign node168 = (inp[8]) ? 1'b1 : 1'b0;
												assign node172 = (inp[11]) ? node174 : 1'b1;
													assign node174 = (inp[14]) ? 1'b0 : node175;
														assign node175 = (inp[8]) ? 1'b0 : 1'b1;
											assign node179 = (inp[8]) ? 1'b1 : node180;
												assign node180 = (inp[14]) ? node182 : 1'b1;
													assign node182 = (inp[0]) ? 1'b1 : node183;
														assign node183 = (inp[2]) ? 1'b1 : node184;
															assign node184 = (inp[11]) ? 1'b1 : 1'b0;
							assign node190 = (inp[0]) ? node212 : node191;
								assign node191 = (inp[8]) ? 1'b0 : node192;
									assign node192 = (inp[1]) ? node194 : 1'b0;
										assign node194 = (inp[2]) ? node206 : node195;
											assign node195 = (inp[14]) ? node201 : node196;
												assign node196 = (inp[11]) ? 1'b1 : node197;
													assign node197 = (inp[13]) ? 1'b0 : 1'b1;
												assign node201 = (inp[11]) ? 1'b0 : node202;
													assign node202 = (inp[13]) ? 1'b1 : 1'b0;
											assign node206 = (inp[13]) ? node208 : 1'b1;
												assign node208 = (inp[11]) ? 1'b1 : 1'b0;
								assign node212 = (inp[4]) ? node240 : node213;
									assign node213 = (inp[8]) ? node227 : node214;
										assign node214 = (inp[1]) ? 1'b0 : node215;
											assign node215 = (inp[14]) ? node219 : node216;
												assign node216 = (inp[5]) ? 1'b0 : 1'b1;
												assign node219 = (inp[2]) ? node221 : 1'b0;
													assign node221 = (inp[13]) ? node223 : 1'b1;
														assign node223 = (inp[5]) ? 1'b1 : 1'b0;
										assign node227 = (inp[2]) ? node235 : node228;
											assign node228 = (inp[14]) ? node232 : node229;
												assign node229 = (inp[3]) ? 1'b0 : 1'b1;
												assign node232 = (inp[13]) ? 1'b1 : 1'b0;
											assign node235 = (inp[11]) ? 1'b1 : node236;
												assign node236 = (inp[13]) ? 1'b0 : 1'b1;
									assign node240 = (inp[1]) ? node242 : 1'b0;
										assign node242 = (inp[8]) ? 1'b0 : node243;
											assign node243 = (inp[11]) ? 1'b1 : node244;
												assign node244 = (inp[13]) ? node250 : node245;
													assign node245 = (inp[14]) ? node247 : 1'b1;
														assign node247 = (inp[2]) ? 1'b1 : 1'b0;
													assign node250 = (inp[2]) ? 1'b0 : node251;
														assign node251 = (inp[14]) ? 1'b1 : 1'b0;
						assign node257 = (inp[7]) ? node381 : node258;
							assign node258 = (inp[3]) ? node318 : node259;
								assign node259 = (inp[1]) ? node279 : node260;
									assign node260 = (inp[0]) ? node262 : 1'b1;
										assign node262 = (inp[4]) ? 1'b1 : node263;
											assign node263 = (inp[11]) ? node273 : node264;
												assign node264 = (inp[2]) ? 1'b1 : node265;
													assign node265 = (inp[14]) ? node269 : node266;
														assign node266 = (inp[13]) ? 1'b1 : 1'b0;
														assign node269 = (inp[13]) ? 1'b0 : 1'b1;
												assign node273 = (inp[14]) ? node275 : 1'b0;
													assign node275 = (inp[2]) ? 1'b0 : 1'b1;
									assign node279 = (inp[8]) ? node305 : node280;
										assign node280 = (inp[4]) ? node294 : node281;
											assign node281 = (inp[0]) ? 1'b1 : node282;
												assign node282 = (inp[2]) ? node288 : node283;
													assign node283 = (inp[5]) ? 1'b0 : node284;
														assign node284 = (inp[14]) ? 1'b1 : 1'b0;
													assign node288 = (inp[13]) ? node290 : 1'b0;
														assign node290 = (inp[5]) ? 1'b1 : 1'b0;
											assign node294 = (inp[13]) ? node296 : 1'b0;
												assign node296 = (inp[2]) ? 1'b0 : node297;
													assign node297 = (inp[0]) ? 1'b1 : node298;
														assign node298 = (inp[14]) ? 1'b0 : node299;
															assign node299 = (inp[11]) ? 1'b0 : 1'b1;
										assign node305 = (inp[14]) ? node311 : node306;
											assign node306 = (inp[0]) ? node308 : 1'b1;
												assign node308 = (inp[4]) ? 1'b1 : 1'b0;
											assign node311 = (inp[4]) ? 1'b1 : node312;
												assign node312 = (inp[13]) ? 1'b1 : node313;
													assign node313 = (inp[11]) ? 1'b0 : 1'b1;
								assign node318 = (inp[8]) ? node364 : node319;
									assign node319 = (inp[1]) ? node333 : node320;
										assign node320 = (inp[0]) ? node322 : 1'b0;
											assign node322 = (inp[4]) ? 1'b0 : node323;
												assign node323 = (inp[13]) ? node329 : node324;
													assign node324 = (inp[11]) ? node326 : 1'b1;
														assign node326 = (inp[2]) ? 1'b1 : 1'b0;
													assign node329 = (inp[2]) ? 1'b0 : 1'b1;
										assign node333 = (inp[0]) ? node355 : node334;
											assign node334 = (inp[13]) ? node340 : node335;
												assign node335 = (inp[2]) ? 1'b1 : node336;
													assign node336 = (inp[14]) ? 1'b0 : 1'b1;
												assign node340 = (inp[5]) ? node346 : node341;
													assign node341 = (inp[14]) ? node343 : 1'b0;
														assign node343 = (inp[4]) ? 1'b1 : 1'b0;
													assign node346 = (inp[2]) ? node352 : node347;
														assign node347 = (inp[11]) ? node349 : 1'b1;
															assign node349 = (inp[14]) ? 1'b0 : 1'b1;
														assign node352 = (inp[11]) ? 1'b1 : 1'b0;
											assign node355 = (inp[4]) ? node357 : 1'b0;
												assign node357 = (inp[11]) ? 1'b1 : node358;
													assign node358 = (inp[14]) ? 1'b0 : node359;
														assign node359 = (inp[13]) ? 1'b0 : 1'b1;
									assign node364 = (inp[0]) ? node366 : 1'b0;
										assign node366 = (inp[4]) ? 1'b0 : node367;
											assign node367 = (inp[5]) ? node375 : node368;
												assign node368 = (inp[11]) ? node370 : 1'b0;
													assign node370 = (inp[14]) ? node372 : 1'b1;
														assign node372 = (inp[2]) ? 1'b1 : 1'b0;
												assign node375 = (inp[11]) ? node377 : 1'b1;
													assign node377 = (inp[13]) ? 1'b1 : 1'b0;
							assign node381 = (inp[4]) ? node431 : node382;
								assign node382 = (inp[0]) ? node398 : node383;
									assign node383 = (inp[8]) ? 1'b1 : node384;
										assign node384 = (inp[1]) ? node386 : 1'b1;
											assign node386 = (inp[11]) ? node392 : node387;
												assign node387 = (inp[13]) ? 1'b1 : node388;
													assign node388 = (inp[2]) ? 1'b0 : 1'b1;
												assign node392 = (inp[2]) ? 1'b0 : node393;
													assign node393 = (inp[14]) ? 1'b1 : 1'b0;
									assign node398 = (inp[1]) ? node420 : node399;
										assign node399 = (inp[11]) ? node415 : node400;
											assign node400 = (inp[13]) ? node406 : node401;
												assign node401 = (inp[14]) ? node403 : 1'b0;
													assign node403 = (inp[2]) ? 1'b0 : 1'b1;
												assign node406 = (inp[8]) ? node408 : 1'b1;
													assign node408 = (inp[3]) ? node410 : 1'b0;
														assign node410 = (inp[5]) ? 1'b1 : node411;
															assign node411 = (inp[14]) ? 1'b0 : 1'b1;
											assign node415 = (inp[2]) ? 1'b0 : node416;
												assign node416 = (inp[14]) ? 1'b1 : 1'b0;
										assign node420 = (inp[8]) ? node422 : 1'b1;
											assign node422 = (inp[2]) ? node426 : node423;
												assign node423 = (inp[14]) ? 1'b1 : 1'b0;
												assign node426 = (inp[13]) ? node428 : 1'b0;
													assign node428 = (inp[11]) ? 1'b0 : 1'b1;
								assign node431 = (inp[8]) ? 1'b1 : node432;
									assign node432 = (inp[1]) ? node434 : 1'b1;
										assign node434 = (inp[11]) ? node452 : node435;
											assign node435 = (inp[5]) ? node445 : node436;
												assign node436 = (inp[14]) ? node438 : 1'b1;
													assign node438 = (inp[0]) ? 1'b0 : node439;
														assign node439 = (inp[13]) ? 1'b0 : node440;
															assign node440 = (inp[2]) ? 1'b0 : 1'b1;
												assign node445 = (inp[13]) ? 1'b1 : node446;
													assign node446 = (inp[14]) ? node448 : 1'b0;
														assign node448 = (inp[2]) ? 1'b0 : 1'b1;
											assign node452 = (inp[5]) ? node454 : 1'b0;
												assign node454 = (inp[13]) ? 1'b1 : 1'b0;
					assign node458 = (inp[3]) ? node552 : node459;
						assign node459 = (inp[0]) ? node481 : node460;
							assign node460 = (inp[1]) ? node462 : 1'b0;
								assign node462 = (inp[8]) ? 1'b0 : node463;
									assign node463 = (inp[11]) ? node475 : node464;
										assign node464 = (inp[13]) ? node470 : node465;
											assign node465 = (inp[2]) ? 1'b1 : node466;
												assign node466 = (inp[14]) ? 1'b0 : 1'b1;
											assign node470 = (inp[14]) ? node472 : 1'b0;
												assign node472 = (inp[2]) ? 1'b0 : 1'b1;
										assign node475 = (inp[14]) ? node477 : 1'b1;
											assign node477 = (inp[2]) ? 1'b1 : 1'b0;
							assign node481 = (inp[4]) ? node533 : node482;
								assign node482 = (inp[14]) ? node496 : node483;
									assign node483 = (inp[11]) ? node491 : node484;
										assign node484 = (inp[13]) ? 1'b0 : node485;
											assign node485 = (inp[1]) ? node487 : 1'b1;
												assign node487 = (inp[8]) ? 1'b1 : 1'b0;
										assign node491 = (inp[8]) ? 1'b1 : node492;
											assign node492 = (inp[1]) ? 1'b0 : 1'b1;
									assign node496 = (inp[8]) ? node522 : node497;
										assign node497 = (inp[1]) ? 1'b0 : node498;
											assign node498 = (inp[5]) ? node506 : node499;
												assign node499 = (inp[13]) ? node501 : 1'b0;
													assign node501 = (inp[2]) ? 1'b0 : node502;
														assign node502 = (inp[11]) ? 1'b0 : 1'b1;
												assign node506 = (inp[7]) ? node512 : node507;
													assign node507 = (inp[9]) ? node509 : 1'b1;
														assign node509 = (inp[2]) ? 1'b0 : 1'b1;
													assign node512 = (inp[11]) ? 1'b0 : node513;
														assign node513 = (inp[2]) ? node517 : node514;
															assign node514 = (inp[13]) ? 1'b1 : 1'b0;
															assign node517 = (inp[13]) ? 1'b0 : 1'b1;
										assign node522 = (inp[2]) ? node528 : node523;
											assign node523 = (inp[11]) ? 1'b0 : node524;
												assign node524 = (inp[13]) ? 1'b1 : 1'b0;
											assign node528 = (inp[13]) ? node530 : 1'b1;
												assign node530 = (inp[11]) ? 1'b1 : 1'b0;
								assign node533 = (inp[1]) ? node535 : 1'b0;
									assign node535 = (inp[8]) ? 1'b0 : node536;
										assign node536 = (inp[11]) ? node546 : node537;
											assign node537 = (inp[5]) ? node539 : 1'b0;
												assign node539 = (inp[13]) ? node543 : node540;
													assign node540 = (inp[2]) ? 1'b1 : 1'b0;
													assign node543 = (inp[2]) ? 1'b0 : 1'b1;
											assign node546 = (inp[2]) ? 1'b1 : node547;
												assign node547 = (inp[14]) ? 1'b0 : 1'b1;
						assign node552 = (inp[7]) ? node622 : node553;
							assign node553 = (inp[1]) ? node575 : node554;
								assign node554 = (inp[0]) ? node556 : 1'b1;
									assign node556 = (inp[4]) ? 1'b1 : node557;
										assign node557 = (inp[13]) ? node563 : node558;
											assign node558 = (inp[2]) ? 1'b0 : node559;
												assign node559 = (inp[14]) ? 1'b1 : 1'b0;
											assign node563 = (inp[11]) ? node569 : node564;
												assign node564 = (inp[14]) ? node566 : 1'b1;
													assign node566 = (inp[2]) ? 1'b1 : 1'b0;
												assign node569 = (inp[14]) ? node571 : 1'b0;
													assign node571 = (inp[2]) ? 1'b0 : 1'b1;
								assign node575 = (inp[8]) ? node605 : node576;
									assign node576 = (inp[0]) ? node592 : node577;
										assign node577 = (inp[11]) ? node587 : node578;
											assign node578 = (inp[14]) ? node582 : node579;
												assign node579 = (inp[13]) ? 1'b1 : 1'b0;
												assign node582 = (inp[13]) ? node584 : 1'b1;
													assign node584 = (inp[2]) ? 1'b1 : 1'b0;
											assign node587 = (inp[2]) ? 1'b0 : node588;
												assign node588 = (inp[14]) ? 1'b1 : 1'b0;
										assign node592 = (inp[4]) ? node594 : 1'b1;
											assign node594 = (inp[11]) ? node600 : node595;
												assign node595 = (inp[2]) ? node597 : 1'b1;
													assign node597 = (inp[13]) ? 1'b1 : 1'b0;
												assign node600 = (inp[2]) ? 1'b0 : node601;
													assign node601 = (inp[14]) ? 1'b1 : 1'b0;
									assign node605 = (inp[4]) ? 1'b1 : node606;
										assign node606 = (inp[0]) ? node608 : 1'b1;
											assign node608 = (inp[13]) ? node610 : 1'b0;
												assign node610 = (inp[11]) ? node616 : node611;
													assign node611 = (inp[5]) ? 1'b1 : node612;
														assign node612 = (inp[2]) ? 1'b1 : 1'b0;
													assign node616 = (inp[2]) ? 1'b0 : node617;
														assign node617 = (inp[14]) ? 1'b1 : 1'b0;
							assign node622 = (inp[1]) ? node646 : node623;
								assign node623 = (inp[4]) ? 1'b0 : node624;
									assign node624 = (inp[0]) ? node626 : 1'b0;
										assign node626 = (inp[2]) ? node638 : node627;
											assign node627 = (inp[14]) ? node633 : node628;
												assign node628 = (inp[13]) ? node630 : 1'b1;
													assign node630 = (inp[11]) ? 1'b1 : 1'b0;
												assign node633 = (inp[11]) ? 1'b0 : node634;
													assign node634 = (inp[13]) ? 1'b1 : 1'b0;
											assign node638 = (inp[9]) ? node640 : 1'b1;
												assign node640 = (inp[13]) ? node642 : 1'b1;
													assign node642 = (inp[11]) ? 1'b1 : 1'b0;
								assign node646 = (inp[8]) ? node684 : node647;
									assign node647 = (inp[0]) ? node665 : node648;
										assign node648 = (inp[14]) ? node654 : node649;
											assign node649 = (inp[13]) ? node651 : 1'b1;
												assign node651 = (inp[11]) ? 1'b1 : 1'b0;
											assign node654 = (inp[2]) ? node660 : node655;
												assign node655 = (inp[13]) ? node657 : 1'b0;
													assign node657 = (inp[11]) ? 1'b0 : 1'b1;
												assign node660 = (inp[13]) ? node662 : 1'b1;
													assign node662 = (inp[11]) ? 1'b1 : 1'b0;
										assign node665 = (inp[4]) ? node667 : 1'b0;
											assign node667 = (inp[11]) ? node679 : node668;
												assign node668 = (inp[13]) ? node674 : node669;
													assign node669 = (inp[9]) ? 1'b1 : node670;
														assign node670 = (inp[2]) ? 1'b1 : 1'b0;
													assign node674 = (inp[14]) ? node676 : 1'b0;
														assign node676 = (inp[2]) ? 1'b0 : 1'b1;
												assign node679 = (inp[14]) ? node681 : 1'b1;
													assign node681 = (inp[2]) ? 1'b1 : 1'b0;
									assign node684 = (inp[4]) ? 1'b0 : node685;
										assign node685 = (inp[0]) ? node687 : 1'b0;
											assign node687 = (inp[9]) ? node689 : 1'b1;
												assign node689 = (inp[13]) ? node695 : node690;
													assign node690 = (inp[14]) ? node692 : 1'b1;
														assign node692 = (inp[2]) ? 1'b1 : 1'b0;
													assign node695 = (inp[11]) ? node701 : node696;
														assign node696 = (inp[2]) ? 1'b0 : node697;
															assign node697 = (inp[14]) ? 1'b1 : 1'b0;
														assign node701 = (inp[5]) ? 1'b1 : 1'b0;
			assign node705 = (inp[0]) ? node727 : node706;
				assign node706 = (inp[1]) ? node708 : 1'b1;
					assign node708 = (inp[8]) ? 1'b1 : node709;
						assign node709 = (inp[11]) ? node721 : node710;
							assign node710 = (inp[13]) ? node716 : node711;
								assign node711 = (inp[2]) ? 1'b0 : node712;
									assign node712 = (inp[14]) ? 1'b1 : 1'b0;
								assign node716 = (inp[14]) ? node718 : 1'b1;
									assign node718 = (inp[2]) ? 1'b1 : 1'b0;
							assign node721 = (inp[14]) ? node723 : 1'b0;
								assign node723 = (inp[2]) ? 1'b0 : 1'b1;
				assign node727 = (inp[4]) ? node765 : node728;
					assign node728 = (inp[1]) ? node746 : node729;
						assign node729 = (inp[2]) ? node741 : node730;
							assign node730 = (inp[14]) ? node736 : node731;
								assign node731 = (inp[11]) ? 1'b0 : node732;
									assign node732 = (inp[13]) ? 1'b1 : 1'b0;
								assign node736 = (inp[11]) ? 1'b1 : node737;
									assign node737 = (inp[13]) ? 1'b0 : 1'b1;
							assign node741 = (inp[11]) ? 1'b0 : node742;
								assign node742 = (inp[13]) ? 1'b1 : 1'b0;
						assign node746 = (inp[8]) ? node748 : 1'b1;
							assign node748 = (inp[2]) ? node760 : node749;
								assign node749 = (inp[14]) ? node755 : node750;
									assign node750 = (inp[11]) ? 1'b0 : node751;
										assign node751 = (inp[13]) ? 1'b1 : 1'b0;
									assign node755 = (inp[13]) ? node757 : 1'b1;
										assign node757 = (inp[11]) ? 1'b1 : 1'b0;
								assign node760 = (inp[13]) ? node762 : 1'b0;
									assign node762 = (inp[11]) ? 1'b0 : 1'b1;
					assign node765 = (inp[8]) ? 1'b1 : node766;
						assign node766 = (inp[1]) ? node768 : 1'b1;
							assign node768 = (inp[11]) ? node780 : node769;
								assign node769 = (inp[13]) ? node775 : node770;
									assign node770 = (inp[14]) ? node772 : 1'b0;
										assign node772 = (inp[2]) ? 1'b0 : 1'b1;
									assign node775 = (inp[2]) ? 1'b1 : node776;
										assign node776 = (inp[14]) ? 1'b0 : 1'b1;
								assign node780 = (inp[14]) ? node782 : 1'b0;
									assign node782 = (inp[2]) ? 1'b0 : 1'b1;
		assign node786 = (inp[5]) ? node1926 : node787;
			assign node787 = (inp[12]) ? node1405 : node788;
				assign node788 = (inp[10]) ? node1174 : node789;
					assign node789 = (inp[9]) ? node995 : node790;
						assign node790 = (inp[3]) ? node876 : node791;
							assign node791 = (inp[0]) ? node809 : node792;
								assign node792 = (inp[1]) ? node794 : 1'b0;
									assign node794 = (inp[8]) ? 1'b0 : node795;
										assign node795 = (inp[14]) ? node801 : node796;
											assign node796 = (inp[11]) ? 1'b1 : node797;
												assign node797 = (inp[13]) ? 1'b0 : 1'b1;
											assign node801 = (inp[2]) ? 1'b1 : node802;
												assign node802 = (inp[13]) ? node804 : 1'b0;
													assign node804 = (inp[15]) ? 1'b0 : 1'b1;
								assign node809 = (inp[13]) ? node835 : node810;
									assign node810 = (inp[4]) ? node826 : node811;
										assign node811 = (inp[1]) ? node819 : node812;
											assign node812 = (inp[7]) ? 1'b1 : node813;
												assign node813 = (inp[14]) ? node815 : 1'b1;
													assign node815 = (inp[11]) ? 1'b0 : 1'b1;
											assign node819 = (inp[8]) ? node821 : 1'b0;
												assign node821 = (inp[14]) ? node823 : 1'b1;
													assign node823 = (inp[2]) ? 1'b1 : 1'b0;
										assign node826 = (inp[1]) ? node828 : 1'b0;
											assign node828 = (inp[8]) ? 1'b0 : node829;
												assign node829 = (inp[14]) ? node831 : 1'b1;
													assign node831 = (inp[15]) ? 1'b1 : 1'b0;
									assign node835 = (inp[11]) ? node845 : node836;
										assign node836 = (inp[14]) ? node838 : 1'b0;
											assign node838 = (inp[2]) ? 1'b0 : node839;
												assign node839 = (inp[1]) ? 1'b0 : node840;
													assign node840 = (inp[4]) ? 1'b0 : 1'b1;
										assign node845 = (inp[14]) ? node863 : node846;
											assign node846 = (inp[2]) ? node854 : node847;
												assign node847 = (inp[15]) ? node849 : 1'b1;
													assign node849 = (inp[1]) ? node851 : 1'b1;
														assign node851 = (inp[8]) ? 1'b1 : 1'b0;
												assign node854 = (inp[15]) ? node856 : 1'b0;
													assign node856 = (inp[4]) ? node860 : node857;
														assign node857 = (inp[7]) ? 1'b1 : 1'b0;
														assign node860 = (inp[8]) ? 1'b0 : 1'b1;
											assign node863 = (inp[2]) ? node865 : 1'b0;
												assign node865 = (inp[4]) ? node871 : node866;
													assign node866 = (inp[8]) ? 1'b1 : node867;
														assign node867 = (inp[1]) ? 1'b0 : 1'b1;
													assign node871 = (inp[8]) ? 1'b0 : node872;
														assign node872 = (inp[1]) ? 1'b1 : 1'b0;
							assign node876 = (inp[7]) ? node940 : node877;
								assign node877 = (inp[2]) ? node909 : node878;
									assign node878 = (inp[0]) ? node890 : node879;
										assign node879 = (inp[4]) ? 1'b1 : node880;
											assign node880 = (inp[15]) ? node882 : 1'b1;
												assign node882 = (inp[11]) ? 1'b1 : node883;
													assign node883 = (inp[13]) ? 1'b1 : node884;
														assign node884 = (inp[14]) ? 1'b1 : 1'b0;
										assign node890 = (inp[1]) ? node896 : node891;
											assign node891 = (inp[15]) ? node893 : 1'b1;
												assign node893 = (inp[8]) ? 1'b0 : 1'b1;
											assign node896 = (inp[15]) ? node904 : node897;
												assign node897 = (inp[8]) ? node901 : node898;
													assign node898 = (inp[4]) ? 1'b0 : 1'b1;
													assign node901 = (inp[4]) ? 1'b1 : 1'b0;
												assign node904 = (inp[14]) ? node906 : 1'b1;
													assign node906 = (inp[8]) ? 1'b0 : 1'b1;
									assign node909 = (inp[8]) ? node931 : node910;
										assign node910 = (inp[1]) ? node916 : node911;
											assign node911 = (inp[0]) ? node913 : 1'b1;
												assign node913 = (inp[4]) ? 1'b1 : 1'b0;
											assign node916 = (inp[0]) ? node924 : node917;
												assign node917 = (inp[14]) ? node919 : 1'b0;
													assign node919 = (inp[11]) ? 1'b0 : node920;
														assign node920 = (inp[13]) ? 1'b1 : 1'b0;
												assign node924 = (inp[4]) ? node926 : 1'b1;
													assign node926 = (inp[14]) ? 1'b0 : node927;
														assign node927 = (inp[13]) ? 1'b1 : 1'b0;
										assign node931 = (inp[4]) ? 1'b1 : node932;
											assign node932 = (inp[0]) ? node934 : 1'b1;
												assign node934 = (inp[13]) ? node936 : 1'b0;
													assign node936 = (inp[11]) ? 1'b0 : 1'b1;
								assign node940 = (inp[8]) ? node976 : node941;
									assign node941 = (inp[1]) ? node955 : node942;
										assign node942 = (inp[4]) ? 1'b0 : node943;
											assign node943 = (inp[0]) ? node945 : 1'b0;
												assign node945 = (inp[15]) ? node951 : node946;
													assign node946 = (inp[14]) ? node948 : 1'b1;
														assign node948 = (inp[2]) ? 1'b1 : 1'b0;
													assign node951 = (inp[14]) ? 1'b1 : 1'b0;
										assign node955 = (inp[0]) ? node969 : node956;
											assign node956 = (inp[14]) ? node962 : node957;
												assign node957 = (inp[13]) ? node959 : 1'b1;
													assign node959 = (inp[11]) ? 1'b1 : 1'b0;
												assign node962 = (inp[2]) ? node966 : node963;
													assign node963 = (inp[4]) ? 1'b0 : 1'b1;
													assign node966 = (inp[4]) ? 1'b1 : 1'b0;
											assign node969 = (inp[4]) ? node971 : 1'b0;
												assign node971 = (inp[15]) ? 1'b1 : node972;
													assign node972 = (inp[11]) ? 1'b1 : 1'b0;
									assign node976 = (inp[4]) ? 1'b0 : node977;
										assign node977 = (inp[0]) ? node979 : 1'b0;
											assign node979 = (inp[2]) ? node989 : node980;
												assign node980 = (inp[15]) ? node984 : node981;
													assign node981 = (inp[14]) ? 1'b0 : 1'b1;
													assign node984 = (inp[1]) ? node986 : 1'b0;
														assign node986 = (inp[13]) ? 1'b1 : 1'b0;
												assign node989 = (inp[11]) ? 1'b1 : node990;
													assign node990 = (inp[13]) ? 1'b0 : 1'b1;
						assign node995 = (inp[7]) ? node1099 : node996;
							assign node996 = (inp[3]) ? node1054 : node997;
								assign node997 = (inp[1]) ? node1015 : node998;
									assign node998 = (inp[0]) ? node1000 : 1'b1;
										assign node1000 = (inp[4]) ? 1'b1 : node1001;
											assign node1001 = (inp[13]) ? node1007 : node1002;
												assign node1002 = (inp[11]) ? node1004 : 1'b0;
													assign node1004 = (inp[14]) ? 1'b1 : 1'b0;
												assign node1007 = (inp[14]) ? node1009 : 1'b1;
													assign node1009 = (inp[11]) ? node1011 : 1'b0;
														assign node1011 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1015 = (inp[8]) ? node1043 : node1016;
										assign node1016 = (inp[4]) ? node1030 : node1017;
											assign node1017 = (inp[0]) ? 1'b1 : node1018;
												assign node1018 = (inp[11]) ? 1'b0 : node1019;
													assign node1019 = (inp[15]) ? node1021 : 1'b1;
														assign node1021 = (inp[13]) ? node1025 : node1022;
															assign node1022 = (inp[14]) ? 1'b1 : 1'b0;
															assign node1025 = (inp[14]) ? 1'b0 : 1'b1;
											assign node1030 = (inp[13]) ? node1036 : node1031;
												assign node1031 = (inp[14]) ? node1033 : 1'b0;
													assign node1033 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1036 = (inp[11]) ? node1040 : node1037;
													assign node1037 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1040 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1043 = (inp[0]) ? node1045 : 1'b1;
											assign node1045 = (inp[4]) ? 1'b1 : node1046;
												assign node1046 = (inp[11]) ? node1050 : node1047;
													assign node1047 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1050 = (inp[14]) ? 1'b1 : 1'b0;
								assign node1054 = (inp[1]) ? node1068 : node1055;
									assign node1055 = (inp[4]) ? 1'b0 : node1056;
										assign node1056 = (inp[0]) ? node1058 : 1'b0;
											assign node1058 = (inp[11]) ? node1062 : node1059;
												assign node1059 = (inp[15]) ? 1'b1 : 1'b0;
												assign node1062 = (inp[14]) ? node1064 : 1'b1;
													assign node1064 = (inp[2]) ? 1'b1 : 1'b0;
									assign node1068 = (inp[14]) ? node1082 : node1069;
										assign node1069 = (inp[8]) ? node1077 : node1070;
											assign node1070 = (inp[4]) ? 1'b1 : node1071;
												assign node1071 = (inp[0]) ? 1'b0 : node1072;
													assign node1072 = (inp[13]) ? 1'b0 : 1'b1;
											assign node1077 = (inp[0]) ? node1079 : 1'b0;
												assign node1079 = (inp[4]) ? 1'b0 : 1'b1;
										assign node1082 = (inp[2]) ? node1084 : 1'b0;
											assign node1084 = (inp[11]) ? node1088 : node1085;
												assign node1085 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1088 = (inp[13]) ? node1090 : 1'b0;
													assign node1090 = (inp[8]) ? node1094 : node1091;
														assign node1091 = (inp[0]) ? 1'b0 : 1'b1;
														assign node1094 = (inp[15]) ? node1096 : 1'b0;
															assign node1096 = (inp[0]) ? 1'b1 : 1'b0;
							assign node1099 = (inp[8]) ? node1155 : node1100;
								assign node1100 = (inp[1]) ? node1116 : node1101;
									assign node1101 = (inp[4]) ? 1'b1 : node1102;
										assign node1102 = (inp[0]) ? node1104 : 1'b1;
											assign node1104 = (inp[11]) ? node1110 : node1105;
												assign node1105 = (inp[13]) ? 1'b1 : node1106;
													assign node1106 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1110 = (inp[14]) ? node1112 : 1'b0;
													assign node1112 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1116 = (inp[4]) ? node1130 : node1117;
										assign node1117 = (inp[0]) ? 1'b1 : node1118;
											assign node1118 = (inp[2]) ? node1124 : node1119;
												assign node1119 = (inp[15]) ? node1121 : 1'b1;
													assign node1121 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1124 = (inp[11]) ? 1'b0 : node1125;
													assign node1125 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1130 = (inp[2]) ? node1150 : node1131;
											assign node1131 = (inp[0]) ? node1141 : node1132;
												assign node1132 = (inp[3]) ? 1'b1 : node1133;
													assign node1133 = (inp[14]) ? node1135 : 1'b0;
														assign node1135 = (inp[15]) ? node1137 : 1'b1;
															assign node1137 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1141 = (inp[13]) ? node1143 : 1'b0;
													assign node1143 = (inp[14]) ? node1147 : node1144;
														assign node1144 = (inp[11]) ? 1'b0 : 1'b1;
														assign node1147 = (inp[11]) ? 1'b1 : 1'b0;
											assign node1150 = (inp[13]) ? node1152 : 1'b0;
												assign node1152 = (inp[0]) ? 1'b1 : 1'b0;
								assign node1155 = (inp[4]) ? 1'b1 : node1156;
									assign node1156 = (inp[0]) ? node1158 : 1'b1;
										assign node1158 = (inp[14]) ? node1164 : node1159;
											assign node1159 = (inp[13]) ? node1161 : 1'b0;
												assign node1161 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1164 = (inp[2]) ? node1170 : node1165;
												assign node1165 = (inp[11]) ? 1'b1 : node1166;
													assign node1166 = (inp[15]) ? 1'b1 : 1'b0;
												assign node1170 = (inp[11]) ? 1'b0 : 1'b1;
					assign node1174 = (inp[3]) ? node1254 : node1175;
						assign node1175 = (inp[4]) ? node1233 : node1176;
							assign node1176 = (inp[0]) ? node1200 : node1177;
								assign node1177 = (inp[8]) ? 1'b0 : node1178;
									assign node1178 = (inp[1]) ? node1180 : 1'b0;
										assign node1180 = (inp[2]) ? node1192 : node1181;
											assign node1181 = (inp[14]) ? node1187 : node1182;
												assign node1182 = (inp[11]) ? 1'b1 : node1183;
													assign node1183 = (inp[13]) ? 1'b0 : 1'b1;
												assign node1187 = (inp[13]) ? node1189 : 1'b0;
													assign node1189 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1192 = (inp[15]) ? 1'b1 : node1193;
												assign node1193 = (inp[13]) ? node1195 : 1'b1;
													assign node1195 = (inp[11]) ? 1'b1 : 1'b0;
								assign node1200 = (inp[8]) ? node1216 : node1201;
									assign node1201 = (inp[1]) ? 1'b0 : node1202;
										assign node1202 = (inp[2]) ? node1210 : node1203;
											assign node1203 = (inp[14]) ? 1'b0 : node1204;
												assign node1204 = (inp[13]) ? node1206 : 1'b1;
													assign node1206 = (inp[11]) ? 1'b1 : 1'b0;
											assign node1210 = (inp[13]) ? node1212 : 1'b1;
												assign node1212 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1216 = (inp[14]) ? node1222 : node1217;
										assign node1217 = (inp[13]) ? node1219 : 1'b1;
											assign node1219 = (inp[11]) ? 1'b1 : 1'b0;
										assign node1222 = (inp[13]) ? node1226 : node1223;
											assign node1223 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1226 = (inp[2]) ? node1230 : node1227;
												assign node1227 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1230 = (inp[11]) ? 1'b1 : 1'b0;
							assign node1233 = (inp[8]) ? 1'b0 : node1234;
								assign node1234 = (inp[1]) ? node1236 : 1'b0;
									assign node1236 = (inp[14]) ? node1242 : node1237;
										assign node1237 = (inp[11]) ? 1'b1 : node1238;
											assign node1238 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1242 = (inp[2]) ? node1248 : node1243;
											assign node1243 = (inp[11]) ? 1'b0 : node1244;
												assign node1244 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1248 = (inp[13]) ? node1250 : 1'b1;
												assign node1250 = (inp[11]) ? 1'b1 : 1'b0;
						assign node1254 = (inp[7]) ? node1340 : node1255;
							assign node1255 = (inp[0]) ? node1275 : node1256;
								assign node1256 = (inp[8]) ? 1'b1 : node1257;
									assign node1257 = (inp[1]) ? node1259 : 1'b1;
										assign node1259 = (inp[11]) ? node1269 : node1260;
											assign node1260 = (inp[13]) ? node1264 : node1261;
												assign node1261 = (inp[4]) ? 1'b1 : 1'b0;
												assign node1264 = (inp[14]) ? node1266 : 1'b1;
													assign node1266 = (inp[15]) ? 1'b1 : 1'b0;
											assign node1269 = (inp[14]) ? node1271 : 1'b0;
												assign node1271 = (inp[2]) ? 1'b0 : 1'b1;
								assign node1275 = (inp[4]) ? node1313 : node1276;
									assign node1276 = (inp[1]) ? node1298 : node1277;
										assign node1277 = (inp[13]) ? node1283 : node1278;
											assign node1278 = (inp[14]) ? node1280 : 1'b0;
												assign node1280 = (inp[2]) ? 1'b0 : 1'b1;
											assign node1283 = (inp[2]) ? node1295 : node1284;
												assign node1284 = (inp[8]) ? node1290 : node1285;
													assign node1285 = (inp[15]) ? node1287 : 1'b1;
														assign node1287 = (inp[14]) ? 1'b1 : 1'b0;
													assign node1290 = (inp[11]) ? 1'b1 : node1291;
														assign node1291 = (inp[14]) ? 1'b0 : 1'b1;
												assign node1295 = (inp[11]) ? 1'b0 : 1'b1;
										assign node1298 = (inp[8]) ? node1300 : 1'b1;
											assign node1300 = (inp[2]) ? node1308 : node1301;
												assign node1301 = (inp[14]) ? node1305 : node1302;
													assign node1302 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1305 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1308 = (inp[14]) ? 1'b0 : node1309;
													assign node1309 = (inp[15]) ? 1'b1 : 1'b0;
									assign node1313 = (inp[1]) ? node1315 : 1'b1;
										assign node1315 = (inp[8]) ? 1'b1 : node1316;
											assign node1316 = (inp[11]) ? node1334 : node1317;
												assign node1317 = (inp[9]) ? node1325 : node1318;
													assign node1318 = (inp[15]) ? node1320 : 1'b1;
														assign node1320 = (inp[2]) ? 1'b1 : node1321;
															assign node1321 = (inp[14]) ? 1'b0 : 1'b0;
													assign node1325 = (inp[13]) ? node1331 : node1326;
														assign node1326 = (inp[14]) ? node1328 : 1'b0;
															assign node1328 = (inp[2]) ? 1'b0 : 1'b1;
														assign node1331 = (inp[2]) ? 1'b1 : 1'b0;
												assign node1334 = (inp[14]) ? node1336 : 1'b0;
													assign node1336 = (inp[2]) ? 1'b0 : 1'b1;
							assign node1340 = (inp[0]) ? node1360 : node1341;
								assign node1341 = (inp[1]) ? node1343 : 1'b0;
									assign node1343 = (inp[8]) ? 1'b0 : node1344;
										assign node1344 = (inp[2]) ? node1354 : node1345;
											assign node1345 = (inp[14]) ? node1349 : node1346;
												assign node1346 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1349 = (inp[11]) ? 1'b0 : node1350;
													assign node1350 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1354 = (inp[11]) ? 1'b1 : node1355;
												assign node1355 = (inp[13]) ? 1'b0 : 1'b1;
								assign node1360 = (inp[4]) ? node1390 : node1361;
									assign node1361 = (inp[2]) ? node1377 : node1362;
										assign node1362 = (inp[1]) ? node1372 : node1363;
											assign node1363 = (inp[11]) ? 1'b1 : node1364;
												assign node1364 = (inp[13]) ? node1368 : node1365;
													assign node1365 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1368 = (inp[14]) ? 1'b1 : 1'b0;
											assign node1372 = (inp[15]) ? 1'b0 : node1373;
												assign node1373 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1377 = (inp[8]) ? node1385 : node1378;
											assign node1378 = (inp[1]) ? 1'b0 : node1379;
												assign node1379 = (inp[13]) ? node1381 : 1'b1;
													assign node1381 = (inp[11]) ? 1'b1 : 1'b0;
											assign node1385 = (inp[13]) ? node1387 : 1'b1;
												assign node1387 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1390 = (inp[8]) ? 1'b0 : node1391;
										assign node1391 = (inp[1]) ? node1393 : 1'b0;
											assign node1393 = (inp[9]) ? node1395 : 1'b1;
												assign node1395 = (inp[14]) ? node1401 : node1396;
													assign node1396 = (inp[11]) ? 1'b1 : node1397;
														assign node1397 = (inp[13]) ? 1'b0 : 1'b1;
													assign node1401 = (inp[11]) ? 1'b0 : 1'b1;
				assign node1405 = (inp[15]) ? node1485 : node1406;
					assign node1406 = (inp[0]) ? node1428 : node1407;
						assign node1407 = (inp[8]) ? 1'b1 : node1408;
							assign node1408 = (inp[1]) ? node1410 : 1'b1;
								assign node1410 = (inp[2]) ? node1422 : node1411;
									assign node1411 = (inp[14]) ? node1417 : node1412;
										assign node1412 = (inp[11]) ? 1'b0 : node1413;
											assign node1413 = (inp[13]) ? 1'b1 : 1'b0;
										assign node1417 = (inp[13]) ? node1419 : 1'b1;
											assign node1419 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1422 = (inp[11]) ? 1'b0 : node1423;
										assign node1423 = (inp[13]) ? 1'b1 : 1'b0;
						assign node1428 = (inp[4]) ? node1464 : node1429;
							assign node1429 = (inp[8]) ? node1447 : node1430;
								assign node1430 = (inp[1]) ? 1'b1 : node1431;
									assign node1431 = (inp[2]) ? node1441 : node1432;
										assign node1432 = (inp[14]) ? node1436 : node1433;
											assign node1433 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1436 = (inp[11]) ? 1'b1 : node1437;
												assign node1437 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1441 = (inp[11]) ? 1'b0 : node1442;
											assign node1442 = (inp[13]) ? 1'b1 : 1'b0;
								assign node1447 = (inp[14]) ? node1453 : node1448;
									assign node1448 = (inp[13]) ? node1450 : 1'b0;
										assign node1450 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1453 = (inp[2]) ? node1459 : node1454;
										assign node1454 = (inp[13]) ? node1456 : 1'b1;
											assign node1456 = (inp[11]) ? 1'b1 : 1'b0;
										assign node1459 = (inp[13]) ? node1461 : 1'b0;
											assign node1461 = (inp[11]) ? 1'b0 : 1'b1;
							assign node1464 = (inp[1]) ? node1466 : 1'b1;
								assign node1466 = (inp[8]) ? 1'b1 : node1467;
									assign node1467 = (inp[2]) ? node1479 : node1468;
										assign node1468 = (inp[14]) ? node1474 : node1469;
											assign node1469 = (inp[11]) ? 1'b0 : node1470;
												assign node1470 = (inp[13]) ? 1'b1 : 1'b0;
											assign node1474 = (inp[11]) ? 1'b1 : node1475;
												assign node1475 = (inp[13]) ? 1'b0 : 1'b1;
										assign node1479 = (inp[11]) ? 1'b0 : node1480;
											assign node1480 = (inp[13]) ? 1'b1 : 1'b0;
					assign node1485 = (inp[10]) ? node1747 : node1486;
						assign node1486 = (inp[9]) ? node1620 : node1487;
							assign node1487 = (inp[7]) ? node1571 : node1488;
								assign node1488 = (inp[3]) ? node1520 : node1489;
									assign node1489 = (inp[0]) ? node1497 : node1490;
										assign node1490 = (inp[1]) ? node1492 : 1'b0;
											assign node1492 = (inp[13]) ? 1'b0 : node1493;
												assign node1493 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1497 = (inp[11]) ? node1507 : node1498;
											assign node1498 = (inp[14]) ? node1504 : node1499;
												assign node1499 = (inp[13]) ? 1'b0 : node1500;
													assign node1500 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1504 = (inp[8]) ? 1'b0 : 1'b1;
											assign node1507 = (inp[8]) ? node1517 : node1508;
												assign node1508 = (inp[1]) ? node1514 : node1509;
													assign node1509 = (inp[4]) ? 1'b0 : node1510;
														assign node1510 = (inp[14]) ? 1'b0 : 1'b1;
													assign node1514 = (inp[4]) ? 1'b1 : 1'b0;
												assign node1517 = (inp[4]) ? 1'b0 : 1'b1;
									assign node1520 = (inp[14]) ? node1544 : node1521;
										assign node1521 = (inp[4]) ? node1539 : node1522;
											assign node1522 = (inp[2]) ? node1534 : node1523;
												assign node1523 = (inp[8]) ? node1529 : node1524;
													assign node1524 = (inp[1]) ? 1'b1 : node1525;
														assign node1525 = (inp[0]) ? 1'b0 : 1'b1;
													assign node1529 = (inp[1]) ? node1531 : 1'b0;
														assign node1531 = (inp[13]) ? 1'b1 : 1'b0;
												assign node1534 = (inp[0]) ? 1'b0 : node1535;
													assign node1535 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1539 = (inp[1]) ? node1541 : 1'b1;
												assign node1541 = (inp[8]) ? 1'b1 : 1'b0;
										assign node1544 = (inp[11]) ? node1560 : node1545;
											assign node1545 = (inp[8]) ? node1555 : node1546;
												assign node1546 = (inp[0]) ? node1548 : 1'b0;
													assign node1548 = (inp[13]) ? node1550 : 1'b1;
														assign node1550 = (inp[2]) ? 1'b1 : node1551;
															assign node1551 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1555 = (inp[0]) ? node1557 : 1'b1;
													assign node1557 = (inp[4]) ? 1'b1 : 1'b0;
											assign node1560 = (inp[13]) ? node1562 : 1'b1;
												assign node1562 = (inp[2]) ? node1564 : 1'b1;
													assign node1564 = (inp[4]) ? node1566 : 1'b1;
														assign node1566 = (inp[8]) ? 1'b1 : node1567;
															assign node1567 = (inp[0]) ? 1'b0 : 1'b1;
								assign node1571 = (inp[0]) ? node1583 : node1572;
									assign node1572 = (inp[1]) ? node1574 : 1'b0;
										assign node1574 = (inp[8]) ? 1'b0 : node1575;
											assign node1575 = (inp[2]) ? 1'b1 : node1576;
												assign node1576 = (inp[14]) ? 1'b0 : node1577;
													assign node1577 = (inp[11]) ? 1'b1 : 1'b0;
									assign node1583 = (inp[13]) ? node1597 : node1584;
										assign node1584 = (inp[4]) ? node1592 : node1585;
											assign node1585 = (inp[14]) ? node1587 : 1'b1;
												assign node1587 = (inp[2]) ? node1589 : 1'b0;
													assign node1589 = (inp[1]) ? 1'b0 : 1'b1;
											assign node1592 = (inp[2]) ? node1594 : 1'b0;
												assign node1594 = (inp[1]) ? 1'b1 : 1'b0;
										assign node1597 = (inp[3]) ? node1611 : node1598;
											assign node1598 = (inp[11]) ? node1604 : node1599;
												assign node1599 = (inp[14]) ? node1601 : 1'b0;
													assign node1601 = (inp[8]) ? 1'b0 : 1'b1;
												assign node1604 = (inp[4]) ? node1608 : node1605;
													assign node1605 = (inp[8]) ? 1'b1 : 1'b0;
													assign node1608 = (inp[1]) ? 1'b1 : 1'b0;
											assign node1611 = (inp[1]) ? node1613 : 1'b0;
												assign node1613 = (inp[14]) ? 1'b0 : node1614;
													assign node1614 = (inp[4]) ? node1616 : 1'b0;
														assign node1616 = (inp[8]) ? 1'b0 : 1'b1;
							assign node1620 = (inp[7]) ? node1678 : node1621;
								assign node1621 = (inp[3]) ? node1647 : node1622;
									assign node1622 = (inp[2]) ? node1630 : node1623;
										assign node1623 = (inp[0]) ? node1625 : 1'b1;
											assign node1625 = (inp[14]) ? 1'b1 : node1626;
												assign node1626 = (inp[13]) ? 1'b1 : 1'b0;
										assign node1630 = (inp[13]) ? node1640 : node1631;
											assign node1631 = (inp[8]) ? node1635 : node1632;
												assign node1632 = (inp[1]) ? 1'b0 : 1'b1;
												assign node1635 = (inp[0]) ? node1637 : 1'b1;
													assign node1637 = (inp[4]) ? 1'b1 : 1'b0;
											assign node1640 = (inp[8]) ? node1642 : 1'b1;
												assign node1642 = (inp[0]) ? node1644 : 1'b1;
													assign node1644 = (inp[4]) ? 1'b1 : 1'b0;
									assign node1647 = (inp[1]) ? node1653 : node1648;
										assign node1648 = (inp[4]) ? 1'b0 : node1649;
											assign node1649 = (inp[0]) ? 1'b1 : 1'b0;
										assign node1653 = (inp[8]) ? node1669 : node1654;
											assign node1654 = (inp[0]) ? node1660 : node1655;
												assign node1655 = (inp[13]) ? node1657 : 1'b1;
													assign node1657 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1660 = (inp[4]) ? node1662 : 1'b0;
													assign node1662 = (inp[2]) ? 1'b1 : node1663;
														assign node1663 = (inp[14]) ? 1'b0 : node1664;
															assign node1664 = (inp[11]) ? 1'b1 : 1'b0;
											assign node1669 = (inp[4]) ? 1'b0 : node1670;
												assign node1670 = (inp[0]) ? node1672 : 1'b0;
													assign node1672 = (inp[13]) ? 1'b1 : node1673;
														assign node1673 = (inp[2]) ? 1'b1 : 1'b0;
								assign node1678 = (inp[1]) ? node1702 : node1679;
									assign node1679 = (inp[0]) ? node1681 : 1'b1;
										assign node1681 = (inp[4]) ? 1'b1 : node1682;
											assign node1682 = (inp[13]) ? node1688 : node1683;
												assign node1683 = (inp[14]) ? node1685 : 1'b0;
													assign node1685 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1688 = (inp[3]) ? node1696 : node1689;
													assign node1689 = (inp[14]) ? node1691 : 1'b1;
														assign node1691 = (inp[2]) ? node1693 : 1'b0;
															assign node1693 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1696 = (inp[2]) ? node1698 : 1'b1;
														assign node1698 = (inp[11]) ? 1'b0 : 1'b1;
									assign node1702 = (inp[2]) ? node1728 : node1703;
										assign node1703 = (inp[3]) ? node1715 : node1704;
											assign node1704 = (inp[11]) ? node1706 : 1'b1;
												assign node1706 = (inp[14]) ? 1'b1 : node1707;
													assign node1707 = (inp[8]) ? node1711 : node1708;
														assign node1708 = (inp[0]) ? 1'b1 : 1'b0;
														assign node1711 = (inp[4]) ? 1'b1 : 1'b0;
											assign node1715 = (inp[14]) ? node1723 : node1716;
												assign node1716 = (inp[8]) ? node1718 : 1'b0;
													assign node1718 = (inp[0]) ? node1720 : 1'b1;
														assign node1720 = (inp[11]) ? 1'b0 : 1'b1;
												assign node1723 = (inp[13]) ? node1725 : 1'b1;
													assign node1725 = (inp[11]) ? 1'b1 : 1'b0;
										assign node1728 = (inp[8]) ? node1742 : node1729;
											assign node1729 = (inp[11]) ? node1737 : node1730;
												assign node1730 = (inp[13]) ? 1'b1 : node1731;
													assign node1731 = (inp[0]) ? node1733 : 1'b0;
														assign node1733 = (inp[4]) ? 1'b0 : 1'b1;
												assign node1737 = (inp[14]) ? 1'b0 : node1738;
													assign node1738 = (inp[4]) ? 1'b0 : 1'b1;
											assign node1742 = (inp[0]) ? node1744 : 1'b1;
												assign node1744 = (inp[4]) ? 1'b1 : 1'b0;
						assign node1747 = (inp[7]) ? node1857 : node1748;
							assign node1748 = (inp[3]) ? node1806 : node1749;
								assign node1749 = (inp[13]) ? node1777 : node1750;
									assign node1750 = (inp[14]) ? node1768 : node1751;
										assign node1751 = (inp[4]) ? node1763 : node1752;
											assign node1752 = (inp[0]) ? node1758 : node1753;
												assign node1753 = (inp[1]) ? node1755 : 1'b0;
													assign node1755 = (inp[8]) ? 1'b0 : 1'b1;
												assign node1758 = (inp[1]) ? node1760 : 1'b1;
													assign node1760 = (inp[8]) ? 1'b1 : 1'b0;
											assign node1763 = (inp[1]) ? node1765 : 1'b0;
												assign node1765 = (inp[8]) ? 1'b0 : 1'b1;
										assign node1768 = (inp[0]) ? node1770 : 1'b0;
											assign node1770 = (inp[11]) ? 1'b1 : node1771;
												assign node1771 = (inp[4]) ? 1'b0 : node1772;
													assign node1772 = (inp[9]) ? 1'b1 : 1'b0;
									assign node1777 = (inp[1]) ? node1779 : 1'b0;
										assign node1779 = (inp[11]) ? node1789 : node1780;
											assign node1780 = (inp[8]) ? 1'b0 : node1781;
												assign node1781 = (inp[2]) ? 1'b0 : node1782;
													assign node1782 = (inp[4]) ? node1784 : 1'b0;
														assign node1784 = (inp[14]) ? 1'b1 : 1'b0;
											assign node1789 = (inp[2]) ? node1795 : node1790;
												assign node1790 = (inp[4]) ? 1'b0 : node1791;
													assign node1791 = (inp[8]) ? 1'b1 : 1'b0;
												assign node1795 = (inp[8]) ? node1801 : node1796;
													assign node1796 = (inp[0]) ? node1798 : 1'b1;
														assign node1798 = (inp[4]) ? 1'b1 : 1'b0;
													assign node1801 = (inp[0]) ? node1803 : 1'b0;
														assign node1803 = (inp[4]) ? 1'b0 : 1'b1;
								assign node1806 = (inp[0]) ? node1824 : node1807;
									assign node1807 = (inp[1]) ? node1809 : 1'b1;
										assign node1809 = (inp[8]) ? 1'b1 : node1810;
											assign node1810 = (inp[11]) ? node1818 : node1811;
												assign node1811 = (inp[13]) ? 1'b1 : node1812;
													assign node1812 = (inp[4]) ? 1'b0 : node1813;
														assign node1813 = (inp[2]) ? 1'b0 : 1'b1;
												assign node1818 = (inp[2]) ? 1'b0 : node1819;
													assign node1819 = (inp[14]) ? 1'b1 : 1'b0;
									assign node1824 = (inp[4]) ? node1844 : node1825;
										assign node1825 = (inp[8]) ? node1833 : node1826;
											assign node1826 = (inp[1]) ? 1'b1 : node1827;
												assign node1827 = (inp[13]) ? node1829 : 1'b0;
													assign node1829 = (inp[11]) ? 1'b0 : 1'b1;
											assign node1833 = (inp[1]) ? node1835 : 1'b0;
												assign node1835 = (inp[14]) ? node1841 : node1836;
													assign node1836 = (inp[11]) ? 1'b0 : node1837;
														assign node1837 = (inp[13]) ? 1'b1 : 1'b0;
													assign node1841 = (inp[2]) ? 1'b0 : 1'b1;
										assign node1844 = (inp[8]) ? 1'b1 : node1845;
											assign node1845 = (inp[1]) ? node1847 : 1'b1;
												assign node1847 = (inp[9]) ? 1'b0 : node1848;
													assign node1848 = (inp[2]) ? node1850 : 1'b1;
														assign node1850 = (inp[14]) ? 1'b0 : node1851;
															assign node1851 = (inp[11]) ? 1'b0 : 1'b1;
							assign node1857 = (inp[1]) ? node1875 : node1858;
								assign node1858 = (inp[0]) ? node1860 : 1'b0;
									assign node1860 = (inp[4]) ? 1'b0 : node1861;
										assign node1861 = (inp[13]) ? node1867 : node1862;
											assign node1862 = (inp[14]) ? node1864 : 1'b1;
												assign node1864 = (inp[2]) ? 1'b1 : 1'b0;
											assign node1867 = (inp[11]) ? 1'b1 : node1868;
												assign node1868 = (inp[14]) ? node1870 : 1'b0;
													assign node1870 = (inp[3]) ? 1'b0 : 1'b1;
								assign node1875 = (inp[8]) ? node1903 : node1876;
									assign node1876 = (inp[0]) ? node1890 : node1877;
										assign node1877 = (inp[14]) ? node1883 : node1878;
											assign node1878 = (inp[13]) ? node1880 : 1'b1;
												assign node1880 = (inp[11]) ? 1'b1 : 1'b0;
											assign node1883 = (inp[2]) ? 1'b1 : node1884;
												assign node1884 = (inp[11]) ? 1'b0 : node1885;
													assign node1885 = (inp[13]) ? 1'b1 : 1'b0;
										assign node1890 = (inp[4]) ? node1892 : 1'b0;
											assign node1892 = (inp[13]) ? node1894 : 1'b1;
												assign node1894 = (inp[3]) ? node1900 : node1895;
													assign node1895 = (inp[2]) ? node1897 : 1'b1;
														assign node1897 = (inp[11]) ? 1'b1 : 1'b0;
													assign node1900 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1903 = (inp[4]) ? 1'b0 : node1904;
										assign node1904 = (inp[0]) ? node1906 : 1'b0;
											assign node1906 = (inp[14]) ? node1912 : node1907;
												assign node1907 = (inp[13]) ? node1909 : 1'b1;
													assign node1909 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1912 = (inp[11]) ? 1'b0 : node1913;
													assign node1913 = (inp[9]) ? node1919 : node1914;
														assign node1914 = (inp[3]) ? 1'b0 : node1915;
															assign node1915 = (inp[13]) ? 1'b0 : 1'b1;
														assign node1919 = (inp[2]) ? 1'b1 : node1920;
															assign node1920 = (inp[13]) ? 1'b1 : 1'b0;
			assign node1926 = (inp[12]) ? node2008 : node1927;
				assign node1927 = (inp[4]) ? node1987 : node1928;
					assign node1928 = (inp[0]) ? node1950 : node1929;
						assign node1929 = (inp[8]) ? 1'b1 : node1930;
							assign node1930 = (inp[1]) ? node1932 : 1'b1;
								assign node1932 = (inp[13]) ? node1938 : node1933;
									assign node1933 = (inp[14]) ? node1935 : 1'b0;
										assign node1935 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1938 = (inp[11]) ? node1944 : node1939;
										assign node1939 = (inp[2]) ? 1'b1 : node1940;
											assign node1940 = (inp[14]) ? 1'b0 : 1'b1;
										assign node1944 = (inp[14]) ? node1946 : 1'b0;
											assign node1946 = (inp[2]) ? 1'b0 : 1'b1;
						assign node1950 = (inp[1]) ? node1968 : node1951;
							assign node1951 = (inp[2]) ? node1963 : node1952;
								assign node1952 = (inp[14]) ? node1958 : node1953;
									assign node1953 = (inp[11]) ? 1'b0 : node1954;
										assign node1954 = (inp[13]) ? 1'b1 : 1'b0;
									assign node1958 = (inp[11]) ? 1'b1 : node1959;
										assign node1959 = (inp[13]) ? 1'b0 : 1'b1;
								assign node1963 = (inp[13]) ? node1965 : 1'b0;
									assign node1965 = (inp[11]) ? 1'b0 : 1'b1;
							assign node1968 = (inp[8]) ? node1970 : 1'b1;
								assign node1970 = (inp[13]) ? node1976 : node1971;
									assign node1971 = (inp[2]) ? 1'b0 : node1972;
										assign node1972 = (inp[14]) ? 1'b1 : 1'b0;
									assign node1976 = (inp[11]) ? node1982 : node1977;
										assign node1977 = (inp[14]) ? node1979 : 1'b1;
											assign node1979 = (inp[2]) ? 1'b1 : 1'b0;
										assign node1982 = (inp[2]) ? 1'b0 : node1983;
											assign node1983 = (inp[14]) ? 1'b1 : 1'b0;
					assign node1987 = (inp[1]) ? node1989 : 1'b1;
						assign node1989 = (inp[8]) ? 1'b1 : node1990;
							assign node1990 = (inp[11]) ? node2002 : node1991;
								assign node1991 = (inp[13]) ? node1997 : node1992;
									assign node1992 = (inp[14]) ? node1994 : 1'b0;
										assign node1994 = (inp[2]) ? 1'b0 : 1'b1;
									assign node1997 = (inp[2]) ? 1'b1 : node1998;
										assign node1998 = (inp[14]) ? 1'b0 : 1'b1;
								assign node2002 = (inp[2]) ? 1'b0 : node2003;
									assign node2003 = (inp[14]) ? 1'b1 : 1'b0;
				assign node2008 = (inp[15]) ? node2430 : node2009;
					assign node2009 = (inp[7]) ? node2241 : node2010;
						assign node2010 = (inp[3]) ? node2138 : node2011;
							assign node2011 = (inp[10]) ? node2099 : node2012;
								assign node2012 = (inp[9]) ? node2058 : node2013;
									assign node2013 = (inp[0]) ? node2023 : node2014;
										assign node2014 = (inp[11]) ? node2016 : 1'b0;
											assign node2016 = (inp[14]) ? 1'b0 : node2017;
												assign node2017 = (inp[1]) ? node2019 : 1'b0;
													assign node2019 = (inp[8]) ? 1'b0 : 1'b1;
										assign node2023 = (inp[4]) ? node2049 : node2024;
											assign node2024 = (inp[14]) ? node2034 : node2025;
												assign node2025 = (inp[2]) ? 1'b1 : node2026;
													assign node2026 = (inp[13]) ? 1'b0 : node2027;
														assign node2027 = (inp[1]) ? node2029 : 1'b1;
															assign node2029 = (inp[8]) ? 1'b1 : 1'b0;
												assign node2034 = (inp[8]) ? node2038 : node2035;
													assign node2035 = (inp[1]) ? 1'b0 : 1'b1;
													assign node2038 = (inp[1]) ? node2044 : node2039;
														assign node2039 = (inp[2]) ? 1'b0 : node2040;
															assign node2040 = (inp[13]) ? 1'b0 : 1'b0;
														assign node2044 = (inp[2]) ? node2046 : 1'b1;
															assign node2046 = (inp[11]) ? 1'b1 : 1'b0;
											assign node2049 = (inp[1]) ? node2051 : 1'b0;
												assign node2051 = (inp[8]) ? 1'b0 : node2052;
													assign node2052 = (inp[13]) ? 1'b1 : node2053;
														assign node2053 = (inp[2]) ? 1'b1 : 1'b0;
									assign node2058 = (inp[2]) ? node2074 : node2059;
										assign node2059 = (inp[1]) ? node2061 : 1'b1;
											assign node2061 = (inp[11]) ? node2069 : node2062;
												assign node2062 = (inp[0]) ? node2064 : 1'b1;
													assign node2064 = (inp[8]) ? node2066 : 1'b0;
														assign node2066 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2069 = (inp[13]) ? 1'b1 : node2070;
													assign node2070 = (inp[8]) ? 1'b1 : 1'b0;
										assign node2074 = (inp[11]) ? node2082 : node2075;
											assign node2075 = (inp[13]) ? 1'b1 : node2076;
												assign node2076 = (inp[1]) ? node2078 : 1'b1;
													assign node2078 = (inp[14]) ? 1'b0 : 1'b1;
											assign node2082 = (inp[0]) ? node2088 : node2083;
												assign node2083 = (inp[1]) ? node2085 : 1'b1;
													assign node2085 = (inp[8]) ? 1'b1 : 1'b0;
												assign node2088 = (inp[8]) ? 1'b0 : node2089;
													assign node2089 = (inp[13]) ? node2093 : node2090;
														assign node2090 = (inp[4]) ? 1'b1 : 1'b0;
														assign node2093 = (inp[1]) ? node2095 : 1'b0;
															assign node2095 = (inp[4]) ? 1'b0 : 1'b1;
								assign node2099 = (inp[0]) ? node2111 : node2100;
									assign node2100 = (inp[8]) ? 1'b0 : node2101;
										assign node2101 = (inp[1]) ? node2103 : 1'b0;
											assign node2103 = (inp[2]) ? 1'b1 : node2104;
												assign node2104 = (inp[11]) ? node2106 : 1'b0;
													assign node2106 = (inp[14]) ? 1'b0 : 1'b1;
									assign node2111 = (inp[4]) ? node2131 : node2112;
										assign node2112 = (inp[1]) ? node2124 : node2113;
											assign node2113 = (inp[9]) ? node2115 : 1'b1;
												assign node2115 = (inp[13]) ? node2117 : 1'b1;
													assign node2117 = (inp[11]) ? node2121 : node2118;
														assign node2118 = (inp[14]) ? 1'b1 : 1'b0;
														assign node2121 = (inp[8]) ? 1'b0 : 1'b1;
											assign node2124 = (inp[8]) ? node2126 : 1'b0;
												assign node2126 = (inp[13]) ? node2128 : 1'b1;
													assign node2128 = (inp[11]) ? 1'b1 : 1'b0;
										assign node2131 = (inp[8]) ? 1'b0 : node2132;
											assign node2132 = (inp[1]) ? node2134 : 1'b0;
												assign node2134 = (inp[11]) ? 1'b1 : 1'b0;
							assign node2138 = (inp[9]) ? node2180 : node2139;
								assign node2139 = (inp[4]) ? node2169 : node2140;
									assign node2140 = (inp[0]) ? node2150 : node2141;
										assign node2141 = (inp[8]) ? 1'b1 : node2142;
											assign node2142 = (inp[1]) ? node2144 : 1'b1;
												assign node2144 = (inp[14]) ? node2146 : 1'b0;
													assign node2146 = (inp[11]) ? 1'b1 : 1'b0;
										assign node2150 = (inp[1]) ? node2162 : node2151;
											assign node2151 = (inp[2]) ? node2157 : node2152;
												assign node2152 = (inp[14]) ? 1'b1 : node2153;
													assign node2153 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2157 = (inp[13]) ? node2159 : 1'b0;
													assign node2159 = (inp[11]) ? 1'b0 : 1'b1;
											assign node2162 = (inp[8]) ? node2164 : 1'b1;
												assign node2164 = (inp[11]) ? node2166 : 1'b1;
													assign node2166 = (inp[10]) ? 1'b1 : 1'b0;
									assign node2169 = (inp[1]) ? node2171 : 1'b1;
										assign node2171 = (inp[8]) ? 1'b1 : node2172;
											assign node2172 = (inp[14]) ? node2174 : 1'b0;
												assign node2174 = (inp[2]) ? node2176 : 1'b1;
													assign node2176 = (inp[11]) ? 1'b0 : 1'b1;
								assign node2180 = (inp[10]) ? node2208 : node2181;
									assign node2181 = (inp[2]) ? node2191 : node2182;
										assign node2182 = (inp[8]) ? 1'b0 : node2183;
											assign node2183 = (inp[1]) ? node2185 : 1'b0;
												assign node2185 = (inp[4]) ? node2187 : 1'b0;
													assign node2187 = (inp[0]) ? 1'b1 : 1'b0;
										assign node2191 = (inp[1]) ? node2197 : node2192;
											assign node2192 = (inp[0]) ? node2194 : 1'b0;
												assign node2194 = (inp[4]) ? 1'b0 : 1'b1;
											assign node2197 = (inp[8]) ? node2203 : node2198;
												assign node2198 = (inp[11]) ? 1'b1 : node2199;
													assign node2199 = (inp[13]) ? 1'b0 : 1'b1;
												assign node2203 = (inp[14]) ? 1'b0 : node2204;
													assign node2204 = (inp[4]) ? 1'b0 : 1'b1;
									assign node2208 = (inp[1]) ? node2220 : node2209;
										assign node2209 = (inp[0]) ? node2211 : 1'b1;
											assign node2211 = (inp[4]) ? 1'b1 : node2212;
												assign node2212 = (inp[11]) ? node2214 : 1'b1;
													assign node2214 = (inp[2]) ? 1'b0 : node2215;
														assign node2215 = (inp[14]) ? 1'b1 : 1'b0;
										assign node2220 = (inp[2]) ? node2230 : node2221;
											assign node2221 = (inp[8]) ? 1'b1 : node2222;
												assign node2222 = (inp[14]) ? 1'b1 : node2223;
													assign node2223 = (inp[11]) ? 1'b0 : node2224;
														assign node2224 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2230 = (inp[13]) ? node2236 : node2231;
												assign node2231 = (inp[11]) ? node2233 : 1'b0;
													assign node2233 = (inp[8]) ? 1'b0 : 1'b1;
												assign node2236 = (inp[4]) ? 1'b1 : node2237;
													assign node2237 = (inp[11]) ? 1'b0 : 1'b1;
						assign node2241 = (inp[9]) ? node2327 : node2242;
							assign node2242 = (inp[4]) ? node2300 : node2243;
								assign node2243 = (inp[0]) ? node2259 : node2244;
									assign node2244 = (inp[1]) ? node2246 : 1'b0;
										assign node2246 = (inp[8]) ? 1'b0 : node2247;
											assign node2247 = (inp[2]) ? node2253 : node2248;
												assign node2248 = (inp[14]) ? 1'b0 : node2249;
													assign node2249 = (inp[10]) ? 1'b1 : 1'b0;
												assign node2253 = (inp[11]) ? 1'b1 : node2254;
													assign node2254 = (inp[13]) ? 1'b0 : 1'b1;
									assign node2259 = (inp[8]) ? node2279 : node2260;
										assign node2260 = (inp[1]) ? 1'b0 : node2261;
											assign node2261 = (inp[11]) ? node2273 : node2262;
												assign node2262 = (inp[13]) ? node2266 : node2263;
													assign node2263 = (inp[2]) ? 1'b1 : 1'b0;
													assign node2266 = (inp[3]) ? node2268 : 1'b0;
														assign node2268 = (inp[14]) ? node2270 : 1'b0;
															assign node2270 = (inp[2]) ? 1'b0 : 1'b1;
												assign node2273 = (inp[14]) ? node2275 : 1'b1;
													assign node2275 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2279 = (inp[13]) ? node2285 : node2280;
											assign node2280 = (inp[14]) ? node2282 : 1'b1;
												assign node2282 = (inp[2]) ? 1'b1 : 1'b0;
											assign node2285 = (inp[1]) ? node2295 : node2286;
												assign node2286 = (inp[10]) ? node2288 : 1'b0;
													assign node2288 = (inp[2]) ? 1'b0 : node2289;
														assign node2289 = (inp[14]) ? node2291 : 1'b1;
															assign node2291 = (inp[11]) ? 1'b0 : 1'b1;
												assign node2295 = (inp[11]) ? 1'b1 : node2296;
													assign node2296 = (inp[2]) ? 1'b0 : 1'b1;
								assign node2300 = (inp[8]) ? 1'b0 : node2301;
									assign node2301 = (inp[1]) ? node2303 : 1'b0;
										assign node2303 = (inp[3]) ? node2311 : node2304;
											assign node2304 = (inp[14]) ? 1'b0 : node2305;
												assign node2305 = (inp[11]) ? 1'b1 : node2306;
													assign node2306 = (inp[13]) ? 1'b0 : 1'b1;
											assign node2311 = (inp[13]) ? node2317 : node2312;
												assign node2312 = (inp[2]) ? 1'b1 : node2313;
													assign node2313 = (inp[14]) ? 1'b0 : 1'b1;
												assign node2317 = (inp[14]) ? node2319 : 1'b0;
													assign node2319 = (inp[0]) ? 1'b0 : node2320;
														assign node2320 = (inp[11]) ? 1'b1 : node2321;
															assign node2321 = (inp[10]) ? 1'b1 : 1'b0;
							assign node2327 = (inp[10]) ? node2377 : node2328;
								assign node2328 = (inp[4]) ? node2362 : node2329;
									assign node2329 = (inp[0]) ? node2343 : node2330;
										assign node2330 = (inp[8]) ? 1'b1 : node2331;
											assign node2331 = (inp[1]) ? node2333 : 1'b1;
												assign node2333 = (inp[3]) ? 1'b0 : node2334;
													assign node2334 = (inp[13]) ? node2336 : 1'b0;
														assign node2336 = (inp[11]) ? 1'b0 : node2337;
															assign node2337 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2343 = (inp[1]) ? node2359 : node2344;
											assign node2344 = (inp[11]) ? node2354 : node2345;
												assign node2345 = (inp[2]) ? node2351 : node2346;
													assign node2346 = (inp[13]) ? node2348 : 1'b0;
														assign node2348 = (inp[14]) ? 1'b0 : 1'b1;
													assign node2351 = (inp[13]) ? 1'b1 : 1'b0;
												assign node2354 = (inp[2]) ? 1'b0 : node2355;
													assign node2355 = (inp[14]) ? 1'b1 : 1'b0;
											assign node2359 = (inp[8]) ? 1'b0 : 1'b1;
									assign node2362 = (inp[1]) ? node2364 : 1'b1;
										assign node2364 = (inp[8]) ? 1'b1 : node2365;
											assign node2365 = (inp[11]) ? node2371 : node2366;
												assign node2366 = (inp[13]) ? 1'b1 : node2367;
													assign node2367 = (inp[14]) ? 1'b1 : 1'b0;
												assign node2371 = (inp[14]) ? node2373 : 1'b0;
													assign node2373 = (inp[2]) ? 1'b0 : 1'b1;
								assign node2377 = (inp[2]) ? node2405 : node2378;
									assign node2378 = (inp[1]) ? node2390 : node2379;
										assign node2379 = (inp[11]) ? 1'b0 : node2380;
											assign node2380 = (inp[0]) ? node2382 : 1'b0;
												assign node2382 = (inp[14]) ? 1'b0 : node2383;
													assign node2383 = (inp[4]) ? 1'b0 : node2384;
														assign node2384 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2390 = (inp[8]) ? node2398 : node2391;
											assign node2391 = (inp[14]) ? node2393 : 1'b1;
												assign node2393 = (inp[11]) ? 1'b0 : node2394;
													assign node2394 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2398 = (inp[4]) ? 1'b0 : node2399;
												assign node2399 = (inp[0]) ? node2401 : 1'b0;
													assign node2401 = (inp[11]) ? 1'b0 : 1'b1;
									assign node2405 = (inp[0]) ? node2415 : node2406;
										assign node2406 = (inp[8]) ? 1'b0 : node2407;
											assign node2407 = (inp[1]) ? node2409 : 1'b0;
												assign node2409 = (inp[4]) ? node2411 : 1'b1;
													assign node2411 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2415 = (inp[4]) ? node2425 : node2416;
											assign node2416 = (inp[1]) ? node2418 : 1'b1;
												assign node2418 = (inp[8]) ? node2420 : 1'b0;
													assign node2420 = (inp[13]) ? node2422 : 1'b1;
														assign node2422 = (inp[11]) ? 1'b1 : 1'b0;
											assign node2425 = (inp[8]) ? 1'b0 : node2426;
												assign node2426 = (inp[1]) ? 1'b1 : 1'b0;
					assign node2430 = (inp[1]) ? node2452 : node2431;
						assign node2431 = (inp[4]) ? 1'b1 : node2432;
							assign node2432 = (inp[0]) ? node2434 : 1'b1;
								assign node2434 = (inp[13]) ? node2440 : node2435;
									assign node2435 = (inp[14]) ? node2437 : 1'b0;
										assign node2437 = (inp[2]) ? 1'b0 : 1'b1;
									assign node2440 = (inp[11]) ? node2446 : node2441;
										assign node2441 = (inp[14]) ? node2443 : 1'b1;
											assign node2443 = (inp[2]) ? 1'b1 : 1'b0;
										assign node2446 = (inp[2]) ? 1'b0 : node2447;
											assign node2447 = (inp[14]) ? 1'b1 : 1'b0;
						assign node2452 = (inp[8]) ? node2490 : node2453;
							assign node2453 = (inp[4]) ? node2473 : node2454;
								assign node2454 = (inp[0]) ? 1'b1 : node2455;
									assign node2455 = (inp[2]) ? node2467 : node2456;
										assign node2456 = (inp[14]) ? node2462 : node2457;
											assign node2457 = (inp[11]) ? 1'b0 : node2458;
												assign node2458 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2462 = (inp[11]) ? 1'b1 : node2463;
												assign node2463 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2467 = (inp[11]) ? 1'b0 : node2468;
											assign node2468 = (inp[13]) ? 1'b1 : 1'b0;
								assign node2473 = (inp[13]) ? node2479 : node2474;
									assign node2474 = (inp[2]) ? 1'b0 : node2475;
										assign node2475 = (inp[14]) ? 1'b1 : 1'b0;
									assign node2479 = (inp[11]) ? node2485 : node2480;
										assign node2480 = (inp[2]) ? 1'b1 : node2481;
											assign node2481 = (inp[14]) ? 1'b0 : 1'b1;
										assign node2485 = (inp[2]) ? 1'b0 : node2486;
											assign node2486 = (inp[14]) ? 1'b1 : 1'b0;
							assign node2490 = (inp[4]) ? 1'b1 : node2491;
								assign node2491 = (inp[0]) ? node2493 : 1'b1;
									assign node2493 = (inp[2]) ? node2505 : node2494;
										assign node2494 = (inp[14]) ? node2500 : node2495;
											assign node2495 = (inp[11]) ? 1'b0 : node2496;
												assign node2496 = (inp[13]) ? 1'b1 : 1'b0;
											assign node2500 = (inp[11]) ? 1'b1 : node2501;
												assign node2501 = (inp[13]) ? 1'b0 : 1'b1;
										assign node2505 = (inp[11]) ? 1'b0 : node2506;
											assign node2506 = (inp[13]) ? 1'b1 : 1'b0;

endmodule