module dtc_split66_bm48 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node6;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node12;
	wire [14-1:0] node13;
	wire [14-1:0] node17;
	wire [14-1:0] node18;
	wire [14-1:0] node19;
	wire [14-1:0] node20;
	wire [14-1:0] node21;
	wire [14-1:0] node25;
	wire [14-1:0] node30;
	wire [14-1:0] node31;
	wire [14-1:0] node32;
	wire [14-1:0] node34;
	wire [14-1:0] node36;
	wire [14-1:0] node38;
	wire [14-1:0] node42;
	wire [14-1:0] node44;
	wire [14-1:0] node46;
	wire [14-1:0] node49;
	wire [14-1:0] node50;
	wire [14-1:0] node51;
	wire [14-1:0] node52;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node56;
	wire [14-1:0] node59;
	wire [14-1:0] node60;
	wire [14-1:0] node62;
	wire [14-1:0] node63;
	wire [14-1:0] node68;
	wire [14-1:0] node69;
	wire [14-1:0] node70;
	wire [14-1:0] node71;
	wire [14-1:0] node74;
	wire [14-1:0] node75;
	wire [14-1:0] node81;
	wire [14-1:0] node82;
	wire [14-1:0] node84;
	wire [14-1:0] node86;
	wire [14-1:0] node87;
	wire [14-1:0] node88;
	wire [14-1:0] node95;
	wire [14-1:0] node96;
	wire [14-1:0] node98;
	wire [14-1:0] node99;
	wire [14-1:0] node100;
	wire [14-1:0] node101;
	wire [14-1:0] node103;
	wire [14-1:0] node106;
	wire [14-1:0] node108;
	wire [14-1:0] node111;
	wire [14-1:0] node112;
	wire [14-1:0] node113;
	wire [14-1:0] node114;
	wire [14-1:0] node121;
	wire [14-1:0] node122;
	wire [14-1:0] node124;
	wire [14-1:0] node125;
	wire [14-1:0] node127;
	wire [14-1:0] node128;
	wire [14-1:0] node129;
	wire [14-1:0] node135;
	wire [14-1:0] node137;
	wire [14-1:0] node140;
	wire [14-1:0] node141;
	wire [14-1:0] node143;
	wire [14-1:0] node145;
	wire [14-1:0] node147;
	wire [14-1:0] node148;
	wire [14-1:0] node151;
	wire [14-1:0] node154;
	wire [14-1:0] node155;
	wire [14-1:0] node156;
	wire [14-1:0] node157;
	wire [14-1:0] node158;
	wire [14-1:0] node160;
	wire [14-1:0] node161;
	wire [14-1:0] node163;
	wire [14-1:0] node167;
	wire [14-1:0] node169;
	wire [14-1:0] node170;
	wire [14-1:0] node174;
	wire [14-1:0] node175;
	wire [14-1:0] node178;
	wire [14-1:0] node179;
	wire [14-1:0] node180;
	wire [14-1:0] node182;
	wire [14-1:0] node187;
	wire [14-1:0] node188;
	wire [14-1:0] node189;
	wire [14-1:0] node190;
	wire [14-1:0] node191;
	wire [14-1:0] node193;
	wire [14-1:0] node196;
	wire [14-1:0] node197;
	wire [14-1:0] node198;
	wire [14-1:0] node201;
	wire [14-1:0] node208;
	wire [14-1:0] node209;
	wire [14-1:0] node210;
	wire [14-1:0] node211;
	wire [14-1:0] node212;
	wire [14-1:0] node214;
	wire [14-1:0] node215;
	wire [14-1:0] node222;
	wire [14-1:0] node223;
	wire [14-1:0] node224;
	wire [14-1:0] node225;
	wire [14-1:0] node226;
	wire [14-1:0] node228;
	wire [14-1:0] node229;
	wire [14-1:0] node232;
	wire [14-1:0] node235;
	wire [14-1:0] node236;
	wire [14-1:0] node239;
	wire [14-1:0] node244;
	wire [14-1:0] node245;
	wire [14-1:0] node247;
	wire [14-1:0] node248;
	wire [14-1:0] node252;
	wire [14-1:0] node253;
	wire [14-1:0] node254;
	wire [14-1:0] node255;
	wire [14-1:0] node256;
	wire [14-1:0] node262;
	wire [14-1:0] node264;
	wire [14-1:0] node267;
	wire [14-1:0] node268;
	wire [14-1:0] node269;
	wire [14-1:0] node270;
	wire [14-1:0] node271;
	wire [14-1:0] node273;
	wire [14-1:0] node274;
	wire [14-1:0] node276;
	wire [14-1:0] node281;
	wire [14-1:0] node283;
	wire [14-1:0] node284;
	wire [14-1:0] node285;
	wire [14-1:0] node287;
	wire [14-1:0] node288;
	wire [14-1:0] node290;
	wire [14-1:0] node296;
	wire [14-1:0] node297;
	wire [14-1:0] node298;
	wire [14-1:0] node299;
	wire [14-1:0] node300;
	wire [14-1:0] node304;
	wire [14-1:0] node306;
	wire [14-1:0] node307;
	wire [14-1:0] node309;
	wire [14-1:0] node311;
	wire [14-1:0] node312;
	wire [14-1:0] node315;
	wire [14-1:0] node319;
	wire [14-1:0] node320;
	wire [14-1:0] node322;
	wire [14-1:0] node323;
	wire [14-1:0] node324;
	wire [14-1:0] node325;
	wire [14-1:0] node326;
	wire [14-1:0] node331;
	wire [14-1:0] node332;
	wire [14-1:0] node333;
	wire [14-1:0] node336;
	wire [14-1:0] node342;
	wire [14-1:0] node343;
	wire [14-1:0] node344;
	wire [14-1:0] node345;
	wire [14-1:0] node346;
	wire [14-1:0] node348;
	wire [14-1:0] node349;
	wire [14-1:0] node353;
	wire [14-1:0] node354;
	wire [14-1:0] node355;
	wire [14-1:0] node360;
	wire [14-1:0] node362;
	wire [14-1:0] node363;
	wire [14-1:0] node364;
	wire [14-1:0] node369;
	wire [14-1:0] node370;
	wire [14-1:0] node372;
	wire [14-1:0] node373;
	wire [14-1:0] node374;
	wire [14-1:0] node377;
	wire [14-1:0] node382;
	wire [14-1:0] node384;
	wire [14-1:0] node386;
	wire [14-1:0] node388;
	wire [14-1:0] node389;
	wire [14-1:0] node392;
	wire [14-1:0] node395;
	wire [14-1:0] node396;
	wire [14-1:0] node397;
	wire [14-1:0] node399;
	wire [14-1:0] node400;
	wire [14-1:0] node401;
	wire [14-1:0] node402;
	wire [14-1:0] node404;
	wire [14-1:0] node405;
	wire [14-1:0] node406;
	wire [14-1:0] node409;
	wire [14-1:0] node413;
	wire [14-1:0] node415;
	wire [14-1:0] node416;
	wire [14-1:0] node420;
	wire [14-1:0] node421;
	wire [14-1:0] node423;
	wire [14-1:0] node424;
	wire [14-1:0] node429;
	wire [14-1:0] node430;
	wire [14-1:0] node431;
	wire [14-1:0] node432;
	wire [14-1:0] node434;
	wire [14-1:0] node440;
	wire [14-1:0] node441;
	wire [14-1:0] node442;
	wire [14-1:0] node443;
	wire [14-1:0] node445;
	wire [14-1:0] node447;
	wire [14-1:0] node448;
	wire [14-1:0] node449;
	wire [14-1:0] node456;
	wire [14-1:0] node457;
	wire [14-1:0] node458;
	wire [14-1:0] node459;
	wire [14-1:0] node460;
	wire [14-1:0] node462;
	wire [14-1:0] node466;
	wire [14-1:0] node467;
	wire [14-1:0] node468;
	wire [14-1:0] node469;
	wire [14-1:0] node474;
	wire [14-1:0] node478;
	wire [14-1:0] node479;
	wire [14-1:0] node482;
	wire [14-1:0] node484;
	wire [14-1:0] node486;
	wire [14-1:0] node489;
	wire [14-1:0] node490;
	wire [14-1:0] node491;
	wire [14-1:0] node493;
	wire [14-1:0] node494;
	wire [14-1:0] node495;
	wire [14-1:0] node496;
	wire [14-1:0] node497;
	wire [14-1:0] node500;
	wire [14-1:0] node503;
	wire [14-1:0] node504;
	wire [14-1:0] node510;
	wire [14-1:0] node511;
	wire [14-1:0] node512;
	wire [14-1:0] node514;
	wire [14-1:0] node515;
	wire [14-1:0] node517;
	wire [14-1:0] node518;
	wire [14-1:0] node521;
	wire [14-1:0] node524;
	wire [14-1:0] node528;
	wire [14-1:0] node530;
	wire [14-1:0] node532;
	wire [14-1:0] node534;
	wire [14-1:0] node538;
	wire [14-1:0] node539;
	wire [14-1:0] node540;
	wire [14-1:0] node541;
	wire [14-1:0] node542;
	wire [14-1:0] node543;
	wire [14-1:0] node548;
	wire [14-1:0] node550;
	wire [14-1:0] node552;
	wire [14-1:0] node555;
	wire [14-1:0] node556;
	wire [14-1:0] node557;
	wire [14-1:0] node558;
	wire [14-1:0] node562;
	wire [14-1:0] node564;
	wire [14-1:0] node565;
	wire [14-1:0] node567;
	wire [14-1:0] node568;
	wire [14-1:0] node569;
	wire [14-1:0] node570;
	wire [14-1:0] node577;
	wire [14-1:0] node578;
	wire [14-1:0] node580;
	wire [14-1:0] node581;
	wire [14-1:0] node582;
	wire [14-1:0] node583;
	wire [14-1:0] node584;
	wire [14-1:0] node585;
	wire [14-1:0] node586;
	wire [14-1:0] node593;
	wire [14-1:0] node596;
	wire [14-1:0] node597;
	wire [14-1:0] node601;
	wire [14-1:0] node602;
	wire [14-1:0] node604;
	wire [14-1:0] node605;
	wire [14-1:0] node606;
	wire [14-1:0] node607;
	wire [14-1:0] node608;
	wire [14-1:0] node609;
	wire [14-1:0] node616;
	wire [14-1:0] node619;
	wire [14-1:0] node620;
	wire [14-1:0] node621;
	wire [14-1:0] node626;
	wire [14-1:0] node627;
	wire [14-1:0] node628;
	wire [14-1:0] node629;
	wire [14-1:0] node630;
	wire [14-1:0] node631;
	wire [14-1:0] node632;
	wire [14-1:0] node635;
	wire [14-1:0] node636;
	wire [14-1:0] node638;
	wire [14-1:0] node641;
	wire [14-1:0] node642;
	wire [14-1:0] node643;
	wire [14-1:0] node647;
	wire [14-1:0] node648;
	wire [14-1:0] node652;
	wire [14-1:0] node653;
	wire [14-1:0] node654;
	wire [14-1:0] node656;
	wire [14-1:0] node658;
	wire [14-1:0] node662;
	wire [14-1:0] node663;
	wire [14-1:0] node665;
	wire [14-1:0] node667;
	wire [14-1:0] node670;
	wire [14-1:0] node671;
	wire [14-1:0] node675;
	wire [14-1:0] node676;
	wire [14-1:0] node677;
	wire [14-1:0] node678;
	wire [14-1:0] node679;
	wire [14-1:0] node681;
	wire [14-1:0] node684;
	wire [14-1:0] node685;
	wire [14-1:0] node689;
	wire [14-1:0] node690;
	wire [14-1:0] node691;
	wire [14-1:0] node693;
	wire [14-1:0] node696;
	wire [14-1:0] node699;
	wire [14-1:0] node700;
	wire [14-1:0] node704;
	wire [14-1:0] node705;
	wire [14-1:0] node707;
	wire [14-1:0] node708;
	wire [14-1:0] node711;
	wire [14-1:0] node715;
	wire [14-1:0] node716;
	wire [14-1:0] node717;
	wire [14-1:0] node718;
	wire [14-1:0] node719;
	wire [14-1:0] node721;
	wire [14-1:0] node725;
	wire [14-1:0] node727;
	wire [14-1:0] node729;
	wire [14-1:0] node732;
	wire [14-1:0] node734;
	wire [14-1:0] node735;
	wire [14-1:0] node736;
	wire [14-1:0] node741;
	wire [14-1:0] node742;
	wire [14-1:0] node743;
	wire [14-1:0] node746;
	wire [14-1:0] node747;
	wire [14-1:0] node752;
	wire [14-1:0] node753;
	wire [14-1:0] node754;
	wire [14-1:0] node755;
	wire [14-1:0] node756;
	wire [14-1:0] node757;
	wire [14-1:0] node759;
	wire [14-1:0] node761;
	wire [14-1:0] node765;
	wire [14-1:0] node766;
	wire [14-1:0] node768;
	wire [14-1:0] node769;
	wire [14-1:0] node772;
	wire [14-1:0] node775;
	wire [14-1:0] node776;
	wire [14-1:0] node777;
	wire [14-1:0] node782;
	wire [14-1:0] node783;
	wire [14-1:0] node784;
	wire [14-1:0] node785;
	wire [14-1:0] node788;
	wire [14-1:0] node789;
	wire [14-1:0] node793;
	wire [14-1:0] node796;
	wire [14-1:0] node797;
	wire [14-1:0] node798;
	wire [14-1:0] node799;
	wire [14-1:0] node804;
	wire [14-1:0] node805;
	wire [14-1:0] node809;
	wire [14-1:0] node810;
	wire [14-1:0] node811;
	wire [14-1:0] node812;
	wire [14-1:0] node817;
	wire [14-1:0] node819;
	wire [14-1:0] node821;
	wire [14-1:0] node824;
	wire [14-1:0] node825;
	wire [14-1:0] node826;
	wire [14-1:0] node827;
	wire [14-1:0] node828;
	wire [14-1:0] node829;
	wire [14-1:0] node834;
	wire [14-1:0] node836;
	wire [14-1:0] node838;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node843;
	wire [14-1:0] node844;
	wire [14-1:0] node849;
	wire [14-1:0] node851;
	wire [14-1:0] node853;
	wire [14-1:0] node856;
	wire [14-1:0] node857;
	wire [14-1:0] node859;
	wire [14-1:0] node861;
	wire [14-1:0] node863;
	wire [14-1:0] node866;
	wire [14-1:0] node867;
	wire [14-1:0] node868;
	wire [14-1:0] node869;
	wire [14-1:0] node875;
	wire [14-1:0] node876;
	wire [14-1:0] node877;
	wire [14-1:0] node878;
	wire [14-1:0] node879;
	wire [14-1:0] node881;
	wire [14-1:0] node883;
	wire [14-1:0] node885;
	wire [14-1:0] node886;
	wire [14-1:0] node891;
	wire [14-1:0] node893;
	wire [14-1:0] node894;
	wire [14-1:0] node895;
	wire [14-1:0] node896;
	wire [14-1:0] node901;
	wire [14-1:0] node904;
	wire [14-1:0] node905;
	wire [14-1:0] node907;
	wire [14-1:0] node909;
	wire [14-1:0] node911;
	wire [14-1:0] node912;
	wire [14-1:0] node916;
	wire [14-1:0] node918;
	wire [14-1:0] node921;
	wire [14-1:0] node922;
	wire [14-1:0] node923;
	wire [14-1:0] node924;
	wire [14-1:0] node925;
	wire [14-1:0] node926;
	wire [14-1:0] node927;
	wire [14-1:0] node928;
	wire [14-1:0] node934;
	wire [14-1:0] node936;
	wire [14-1:0] node938;
	wire [14-1:0] node941;
	wire [14-1:0] node942;
	wire [14-1:0] node943;
	wire [14-1:0] node944;
	wire [14-1:0] node949;
	wire [14-1:0] node951;
	wire [14-1:0] node953;
	wire [14-1:0] node956;
	wire [14-1:0] node957;
	wire [14-1:0] node958;
	wire [14-1:0] node959;
	wire [14-1:0] node964;
	wire [14-1:0] node966;
	wire [14-1:0] node968;
	wire [14-1:0] node971;
	wire [14-1:0] node972;
	wire [14-1:0] node973;
	wire [14-1:0] node974;
	wire [14-1:0] node976;
	wire [14-1:0] node978;
	wire [14-1:0] node979;
	wire [14-1:0] node983;
	wire [14-1:0] node984;
	wire [14-1:0] node986;
	wire [14-1:0] node987;
	wire [14-1:0] node992;
	wire [14-1:0] node994;
	wire [14-1:0] node995;
	wire [14-1:0] node996;
	wire [14-1:0] node1000;
	wire [14-1:0] node1002;
	wire [14-1:0] node1005;
	wire [14-1:0] node1006;
	wire [14-1:0] node1007;
	wire [14-1:0] node1008;
	wire [14-1:0] node1010;
	wire [14-1:0] node1013;
	wire [14-1:0] node1014;
	wire [14-1:0] node1015;
	wire [14-1:0] node1020;
	wire [14-1:0] node1021;
	wire [14-1:0] node1025;
	wire [14-1:0] node1026;
	wire [14-1:0] node1028;
	wire [14-1:0] node1029;
	wire [14-1:0] node1030;
	wire [14-1:0] node1034;
	wire [14-1:0] node1037;
	wire [14-1:0] node1038;
	wire [14-1:0] node1040;
	wire [14-1:0] node1044;
	wire [14-1:0] node1045;
	wire [14-1:0] node1046;
	wire [14-1:0] node1047;
	wire [14-1:0] node1049;
	wire [14-1:0] node1050;
	wire [14-1:0] node1051;
	wire [14-1:0] node1052;
	wire [14-1:0] node1053;
	wire [14-1:0] node1056;
	wire [14-1:0] node1061;
	wire [14-1:0] node1063;
	wire [14-1:0] node1065;
	wire [14-1:0] node1067;
	wire [14-1:0] node1068;
	wire [14-1:0] node1072;
	wire [14-1:0] node1073;
	wire [14-1:0] node1074;
	wire [14-1:0] node1075;
	wire [14-1:0] node1076;
	wire [14-1:0] node1077;
	wire [14-1:0] node1079;
	wire [14-1:0] node1082;
	wire [14-1:0] node1083;
	wire [14-1:0] node1090;
	wire [14-1:0] node1091;
	wire [14-1:0] node1092;
	wire [14-1:0] node1093;
	wire [14-1:0] node1095;
	wire [14-1:0] node1099;
	wire [14-1:0] node1101;
	wire [14-1:0] node1103;
	wire [14-1:0] node1106;
	wire [14-1:0] node1107;
	wire [14-1:0] node1108;
	wire [14-1:0] node1109;
	wire [14-1:0] node1110;
	wire [14-1:0] node1114;
	wire [14-1:0] node1115;
	wire [14-1:0] node1120;
	wire [14-1:0] node1122;
	wire [14-1:0] node1123;
	wire [14-1:0] node1125;
	wire [14-1:0] node1129;
	wire [14-1:0] node1130;
	wire [14-1:0] node1131;
	wire [14-1:0] node1133;
	wire [14-1:0] node1134;
	wire [14-1:0] node1136;
	wire [14-1:0] node1137;
	wire [14-1:0] node1138;
	wire [14-1:0] node1145;
	wire [14-1:0] node1146;
	wire [14-1:0] node1147;
	wire [14-1:0] node1148;
	wire [14-1:0] node1149;
	wire [14-1:0] node1150;
	wire [14-1:0] node1151;
	wire [14-1:0] node1159;
	wire [14-1:0] node1161;
	wire [14-1:0] node1163;
	wire [14-1:0] node1164;
	wire [14-1:0] node1165;
	wire [14-1:0] node1169;
	wire [14-1:0] node1171;
	wire [14-1:0] node1174;
	wire [14-1:0] node1175;
	wire [14-1:0] node1177;
	wire [14-1:0] node1178;
	wire [14-1:0] node1179;
	wire [14-1:0] node1180;
	wire [14-1:0] node1181;
	wire [14-1:0] node1182;
	wire [14-1:0] node1184;
	wire [14-1:0] node1187;
	wire [14-1:0] node1188;
	wire [14-1:0] node1195;
	wire [14-1:0] node1196;
	wire [14-1:0] node1197;
	wire [14-1:0] node1198;
	wire [14-1:0] node1199;
	wire [14-1:0] node1200;
	wire [14-1:0] node1204;
	wire [14-1:0] node1205;
	wire [14-1:0] node1211;
	wire [14-1:0] node1213;
	wire [14-1:0] node1215;
	wire [14-1:0] node1216;
	wire [14-1:0] node1217;
	wire [14-1:0] node1221;
	wire [14-1:0] node1224;
	wire [14-1:0] node1225;
	wire [14-1:0] node1226;
	wire [14-1:0] node1227;
	wire [14-1:0] node1228;
	wire [14-1:0] node1232;
	wire [14-1:0] node1234;
	wire [14-1:0] node1236;
	wire [14-1:0] node1237;
	wire [14-1:0] node1241;
	wire [14-1:0] node1243;
	wire [14-1:0] node1245;
	wire [14-1:0] node1247;
	wire [14-1:0] node1248;
	wire [14-1:0] node1252;
	wire [14-1:0] node1253;
	wire [14-1:0] node1254;
	wire [14-1:0] node1255;
	wire [14-1:0] node1259;
	wire [14-1:0] node1261;
	wire [14-1:0] node1263;
	wire [14-1:0] node1265;

	assign outp = (inp[10]) ? node538 : node1;
		assign node1 = (inp[13]) ? node267 : node2;
			assign node2 = (inp[11]) ? node140 : node3;
				assign node3 = (inp[12]) ? node49 : node4;
					assign node4 = (inp[8]) ? node6 : 14'b00000100000011;
						assign node6 = (inp[1]) ? node8 : 14'b00000000000000;
							assign node8 = (inp[6]) ? node30 : node9;
								assign node9 = (inp[0]) ? node17 : node10;
									assign node10 = (inp[3]) ? node12 : 14'b00000000000000;
										assign node12 = (inp[2]) ? 14'b00000000000000 : node13;
											assign node13 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
									assign node17 = (inp[4]) ? 14'b00000000000000 : node18;
										assign node18 = (inp[3]) ? 14'b00000000000000 : node19;
											assign node19 = (inp[2]) ? node25 : node20;
												assign node20 = (inp[5]) ? 14'b00000000000000 : node21;
													assign node21 = (inp[9]) ? 14'b00000000000000 : 14'b00100100001100;
												assign node25 = (inp[9]) ? 14'b00000000000000 : 14'b10000000011010;
								assign node30 = (inp[5]) ? node42 : node31;
									assign node31 = (inp[0]) ? 14'b00000000000000 : node32;
										assign node32 = (inp[3]) ? node34 : 14'b00000000000000;
											assign node34 = (inp[9]) ? node36 : 14'b00000000000000;
												assign node36 = (inp[7]) ? node38 : 14'b00000000000000;
													assign node38 = (inp[4]) ? 14'b00000000000000 : 14'b01000000000000;
									assign node42 = (inp[3]) ? node44 : 14'b00000000000000;
										assign node44 = (inp[7]) ? node46 : 14'b00000000000000;
											assign node46 = (inp[9]) ? 14'b00000000011100 : 14'b00000000000000;
					assign node49 = (inp[8]) ? node95 : node50;
						assign node50 = (inp[9]) ? 14'b00000000000000 : node51;
							assign node51 = (inp[2]) ? node81 : node52;
								assign node52 = (inp[7]) ? node68 : node53;
									assign node53 = (inp[1]) ? node59 : node54;
										assign node54 = (inp[3]) ? node56 : 14'b00000000000000;
											assign node56 = (inp[0]) ? 14'b00000000000000 : 14'b00100000000011;
										assign node59 = (inp[3]) ? 14'b00000000000000 : node60;
											assign node60 = (inp[0]) ? node62 : 14'b00000000000000;
												assign node62 = (inp[6]) ? 14'b00000000000000 : node63;
													assign node63 = (inp[5]) ? 14'b00000000000000 : 14'b00100000000011;
									assign node68 = (inp[3]) ? 14'b00000000000000 : node69;
										assign node69 = (inp[4]) ? 14'b00000000000000 : node70;
											assign node70 = (inp[0]) ? node74 : node71;
												assign node71 = (inp[6]) ? 14'b00001000000101 : 14'b00000000000000;
												assign node74 = (inp[6]) ? 14'b00000000000000 : node75;
													assign node75 = (inp[5]) ? 14'b00000000000000 : 14'b00100000000011;
								assign node81 = (inp[6]) ? 14'b00000000000000 : node82;
									assign node82 = (inp[1]) ? node84 : 14'b00000000000000;
										assign node84 = (inp[0]) ? node86 : 14'b00000000000000;
											assign node86 = (inp[3]) ? 14'b00000000000000 : node87;
												assign node87 = (inp[7]) ? 14'b00100000000011 : node88;
													assign node88 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node95 = (inp[6]) ? node121 : node96;
							assign node96 = (inp[1]) ? node98 : 14'b00000000000000;
								assign node98 = (inp[2]) ? 14'b00000000000000 : node99;
									assign node99 = (inp[0]) ? node111 : node100;
										assign node100 = (inp[9]) ? node106 : node101;
											assign node101 = (inp[3]) ? node103 : 14'b00100000000011;
												assign node103 = (inp[7]) ? 14'b00000000000000 : 14'b00001000000000;
											assign node106 = (inp[3]) ? node108 : 14'b00000000000000;
												assign node108 = (inp[7]) ? 14'b00000000000000 : 14'b00001000000101;
										assign node111 = (inp[9]) ? 14'b00000000000000 : node112;
											assign node112 = (inp[3]) ? 14'b00000000000000 : node113;
												assign node113 = (inp[5]) ? 14'b00000000000000 : node114;
													assign node114 = (inp[4]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node121 = (inp[9]) ? node135 : node122;
								assign node122 = (inp[7]) ? node124 : 14'b00000000000000;
									assign node124 = (inp[3]) ? 14'b00000000000000 : node125;
										assign node125 = (inp[1]) ? node127 : 14'b00000000000000;
											assign node127 = (inp[2]) ? 14'b00000000000000 : node128;
												assign node128 = (inp[0]) ? 14'b00000000000000 : node129;
													assign node129 = (inp[4]) ? 14'b10100100111111 : 14'b00000000000000;
								assign node135 = (inp[3]) ? node137 : 14'b00000000000000;
									assign node137 = (inp[1]) ? 14'b00000000000000 : 14'b11110111110010;
				assign node140 = (inp[1]) ? node154 : node141;
					assign node141 = (inp[3]) ? node143 : 14'b00000000000000;
						assign node143 = (inp[6]) ? node145 : 14'b00000000000000;
							assign node145 = (inp[12]) ? node147 : 14'b00000000000000;
								assign node147 = (inp[8]) ? node151 : node148;
									assign node148 = (inp[9]) ? 14'b00000000000000 : 14'b01100000001010;
									assign node151 = (inp[9]) ? 14'b10100010001100 : 14'b00000000000000;
					assign node154 = (inp[9]) ? node208 : node155;
						assign node155 = (inp[3]) ? node187 : node156;
							assign node156 = (inp[12]) ? node174 : node157;
								assign node157 = (inp[8]) ? node167 : node158;
									assign node158 = (inp[2]) ? node160 : 14'b00000000000000;
										assign node160 = (inp[6]) ? 14'b00000000000000 : node161;
											assign node161 = (inp[0]) ? node163 : 14'b00000000000000;
												assign node163 = (inp[4]) ? 14'b00000000000000 : 14'b00100000000011;
									assign node167 = (inp[6]) ? node169 : 14'b01001000000100;
										assign node169 = (inp[5]) ? 14'b00000000000000 : node170;
											assign node170 = (inp[7]) ? 14'b00000000000000 : 14'b11000000000100;
								assign node174 = (inp[6]) ? node178 : node175;
									assign node175 = (inp[8]) ? 14'b00100100011111 : 14'b10000100011000;
									assign node178 = (inp[8]) ? 14'b01000100000100 : node179;
										assign node179 = (inp[2]) ? 14'b00000000000000 : node180;
											assign node180 = (inp[5]) ? node182 : 14'b00000000000000;
												assign node182 = (inp[0]) ? 14'b00000000000000 : 14'b10100000001000;
							assign node187 = (inp[6]) ? 14'b00000000000000 : node188;
								assign node188 = (inp[2]) ? 14'b00000000000000 : node189;
									assign node189 = (inp[0]) ? 14'b00000000000000 : node190;
										assign node190 = (inp[7]) ? node196 : node191;
											assign node191 = (inp[8]) ? node193 : 14'b00000000000000;
												assign node193 = (inp[12]) ? 14'b00000000000000 : 14'b00000100000001;
											assign node196 = (inp[8]) ? 14'b00000000000000 : node197;
												assign node197 = (inp[12]) ? node201 : node198;
													assign node198 = (inp[5]) ? 14'b10010000001101 : 14'b00000000000000;
													assign node201 = (inp[5]) ? 14'b01001000000100 : 14'b01001000000101;
						assign node208 = (inp[3]) ? node222 : node209;
							assign node209 = (inp[6]) ? 14'b00000000000000 : node210;
								assign node210 = (inp[2]) ? 14'b00000000000000 : node211;
									assign node211 = (inp[8]) ? 14'b00000000000000 : node212;
										assign node212 = (inp[7]) ? node214 : 14'b00000000000000;
											assign node214 = (inp[0]) ? 14'b00000000000000 : node215;
												assign node215 = (inp[12]) ? 14'b01001000000100 : 14'b10010000001101;
							assign node222 = (inp[6]) ? node244 : node223;
								assign node223 = (inp[2]) ? 14'b00000000000000 : node224;
									assign node224 = (inp[0]) ? 14'b00000000000000 : node225;
										assign node225 = (inp[7]) ? node235 : node226;
											assign node226 = (inp[8]) ? node228 : 14'b00000000000000;
												assign node228 = (inp[5]) ? node232 : node229;
													assign node229 = (inp[12]) ? 14'b00000000000000 : 14'b00000100000001;
													assign node232 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
											assign node235 = (inp[12]) ? node239 : node236;
												assign node236 = (inp[8]) ? 14'b00000000000000 : 14'b10010000001101;
												assign node239 = (inp[8]) ? 14'b00000000000000 : 14'b01001000000100;
								assign node244 = (inp[7]) ? node252 : node245;
									assign node245 = (inp[12]) ? node247 : 14'b00000000000000;
										assign node247 = (inp[8]) ? 14'b00000000000000 : node248;
											assign node248 = (inp[5]) ? 14'b01001000001100 : 14'b00000000000000;
									assign node252 = (inp[12]) ? node262 : node253;
										assign node253 = (inp[5]) ? 14'b00000000000000 : node254;
											assign node254 = (inp[8]) ? 14'b01100000001010 : node255;
												assign node255 = (inp[0]) ? 14'b01001000000100 : node256;
													assign node256 = (inp[4]) ? 14'b10100000101010 : 14'b10100000111010;
										assign node262 = (inp[5]) ? node264 : 14'b00000000000000;
											assign node264 = (inp[8]) ? 14'b10000000011010 : 14'b00000000000000;
			assign node267 = (inp[12]) ? node395 : node268;
				assign node268 = (inp[1]) ? node296 : node269;
					assign node269 = (inp[8]) ? node281 : node270;
						assign node270 = (inp[7]) ? 14'b00000000000000 : node271;
							assign node271 = (inp[6]) ? node273 : 14'b00000000000000;
								assign node273 = (inp[11]) ? 14'b00000000000000 : node274;
									assign node274 = (inp[3]) ? node276 : 14'b00000000000000;
										assign node276 = (inp[9]) ? 14'b00000000000000 : 14'b11000000000100;
						assign node281 = (inp[6]) ? node283 : 14'b00000000000000;
							assign node283 = (inp[0]) ? 14'b00000000000000 : node284;
								assign node284 = (inp[2]) ? 14'b00000000000000 : node285;
									assign node285 = (inp[11]) ? node287 : 14'b00000000000000;
										assign node287 = (inp[7]) ? 14'b00000000000000 : node288;
											assign node288 = (inp[3]) ? node290 : 14'b00000000000000;
												assign node290 = (inp[9]) ? 14'b00000000000000 : 14'b00100000000011;
					assign node296 = (inp[11]) ? node342 : node297;
						assign node297 = (inp[8]) ? node319 : node298;
							assign node298 = (inp[9]) ? node304 : node299;
								assign node299 = (inp[6]) ? 14'b00000000000000 : node300;
									assign node300 = (inp[3]) ? 14'b00000000000000 : 14'b11000000000100;
								assign node304 = (inp[7]) ? node306 : 14'b00000000000000;
									assign node306 = (inp[5]) ? 14'b00000000000000 : node307;
										assign node307 = (inp[6]) ? node309 : 14'b00000000000000;
											assign node309 = (inp[3]) ? node311 : 14'b00000000000000;
												assign node311 = (inp[2]) ? node315 : node312;
													assign node312 = (inp[0]) ? 14'b01100000000110 : 14'b00001000000101;
													assign node315 = (inp[4]) ? 14'b00000000000000 : 14'b01100000000110;
							assign node319 = (inp[4]) ? 14'b00000000000000 : node320;
								assign node320 = (inp[7]) ? node322 : 14'b00000000000000;
									assign node322 = (inp[2]) ? 14'b00000000000000 : node323;
										assign node323 = (inp[3]) ? node331 : node324;
											assign node324 = (inp[9]) ? 14'b00000000000000 : node325;
												assign node325 = (inp[6]) ? 14'b00000000000000 : node326;
													assign node326 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
											assign node331 = (inp[0]) ? 14'b00000000000000 : node332;
												assign node332 = (inp[5]) ? node336 : node333;
													assign node333 = (inp[9]) ? 14'b00000000011100 : 14'b00000000000000;
													assign node336 = (inp[6]) ? 14'b00000000000000 : 14'b10000000111000;
						assign node342 = (inp[6]) ? node382 : node343;
							assign node343 = (inp[9]) ? node369 : node344;
								assign node344 = (inp[8]) ? node360 : node345;
									assign node345 = (inp[3]) ? node353 : node346;
										assign node346 = (inp[0]) ? node348 : 14'b00000000000000;
											assign node348 = (inp[4]) ? 14'b00000000000000 : node349;
												assign node349 = (inp[5]) ? 14'b00000000000000 : 14'b01001000000100;
										assign node353 = (inp[2]) ? 14'b00000000000000 : node354;
											assign node354 = (inp[0]) ? 14'b00000000000000 : node355;
												assign node355 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
									assign node360 = (inp[3]) ? node362 : 14'b00000000011100;
										assign node362 = (inp[2]) ? 14'b00000000000000 : node363;
											assign node363 = (inp[7]) ? 14'b00000000000000 : node364;
												assign node364 = (inp[0]) ? 14'b00000000000000 : 14'b00000000011100;
								assign node369 = (inp[2]) ? 14'b00000000000000 : node370;
									assign node370 = (inp[3]) ? node372 : 14'b00000000000000;
										assign node372 = (inp[0]) ? 14'b00000000000000 : node373;
											assign node373 = (inp[8]) ? node377 : node374;
												assign node374 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
												assign node377 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node382 = (inp[7]) ? node384 : 14'b00000000000000;
								assign node384 = (inp[3]) ? node386 : 14'b00000000000000;
									assign node386 = (inp[9]) ? node388 : 14'b00000000000000;
										assign node388 = (inp[5]) ? node392 : node389;
											assign node389 = (inp[8]) ? 14'b10100010001100 : 14'b10000010001100;
											assign node392 = (inp[8]) ? 14'b00000000000000 : 14'b01001000000101;
				assign node395 = (inp[8]) ? node489 : node396;
					assign node396 = (inp[3]) ? node440 : node397;
						assign node397 = (inp[1]) ? node399 : 14'b00000000000000;
							assign node399 = (inp[6]) ? node429 : node400;
								assign node400 = (inp[2]) ? node420 : node401;
									assign node401 = (inp[7]) ? node413 : node402;
										assign node402 = (inp[0]) ? node404 : 14'b00000000000000;
											assign node404 = (inp[5]) ? 14'b00000000000000 : node405;
												assign node405 = (inp[11]) ? node409 : node406;
													assign node406 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
													assign node409 = (inp[4]) ? 14'b00000000000000 : 14'b01001000000101;
										assign node413 = (inp[9]) ? node415 : 14'b00000000000000;
											assign node415 = (inp[0]) ? 14'b00000000000000 : node416;
												assign node416 = (inp[11]) ? 14'b10100010001100 : 14'b11110111110010;
									assign node420 = (inp[11]) ? 14'b00000000000000 : node421;
										assign node421 = (inp[0]) ? node423 : 14'b00000000000000;
											assign node423 = (inp[4]) ? 14'b00000000000000 : node424;
												assign node424 = (inp[9]) ? 14'b00000000000000 : 14'b10000000101100;
								assign node429 = (inp[0]) ? 14'b00000000000000 : node430;
									assign node430 = (inp[9]) ? 14'b00000000000000 : node431;
										assign node431 = (inp[2]) ? 14'b00000000000000 : node432;
											assign node432 = (inp[5]) ? node434 : 14'b00000000000000;
												assign node434 = (inp[11]) ? 14'b00001000000001 : 14'b01001000000101;
						assign node440 = (inp[6]) ? node456 : node441;
							assign node441 = (inp[2]) ? 14'b00000000000000 : node442;
								assign node442 = (inp[0]) ? 14'b00000000000000 : node443;
									assign node443 = (inp[7]) ? node445 : 14'b00000000000000;
										assign node445 = (inp[1]) ? node447 : 14'b00000000000000;
											assign node447 = (inp[11]) ? 14'b10100010001100 : node448;
												assign node448 = (inp[9]) ? 14'b11110111110010 : node449;
													assign node449 = (inp[4]) ? 14'b11110111110010 : 14'b00000000000000;
							assign node456 = (inp[11]) ? node478 : node457;
								assign node457 = (inp[7]) ? 14'b00000000000000 : node458;
									assign node458 = (inp[5]) ? node466 : node459;
										assign node459 = (inp[2]) ? 14'b00000000000000 : node460;
											assign node460 = (inp[4]) ? node462 : 14'b00000000000000;
												assign node462 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
										assign node466 = (inp[9]) ? node474 : node467;
											assign node467 = (inp[2]) ? 14'b00000000000000 : node468;
												assign node468 = (inp[0]) ? 14'b00000000000000 : node469;
													assign node469 = (inp[1]) ? 14'b00000000000000 : 14'b00000000011100;
											assign node474 = (inp[1]) ? 14'b00000000011101 : 14'b00000000000000;
								assign node478 = (inp[9]) ? node482 : node479;
									assign node479 = (inp[1]) ? 14'b00000000000000 : 14'b00100100001101;
									assign node482 = (inp[5]) ? node484 : 14'b00000000000000;
										assign node484 = (inp[1]) ? node486 : 14'b00000000000000;
											assign node486 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
					assign node489 = (inp[11]) ? 14'b01000000010100 : node490;
						assign node490 = (inp[6]) ? node510 : node491;
							assign node491 = (inp[1]) ? node493 : 14'b00000000000000;
								assign node493 = (inp[0]) ? 14'b00000000000000 : node494;
									assign node494 = (inp[2]) ? 14'b00000000000000 : node495;
										assign node495 = (inp[7]) ? node503 : node496;
											assign node496 = (inp[3]) ? node500 : node497;
												assign node497 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
												assign node500 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
											assign node503 = (inp[9]) ? 14'b00000000000000 : node504;
												assign node504 = (inp[3]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node510 = (inp[3]) ? node528 : node511;
								assign node511 = (inp[9]) ? 14'b00000000000000 : node512;
									assign node512 = (inp[1]) ? node514 : 14'b00000000000000;
										assign node514 = (inp[5]) ? node524 : node515;
											assign node515 = (inp[7]) ? node517 : 14'b10010100011100;
												assign node517 = (inp[0]) ? node521 : node518;
													assign node518 = (inp[2]) ? 14'b00000000000000 : 14'b10010010001100;
													assign node521 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
											assign node524 = (inp[7]) ? 14'b11100100010100 : 14'b11100100000100;
								assign node528 = (inp[9]) ? node530 : 14'b00000000000000;
									assign node530 = (inp[1]) ? node532 : 14'b01001000000100;
										assign node532 = (inp[7]) ? node534 : 14'b00000000000000;
											assign node534 = (inp[5]) ? 14'b01001000001001 : 14'b00000000000000;
		assign node538 = (inp[1]) ? node626 : node539;
			assign node539 = (inp[6]) ? node555 : node540;
				assign node540 = (inp[11]) ? node548 : node541;
					assign node541 = (inp[12]) ? 14'b00000000000000 : node542;
						assign node542 = (inp[13]) ? 14'b00000000000000 : node543;
							assign node543 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
					assign node548 = (inp[8]) ? node550 : 14'b00000000000000;
						assign node550 = (inp[13]) ? node552 : 14'b00000000000000;
							assign node552 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
				assign node555 = (inp[12]) ? node577 : node556;
					assign node556 = (inp[8]) ? node562 : node557;
						assign node557 = (inp[11]) ? 14'b00000000000000 : node558;
							assign node558 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
						assign node562 = (inp[13]) ? node564 : 14'b00000000000000;
							assign node564 = (inp[7]) ? 14'b00000000000000 : node565;
								assign node565 = (inp[3]) ? node567 : 14'b00000000000000;
									assign node567 = (inp[9]) ? 14'b00000000000000 : node568;
										assign node568 = (inp[2]) ? 14'b00000000000000 : node569;
											assign node569 = (inp[0]) ? 14'b00000000000000 : node570;
												assign node570 = (inp[5]) ? 14'b10000100111010 : 14'b10000100101010;
					assign node577 = (inp[13]) ? node601 : node578;
						assign node578 = (inp[3]) ? node580 : 14'b00000000000000;
							assign node580 = (inp[11]) ? node596 : node581;
								assign node581 = (inp[8]) ? node593 : node582;
									assign node582 = (inp[7]) ? 14'b00000000000000 : node583;
										assign node583 = (inp[0]) ? 14'b00000000000000 : node584;
											assign node584 = (inp[9]) ? 14'b00000000000000 : node585;
												assign node585 = (inp[2]) ? 14'b00000000000000 : node586;
													assign node586 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
									assign node593 = (inp[9]) ? 14'b01100000001010 : 14'b00000000000000;
								assign node596 = (inp[8]) ? 14'b00000000000000 : node597;
									assign node597 = (inp[9]) ? 14'b00000000000000 : 14'b01001000000101;
						assign node601 = (inp[11]) ? node619 : node602;
							assign node602 = (inp[3]) ? node604 : 14'b00000000000000;
								assign node604 = (inp[9]) ? node616 : node605;
									assign node605 = (inp[8]) ? 14'b00000000000000 : node606;
										assign node606 = (inp[0]) ? 14'b00000000000000 : node607;
											assign node607 = (inp[2]) ? 14'b00000000000000 : node608;
												assign node608 = (inp[7]) ? 14'b00000000000000 : node609;
													assign node609 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
									assign node616 = (inp[8]) ? 14'b00100100001101 : 14'b00000000000000;
							assign node619 = (inp[8]) ? 14'b10000100001000 : node620;
								assign node620 = (inp[9]) ? 14'b00000000000000 : node621;
									assign node621 = (inp[3]) ? 14'b10010101111110 : 14'b00000000000000;
			assign node626 = (inp[2]) ? node1044 : node627;
				assign node627 = (inp[6]) ? node875 : node628;
					assign node628 = (inp[0]) ? node752 : node629;
						assign node629 = (inp[8]) ? node675 : node630;
							assign node630 = (inp[11]) ? node652 : node631;
								assign node631 = (inp[13]) ? node635 : node632;
									assign node632 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node635 = (inp[12]) ? node641 : node636;
										assign node636 = (inp[9]) ? node638 : 14'b00000000000000;
											assign node638 = (inp[7]) ? 14'b00001000000100 : 14'b00000000000000;
										assign node641 = (inp[7]) ? node647 : node642;
											assign node642 = (inp[3]) ? 14'b00000000000000 : node643;
												assign node643 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011101;
											assign node647 = (inp[3]) ? 14'b01100000001010 : node648;
												assign node648 = (inp[9]) ? 14'b01100000001010 : 14'b00000000011101;
								assign node652 = (inp[3]) ? node662 : node653;
									assign node653 = (inp[13]) ? 14'b00000000000000 : node654;
										assign node654 = (inp[9]) ? node656 : 14'b00000000000000;
											assign node656 = (inp[7]) ? node658 : 14'b00000000000000;
												assign node658 = (inp[12]) ? 14'b00100100001101 : 14'b00000000000000;
									assign node662 = (inp[12]) ? node670 : node663;
										assign node663 = (inp[7]) ? node665 : 14'b00100000000011;
											assign node665 = (inp[5]) ? node667 : 14'b00000000000000;
												assign node667 = (inp[9]) ? 14'b00000000000000 : 14'b00100000000011;
										assign node670 = (inp[13]) ? 14'b00000000000000 : node671;
											assign node671 = (inp[7]) ? 14'b00100100001101 : 14'b00000000000000;
							assign node675 = (inp[13]) ? node715 : node676;
								assign node676 = (inp[9]) ? node704 : node677;
									assign node677 = (inp[3]) ? node689 : node678;
										assign node678 = (inp[11]) ? node684 : node679;
											assign node679 = (inp[12]) ? node681 : 14'b00100000000011;
												assign node681 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
											assign node684 = (inp[12]) ? 14'b00000000000000 : node685;
												assign node685 = (inp[4]) ? 14'b10000010001101 : 14'b10000001001101;
										assign node689 = (inp[11]) ? node699 : node690;
											assign node690 = (inp[12]) ? node696 : node691;
												assign node691 = (inp[7]) ? node693 : 14'b00000000000000;
													assign node693 = (inp[5]) ? 14'b00000000011100 : 14'b00000000000000;
												assign node696 = (inp[7]) ? 14'b00000000000000 : 14'b00000000011100;
											assign node699 = (inp[7]) ? 14'b00000000000000 : node700;
												assign node700 = (inp[12]) ? 14'b00000000000000 : 14'b00100000001010;
									assign node704 = (inp[7]) ? 14'b00000000000000 : node705;
										assign node705 = (inp[3]) ? node707 : 14'b00000000000000;
											assign node707 = (inp[11]) ? node711 : node708;
												assign node708 = (inp[12]) ? 14'b00000000011100 : 14'b00000000000000;
												assign node711 = (inp[12]) ? 14'b00000000000000 : 14'b00100000001010;
								assign node715 = (inp[11]) ? node741 : node716;
									assign node716 = (inp[7]) ? node732 : node717;
										assign node717 = (inp[3]) ? node725 : node718;
											assign node718 = (inp[9]) ? 14'b00000000000000 : node719;
												assign node719 = (inp[12]) ? node721 : 14'b00000000000000;
													assign node721 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
											assign node725 = (inp[12]) ? node727 : 14'b00001000001001;
												assign node727 = (inp[9]) ? node729 : 14'b00000000000000;
													assign node729 = (inp[5]) ? 14'b00000000011101 : 14'b00000000000000;
										assign node732 = (inp[12]) ? node734 : 14'b00000000000000;
											assign node734 = (inp[3]) ? 14'b00000000000000 : node735;
												assign node735 = (inp[9]) ? 14'b00000000000000 : node736;
													assign node736 = (inp[5]) ? 14'b10000000101000 : 14'b10000000111000;
									assign node741 = (inp[12]) ? 14'b10000100001000 : node742;
										assign node742 = (inp[3]) ? node746 : node743;
											assign node743 = (inp[9]) ? 14'b00000000000000 : 14'b10000000001010;
											assign node746 = (inp[7]) ? 14'b00000000000000 : node747;
												assign node747 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
						assign node752 = (inp[3]) ? node824 : node753;
							assign node753 = (inp[9]) ? node809 : node754;
								assign node754 = (inp[12]) ? node782 : node755;
									assign node755 = (inp[8]) ? node765 : node756;
										assign node756 = (inp[13]) ? 14'b00000000000000 : node757;
											assign node757 = (inp[11]) ? node759 : 14'b10000100001000;
												assign node759 = (inp[7]) ? node761 : 14'b00000000000000;
													assign node761 = (inp[5]) ? 14'b00000000000000 : 14'b01100000001010;
										assign node765 = (inp[11]) ? node775 : node766;
											assign node766 = (inp[7]) ? node768 : 14'b00000000000000;
												assign node768 = (inp[13]) ? node772 : node769;
													assign node769 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
													assign node772 = (inp[5]) ? 14'b00000000000000 : 14'b10110111101111;
											assign node775 = (inp[13]) ? 14'b10100100011000 : node776;
												assign node776 = (inp[4]) ? 14'b10000000011101 : node777;
													assign node777 = (inp[5]) ? 14'b00000000000000 : 14'b10100000001101;
									assign node782 = (inp[11]) ? node796 : node783;
										assign node783 = (inp[13]) ? node793 : node784;
											assign node784 = (inp[8]) ? node788 : node785;
												assign node785 = (inp[4]) ? 14'b00000000000000 : 14'b01001000000100;
												assign node788 = (inp[4]) ? 14'b00000000000000 : node789;
													assign node789 = (inp[5]) ? 14'b00000000000000 : 14'b10000100011000;
											assign node793 = (inp[8]) ? 14'b00001000000100 : 14'b00000000011101;
										assign node796 = (inp[13]) ? node804 : node797;
											assign node797 = (inp[4]) ? 14'b00000000000000 : node798;
												assign node798 = (inp[8]) ? 14'b00000000000000 : node799;
													assign node799 = (inp[5]) ? 14'b00000000000000 : 14'b00001000000101;
											assign node804 = (inp[8]) ? 14'b10000100001000 : node805;
												assign node805 = (inp[4]) ? 14'b00000000000000 : 14'b10000000001111;
								assign node809 = (inp[13]) ? node817 : node810;
									assign node810 = (inp[8]) ? 14'b00000000000000 : node811;
										assign node811 = (inp[11]) ? 14'b00000000000000 : node812;
											assign node812 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node817 = (inp[11]) ? node819 : 14'b00000000000000;
										assign node819 = (inp[8]) ? node821 : 14'b00000000000000;
											assign node821 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node824 = (inp[4]) ? node856 : node825;
								assign node825 = (inp[7]) ? node841 : node826;
									assign node826 = (inp[11]) ? node834 : node827;
										assign node827 = (inp[8]) ? 14'b00000000000000 : node828;
											assign node828 = (inp[13]) ? 14'b00000000000000 : node829;
												assign node829 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node834 = (inp[13]) ? node836 : 14'b00000000000000;
											assign node836 = (inp[12]) ? node838 : 14'b00000000000000;
												assign node838 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node841 = (inp[11]) ? node849 : node842;
										assign node842 = (inp[13]) ? 14'b00000000000000 : node843;
											assign node843 = (inp[8]) ? 14'b00000000000000 : node844;
												assign node844 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node849 = (inp[13]) ? node851 : 14'b00000000000000;
											assign node851 = (inp[8]) ? node853 : 14'b00000000000000;
												assign node853 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node856 = (inp[9]) ? node866 : node857;
									assign node857 = (inp[8]) ? node859 : 14'b00000000000000;
										assign node859 = (inp[11]) ? node861 : 14'b00000000000000;
											assign node861 = (inp[12]) ? node863 : 14'b00000000000000;
												assign node863 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node866 = (inp[13]) ? 14'b00000000000000 : node867;
										assign node867 = (inp[8]) ? 14'b00000000000000 : node868;
											assign node868 = (inp[11]) ? 14'b00000000000000 : node869;
												assign node869 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
					assign node875 = (inp[3]) ? node921 : node876;
						assign node876 = (inp[11]) ? node904 : node877;
							assign node877 = (inp[13]) ? node891 : node878;
								assign node878 = (inp[8]) ? 14'b00000000000000 : node879;
									assign node879 = (inp[12]) ? node881 : 14'b10000100001000;
										assign node881 = (inp[5]) ? node883 : 14'b00000000000000;
											assign node883 = (inp[7]) ? node885 : 14'b00000000000000;
												assign node885 = (inp[9]) ? 14'b00000000000000 : node886;
													assign node886 = (inp[0]) ? 14'b00000000000000 : 14'b00000100001101;
								assign node891 = (inp[12]) ? node893 : 14'b00000000000000;
									assign node893 = (inp[8]) ? node901 : node894;
										assign node894 = (inp[9]) ? 14'b00000000000000 : node895;
											assign node895 = (inp[4]) ? 14'b00000000000000 : node896;
												assign node896 = (inp[7]) ? 14'b00000000011100 : 14'b00000000000000;
										assign node901 = (inp[9]) ? 14'b00000000000000 : 14'b00000100001110;
							assign node904 = (inp[8]) ? node916 : node905;
								assign node905 = (inp[7]) ? node907 : 14'b00000000000000;
									assign node907 = (inp[12]) ? node909 : 14'b00000000000000;
										assign node909 = (inp[5]) ? node911 : 14'b00000000000000;
											assign node911 = (inp[0]) ? 14'b00000000000000 : node912;
												assign node912 = (inp[9]) ? 14'b00000000000000 : 14'b01001000000101;
								assign node916 = (inp[13]) ? node918 : 14'b00000000000000;
									assign node918 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node921 = (inp[9]) ? node971 : node922;
							assign node922 = (inp[5]) ? node956 : node923;
								assign node923 = (inp[4]) ? node941 : node924;
									assign node924 = (inp[7]) ? node934 : node925;
										assign node925 = (inp[8]) ? 14'b00000000000000 : node926;
											assign node926 = (inp[11]) ? 14'b00000000000000 : node927;
												assign node927 = (inp[12]) ? 14'b00000000000000 : node928;
													assign node928 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node934 = (inp[8]) ? node936 : 14'b00000000000000;
											assign node936 = (inp[11]) ? node938 : 14'b00000000000000;
												assign node938 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node941 = (inp[13]) ? node949 : node942;
										assign node942 = (inp[8]) ? 14'b00000000000000 : node943;
											assign node943 = (inp[11]) ? 14'b00000000000000 : node944;
												assign node944 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node949 = (inp[8]) ? node951 : 14'b00000000000000;
											assign node951 = (inp[12]) ? node953 : 14'b00000000000000;
												assign node953 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node956 = (inp[8]) ? node964 : node957;
									assign node957 = (inp[12]) ? 14'b00000000000000 : node958;
										assign node958 = (inp[11]) ? 14'b00000000000000 : node959;
											assign node959 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node964 = (inp[11]) ? node966 : 14'b00000000000000;
										assign node966 = (inp[12]) ? node968 : 14'b00000000000000;
											assign node968 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node971 = (inp[11]) ? node1005 : node972;
								assign node972 = (inp[12]) ? node992 : node973;
									assign node973 = (inp[13]) ? node983 : node974;
										assign node974 = (inp[8]) ? node976 : 14'b10000100001000;
											assign node976 = (inp[7]) ? node978 : 14'b00000000000000;
												assign node978 = (inp[5]) ? 14'b10100000001000 : node979;
													assign node979 = (inp[0]) ? 14'b00000000000000 : 14'b00100000001010;
										assign node983 = (inp[5]) ? 14'b00000000000000 : node984;
											assign node984 = (inp[7]) ? node986 : 14'b00000000000000;
												assign node986 = (inp[0]) ? 14'b00000000000000 : node987;
													assign node987 = (inp[8]) ? 14'b10000100111000 : 14'b00000000011101;
									assign node992 = (inp[5]) ? node994 : 14'b00000000000000;
										assign node994 = (inp[8]) ? node1000 : node995;
											assign node995 = (inp[7]) ? 14'b00000000000000 : node996;
												assign node996 = (inp[13]) ? 14'b10100000001000 : 14'b00001000001100;
											assign node1000 = (inp[7]) ? node1002 : 14'b00000000000000;
												assign node1002 = (inp[13]) ? 14'b00000000011100 : 14'b01100000000110;
								assign node1005 = (inp[13]) ? node1025 : node1006;
									assign node1006 = (inp[8]) ? node1020 : node1007;
										assign node1007 = (inp[7]) ? node1013 : node1008;
											assign node1008 = (inp[12]) ? node1010 : 14'b00000000000000;
												assign node1010 = (inp[5]) ? 14'b00000100001111 : 14'b00000000000000;
											assign node1013 = (inp[12]) ? 14'b00000000000000 : node1014;
												assign node1014 = (inp[5]) ? 14'b00000000000000 : node1015;
													assign node1015 = (inp[0]) ? 14'b00000100001111 : 14'b00100000000011;
										assign node1020 = (inp[5]) ? 14'b00000000000000 : node1021;
											assign node1021 = (inp[7]) ? 14'b01001000000100 : 14'b00000000000000;
									assign node1025 = (inp[12]) ? node1037 : node1026;
										assign node1026 = (inp[7]) ? node1028 : 14'b00000000000000;
											assign node1028 = (inp[8]) ? node1034 : node1029;
												assign node1029 = (inp[5]) ? 14'b10100101111111 : node1030;
													assign node1030 = (inp[0]) ? 14'b01000100000010 : 14'b00001000001001;
												assign node1034 = (inp[5]) ? 14'b00000000000000 : 14'b00100100001101;
										assign node1037 = (inp[8]) ? 14'b10000100001000 : node1038;
											assign node1038 = (inp[5]) ? node1040 : 14'b00000000000000;
												assign node1040 = (inp[7]) ? 14'b00000000000000 : 14'b10100100001000;
				assign node1044 = (inp[13]) ? node1174 : node1045;
					assign node1045 = (inp[12]) ? node1129 : node1046;
						assign node1046 = (inp[11]) ? node1072 : node1047;
							assign node1047 = (inp[8]) ? node1049 : 14'b10000100001000;
								assign node1049 = (inp[9]) ? node1061 : node1050;
									assign node1050 = (inp[6]) ? 14'b00000000000000 : node1051;
										assign node1051 = (inp[3]) ? 14'b00000000000000 : node1052;
											assign node1052 = (inp[4]) ? node1056 : node1053;
												assign node1053 = (inp[0]) ? 14'b00100000000011 : 14'b00000000000000;
												assign node1056 = (inp[0]) ? 14'b00000000000000 : 14'b00100000000011;
									assign node1061 = (inp[3]) ? node1063 : 14'b00000000000000;
										assign node1063 = (inp[6]) ? node1065 : 14'b00000000000000;
											assign node1065 = (inp[7]) ? node1067 : 14'b00000000000000;
												assign node1067 = (inp[5]) ? 14'b10100000001000 : node1068;
													assign node1068 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
							assign node1072 = (inp[7]) ? node1090 : node1073;
								assign node1073 = (inp[6]) ? 14'b00000000000000 : node1074;
									assign node1074 = (inp[3]) ? 14'b00000000000000 : node1075;
										assign node1075 = (inp[9]) ? 14'b00000000000000 : node1076;
											assign node1076 = (inp[0]) ? node1082 : node1077;
												assign node1077 = (inp[4]) ? node1079 : 14'b00000000000000;
													assign node1079 = (inp[8]) ? 14'b10000100001101 : 14'b00000000000000;
												assign node1082 = (inp[4]) ? 14'b00000000000000 : node1083;
													assign node1083 = (inp[8]) ? 14'b10010000001101 : 14'b01001000000101;
								assign node1090 = (inp[5]) ? node1106 : node1091;
									assign node1091 = (inp[3]) ? node1099 : node1092;
										assign node1092 = (inp[9]) ? 14'b00000000000000 : node1093;
											assign node1093 = (inp[8]) ? node1095 : 14'b00000000000000;
												assign node1095 = (inp[4]) ? 14'b00000000000000 : 14'b10010000001101;
										assign node1099 = (inp[9]) ? node1101 : 14'b00000000000000;
											assign node1101 = (inp[6]) ? node1103 : 14'b00000000000000;
												assign node1103 = (inp[8]) ? 14'b01001000000100 : 14'b00000100001111;
									assign node1106 = (inp[9]) ? node1120 : node1107;
										assign node1107 = (inp[6]) ? 14'b00000000000000 : node1108;
											assign node1108 = (inp[8]) ? node1114 : node1109;
												assign node1109 = (inp[3]) ? 14'b00000000000000 : node1110;
													assign node1110 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
												assign node1114 = (inp[4]) ? 14'b10000100001101 : node1115;
													assign node1115 = (inp[0]) ? 14'b10010000001101 : 14'b00000000000000;
										assign node1120 = (inp[4]) ? node1122 : 14'b00000000000000;
											assign node1122 = (inp[8]) ? 14'b00000000000000 : node1123;
												assign node1123 = (inp[3]) ? node1125 : 14'b00000000000000;
													assign node1125 = (inp[0]) ? 14'b00100000000011 : 14'b00000000000000;
						assign node1129 = (inp[5]) ? node1145 : node1130;
							assign node1130 = (inp[11]) ? 14'b00000000000000 : node1131;
								assign node1131 = (inp[7]) ? node1133 : 14'b00000000000000;
									assign node1133 = (inp[9]) ? 14'b00000000000000 : node1134;
										assign node1134 = (inp[0]) ? node1136 : 14'b00000000000000;
											assign node1136 = (inp[8]) ? 14'b00000000000000 : node1137;
												assign node1137 = (inp[3]) ? 14'b00000000000000 : node1138;
													assign node1138 = (inp[6]) ? 14'b00000000000000 : 14'b01001000000100;
							assign node1145 = (inp[3]) ? node1159 : node1146;
								assign node1146 = (inp[9]) ? 14'b00000000000000 : node1147;
									assign node1147 = (inp[4]) ? 14'b00000000000000 : node1148;
										assign node1148 = (inp[8]) ? 14'b00000000000000 : node1149;
											assign node1149 = (inp[6]) ? 14'b00000000000000 : node1150;
												assign node1150 = (inp[11]) ? 14'b00000000000000 : node1151;
													assign node1151 = (inp[0]) ? 14'b01001000000100 : 14'b00000000000000;
								assign node1159 = (inp[9]) ? node1161 : 14'b00000000000000;
									assign node1161 = (inp[6]) ? node1163 : 14'b00000000000000;
										assign node1163 = (inp[8]) ? node1169 : node1164;
											assign node1164 = (inp[7]) ? 14'b00000000000000 : node1165;
												assign node1165 = (inp[11]) ? 14'b00000100001111 : 14'b00001000001100;
											assign node1169 = (inp[7]) ? node1171 : 14'b00000000000000;
												assign node1171 = (inp[11]) ? 14'b00000000000000 : 14'b01100000000110;
					assign node1174 = (inp[12]) ? node1224 : node1175;
						assign node1175 = (inp[11]) ? node1177 : 14'b00000000000000;
							assign node1177 = (inp[7]) ? node1195 : node1178;
								assign node1178 = (inp[9]) ? 14'b00000000000000 : node1179;
									assign node1179 = (inp[3]) ? 14'b00000000000000 : node1180;
										assign node1180 = (inp[6]) ? 14'b00000000000000 : node1181;
											assign node1181 = (inp[8]) ? node1187 : node1182;
												assign node1182 = (inp[0]) ? node1184 : 14'b00000000000000;
													assign node1184 = (inp[4]) ? 14'b00000000000000 : 14'b00000000011100;
												assign node1187 = (inp[4]) ? 14'b10100100011000 : node1188;
													assign node1188 = (inp[0]) ? 14'b10100100011000 : 14'b00000000000000;
								assign node1195 = (inp[3]) ? node1211 : node1196;
									assign node1196 = (inp[9]) ? 14'b00000000000000 : node1197;
										assign node1197 = (inp[6]) ? 14'b00000000000000 : node1198;
											assign node1198 = (inp[8]) ? node1204 : node1199;
												assign node1199 = (inp[4]) ? 14'b00000000000000 : node1200;
													assign node1200 = (inp[0]) ? 14'b00000000011100 : 14'b00000000000000;
												assign node1204 = (inp[4]) ? 14'b10100100011000 : node1205;
													assign node1205 = (inp[5]) ? 14'b00000000000000 : 14'b10100100011000;
									assign node1211 = (inp[9]) ? node1213 : 14'b00000000000000;
										assign node1213 = (inp[6]) ? node1215 : 14'b00000000000000;
											assign node1215 = (inp[8]) ? node1221 : node1216;
												assign node1216 = (inp[5]) ? 14'b10100101111111 : node1217;
													assign node1217 = (inp[4]) ? 14'b01000100000010 : 14'b01100000000010;
												assign node1221 = (inp[5]) ? 14'b00000000000000 : 14'b00100100001101;
						assign node1224 = (inp[8]) ? node1252 : node1225;
							assign node1225 = (inp[11]) ? node1241 : node1226;
								assign node1226 = (inp[6]) ? node1232 : node1227;
									assign node1227 = (inp[3]) ? 14'b00000000000000 : node1228;
										assign node1228 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011101;
									assign node1232 = (inp[9]) ? node1234 : 14'b00000000000000;
										assign node1234 = (inp[5]) ? node1236 : 14'b00000000000000;
											assign node1236 = (inp[7]) ? 14'b00000000000000 : node1237;
												assign node1237 = (inp[3]) ? 14'b10100000001000 : 14'b00000000000000;
								assign node1241 = (inp[5]) ? node1243 : 14'b00000000000000;
									assign node1243 = (inp[6]) ? node1245 : 14'b00000000000000;
										assign node1245 = (inp[9]) ? node1247 : 14'b00000000000000;
											assign node1247 = (inp[7]) ? 14'b00000000000000 : node1248;
												assign node1248 = (inp[3]) ? 14'b10100100001000 : 14'b00000000000000;
							assign node1252 = (inp[11]) ? 14'b10000100001000 : node1253;
								assign node1253 = (inp[3]) ? node1259 : node1254;
									assign node1254 = (inp[9]) ? 14'b00000000000000 : node1255;
										assign node1255 = (inp[6]) ? 14'b00000100001110 : 14'b00001000000100;
									assign node1259 = (inp[5]) ? node1261 : 14'b00000000000000;
										assign node1261 = (inp[9]) ? node1263 : 14'b00000000000000;
											assign node1263 = (inp[7]) ? node1265 : 14'b00000000000000;
												assign node1265 = (inp[6]) ? 14'b00000000011100 : 14'b00000000000000;

endmodule