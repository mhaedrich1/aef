module dtc_split66_bm81 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node317;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node390;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node463;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node548;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node567;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node627;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node655;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node670;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node707;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node722;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node729;
	wire [3-1:0] node731;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node770;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node783;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node795;
	wire [3-1:0] node799;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node823;
	wire [3-1:0] node827;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node845;
	wire [3-1:0] node846;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node853;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node865;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node879;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node901;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node932;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node939;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node945;
	wire [3-1:0] node948;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node969;
	wire [3-1:0] node970;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node980;
	wire [3-1:0] node982;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1002;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1017;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1036;
	wire [3-1:0] node1038;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1069;
	wire [3-1:0] node1071;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1078;
	wire [3-1:0] node1081;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1087;
	wire [3-1:0] node1090;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1103;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1108;
	wire [3-1:0] node1111;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1118;
	wire [3-1:0] node1120;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1130;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1141;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1153;
	wire [3-1:0] node1155;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1162;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1167;
	wire [3-1:0] node1168;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1175;
	wire [3-1:0] node1177;
	wire [3-1:0] node1178;
	wire [3-1:0] node1182;
	wire [3-1:0] node1183;
	wire [3-1:0] node1185;
	wire [3-1:0] node1188;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1195;
	wire [3-1:0] node1196;
	wire [3-1:0] node1200;
	wire [3-1:0] node1202;
	wire [3-1:0] node1205;
	wire [3-1:0] node1206;
	wire [3-1:0] node1209;
	wire [3-1:0] node1211;
	wire [3-1:0] node1213;
	wire [3-1:0] node1216;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1242;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1249;
	wire [3-1:0] node1252;
	wire [3-1:0] node1255;
	wire [3-1:0] node1256;
	wire [3-1:0] node1257;
	wire [3-1:0] node1259;
	wire [3-1:0] node1263;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1269;
	wire [3-1:0] node1270;
	wire [3-1:0] node1275;
	wire [3-1:0] node1276;
	wire [3-1:0] node1278;
	wire [3-1:0] node1279;
	wire [3-1:0] node1280;
	wire [3-1:0] node1286;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1292;
	wire [3-1:0] node1295;
	wire [3-1:0] node1298;
	wire [3-1:0] node1300;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1308;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1315;
	wire [3-1:0] node1318;
	wire [3-1:0] node1319;
	wire [3-1:0] node1320;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1327;
	wire [3-1:0] node1329;
	wire [3-1:0] node1332;
	wire [3-1:0] node1333;
	wire [3-1:0] node1335;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1341;
	wire [3-1:0] node1342;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1350;
	wire [3-1:0] node1351;
	wire [3-1:0] node1353;
	wire [3-1:0] node1357;
	wire [3-1:0] node1358;
	wire [3-1:0] node1360;
	wire [3-1:0] node1362;
	wire [3-1:0] node1365;
	wire [3-1:0] node1366;
	wire [3-1:0] node1368;
	wire [3-1:0] node1372;
	wire [3-1:0] node1373;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1379;
	wire [3-1:0] node1382;
	wire [3-1:0] node1383;
	wire [3-1:0] node1385;
	wire [3-1:0] node1389;
	wire [3-1:0] node1390;
	wire [3-1:0] node1391;
	wire [3-1:0] node1393;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1401;
	wire [3-1:0] node1403;
	wire [3-1:0] node1406;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;

	assign outp = (inp[9]) ? node416 : node1;
		assign node1 = (inp[3]) ? node339 : node2;
			assign node2 = (inp[6]) ? node224 : node3;
				assign node3 = (inp[4]) ? node91 : node4;
					assign node4 = (inp[7]) ? node18 : node5;
						assign node5 = (inp[11]) ? 3'b001 : node6;
							assign node6 = (inp[10]) ? 3'b001 : node7;
								assign node7 = (inp[8]) ? node9 : 3'b001;
									assign node9 = (inp[5]) ? node11 : 3'b001;
										assign node11 = (inp[1]) ? 3'b000 : node12;
											assign node12 = (inp[2]) ? 3'b000 : 3'b001;
						assign node18 = (inp[10]) ? node52 : node19;
							assign node19 = (inp[5]) ? node39 : node20;
								assign node20 = (inp[8]) ? node32 : node21;
									assign node21 = (inp[11]) ? node27 : node22;
										assign node22 = (inp[0]) ? node24 : 3'b100;
											assign node24 = (inp[1]) ? 3'b000 : 3'b100;
										assign node27 = (inp[0]) ? node29 : 3'b101;
											assign node29 = (inp[1]) ? 3'b001 : 3'b101;
									assign node32 = (inp[2]) ? node34 : 3'b000;
										assign node34 = (inp[0]) ? node36 : 3'b000;
											assign node36 = (inp[1]) ? 3'b100 : 3'b000;
								assign node39 = (inp[8]) ? node45 : node40;
									assign node40 = (inp[0]) ? node42 : 3'b000;
										assign node42 = (inp[1]) ? 3'b100 : 3'b000;
									assign node45 = (inp[0]) ? node47 : 3'b100;
										assign node47 = (inp[2]) ? node49 : 3'b100;
											assign node49 = (inp[1]) ? 3'b000 : 3'b100;
							assign node52 = (inp[5]) ? node78 : node53;
								assign node53 = (inp[11]) ? node67 : node54;
									assign node54 = (inp[8]) ? node60 : node55;
										assign node55 = (inp[1]) ? node57 : 3'b101;
											assign node57 = (inp[0]) ? 3'b001 : 3'b101;
										assign node60 = (inp[2]) ? node62 : 3'b001;
											assign node62 = (inp[1]) ? node64 : 3'b001;
												assign node64 = (inp[0]) ? 3'b101 : 3'b001;
									assign node67 = (inp[8]) ? node73 : node68;
										assign node68 = (inp[0]) ? node70 : 3'b100;
											assign node70 = (inp[1]) ? 3'b000 : 3'b100;
										assign node73 = (inp[1]) ? 3'b001 : node74;
											assign node74 = (inp[0]) ? 3'b001 : 3'b000;
								assign node78 = (inp[8]) ? node84 : node79;
									assign node79 = (inp[0]) ? node81 : 3'b001;
										assign node81 = (inp[1]) ? 3'b101 : 3'b001;
									assign node84 = (inp[11]) ? node86 : 3'b100;
										assign node86 = (inp[1]) ? node88 : 3'b101;
											assign node88 = (inp[0]) ? 3'b001 : 3'b101;
					assign node91 = (inp[10]) ? node157 : node92;
						assign node92 = (inp[7]) ? node144 : node93;
							assign node93 = (inp[11]) ? node117 : node94;
								assign node94 = (inp[1]) ? node112 : node95;
									assign node95 = (inp[0]) ? node107 : node96;
										assign node96 = (inp[8]) ? node100 : node97;
											assign node97 = (inp[5]) ? 3'b110 : 3'b100;
											assign node100 = (inp[5]) ? node104 : node101;
												assign node101 = (inp[2]) ? 3'b010 : 3'b110;
												assign node104 = (inp[2]) ? 3'b110 : 3'b010;
										assign node107 = (inp[5]) ? node109 : 3'b010;
											assign node109 = (inp[8]) ? 3'b100 : 3'b010;
									assign node112 = (inp[8]) ? 3'b010 : node113;
										assign node113 = (inp[0]) ? 3'b110 : 3'b010;
								assign node117 = (inp[5]) ? node135 : node118;
									assign node118 = (inp[0]) ? node128 : node119;
										assign node119 = (inp[1]) ? node125 : node120;
											assign node120 = (inp[8]) ? 3'b001 : node121;
												assign node121 = (inp[2]) ? 3'b101 : 3'b100;
											assign node125 = (inp[8]) ? 3'b100 : 3'b001;
										assign node128 = (inp[8]) ? node130 : 3'b001;
											assign node130 = (inp[2]) ? 3'b110 : node131;
												assign node131 = (inp[1]) ? 3'b110 : 3'b100;
									assign node135 = (inp[8]) ? node139 : node136;
										assign node136 = (inp[0]) ? 3'b110 : 3'b000;
										assign node139 = (inp[0]) ? 3'b010 : node140;
											assign node140 = (inp[2]) ? 3'b010 : 3'b110;
							assign node144 = (inp[5]) ? node152 : node145;
								assign node145 = (inp[11]) ? node149 : node146;
									assign node146 = (inp[8]) ? 3'b000 : 3'b100;
									assign node149 = (inp[8]) ? 3'b100 : 3'b010;
								assign node152 = (inp[11]) ? node154 : 3'b000;
									assign node154 = (inp[8]) ? 3'b000 : 3'b100;
						assign node157 = (inp[7]) ? node195 : node158;
							assign node158 = (inp[11]) ? node172 : node159;
								assign node159 = (inp[8]) ? node163 : node160;
									assign node160 = (inp[5]) ? 3'b001 : 3'b101;
									assign node163 = (inp[5]) ? node169 : node164;
										assign node164 = (inp[0]) ? 3'b001 : node165;
											assign node165 = (inp[1]) ? 3'b001 : 3'b000;
										assign node169 = (inp[2]) ? 3'b110 : 3'b001;
								assign node172 = (inp[5]) ? node182 : node173;
									assign node173 = (inp[8]) ? node179 : node174;
										assign node174 = (inp[0]) ? 3'b011 : node175;
											assign node175 = (inp[1]) ? 3'b011 : 3'b111;
										assign node179 = (inp[0]) ? 3'b101 : 3'b011;
									assign node182 = (inp[8]) ? node188 : node183;
										assign node183 = (inp[0]) ? 3'b101 : node184;
											assign node184 = (inp[1]) ? 3'b101 : 3'b001;
										assign node188 = (inp[0]) ? 3'b001 : node189;
											assign node189 = (inp[2]) ? node191 : 3'b101;
												assign node191 = (inp[1]) ? 3'b001 : 3'b101;
							assign node195 = (inp[11]) ? node207 : node196;
								assign node196 = (inp[8]) ? node200 : node197;
									assign node197 = (inp[5]) ? 3'b010 : 3'b110;
									assign node200 = (inp[5]) ? node202 : 3'b010;
										assign node202 = (inp[1]) ? 3'b100 : node203;
											assign node203 = (inp[2]) ? 3'b100 : 3'b110;
								assign node207 = (inp[5]) ? node215 : node208;
									assign node208 = (inp[8]) ? node210 : 3'b001;
										assign node210 = (inp[1]) ? 3'b110 : node211;
											assign node211 = (inp[0]) ? 3'b110 : 3'b100;
									assign node215 = (inp[8]) ? 3'b010 : node216;
										assign node216 = (inp[0]) ? 3'b110 : node217;
											assign node217 = (inp[1]) ? 3'b110 : node218;
												assign node218 = (inp[2]) ? 3'b110 : 3'b010;
				assign node224 = (inp[7]) ? node322 : node225;
					assign node225 = (inp[4]) ? node301 : node226;
						assign node226 = (inp[10]) ? node254 : node227;
							assign node227 = (inp[11]) ? node241 : node228;
								assign node228 = (inp[5]) ? 3'b000 : node229;
									assign node229 = (inp[8]) ? node235 : node230;
										assign node230 = (inp[1]) ? 3'b100 : node231;
											assign node231 = (inp[0]) ? 3'b100 : 3'b000;
										assign node235 = (inp[2]) ? 3'b000 : node236;
											assign node236 = (inp[0]) ? 3'b000 : 3'b100;
								assign node241 = (inp[5]) ? node249 : node242;
									assign node242 = (inp[8]) ? node244 : 3'b010;
										assign node244 = (inp[1]) ? 3'b100 : node245;
											assign node245 = (inp[0]) ? 3'b100 : 3'b000;
									assign node249 = (inp[0]) ? node251 : 3'b100;
										assign node251 = (inp[8]) ? 3'b000 : 3'b100;
							assign node254 = (inp[8]) ? node272 : node255;
								assign node255 = (inp[11]) ? node261 : node256;
									assign node256 = (inp[5]) ? 3'b110 : node257;
										assign node257 = (inp[0]) ? 3'b110 : 3'b011;
									assign node261 = (inp[5]) ? node267 : node262;
										assign node262 = (inp[0]) ? node264 : 3'b101;
											assign node264 = (inp[1]) ? 3'b001 : 3'b101;
										assign node267 = (inp[1]) ? node269 : 3'b011;
											assign node269 = (inp[0]) ? 3'b110 : 3'b011;
								assign node272 = (inp[11]) ? node288 : node273;
									assign node273 = (inp[5]) ? node277 : node274;
										assign node274 = (inp[0]) ? 3'b010 : 3'b110;
										assign node277 = (inp[0]) ? node283 : node278;
											assign node278 = (inp[2]) ? 3'b000 : node279;
												assign node279 = (inp[1]) ? 3'b000 : 3'b010;
											assign node283 = (inp[1]) ? 3'b100 : node284;
												assign node284 = (inp[2]) ? 3'b100 : 3'b000;
									assign node288 = (inp[5]) ? node296 : node289;
										assign node289 = (inp[0]) ? node293 : node290;
											assign node290 = (inp[1]) ? 3'b011 : 3'b001;
											assign node293 = (inp[1]) ? 3'b110 : 3'b011;
										assign node296 = (inp[0]) ? node298 : 3'b110;
											assign node298 = (inp[1]) ? 3'b010 : 3'b110;
						assign node301 = (inp[10]) ? node303 : 3'b000;
							assign node303 = (inp[5]) ? node317 : node304;
								assign node304 = (inp[8]) ? node308 : node305;
									assign node305 = (inp[11]) ? 3'b010 : 3'b100;
									assign node308 = (inp[11]) ? node310 : 3'b000;
										assign node310 = (inp[2]) ? 3'b100 : node311;
											assign node311 = (inp[1]) ? 3'b100 : node312;
												assign node312 = (inp[0]) ? 3'b100 : 3'b000;
								assign node317 = (inp[11]) ? node319 : 3'b000;
									assign node319 = (inp[8]) ? 3'b000 : 3'b100;
					assign node322 = (inp[4]) ? 3'b000 : node323;
						assign node323 = (inp[10]) ? node325 : 3'b000;
							assign node325 = (inp[8]) ? node333 : node326;
								assign node326 = (inp[11]) ? node330 : node327;
									assign node327 = (inp[5]) ? 3'b000 : 3'b100;
									assign node330 = (inp[5]) ? 3'b100 : 3'b010;
								assign node333 = (inp[11]) ? node335 : 3'b000;
									assign node335 = (inp[5]) ? 3'b000 : 3'b100;
			assign node339 = (inp[6]) ? 3'b000 : node340;
				assign node340 = (inp[7]) ? node398 : node341;
					assign node341 = (inp[4]) ? node383 : node342;
						assign node342 = (inp[10]) ? node356 : node343;
							assign node343 = (inp[5]) ? node351 : node344;
								assign node344 = (inp[8]) ? node348 : node345;
									assign node345 = (inp[11]) ? 3'b010 : 3'b100;
									assign node348 = (inp[11]) ? 3'b100 : 3'b000;
								assign node351 = (inp[8]) ? 3'b000 : node352;
									assign node352 = (inp[11]) ? 3'b100 : 3'b000;
							assign node356 = (inp[11]) ? node368 : node357;
								assign node357 = (inp[5]) ? node361 : node358;
									assign node358 = (inp[8]) ? 3'b010 : 3'b110;
									assign node361 = (inp[8]) ? node363 : 3'b010;
										assign node363 = (inp[1]) ? 3'b100 : node364;
											assign node364 = (inp[0]) ? 3'b100 : 3'b110;
								assign node368 = (inp[5]) ? node376 : node369;
									assign node369 = (inp[8]) ? node371 : 3'b001;
										assign node371 = (inp[1]) ? 3'b110 : node372;
											assign node372 = (inp[0]) ? 3'b110 : 3'b100;
									assign node376 = (inp[8]) ? 3'b010 : node377;
										assign node377 = (inp[0]) ? 3'b110 : node378;
											assign node378 = (inp[1]) ? 3'b110 : 3'b010;
						assign node383 = (inp[10]) ? node385 : 3'b000;
							assign node385 = (inp[8]) ? node393 : node386;
								assign node386 = (inp[5]) ? node390 : node387;
									assign node387 = (inp[11]) ? 3'b010 : 3'b100;
									assign node390 = (inp[11]) ? 3'b100 : 3'b000;
								assign node393 = (inp[5]) ? 3'b000 : node394;
									assign node394 = (inp[11]) ? 3'b100 : 3'b000;
					assign node398 = (inp[4]) ? 3'b000 : node399;
						assign node399 = (inp[10]) ? node401 : 3'b000;
							assign node401 = (inp[8]) ? node409 : node402;
								assign node402 = (inp[5]) ? node406 : node403;
									assign node403 = (inp[11]) ? 3'b010 : 3'b100;
									assign node406 = (inp[11]) ? 3'b100 : 3'b000;
								assign node409 = (inp[11]) ? node411 : 3'b000;
									assign node411 = (inp[5]) ? 3'b000 : 3'b100;
		assign node416 = (inp[6]) ? node868 : node417;
			assign node417 = (inp[3]) ? node559 : node418;
				assign node418 = (inp[10]) ? node524 : node419;
					assign node419 = (inp[7]) ? node473 : node420;
						assign node420 = (inp[4]) ? node422 : 3'b111;
							assign node422 = (inp[0]) ? node452 : node423;
								assign node423 = (inp[8]) ? node437 : node424;
									assign node424 = (inp[11]) ? node432 : node425;
										assign node425 = (inp[5]) ? node427 : 3'b111;
											assign node427 = (inp[2]) ? 3'b011 : node428;
												assign node428 = (inp[1]) ? 3'b011 : 3'b111;
										assign node432 = (inp[5]) ? 3'b111 : node433;
											assign node433 = (inp[2]) ? 3'b001 : 3'b101;
									assign node437 = (inp[1]) ? node447 : node438;
										assign node438 = (inp[11]) ? node444 : node439;
											assign node439 = (inp[2]) ? 3'b011 : node440;
												assign node440 = (inp[5]) ? 3'b011 : 3'b111;
											assign node444 = (inp[2]) ? 3'b111 : 3'b001;
										assign node447 = (inp[11]) ? node449 : 3'b101;
											assign node449 = (inp[5]) ? 3'b011 : 3'b111;
								assign node452 = (inp[5]) ? node466 : node453;
									assign node453 = (inp[1]) ? node459 : node454;
										assign node454 = (inp[11]) ? 3'b111 : node455;
											assign node455 = (inp[8]) ? 3'b011 : 3'b111;
										assign node459 = (inp[11]) ? node463 : node460;
											assign node460 = (inp[8]) ? 3'b011 : 3'b111;
											assign node463 = (inp[8]) ? 3'b111 : 3'b001;
									assign node466 = (inp[11]) ? node470 : node467;
										assign node467 = (inp[8]) ? 3'b101 : 3'b011;
										assign node470 = (inp[8]) ? 3'b011 : 3'b111;
						assign node473 = (inp[4]) ? node503 : node474;
							assign node474 = (inp[5]) ? node492 : node475;
								assign node475 = (inp[0]) ? node483 : node476;
									assign node476 = (inp[8]) ? node480 : node477;
										assign node477 = (inp[11]) ? 3'b101 : 3'b001;
										assign node480 = (inp[11]) ? 3'b001 : 3'b111;
									assign node483 = (inp[11]) ? node487 : node484;
										assign node484 = (inp[8]) ? 3'b011 : 3'b111;
										assign node487 = (inp[8]) ? node489 : 3'b001;
											assign node489 = (inp[1]) ? 3'b111 : 3'b001;
								assign node492 = (inp[11]) ? node498 : node493;
									assign node493 = (inp[8]) ? 3'b011 : node494;
										assign node494 = (inp[0]) ? 3'b011 : 3'b111;
									assign node498 = (inp[8]) ? 3'b111 : node499;
										assign node499 = (inp[1]) ? 3'b111 : 3'b001;
							assign node503 = (inp[8]) ? node511 : node504;
								assign node504 = (inp[11]) ? node508 : node505;
									assign node505 = (inp[5]) ? 3'b001 : 3'b101;
									assign node508 = (inp[5]) ? 3'b101 : 3'b011;
								assign node511 = (inp[5]) ? node515 : node512;
									assign node512 = (inp[11]) ? 3'b101 : 3'b001;
									assign node515 = (inp[11]) ? 3'b001 : node516;
										assign node516 = (inp[0]) ? 3'b110 : node517;
											assign node517 = (inp[2]) ? 3'b110 : node518;
												assign node518 = (inp[1]) ? 3'b110 : 3'b101;
					assign node524 = (inp[4]) ? node526 : 3'b111;
						assign node526 = (inp[7]) ? node528 : 3'b111;
							assign node528 = (inp[11]) ? node552 : node529;
								assign node529 = (inp[8]) ? node537 : node530;
									assign node530 = (inp[5]) ? node532 : 3'b111;
										assign node532 = (inp[0]) ? 3'b011 : node533;
											assign node533 = (inp[1]) ? 3'b011 : 3'b111;
									assign node537 = (inp[1]) ? node545 : node538;
										assign node538 = (inp[5]) ? 3'b011 : node539;
											assign node539 = (inp[0]) ? 3'b011 : node540;
												assign node540 = (inp[2]) ? 3'b101 : 3'b111;
										assign node545 = (inp[0]) ? 3'b101 : node546;
											assign node546 = (inp[2]) ? node548 : 3'b011;
												assign node548 = (inp[5]) ? 3'b101 : 3'b011;
								assign node552 = (inp[5]) ? node554 : 3'b111;
									assign node554 = (inp[8]) ? node556 : 3'b111;
										assign node556 = (inp[0]) ? 3'b011 : 3'b111;
				assign node559 = (inp[10]) ? node711 : node560;
					assign node560 = (inp[4]) ? node630 : node561;
						assign node561 = (inp[7]) ? node593 : node562;
							assign node562 = (inp[11]) ? node572 : node563;
								assign node563 = (inp[8]) ? node567 : node564;
									assign node564 = (inp[5]) ? 3'b001 : 3'b101;
									assign node567 = (inp[5]) ? node569 : 3'b001;
										assign node569 = (inp[1]) ? 3'b110 : 3'b101;
								assign node572 = (inp[5]) ? node580 : node573;
									assign node573 = (inp[8]) ? node575 : 3'b011;
										assign node575 = (inp[2]) ? 3'b101 : node576;
											assign node576 = (inp[1]) ? 3'b101 : 3'b001;
									assign node580 = (inp[8]) ? node588 : node581;
										assign node581 = (inp[0]) ? 3'b101 : node582;
											assign node582 = (inp[2]) ? 3'b101 : node583;
												assign node583 = (inp[1]) ? 3'b101 : 3'b001;
										assign node588 = (inp[0]) ? 3'b001 : node589;
											assign node589 = (inp[2]) ? 3'b001 : 3'b101;
							assign node593 = (inp[11]) ? node609 : node594;
								assign node594 = (inp[5]) ? node598 : node595;
									assign node595 = (inp[8]) ? 3'b010 : 3'b110;
									assign node598 = (inp[8]) ? node602 : node599;
										assign node599 = (inp[2]) ? 3'b010 : 3'b110;
										assign node602 = (inp[1]) ? 3'b100 : node603;
											assign node603 = (inp[2]) ? 3'b100 : node604;
												assign node604 = (inp[0]) ? 3'b100 : 3'b010;
								assign node609 = (inp[5]) ? node621 : node610;
									assign node610 = (inp[8]) ? node616 : node611;
										assign node611 = (inp[1]) ? 3'b001 : node612;
											assign node612 = (inp[0]) ? 3'b001 : 3'b101;
										assign node616 = (inp[0]) ? 3'b110 : node617;
											assign node617 = (inp[1]) ? 3'b110 : 3'b001;
									assign node621 = (inp[0]) ? node627 : node622;
										assign node622 = (inp[1]) ? 3'b110 : node623;
											assign node623 = (inp[8]) ? 3'b110 : 3'b010;
										assign node627 = (inp[8]) ? 3'b010 : 3'b110;
						assign node630 = (inp[7]) ? node662 : node631;
							assign node631 = (inp[11]) ? node643 : node632;
								assign node632 = (inp[8]) ? node636 : node633;
									assign node633 = (inp[5]) ? 3'b010 : 3'b110;
									assign node636 = (inp[5]) ? node638 : 3'b010;
										assign node638 = (inp[1]) ? 3'b100 : node639;
											assign node639 = (inp[0]) ? 3'b100 : 3'b010;
								assign node643 = (inp[5]) ? node655 : node644;
									assign node644 = (inp[8]) ? node650 : node645;
										assign node645 = (inp[1]) ? 3'b001 : node646;
											assign node646 = (inp[2]) ? 3'b001 : 3'b110;
										assign node650 = (inp[0]) ? 3'b110 : node651;
											assign node651 = (inp[2]) ? 3'b001 : 3'b110;
									assign node655 = (inp[8]) ? node657 : 3'b110;
										assign node657 = (inp[0]) ? 3'b010 : node658;
											assign node658 = (inp[1]) ? 3'b010 : 3'b110;
							assign node662 = (inp[11]) ? node680 : node663;
								assign node663 = (inp[5]) ? node673 : node664;
									assign node664 = (inp[8]) ? node670 : node665;
										assign node665 = (inp[2]) ? 3'b100 : node666;
											assign node666 = (inp[0]) ? 3'b100 : 3'b000;
										assign node670 = (inp[0]) ? 3'b000 : 3'b100;
									assign node673 = (inp[2]) ? 3'b000 : node674;
										assign node674 = (inp[1]) ? 3'b000 : node675;
											assign node675 = (inp[8]) ? 3'b000 : 3'b100;
								assign node680 = (inp[8]) ? node698 : node681;
									assign node681 = (inp[2]) ? node687 : node682;
										assign node682 = (inp[0]) ? 3'b010 : node683;
											assign node683 = (inp[5]) ? 3'b010 : 3'b110;
										assign node687 = (inp[5]) ? node693 : node688;
											assign node688 = (inp[0]) ? 3'b010 : node689;
												assign node689 = (inp[1]) ? 3'b010 : 3'b100;
											assign node693 = (inp[0]) ? 3'b100 : node694;
												assign node694 = (inp[1]) ? 3'b100 : 3'b010;
									assign node698 = (inp[5]) ? node704 : node699;
										assign node699 = (inp[2]) ? 3'b100 : node700;
											assign node700 = (inp[0]) ? 3'b100 : 3'b010;
										assign node704 = (inp[0]) ? 3'b000 : node705;
											assign node705 = (inp[2]) ? node707 : 3'b100;
												assign node707 = (inp[1]) ? 3'b000 : 3'b100;
					assign node711 = (inp[4]) ? node777 : node712;
						assign node712 = (inp[7]) ? node736 : node713;
							assign node713 = (inp[11]) ? node729 : node714;
								assign node714 = (inp[5]) ? node722 : node715;
									assign node715 = (inp[8]) ? node717 : 3'b111;
										assign node717 = (inp[0]) ? 3'b011 : node718;
											assign node718 = (inp[2]) ? 3'b011 : 3'b111;
									assign node722 = (inp[8]) ? node724 : 3'b011;
										assign node724 = (inp[0]) ? 3'b101 : node725;
											assign node725 = (inp[2]) ? 3'b101 : 3'b011;
								assign node729 = (inp[0]) ? node731 : 3'b111;
									assign node731 = (inp[5]) ? node733 : 3'b111;
										assign node733 = (inp[8]) ? 3'b011 : 3'b111;
							assign node736 = (inp[8]) ? node754 : node737;
								assign node737 = (inp[5]) ? node747 : node738;
									assign node738 = (inp[0]) ? node744 : node739;
										assign node739 = (inp[11]) ? 3'b111 : node740;
											assign node740 = (inp[2]) ? 3'b111 : 3'b011;
										assign node744 = (inp[11]) ? 3'b011 : 3'b101;
									assign node747 = (inp[0]) ? node751 : node748;
										assign node748 = (inp[11]) ? 3'b011 : 3'b101;
										assign node751 = (inp[11]) ? 3'b101 : 3'b001;
								assign node754 = (inp[11]) ? node764 : node755;
									assign node755 = (inp[5]) ? node761 : node756;
										assign node756 = (inp[1]) ? 3'b001 : node757;
											assign node757 = (inp[0]) ? 3'b001 : 3'b101;
										assign node761 = (inp[0]) ? 3'b110 : 3'b001;
									assign node764 = (inp[5]) ? node770 : node765;
										assign node765 = (inp[2]) ? 3'b101 : node766;
											assign node766 = (inp[1]) ? 3'b101 : 3'b011;
										assign node770 = (inp[0]) ? node772 : 3'b101;
											assign node772 = (inp[2]) ? 3'b001 : node773;
												assign node773 = (inp[1]) ? 3'b001 : 3'b101;
						assign node777 = (inp[7]) ? node817 : node778;
							assign node778 = (inp[0]) ? node802 : node779;
								assign node779 = (inp[11]) ? node791 : node780;
									assign node780 = (inp[5]) ? node786 : node781;
										assign node781 = (inp[8]) ? node783 : 3'b001;
											assign node783 = (inp[2]) ? 3'b110 : 3'b111;
										assign node786 = (inp[8]) ? 3'b001 : node787;
											assign node787 = (inp[2]) ? 3'b001 : 3'b101;
									assign node791 = (inp[8]) ? node799 : node792;
										assign node792 = (inp[5]) ? 3'b011 : node793;
											assign node793 = (inp[1]) ? node795 : 3'b111;
												assign node795 = (inp[2]) ? 3'b011 : 3'b111;
										assign node799 = (inp[5]) ? 3'b101 : 3'b011;
								assign node802 = (inp[11]) ? node810 : node803;
									assign node803 = (inp[8]) ? node807 : node804;
										assign node804 = (inp[5]) ? 3'b001 : 3'b101;
										assign node807 = (inp[5]) ? 3'b110 : 3'b001;
									assign node810 = (inp[8]) ? node814 : node811;
										assign node811 = (inp[5]) ? 3'b101 : 3'b011;
										assign node814 = (inp[5]) ? 3'b001 : 3'b101;
							assign node817 = (inp[5]) ? node843 : node818;
								assign node818 = (inp[0]) ? node830 : node819;
									assign node819 = (inp[11]) ? node827 : node820;
										assign node820 = (inp[8]) ? 3'b100 : node821;
											assign node821 = (inp[2]) ? node823 : 3'b001;
												assign node823 = (inp[1]) ? 3'b110 : 3'b001;
										assign node827 = (inp[8]) ? 3'b001 : 3'b101;
									assign node830 = (inp[11]) ? node834 : node831;
										assign node831 = (inp[8]) ? 3'b010 : 3'b110;
										assign node834 = (inp[8]) ? node838 : node835;
											assign node835 = (inp[2]) ? 3'b001 : 3'b101;
											assign node838 = (inp[1]) ? 3'b110 : node839;
												assign node839 = (inp[2]) ? 3'b110 : 3'b001;
								assign node843 = (inp[2]) ? node851 : node844;
									assign node844 = (inp[8]) ? 3'b010 : node845;
										assign node845 = (inp[11]) ? 3'b110 : node846;
											assign node846 = (inp[0]) ? 3'b010 : 3'b110;
									assign node851 = (inp[8]) ? node859 : node852;
										assign node852 = (inp[0]) ? node856 : node853;
											assign node853 = (inp[11]) ? 3'b001 : 3'b110;
											assign node856 = (inp[11]) ? 3'b110 : 3'b010;
										assign node859 = (inp[11]) ? node863 : node860;
											assign node860 = (inp[0]) ? 3'b100 : 3'b010;
											assign node863 = (inp[1]) ? node865 : 3'b110;
												assign node865 = (inp[0]) ? 3'b010 : 3'b110;
			assign node868 = (inp[3]) ? node1216 : node869;
				assign node869 = (inp[10]) ? node1041 : node870;
					assign node870 = (inp[4]) ? node958 : node871;
						assign node871 = (inp[7]) ? node919 : node872;
							assign node872 = (inp[11]) ? node896 : node873;
								assign node873 = (inp[5]) ? node883 : node874;
									assign node874 = (inp[8]) ? node876 : 3'b101;
										assign node876 = (inp[0]) ? 3'b001 : node877;
											assign node877 = (inp[1]) ? node879 : 3'b101;
												assign node879 = (inp[2]) ? 3'b001 : 3'b101;
									assign node883 = (inp[8]) ? node889 : node884;
										assign node884 = (inp[0]) ? 3'b001 : node885;
											assign node885 = (inp[2]) ? 3'b001 : 3'b101;
										assign node889 = (inp[0]) ? 3'b111 : node890;
											assign node890 = (inp[1]) ? 3'b011 : node891;
												assign node891 = (inp[2]) ? 3'b011 : 3'b001;
								assign node896 = (inp[5]) ? node908 : node897;
									assign node897 = (inp[8]) ? node901 : node898;
										assign node898 = (inp[0]) ? 3'b010 : 3'b110;
										assign node901 = (inp[0]) ? node903 : 3'b000;
											assign node903 = (inp[1]) ? 3'b101 : node904;
												assign node904 = (inp[2]) ? 3'b100 : 3'b000;
									assign node908 = (inp[8]) ? node914 : node909;
										assign node909 = (inp[0]) ? node911 : 3'b000;
											assign node911 = (inp[1]) ? 3'b101 : 3'b100;
										assign node914 = (inp[2]) ? node916 : 3'b101;
											assign node916 = (inp[1]) ? 3'b001 : 3'b101;
							assign node919 = (inp[11]) ? node943 : node920;
								assign node920 = (inp[8]) ? node932 : node921;
									assign node921 = (inp[5]) ? node927 : node922;
										assign node922 = (inp[1]) ? 3'b110 : node923;
											assign node923 = (inp[0]) ? 3'b110 : 3'b010;
										assign node927 = (inp[0]) ? 3'b010 : node928;
											assign node928 = (inp[1]) ? 3'b010 : 3'b110;
									assign node932 = (inp[2]) ? node934 : 3'b010;
										assign node934 = (inp[0]) ? 3'b010 : node935;
											assign node935 = (inp[1]) ? node939 : node936;
												assign node936 = (inp[5]) ? 3'b010 : 3'b100;
												assign node939 = (inp[5]) ? 3'b100 : 3'b010;
								assign node943 = (inp[8]) ? node951 : node944;
									assign node944 = (inp[0]) ? node948 : node945;
										assign node945 = (inp[5]) ? 3'b001 : 3'b101;
										assign node948 = (inp[5]) ? 3'b110 : 3'b001;
									assign node951 = (inp[0]) ? node955 : node952;
										assign node952 = (inp[5]) ? 3'b110 : 3'b001;
										assign node955 = (inp[5]) ? 3'b010 : 3'b110;
						assign node958 = (inp[7]) ? node1006 : node959;
							assign node959 = (inp[11]) ? node985 : node960;
								assign node960 = (inp[8]) ? node974 : node961;
									assign node961 = (inp[5]) ? node969 : node962;
										assign node962 = (inp[2]) ? 3'b110 : node963;
											assign node963 = (inp[1]) ? 3'b110 : node964;
												assign node964 = (inp[0]) ? 3'b110 : 3'b010;
										assign node969 = (inp[0]) ? 3'b010 : node970;
											assign node970 = (inp[1]) ? 3'b010 : 3'b110;
									assign node974 = (inp[5]) ? node980 : node975;
										assign node975 = (inp[1]) ? 3'b010 : node976;
											assign node976 = (inp[0]) ? 3'b010 : 3'b100;
										assign node980 = (inp[2]) ? node982 : 3'b100;
											assign node982 = (inp[1]) ? 3'b100 : 3'b010;
								assign node985 = (inp[5]) ? node993 : node986;
									assign node986 = (inp[0]) ? node990 : node987;
										assign node987 = (inp[8]) ? 3'b001 : 3'b111;
										assign node990 = (inp[8]) ? 3'b110 : 3'b001;
									assign node993 = (inp[8]) ? node999 : node994;
										assign node994 = (inp[0]) ? 3'b110 : node995;
											assign node995 = (inp[1]) ? 3'b110 : 3'b001;
										assign node999 = (inp[0]) ? 3'b010 : node1000;
											assign node1000 = (inp[1]) ? node1002 : 3'b110;
												assign node1002 = (inp[2]) ? 3'b010 : 3'b110;
							assign node1006 = (inp[11]) ? node1028 : node1007;
								assign node1007 = (inp[5]) ? node1021 : node1008;
									assign node1008 = (inp[8]) ? node1014 : node1009;
										assign node1009 = (inp[0]) ? 3'b100 : node1010;
											assign node1010 = (inp[1]) ? 3'b100 : 3'b000;
										assign node1014 = (inp[0]) ? 3'b000 : node1015;
											assign node1015 = (inp[1]) ? node1017 : 3'b100;
												assign node1017 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1021 = (inp[8]) ? 3'b000 : node1022;
										assign node1022 = (inp[0]) ? 3'b000 : node1023;
											assign node1023 = (inp[1]) ? 3'b000 : 3'b100;
								assign node1028 = (inp[5]) ? node1036 : node1029;
									assign node1029 = (inp[1]) ? 3'b010 : node1030;
										assign node1030 = (inp[0]) ? 3'b010 : node1031;
											assign node1031 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1036 = (inp[0]) ? node1038 : 3'b100;
										assign node1038 = (inp[8]) ? 3'b000 : 3'b100;
					assign node1041 = (inp[7]) ? node1123 : node1042;
						assign node1042 = (inp[4]) ? node1074 : node1043;
							assign node1043 = (inp[11]) ? node1067 : node1044;
								assign node1044 = (inp[5]) ? node1060 : node1045;
									assign node1045 = (inp[2]) ? node1055 : node1046;
										assign node1046 = (inp[8]) ? node1052 : node1047;
											assign node1047 = (inp[0]) ? node1049 : 3'b011;
												assign node1049 = (inp[1]) ? 3'b111 : 3'b011;
											assign node1052 = (inp[1]) ? 3'b011 : 3'b111;
										assign node1055 = (inp[0]) ? 3'b111 : node1056;
											assign node1056 = (inp[1]) ? 3'b111 : 3'b101;
									assign node1060 = (inp[8]) ? node1064 : node1061;
										assign node1061 = (inp[1]) ? 3'b011 : 3'b111;
										assign node1064 = (inp[0]) ? 3'b001 : 3'b011;
								assign node1067 = (inp[8]) ? node1069 : 3'b111;
									assign node1069 = (inp[0]) ? node1071 : 3'b111;
										assign node1071 = (inp[2]) ? 3'b011 : 3'b111;
							assign node1074 = (inp[5]) ? node1106 : node1075;
								assign node1075 = (inp[0]) ? node1093 : node1076;
									assign node1076 = (inp[2]) ? node1084 : node1077;
										assign node1077 = (inp[8]) ? node1081 : node1078;
											assign node1078 = (inp[11]) ? 3'b111 : 3'b011;
											assign node1081 = (inp[1]) ? 3'b101 : 3'b111;
										assign node1084 = (inp[1]) ? node1090 : node1085;
											assign node1085 = (inp[8]) ? node1087 : 3'b011;
												assign node1087 = (inp[11]) ? 3'b011 : 3'b111;
											assign node1090 = (inp[8]) ? 3'b011 : 3'b111;
									assign node1093 = (inp[11]) ? node1097 : node1094;
										assign node1094 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1097 = (inp[8]) ? node1103 : node1098;
											assign node1098 = (inp[1]) ? 3'b011 : node1099;
												assign node1099 = (inp[2]) ? 3'b011 : 3'b111;
											assign node1103 = (inp[2]) ? 3'b101 : 3'b011;
								assign node1106 = (inp[0]) ? node1114 : node1107;
									assign node1107 = (inp[11]) ? node1111 : node1108;
										assign node1108 = (inp[8]) ? 3'b001 : 3'b101;
										assign node1111 = (inp[8]) ? 3'b101 : 3'b011;
									assign node1114 = (inp[11]) ? node1118 : node1115;
										assign node1115 = (inp[8]) ? 3'b110 : 3'b001;
										assign node1118 = (inp[8]) ? node1120 : 3'b101;
											assign node1120 = (inp[1]) ? 3'b001 : 3'b101;
						assign node1123 = (inp[4]) ? node1165 : node1124;
							assign node1124 = (inp[11]) ? node1144 : node1125;
								assign node1125 = (inp[0]) ? node1133 : node1126;
									assign node1126 = (inp[8]) ? node1130 : node1127;
										assign node1127 = (inp[5]) ? 3'b101 : 3'b010;
										assign node1130 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1133 = (inp[5]) ? node1141 : node1134;
										assign node1134 = (inp[8]) ? node1136 : 3'b101;
											assign node1136 = (inp[2]) ? 3'b001 : node1137;
												assign node1137 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1141 = (inp[1]) ? 3'b110 : 3'b001;
								assign node1144 = (inp[5]) ? node1158 : node1145;
									assign node1145 = (inp[8]) ? node1153 : node1146;
										assign node1146 = (inp[0]) ? node1148 : 3'b111;
											assign node1148 = (inp[2]) ? 3'b011 : node1149;
												assign node1149 = (inp[1]) ? 3'b011 : 3'b111;
										assign node1153 = (inp[1]) ? node1155 : 3'b011;
											assign node1155 = (inp[2]) ? 3'b101 : 3'b011;
									assign node1158 = (inp[8]) ? node1162 : node1159;
										assign node1159 = (inp[0]) ? 3'b101 : 3'b011;
										assign node1162 = (inp[0]) ? 3'b001 : 3'b101;
							assign node1165 = (inp[5]) ? node1191 : node1166;
								assign node1166 = (inp[11]) ? node1182 : node1167;
									assign node1167 = (inp[8]) ? node1175 : node1168;
										assign node1168 = (inp[0]) ? node1170 : 3'b001;
											assign node1170 = (inp[2]) ? 3'b110 : node1171;
												assign node1171 = (inp[1]) ? 3'b110 : 3'b001;
										assign node1175 = (inp[0]) ? node1177 : 3'b110;
											assign node1177 = (inp[2]) ? 3'b010 : node1178;
												assign node1178 = (inp[1]) ? 3'b010 : 3'b110;
									assign node1182 = (inp[8]) ? node1188 : node1183;
										assign node1183 = (inp[0]) ? node1185 : 3'b101;
											assign node1185 = (inp[1]) ? 3'b001 : 3'b101;
										assign node1188 = (inp[1]) ? 3'b110 : 3'b001;
								assign node1191 = (inp[11]) ? node1205 : node1192;
									assign node1192 = (inp[8]) ? node1200 : node1193;
										assign node1193 = (inp[0]) ? node1195 : 3'b110;
											assign node1195 = (inp[2]) ? 3'b010 : node1196;
												assign node1196 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1200 = (inp[1]) ? node1202 : 3'b010;
											assign node1202 = (inp[0]) ? 3'b100 : 3'b010;
									assign node1205 = (inp[8]) ? node1209 : node1206;
										assign node1206 = (inp[0]) ? 3'b110 : 3'b001;
										assign node1209 = (inp[2]) ? node1211 : 3'b110;
											assign node1211 = (inp[1]) ? node1213 : 3'b110;
												assign node1213 = (inp[0]) ? 3'b010 : 3'b110;
				assign node1216 = (inp[10]) ? node1286 : node1217;
					assign node1217 = (inp[7]) ? node1275 : node1218;
						assign node1218 = (inp[4]) ? node1266 : node1219;
							assign node1219 = (inp[11]) ? node1237 : node1220;
								assign node1220 = (inp[5]) ? node1232 : node1221;
									assign node1221 = (inp[8]) ? node1227 : node1222;
										assign node1222 = (inp[0]) ? 3'b100 : node1223;
											assign node1223 = (inp[1]) ? 3'b100 : 3'b010;
										assign node1227 = (inp[0]) ? 3'b000 : node1228;
											assign node1228 = (inp[1]) ? 3'b000 : 3'b100;
									assign node1232 = (inp[0]) ? 3'b000 : node1233;
										assign node1233 = (inp[1]) ? 3'b000 : 3'b100;
								assign node1237 = (inp[8]) ? node1255 : node1238;
									assign node1238 = (inp[5]) ? node1246 : node1239;
										assign node1239 = (inp[0]) ? 3'b010 : node1240;
											assign node1240 = (inp[1]) ? node1242 : 3'b110;
												assign node1242 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1246 = (inp[0]) ? node1252 : node1247;
											assign node1247 = (inp[2]) ? node1249 : 3'b010;
												assign node1249 = (inp[1]) ? 3'b100 : 3'b010;
											assign node1252 = (inp[2]) ? 3'b110 : 3'b100;
									assign node1255 = (inp[0]) ? node1263 : node1256;
										assign node1256 = (inp[5]) ? 3'b100 : node1257;
											assign node1257 = (inp[2]) ? node1259 : 3'b010;
												assign node1259 = (inp[1]) ? 3'b100 : 3'b010;
										assign node1263 = (inp[5]) ? 3'b000 : 3'b100;
							assign node1266 = (inp[5]) ? 3'b000 : node1267;
								assign node1267 = (inp[11]) ? node1269 : 3'b000;
									assign node1269 = (inp[1]) ? 3'b000 : node1270;
										assign node1270 = (inp[0]) ? 3'b000 : 3'b100;
						assign node1275 = (inp[5]) ? 3'b000 : node1276;
							assign node1276 = (inp[11]) ? node1278 : 3'b000;
								assign node1278 = (inp[4]) ? 3'b000 : node1279;
									assign node1279 = (inp[8]) ? 3'b000 : node1280;
										assign node1280 = (inp[0]) ? 3'b000 : 3'b100;
					assign node1286 = (inp[4]) ? node1372 : node1287;
						assign node1287 = (inp[7]) ? node1339 : node1288;
							assign node1288 = (inp[11]) ? node1318 : node1289;
								assign node1289 = (inp[2]) ? node1303 : node1290;
									assign node1290 = (inp[8]) ? node1298 : node1291;
										assign node1291 = (inp[5]) ? node1295 : node1292;
											assign node1292 = (inp[0]) ? 3'b110 : 3'b001;
											assign node1295 = (inp[0]) ? 3'b010 : 3'b110;
										assign node1298 = (inp[5]) ? node1300 : 3'b110;
											assign node1300 = (inp[1]) ? 3'b100 : 3'b010;
									assign node1303 = (inp[8]) ? node1311 : node1304;
										assign node1304 = (inp[5]) ? node1308 : node1305;
											assign node1305 = (inp[1]) ? 3'b110 : 3'b001;
											assign node1308 = (inp[0]) ? 3'b010 : 3'b110;
										assign node1311 = (inp[0]) ? node1315 : node1312;
											assign node1312 = (inp[5]) ? 3'b010 : 3'b110;
											assign node1315 = (inp[5]) ? 3'b100 : 3'b010;
								assign node1318 = (inp[8]) ? node1332 : node1319;
									assign node1319 = (inp[5]) ? node1327 : node1320;
										assign node1320 = (inp[0]) ? node1322 : 3'b101;
											assign node1322 = (inp[1]) ? 3'b001 : node1323;
												assign node1323 = (inp[2]) ? 3'b001 : 3'b101;
										assign node1327 = (inp[0]) ? node1329 : 3'b001;
											assign node1329 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1332 = (inp[5]) ? 3'b110 : node1333;
										assign node1333 = (inp[0]) ? node1335 : 3'b001;
											assign node1335 = (inp[1]) ? 3'b110 : 3'b001;
							assign node1339 = (inp[11]) ? node1357 : node1340;
								assign node1340 = (inp[8]) ? node1350 : node1341;
									assign node1341 = (inp[5]) ? 3'b100 : node1342;
										assign node1342 = (inp[0]) ? node1344 : 3'b010;
											assign node1344 = (inp[1]) ? 3'b100 : node1345;
												assign node1345 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1350 = (inp[5]) ? 3'b000 : node1351;
										assign node1351 = (inp[1]) ? node1353 : 3'b100;
											assign node1353 = (inp[0]) ? 3'b000 : 3'b100;
								assign node1357 = (inp[5]) ? node1365 : node1358;
									assign node1358 = (inp[8]) ? node1360 : 3'b110;
										assign node1360 = (inp[2]) ? node1362 : 3'b010;
											assign node1362 = (inp[1]) ? 3'b100 : 3'b010;
									assign node1365 = (inp[8]) ? 3'b100 : node1366;
										assign node1366 = (inp[2]) ? node1368 : 3'b010;
											assign node1368 = (inp[1]) ? 3'b100 : 3'b010;
						assign node1372 = (inp[7]) ? node1406 : node1373;
							assign node1373 = (inp[5]) ? node1389 : node1374;
								assign node1374 = (inp[11]) ? node1382 : node1375;
									assign node1375 = (inp[8]) ? node1379 : node1376;
										assign node1376 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1379 = (inp[0]) ? 3'b000 : 3'b100;
									assign node1382 = (inp[8]) ? 3'b010 : node1383;
										assign node1383 = (inp[0]) ? node1385 : 3'b110;
											assign node1385 = (inp[1]) ? 3'b010 : 3'b110;
								assign node1389 = (inp[11]) ? node1397 : node1390;
									assign node1390 = (inp[8]) ? 3'b000 : node1391;
										assign node1391 = (inp[0]) ? node1393 : 3'b100;
											assign node1393 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1397 = (inp[8]) ? node1401 : node1398;
										assign node1398 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1401 = (inp[1]) ? node1403 : 3'b100;
											assign node1403 = (inp[2]) ? 3'b000 : 3'b100;
							assign node1406 = (inp[11]) ? node1408 : 3'b000;
								assign node1408 = (inp[8]) ? 3'b000 : node1409;
									assign node1409 = (inp[5]) ? 3'b000 : 3'b100;

endmodule