module dtc_split5_bm91 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node361;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node369;
	wire [3-1:0] node370;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node390;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node405;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node416;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node464;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node496;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node521;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node533;
	wire [3-1:0] node534;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node547;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node580;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node628;
	wire [3-1:0] node631;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node637;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node651;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node663;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node676;
	wire [3-1:0] node678;
	wire [3-1:0] node680;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node705;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node716;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node746;
	wire [3-1:0] node748;
	wire [3-1:0] node750;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node787;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node813;
	wire [3-1:0] node815;
	wire [3-1:0] node818;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node824;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node832;
	wire [3-1:0] node835;
	wire [3-1:0] node837;
	wire [3-1:0] node840;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node852;
	wire [3-1:0] node854;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node861;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node867;

	assign outp = (inp[3]) ? node634 : node1;
		assign node1 = (inp[9]) ? node293 : node2;
			assign node2 = (inp[1]) ? node104 : node3;
				assign node3 = (inp[5]) ? node57 : node4;
					assign node4 = (inp[6]) ? node24 : node5;
						assign node5 = (inp[0]) ? node9 : node6;
							assign node6 = (inp[4]) ? 3'b000 : 3'b001;
							assign node9 = (inp[4]) ? node17 : node10;
								assign node10 = (inp[2]) ? 3'b000 : node11;
									assign node11 = (inp[8]) ? 3'b000 : node12;
										assign node12 = (inp[7]) ? 3'b000 : 3'b001;
								assign node17 = (inp[8]) ? 3'b001 : node18;
									assign node18 = (inp[2]) ? 3'b001 : node19;
										assign node19 = (inp[7]) ? 3'b001 : 3'b000;
						assign node24 = (inp[10]) ? node34 : node25;
							assign node25 = (inp[7]) ? 3'b000 : node26;
								assign node26 = (inp[2]) ? node28 : 3'b000;
									assign node28 = (inp[11]) ? 3'b000 : node29;
										assign node29 = (inp[4]) ? 3'b001 : 3'b000;
							assign node34 = (inp[7]) ? node42 : node35;
								assign node35 = (inp[8]) ? node37 : 3'b000;
									assign node37 = (inp[11]) ? 3'b000 : node38;
										assign node38 = (inp[0]) ? 3'b000 : 3'b001;
								assign node42 = (inp[11]) ? node50 : node43;
									assign node43 = (inp[8]) ? 3'b000 : node44;
										assign node44 = (inp[0]) ? node46 : 3'b000;
											assign node46 = (inp[4]) ? 3'b000 : 3'b001;
									assign node50 = (inp[4]) ? node54 : node51;
										assign node51 = (inp[0]) ? 3'b001 : 3'b000;
										assign node54 = (inp[0]) ? 3'b000 : 3'b001;
					assign node57 = (inp[4]) ? node77 : node58;
						assign node58 = (inp[6]) ? node64 : node59;
							assign node59 = (inp[7]) ? 3'b001 : node60;
								assign node60 = (inp[0]) ? 3'b001 : 3'b000;
							assign node64 = (inp[0]) ? node70 : node65;
								assign node65 = (inp[8]) ? node67 : 3'b001;
									assign node67 = (inp[7]) ? 3'b000 : 3'b001;
								assign node70 = (inp[2]) ? node72 : 3'b000;
									assign node72 = (inp[10]) ? node74 : 3'b000;
										assign node74 = (inp[7]) ? 3'b001 : 3'b000;
						assign node77 = (inp[6]) ? node89 : node78;
							assign node78 = (inp[8]) ? node80 : 3'b000;
								assign node80 = (inp[0]) ? node82 : 3'b000;
									assign node82 = (inp[2]) ? 3'b000 : node83;
										assign node83 = (inp[10]) ? 3'b000 : node84;
											assign node84 = (inp[7]) ? 3'b000 : 3'b001;
							assign node89 = (inp[0]) ? 3'b001 : node90;
								assign node90 = (inp[8]) ? node92 : 3'b000;
									assign node92 = (inp[10]) ? node96 : node93;
										assign node93 = (inp[7]) ? 3'b000 : 3'b001;
										assign node96 = (inp[2]) ? node98 : 3'b001;
											assign node98 = (inp[11]) ? node100 : 3'b001;
												assign node100 = (inp[7]) ? 3'b001 : 3'b000;
				assign node104 = (inp[6]) ? node212 : node105;
					assign node105 = (inp[5]) ? node149 : node106;
						assign node106 = (inp[7]) ? node124 : node107;
							assign node107 = (inp[0]) ? node119 : node108;
								assign node108 = (inp[4]) ? node116 : node109;
									assign node109 = (inp[10]) ? 3'b001 : node110;
										assign node110 = (inp[8]) ? 3'b000 : node111;
											assign node111 = (inp[11]) ? 3'b000 : 3'b001;
									assign node116 = (inp[10]) ? 3'b000 : 3'b001;
								assign node119 = (inp[8]) ? 3'b000 : node120;
									assign node120 = (inp[4]) ? 3'b001 : 3'b000;
							assign node124 = (inp[4]) ? node138 : node125;
								assign node125 = (inp[8]) ? node133 : node126;
									assign node126 = (inp[0]) ? 3'b000 : node127;
										assign node127 = (inp[10]) ? node129 : 3'b001;
											assign node129 = (inp[2]) ? 3'b000 : 3'b001;
									assign node133 = (inp[0]) ? 3'b001 : node134;
										assign node134 = (inp[2]) ? 3'b000 : 3'b001;
								assign node138 = (inp[0]) ? 3'b001 : node139;
									assign node139 = (inp[11]) ? node141 : 3'b001;
										assign node141 = (inp[10]) ? node143 : 3'b000;
											assign node143 = (inp[8]) ? 3'b001 : node144;
												assign node144 = (inp[2]) ? 3'b001 : 3'b000;
						assign node149 = (inp[0]) ? node189 : node150;
							assign node150 = (inp[4]) ? node170 : node151;
								assign node151 = (inp[7]) ? node157 : node152;
									assign node152 = (inp[10]) ? 3'b001 : node153;
										assign node153 = (inp[8]) ? 3'b000 : 3'b001;
									assign node157 = (inp[2]) ? node165 : node158;
										assign node158 = (inp[10]) ? node162 : node159;
											assign node159 = (inp[11]) ? 3'b000 : 3'b001;
											assign node162 = (inp[8]) ? 3'b000 : 3'b001;
										assign node165 = (inp[11]) ? node167 : 3'b000;
											assign node167 = (inp[8]) ? 3'b001 : 3'b000;
								assign node170 = (inp[10]) ? node182 : node171;
									assign node171 = (inp[8]) ? node177 : node172;
										assign node172 = (inp[7]) ? node174 : 3'b000;
											assign node174 = (inp[11]) ? 3'b001 : 3'b000;
										assign node177 = (inp[11]) ? 3'b001 : node178;
											assign node178 = (inp[7]) ? 3'b000 : 3'b001;
									assign node182 = (inp[7]) ? node184 : 3'b000;
										assign node184 = (inp[8]) ? node186 : 3'b000;
											assign node186 = (inp[11]) ? 3'b000 : 3'b001;
							assign node189 = (inp[8]) ? 3'b001 : node190;
								assign node190 = (inp[10]) ? node200 : node191;
									assign node191 = (inp[4]) ? node195 : node192;
										assign node192 = (inp[7]) ? 3'b000 : 3'b001;
										assign node195 = (inp[7]) ? 3'b001 : node196;
											assign node196 = (inp[11]) ? 3'b000 : 3'b001;
									assign node200 = (inp[11]) ? node206 : node201;
										assign node201 = (inp[2]) ? node203 : 3'b001;
											assign node203 = (inp[4]) ? 3'b001 : 3'b000;
										assign node206 = (inp[7]) ? node208 : 3'b000;
											assign node208 = (inp[4]) ? 3'b001 : 3'b000;
					assign node212 = (inp[8]) ? node250 : node213;
						assign node213 = (inp[5]) ? node225 : node214;
							assign node214 = (inp[0]) ? node222 : node215;
								assign node215 = (inp[4]) ? 3'b001 : node216;
									assign node216 = (inp[10]) ? 3'b000 : node217;
										assign node217 = (inp[7]) ? 3'b001 : 3'b000;
								assign node222 = (inp[4]) ? 3'b000 : 3'b001;
							assign node225 = (inp[11]) ? node233 : node226;
								assign node226 = (inp[4]) ? node228 : 3'b000;
									assign node228 = (inp[7]) ? 3'b000 : node229;
										assign node229 = (inp[0]) ? 3'b001 : 3'b000;
								assign node233 = (inp[10]) ? node245 : node234;
									assign node234 = (inp[0]) ? node242 : node235;
										assign node235 = (inp[7]) ? node237 : 3'b000;
											assign node237 = (inp[2]) ? node239 : 3'b001;
												assign node239 = (inp[4]) ? 3'b000 : 3'b001;
										assign node242 = (inp[7]) ? 3'b000 : 3'b001;
									assign node245 = (inp[2]) ? 3'b000 : node246;
										assign node246 = (inp[7]) ? 3'b001 : 3'b000;
						assign node250 = (inp[4]) ? node268 : node251;
							assign node251 = (inp[0]) ? 3'b001 : node252;
								assign node252 = (inp[7]) ? node258 : node253;
									assign node253 = (inp[10]) ? 3'b000 : node254;
										assign node254 = (inp[5]) ? 3'b000 : 3'b001;
									assign node258 = (inp[5]) ? node262 : node259;
										assign node259 = (inp[10]) ? 3'b001 : 3'b000;
										assign node262 = (inp[10]) ? node264 : 3'b001;
											assign node264 = (inp[11]) ? 3'b000 : 3'b001;
							assign node268 = (inp[5]) ? node276 : node269;
								assign node269 = (inp[0]) ? 3'b000 : node270;
									assign node270 = (inp[2]) ? node272 : 3'b001;
										assign node272 = (inp[7]) ? 3'b000 : 3'b001;
								assign node276 = (inp[10]) ? node284 : node277;
									assign node277 = (inp[0]) ? node281 : node278;
										assign node278 = (inp[7]) ? 3'b001 : 3'b000;
										assign node281 = (inp[7]) ? 3'b000 : 3'b001;
									assign node284 = (inp[11]) ? 3'b000 : node285;
										assign node285 = (inp[2]) ? 3'b001 : node286;
											assign node286 = (inp[7]) ? node288 : 3'b000;
												assign node288 = (inp[0]) ? 3'b000 : 3'b001;
			assign node293 = (inp[4]) ? node485 : node294;
				assign node294 = (inp[6]) ? node380 : node295;
					assign node295 = (inp[0]) ? node327 : node296;
						assign node296 = (inp[1]) ? node304 : node297;
							assign node297 = (inp[5]) ? node301 : node298;
								assign node298 = (inp[7]) ? 3'b110 : 3'b010;
								assign node301 = (inp[7]) ? 3'b010 : 3'b100;
							assign node304 = (inp[7]) ? node312 : node305;
								assign node305 = (inp[5]) ? 3'b010 : node306;
									assign node306 = (inp[2]) ? 3'b110 : node307;
										assign node307 = (inp[10]) ? 3'b110 : 3'b101;
								assign node312 = (inp[11]) ? node318 : node313;
									assign node313 = (inp[5]) ? node315 : 3'b001;
										assign node315 = (inp[2]) ? 3'b110 : 3'b001;
									assign node318 = (inp[10]) ? node324 : node319;
										assign node319 = (inp[8]) ? node321 : 3'b101;
											assign node321 = (inp[2]) ? 3'b110 : 3'b101;
										assign node324 = (inp[8]) ? 3'b001 : 3'b110;
						assign node327 = (inp[5]) ? node351 : node328;
							assign node328 = (inp[8]) ? node344 : node329;
								assign node329 = (inp[1]) ? node339 : node330;
									assign node330 = (inp[7]) ? node336 : node331;
										assign node331 = (inp[2]) ? 3'b001 : node332;
											assign node332 = (inp[11]) ? 3'b110 : 3'b010;
										assign node336 = (inp[2]) ? 3'b101 : 3'b001;
									assign node339 = (inp[7]) ? 3'b101 : node340;
										assign node340 = (inp[11]) ? 3'b001 : 3'b101;
								assign node344 = (inp[1]) ? node346 : 3'b001;
									assign node346 = (inp[7]) ? 3'b011 : node347;
										assign node347 = (inp[11]) ? 3'b000 : 3'b100;
							assign node351 = (inp[1]) ? node369 : node352;
								assign node352 = (inp[8]) ? node358 : node353;
									assign node353 = (inp[7]) ? 3'b110 : node354;
										assign node354 = (inp[2]) ? 3'b110 : 3'b010;
									assign node358 = (inp[10]) ? node366 : node359;
										assign node359 = (inp[7]) ? node361 : 3'b110;
											assign node361 = (inp[2]) ? node363 : 3'b110;
												assign node363 = (inp[11]) ? 3'b110 : 3'b010;
										assign node366 = (inp[11]) ? 3'b110 : 3'b101;
								assign node369 = (inp[7]) ? node375 : node370;
									assign node370 = (inp[11]) ? node372 : 3'b111;
										assign node372 = (inp[8]) ? 3'b111 : 3'b110;
									assign node375 = (inp[8]) ? node377 : 3'b001;
										assign node377 = (inp[11]) ? 3'b101 : 3'b111;
					assign node380 = (inp[1]) ? node438 : node381;
						assign node381 = (inp[7]) ? node395 : node382;
							assign node382 = (inp[0]) ? 3'b101 : node383;
								assign node383 = (inp[5]) ? node387 : node384;
									assign node384 = (inp[10]) ? 3'b001 : 3'b101;
									assign node387 = (inp[2]) ? 3'b110 : node388;
										assign node388 = (inp[10]) ? node390 : 3'b110;
											assign node390 = (inp[8]) ? 3'b110 : 3'b010;
							assign node395 = (inp[8]) ? node421 : node396;
								assign node396 = (inp[5]) ? node408 : node397;
									assign node397 = (inp[0]) ? node405 : node398;
										assign node398 = (inp[10]) ? node400 : 3'b001;
											assign node400 = (inp[2]) ? 3'b101 : node401;
												assign node401 = (inp[11]) ? 3'b001 : 3'b101;
										assign node405 = (inp[10]) ? 3'b011 : 3'b001;
									assign node408 = (inp[0]) ? node416 : node409;
										assign node409 = (inp[11]) ? node411 : 3'b010;
											assign node411 = (inp[2]) ? 3'b010 : node412;
												assign node412 = (inp[10]) ? 3'b110 : 3'b010;
										assign node416 = (inp[2]) ? node418 : 3'b101;
											assign node418 = (inp[10]) ? 3'b011 : 3'b001;
								assign node421 = (inp[0]) ? node427 : node422;
									assign node422 = (inp[5]) ? 3'b001 : node423;
										assign node423 = (inp[10]) ? 3'b101 : 3'b001;
									assign node427 = (inp[5]) ? node433 : node428;
										assign node428 = (inp[2]) ? 3'b111 : node429;
											assign node429 = (inp[10]) ? 3'b011 : 3'b001;
										assign node433 = (inp[11]) ? node435 : 3'b101;
											assign node435 = (inp[2]) ? 3'b001 : 3'b101;
						assign node438 = (inp[5]) ? node468 : node439;
							assign node439 = (inp[0]) ? node459 : node440;
								assign node440 = (inp[10]) ? node450 : node441;
									assign node441 = (inp[7]) ? node447 : node442;
										assign node442 = (inp[2]) ? node444 : 3'b011;
											assign node444 = (inp[8]) ? 3'b011 : 3'b001;
										assign node447 = (inp[8]) ? 3'b001 : 3'b011;
									assign node450 = (inp[7]) ? node454 : node451;
										assign node451 = (inp[8]) ? 3'b101 : 3'b001;
										assign node454 = (inp[2]) ? node456 : 3'b011;
											assign node456 = (inp[8]) ? 3'b011 : 3'b001;
								assign node459 = (inp[7]) ? 3'b111 : node460;
									assign node460 = (inp[10]) ? node462 : 3'b011;
										assign node462 = (inp[2]) ? node464 : 3'b011;
											assign node464 = (inp[8]) ? 3'b111 : 3'b011;
							assign node468 = (inp[8]) ? node480 : node469;
								assign node469 = (inp[0]) ? node473 : node470;
									assign node470 = (inp[7]) ? 3'b011 : 3'b001;
									assign node473 = (inp[7]) ? 3'b001 : node474;
										assign node474 = (inp[2]) ? node476 : 3'b001;
											assign node476 = (inp[10]) ? 3'b101 : 3'b001;
								assign node480 = (inp[0]) ? 3'b011 : node481;
									assign node481 = (inp[10]) ? 3'b001 : 3'b011;
				assign node485 = (inp[0]) ? node583 : node486;
					assign node486 = (inp[6]) ? node538 : node487;
						assign node487 = (inp[5]) ? node521 : node488;
							assign node488 = (inp[1]) ? node500 : node489;
								assign node489 = (inp[10]) ? node491 : 3'b100;
									assign node491 = (inp[7]) ? 3'b100 : node492;
										assign node492 = (inp[2]) ? node494 : 3'b000;
											assign node494 = (inp[11]) ? node496 : 3'b100;
												assign node496 = (inp[8]) ? 3'b100 : 3'b000;
								assign node500 = (inp[7]) ? node510 : node501;
									assign node501 = (inp[10]) ? node505 : node502;
										assign node502 = (inp[8]) ? 3'b110 : 3'b010;
										assign node505 = (inp[8]) ? 3'b100 : node506;
											assign node506 = (inp[2]) ? 3'b100 : 3'b000;
									assign node510 = (inp[10]) ? 3'b010 : node511;
										assign node511 = (inp[11]) ? node513 : 3'b010;
											assign node513 = (inp[8]) ? node517 : node514;
												assign node514 = (inp[2]) ? 3'b000 : 3'b110;
												assign node517 = (inp[2]) ? 3'b010 : 3'b000;
							assign node521 = (inp[1]) ? node523 : 3'b000;
								assign node523 = (inp[7]) ? node529 : node524;
									assign node524 = (inp[11]) ? 3'b000 : node525;
										assign node525 = (inp[8]) ? 3'b010 : 3'b000;
									assign node529 = (inp[8]) ? node531 : 3'b100;
										assign node531 = (inp[11]) ? node533 : 3'b110;
											assign node533 = (inp[10]) ? 3'b100 : node534;
												assign node534 = (inp[2]) ? 3'b100 : 3'b110;
						assign node538 = (inp[8]) ? node554 : node539;
							assign node539 = (inp[1]) ? node547 : node540;
								assign node540 = (inp[7]) ? node542 : 3'b100;
									assign node542 = (inp[11]) ? 3'b100 : node543;
										assign node543 = (inp[10]) ? 3'b010 : 3'b000;
								assign node547 = (inp[5]) ? node549 : 3'b110;
									assign node549 = (inp[7]) ? node551 : 3'b100;
										assign node551 = (inp[10]) ? 3'b101 : 3'b010;
							assign node554 = (inp[1]) ? node572 : node555;
								assign node555 = (inp[5]) ? node561 : node556;
									assign node556 = (inp[7]) ? node558 : 3'b010;
										assign node558 = (inp[10]) ? 3'b110 : 3'b100;
									assign node561 = (inp[11]) ? node567 : node562;
										assign node562 = (inp[10]) ? 3'b010 : node563;
											assign node563 = (inp[7]) ? 3'b000 : 3'b010;
										assign node567 = (inp[2]) ? 3'b010 : node568;
											assign node568 = (inp[10]) ? 3'b100 : 3'b000;
								assign node572 = (inp[7]) ? node576 : node573;
									assign node573 = (inp[5]) ? 3'b100 : 3'b110;
									assign node576 = (inp[10]) ? node580 : node577;
										assign node577 = (inp[2]) ? 3'b010 : 3'b110;
										assign node580 = (inp[5]) ? 3'b110 : 3'b001;
					assign node583 = (inp[6]) ? node615 : node584;
						assign node584 = (inp[1]) ? node602 : node585;
							assign node585 = (inp[5]) ? node591 : node586;
								assign node586 = (inp[2]) ? 3'b010 : node587;
									assign node587 = (inp[7]) ? 3'b010 : 3'b100;
								assign node591 = (inp[7]) ? 3'b100 : node592;
									assign node592 = (inp[8]) ? node596 : node593;
										assign node593 = (inp[2]) ? 3'b100 : 3'b000;
										assign node596 = (inp[2]) ? 3'b100 : node597;
											assign node597 = (inp[11]) ? 3'b100 : 3'b110;
							assign node602 = (inp[5]) ? node608 : node603;
								assign node603 = (inp[7]) ? 3'b110 : node604;
									assign node604 = (inp[8]) ? 3'b100 : 3'b010;
								assign node608 = (inp[7]) ? 3'b010 : node609;
									assign node609 = (inp[8]) ? 3'b010 : node610;
										assign node610 = (inp[11]) ? 3'b100 : 3'b010;
						assign node615 = (inp[5]) ? node625 : node616;
							assign node616 = (inp[7]) ? node618 : 3'b001;
								assign node618 = (inp[1]) ? 3'b101 : node619;
									assign node619 = (inp[10]) ? node621 : 3'b001;
										assign node621 = (inp[2]) ? 3'b101 : 3'b001;
							assign node625 = (inp[1]) ? node631 : node626;
								assign node626 = (inp[7]) ? node628 : 3'b010;
									assign node628 = (inp[10]) ? 3'b110 : 3'b010;
								assign node631 = (inp[7]) ? 3'b001 : 3'b110;
		assign node634 = (inp[6]) ? node656 : node635;
			assign node635 = (inp[9]) ? node637 : 3'b000;
				assign node637 = (inp[0]) ? node639 : 3'b000;
					assign node639 = (inp[4]) ? 3'b000 : node640;
						assign node640 = (inp[1]) ? node642 : 3'b000;
							assign node642 = (inp[5]) ? node648 : node643;
								assign node643 = (inp[7]) ? 3'b100 : node644;
									assign node644 = (inp[8]) ? 3'b100 : 3'b000;
								assign node648 = (inp[7]) ? 3'b000 : node649;
									assign node649 = (inp[10]) ? node651 : 3'b000;
										assign node651 = (inp[2]) ? 3'b100 : 3'b000;
			assign node656 = (inp[9]) ? node794 : node657;
				assign node657 = (inp[4]) ? node683 : node658;
					assign node658 = (inp[0]) ? node676 : node659;
						assign node659 = (inp[7]) ? node661 : 3'b010;
							assign node661 = (inp[1]) ? node663 : 3'b010;
								assign node663 = (inp[2]) ? node665 : 3'b010;
									assign node665 = (inp[11]) ? node671 : node666;
										assign node666 = (inp[5]) ? 3'b010 : node667;
											assign node667 = (inp[8]) ? 3'b011 : 3'b010;
										assign node671 = (inp[5]) ? 3'b011 : node672;
											assign node672 = (inp[8]) ? 3'b011 : 3'b010;
						assign node676 = (inp[5]) ? node678 : 3'b011;
							assign node678 = (inp[1]) ? node680 : 3'b010;
								assign node680 = (inp[7]) ? 3'b011 : 3'b010;
					assign node683 = (inp[0]) ? node731 : node684;
						assign node684 = (inp[10]) ? node714 : node685;
							assign node685 = (inp[7]) ? node699 : node686;
								assign node686 = (inp[1]) ? node694 : node687;
									assign node687 = (inp[5]) ? node691 : node688;
										assign node688 = (inp[11]) ? 3'b010 : 3'b000;
										assign node691 = (inp[11]) ? 3'b000 : 3'b010;
									assign node694 = (inp[11]) ? node696 : 3'b000;
										assign node696 = (inp[5]) ? 3'b100 : 3'b000;
								assign node699 = (inp[1]) ? node703 : node700;
									assign node700 = (inp[8]) ? 3'b010 : 3'b100;
									assign node703 = (inp[8]) ? node705 : 3'b010;
										assign node705 = (inp[11]) ? node707 : 3'b010;
											assign node707 = (inp[5]) ? node711 : node708;
												assign node708 = (inp[2]) ? 3'b100 : 3'b010;
												assign node711 = (inp[2]) ? 3'b010 : 3'b100;
							assign node714 = (inp[5]) ? node716 : 3'b000;
								assign node716 = (inp[1]) ? node718 : 3'b000;
									assign node718 = (inp[11]) ? node726 : node719;
										assign node719 = (inp[7]) ? node721 : 3'b000;
											assign node721 = (inp[2]) ? 3'b100 : node722;
												assign node722 = (inp[8]) ? 3'b100 : 3'b000;
										assign node726 = (inp[8]) ? 3'b100 : node727;
											assign node727 = (inp[7]) ? 3'b000 : 3'b100;
						assign node731 = (inp[7]) ? node753 : node732;
							assign node732 = (inp[10]) ? node744 : node733;
								assign node733 = (inp[1]) ? node739 : node734;
									assign node734 = (inp[8]) ? node736 : 3'b100;
										assign node736 = (inp[2]) ? 3'b010 : 3'b100;
									assign node739 = (inp[5]) ? node741 : 3'b110;
										assign node741 = (inp[2]) ? 3'b110 : 3'b010;
								assign node744 = (inp[1]) ? node746 : 3'b100;
									assign node746 = (inp[8]) ? node748 : 3'b100;
										assign node748 = (inp[5]) ? node750 : 3'b010;
											assign node750 = (inp[11]) ? 3'b100 : 3'b010;
							assign node753 = (inp[1]) ? node771 : node754;
								assign node754 = (inp[10]) ? node764 : node755;
									assign node755 = (inp[2]) ? node759 : node756;
										assign node756 = (inp[8]) ? 3'b110 : 3'b010;
										assign node759 = (inp[8]) ? 3'b010 : node760;
											assign node760 = (inp[5]) ? 3'b010 : 3'b110;
									assign node764 = (inp[8]) ? 3'b010 : node765;
										assign node765 = (inp[11]) ? 3'b100 : node766;
											assign node766 = (inp[2]) ? 3'b010 : 3'b100;
								assign node771 = (inp[10]) ? node787 : node772;
									assign node772 = (inp[8]) ? node782 : node773;
										assign node773 = (inp[5]) ? node777 : node774;
											assign node774 = (inp[2]) ? 3'b110 : 3'b101;
											assign node777 = (inp[11]) ? node779 : 3'b110;
												assign node779 = (inp[2]) ? 3'b110 : 3'b010;
										assign node782 = (inp[11]) ? 3'b001 : node783;
											assign node783 = (inp[2]) ? 3'b001 : 3'b101;
									assign node787 = (inp[5]) ? node789 : 3'b110;
										assign node789 = (inp[11]) ? 3'b010 : node790;
											assign node790 = (inp[2]) ? 3'b110 : 3'b010;
				assign node794 = (inp[0]) ? node828 : node795;
					assign node795 = (inp[4]) ? 3'b000 : node796;
						assign node796 = (inp[10]) ? node810 : node797;
							assign node797 = (inp[2]) ? node799 : 3'b000;
								assign node799 = (inp[1]) ? node801 : 3'b000;
									assign node801 = (inp[7]) ? node803 : 3'b000;
										assign node803 = (inp[11]) ? 3'b010 : node804;
											assign node804 = (inp[5]) ? 3'b000 : node805;
												assign node805 = (inp[8]) ? 3'b010 : 3'b000;
							assign node810 = (inp[1]) ? node818 : node811;
								assign node811 = (inp[7]) ? node813 : 3'b000;
									assign node813 = (inp[8]) ? node815 : 3'b000;
										assign node815 = (inp[5]) ? 3'b000 : 3'b100;
								assign node818 = (inp[2]) ? node822 : node819;
									assign node819 = (inp[7]) ? 3'b100 : 3'b000;
									assign node822 = (inp[7]) ? node824 : 3'b100;
										assign node824 = (inp[11]) ? 3'b010 : 3'b100;
					assign node828 = (inp[4]) ? node840 : node829;
						assign node829 = (inp[5]) ? node835 : node830;
							assign node830 = (inp[1]) ? node832 : 3'b010;
								assign node832 = (inp[7]) ? 3'b110 : 3'b010;
							assign node835 = (inp[7]) ? node837 : 3'b100;
								assign node837 = (inp[1]) ? 3'b010 : 3'b100;
						assign node840 = (inp[7]) ? node848 : node841;
							assign node841 = (inp[10]) ? 3'b000 : node842;
								assign node842 = (inp[5]) ? 3'b000 : node843;
									assign node843 = (inp[11]) ? 3'b000 : 3'b100;
							assign node848 = (inp[1]) ? node858 : node849;
								assign node849 = (inp[10]) ? 3'b000 : node850;
									assign node850 = (inp[8]) ? node852 : 3'b000;
										assign node852 = (inp[5]) ? node854 : 3'b100;
											assign node854 = (inp[11]) ? 3'b000 : 3'b100;
								assign node858 = (inp[5]) ? node864 : node859;
									assign node859 = (inp[8]) ? node861 : 3'b100;
										assign node861 = (inp[10]) ? 3'b100 : 3'b010;
									assign node864 = (inp[10]) ? 3'b000 : node865;
										assign node865 = (inp[8]) ? 3'b100 : node866;
											assign node866 = (inp[2]) ? 3'b100 : node867;
												assign node867 = (inp[11]) ? 3'b000 : 3'b100;

endmodule