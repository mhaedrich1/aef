module dtc_split5_bm60 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node88;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node234;

	assign outp = (inp[2]) ? node92 : node1;
		assign node1 = (inp[4]) ? node35 : node2;
			assign node2 = (inp[10]) ? node24 : node3;
				assign node3 = (inp[5]) ? node5 : 3'b111;
					assign node5 = (inp[9]) ? node7 : 3'b111;
						assign node7 = (inp[3]) ? node17 : node8;
							assign node8 = (inp[7]) ? node10 : 3'b111;
								assign node10 = (inp[6]) ? node12 : 3'b111;
									assign node12 = (inp[8]) ? node14 : 3'b111;
										assign node14 = (inp[11]) ? 3'b110 : 3'b111;
							assign node17 = (inp[7]) ? 3'b110 : node18;
								assign node18 = (inp[6]) ? node20 : 3'b111;
									assign node20 = (inp[8]) ? 3'b110 : 3'b111;
				assign node24 = (inp[5]) ? node26 : 3'b110;
					assign node26 = (inp[9]) ? node28 : 3'b110;
						assign node28 = (inp[3]) ? 3'b011 : node29;
							assign node29 = (inp[7]) ? node31 : 3'b110;
								assign node31 = (inp[8]) ? 3'b111 : 3'b110;
			assign node35 = (inp[3]) ? node61 : node36;
				assign node36 = (inp[5]) ? node56 : node37;
					assign node37 = (inp[10]) ? node45 : node38;
						assign node38 = (inp[7]) ? node40 : 3'b110;
							assign node40 = (inp[9]) ? node42 : 3'b110;
								assign node42 = (inp[8]) ? 3'b111 : 3'b110;
						assign node45 = (inp[9]) ? 3'b110 : node46;
							assign node46 = (inp[7]) ? 3'b110 : node47;
								assign node47 = (inp[8]) ? node49 : 3'b111;
									assign node49 = (inp[11]) ? node51 : 3'b111;
										assign node51 = (inp[6]) ? 3'b110 : 3'b111;
					assign node56 = (inp[10]) ? node58 : 3'b111;
						assign node58 = (inp[9]) ? 3'b011 : 3'b110;
				assign node61 = (inp[5]) ? node83 : node62;
					assign node62 = (inp[9]) ? node64 : 3'b011;
						assign node64 = (inp[7]) ? node74 : node65;
							assign node65 = (inp[11]) ? node67 : 3'b011;
								assign node67 = (inp[8]) ? node69 : 3'b011;
									assign node69 = (inp[6]) ? node71 : 3'b011;
										assign node71 = (inp[10]) ? 3'b011 : 3'b010;
							assign node74 = (inp[10]) ? node76 : 3'b010;
								assign node76 = (inp[6]) ? node78 : 3'b011;
									assign node78 = (inp[11]) ? node80 : 3'b011;
										assign node80 = (inp[8]) ? 3'b010 : 3'b011;
					assign node83 = (inp[8]) ? node85 : 3'b010;
						assign node85 = (inp[10]) ? 3'b010 : node86;
							assign node86 = (inp[9]) ? node88 : 3'b010;
								assign node88 = (inp[7]) ? 3'b011 : 3'b010;
		assign node92 = (inp[4]) ? node144 : node93;
			assign node93 = (inp[10]) ? node121 : node94;
				assign node94 = (inp[5]) ? node108 : node95;
					assign node95 = (inp[3]) ? node97 : 3'b011;
						assign node97 = (inp[9]) ? 3'b010 : node98;
							assign node98 = (inp[8]) ? node100 : 3'b011;
								assign node100 = (inp[6]) ? node102 : 3'b011;
									assign node102 = (inp[11]) ? node104 : 3'b011;
										assign node104 = (inp[7]) ? 3'b010 : 3'b011;
					assign node108 = (inp[3]) ? 3'b010 : node109;
						assign node109 = (inp[7]) ? 3'b010 : node110;
							assign node110 = (inp[9]) ? 3'b010 : node111;
								assign node111 = (inp[6]) ? node113 : 3'b011;
									assign node113 = (inp[8]) ? node115 : 3'b011;
										assign node115 = (inp[11]) ? 3'b010 : 3'b011;
				assign node121 = (inp[3]) ? node131 : node122;
					assign node122 = (inp[5]) ? 3'b011 : node123;
						assign node123 = (inp[7]) ? node125 : 3'b010;
							assign node125 = (inp[9]) ? node127 : 3'b010;
								assign node127 = (inp[8]) ? 3'b011 : 3'b010;
					assign node131 = (inp[5]) ? node133 : 3'b111;
						assign node133 = (inp[9]) ? 3'b110 : node134;
							assign node134 = (inp[11]) ? node136 : 3'b111;
								assign node136 = (inp[8]) ? node138 : 3'b111;
									assign node138 = (inp[7]) ? node140 : 3'b111;
										assign node140 = (inp[6]) ? 3'b110 : 3'b111;
			assign node144 = (inp[3]) ? node176 : node145;
				assign node145 = (inp[5]) ? node167 : node146;
					assign node146 = (inp[9]) ? node148 : 3'b101;
						assign node148 = (inp[7]) ? node158 : node149;
							assign node149 = (inp[6]) ? node151 : 3'b101;
								assign node151 = (inp[0]) ? 3'b101 : node152;
									assign node152 = (inp[8]) ? node154 : 3'b101;
										assign node154 = (inp[11]) ? 3'b100 : 3'b101;
							assign node158 = (inp[10]) ? 3'b100 : node159;
								assign node159 = (inp[11]) ? node161 : 3'b101;
									assign node161 = (inp[8]) ? node163 : 3'b101;
										assign node163 = (inp[6]) ? 3'b100 : 3'b101;
					assign node167 = (inp[9]) ? node169 : 3'b100;
						assign node169 = (inp[10]) ? 3'b001 : node170;
							assign node170 = (inp[7]) ? node172 : 3'b100;
								assign node172 = (inp[8]) ? 3'b101 : 3'b100;
				assign node176 = (inp[10]) ? node204 : node177;
					assign node177 = (inp[9]) ? node197 : node178;
						assign node178 = (inp[7]) ? node188 : node179;
							assign node179 = (inp[11]) ? node181 : 3'b001;
								assign node181 = (inp[6]) ? node183 : 3'b001;
									assign node183 = (inp[1]) ? node185 : 3'b001;
										assign node185 = (inp[8]) ? 3'b000 : 3'b001;
							assign node188 = (inp[5]) ? node190 : 3'b000;
								assign node190 = (inp[1]) ? node192 : 3'b001;
									assign node192 = (inp[8]) ? node194 : 3'b001;
										assign node194 = (inp[6]) ? 3'b000 : 3'b001;
						assign node197 = (inp[5]) ? 3'b000 : node198;
							assign node198 = (inp[7]) ? node200 : 3'b000;
								assign node200 = (inp[8]) ? 3'b001 : 3'b000;
					assign node204 = (inp[9]) ? node222 : node205;
						assign node205 = (inp[5]) ? node215 : node206;
							assign node206 = (inp[8]) ? node208 : 3'b101;
								assign node208 = (inp[1]) ? 3'b101 : node209;
									assign node209 = (inp[6]) ? node211 : 3'b101;
										assign node211 = (inp[11]) ? 3'b100 : 3'b101;
							assign node215 = (inp[7]) ? 3'b100 : node216;
								assign node216 = (inp[8]) ? node218 : 3'b101;
									assign node218 = (inp[11]) ? 3'b100 : 3'b101;
						assign node222 = (inp[5]) ? node228 : node223;
							assign node223 = (inp[8]) ? node225 : 3'b100;
								assign node225 = (inp[7]) ? 3'b101 : 3'b100;
							assign node228 = (inp[7]) ? node230 : 3'b001;
								assign node230 = (inp[8]) ? node232 : 3'b000;
									assign node232 = (inp[6]) ? node234 : 3'b001;
										assign node234 = (inp[11]) ? 3'b000 : 3'b001;

endmodule