module dtc_split75_bm97 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node61;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node205;

	assign outp = (inp[3]) ? node50 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b000;
			assign node3 = (inp[9]) ? node5 : 3'b000;
				assign node5 = (inp[7]) ? node7 : 3'b001;
					assign node7 = (inp[10]) ? node9 : 3'b000;
						assign node9 = (inp[4]) ? node29 : node10;
							assign node10 = (inp[11]) ? node12 : 3'b000;
								assign node12 = (inp[5]) ? node16 : node13;
									assign node13 = (inp[8]) ? 3'b100 : 3'b000;
									assign node16 = (inp[8]) ? node20 : node17;
										assign node17 = (inp[1]) ? 3'b101 : 3'b001;
										assign node20 = (inp[0]) ? node24 : node21;
											assign node21 = (inp[2]) ? 3'b100 : 3'b101;
											assign node24 = (inp[1]) ? node26 : 3'b101;
												assign node26 = (inp[2]) ? 3'b001 : 3'b101;
							assign node29 = (inp[11]) ? node31 : 3'b100;
								assign node31 = (inp[5]) ? node39 : node32;
									assign node32 = (inp[8]) ? node34 : 3'b000;
										assign node34 = (inp[1]) ? node36 : 3'b100;
											assign node36 = (inp[2]) ? 3'b110 : 3'b100;
									assign node39 = (inp[8]) ? node45 : node40;
										assign node40 = (inp[1]) ? node42 : 3'b010;
											assign node42 = (inp[0]) ? 3'b110 : 3'b010;
										assign node45 = (inp[2]) ? node47 : 3'b110;
											assign node47 = (inp[1]) ? 3'b010 : 3'b110;
		assign node50 = (inp[9]) ? node94 : node51;
			assign node51 = (inp[6]) ? 3'b000 : node52;
				assign node52 = (inp[7]) ? 3'b000 : node53;
					assign node53 = (inp[4]) ? node55 : 3'b100;
						assign node55 = (inp[11]) ? node65 : node56;
							assign node56 = (inp[8]) ? 3'b100 : node57;
								assign node57 = (inp[10]) ? node59 : 3'b100;
									assign node59 = (inp[1]) ? node61 : 3'b000;
										assign node61 = (inp[2]) ? 3'b100 : 3'b000;
							assign node65 = (inp[5]) ? node81 : node66;
								assign node66 = (inp[10]) ? node74 : node67;
									assign node67 = (inp[1]) ? node69 : 3'b100;
										assign node69 = (inp[0]) ? node71 : 3'b100;
											assign node71 = (inp[8]) ? 3'b000 : 3'b100;
									assign node74 = (inp[8]) ? 3'b000 : node75;
										assign node75 = (inp[1]) ? node77 : 3'b100;
											assign node77 = (inp[0]) ? 3'b000 : 3'b100;
								assign node81 = (inp[0]) ? 3'b000 : node82;
									assign node82 = (inp[10]) ? node88 : node83;
										assign node83 = (inp[8]) ? node85 : 3'b000;
											assign node85 = (inp[2]) ? 3'b100 : 3'b000;
										assign node88 = (inp[8]) ? 3'b000 : 3'b100;
			assign node94 = (inp[4]) ? node130 : node95;
				assign node95 = (inp[6]) ? node99 : node96;
					assign node96 = (inp[7]) ? 3'b110 : 3'b000;
					assign node99 = (inp[7]) ? node101 : 3'b110;
						assign node101 = (inp[10]) ? node103 : 3'b000;
							assign node103 = (inp[5]) ? node115 : node104;
								assign node104 = (inp[0]) ? node106 : 3'b010;
									assign node106 = (inp[1]) ? node108 : 3'b010;
										assign node108 = (inp[2]) ? node110 : 3'b010;
											assign node110 = (inp[8]) ? node112 : 3'b010;
												assign node112 = (inp[11]) ? 3'b100 : 3'b000;
								assign node115 = (inp[11]) ? node123 : node116;
									assign node116 = (inp[8]) ? node118 : 3'b000;
										assign node118 = (inp[0]) ? 3'b000 : node119;
											assign node119 = (inp[2]) ? 3'b010 : 3'b000;
									assign node123 = (inp[0]) ? 3'b100 : node124;
										assign node124 = (inp[2]) ? node126 : 3'b100;
											assign node126 = (inp[8]) ? 3'b010 : 3'b100;
				assign node130 = (inp[6]) ? node186 : node131;
					assign node131 = (inp[7]) ? node167 : node132;
						assign node132 = (inp[10]) ? node150 : node133;
							assign node133 = (inp[11]) ? node135 : 3'b010;
								assign node135 = (inp[5]) ? node143 : node136;
									assign node136 = (inp[1]) ? node138 : 3'b010;
										assign node138 = (inp[0]) ? node140 : 3'b010;
											assign node140 = (inp[8]) ? 3'b110 : 3'b010;
									assign node143 = (inp[2]) ? node145 : 3'b110;
										assign node145 = (inp[0]) ? 3'b110 : node146;
											assign node146 = (inp[8]) ? 3'b010 : 3'b110;
							assign node150 = (inp[11]) ? node158 : node151;
								assign node151 = (inp[8]) ? 3'b001 : node152;
									assign node152 = (inp[2]) ? node154 : 3'b101;
										assign node154 = (inp[1]) ? 3'b001 : 3'b101;
								assign node158 = (inp[8]) ? 3'b101 : node159;
									assign node159 = (inp[0]) ? node161 : 3'b011;
										assign node161 = (inp[1]) ? 3'b101 : node162;
											assign node162 = (inp[5]) ? 3'b101 : 3'b011;
						assign node167 = (inp[10]) ? node169 : 3'b001;
							assign node169 = (inp[11]) ? node171 : 3'b001;
								assign node171 = (inp[8]) ? node177 : node172;
									assign node172 = (inp[0]) ? node174 : 3'b001;
										assign node174 = (inp[5]) ? 3'b110 : 3'b001;
									assign node177 = (inp[0]) ? node179 : 3'b110;
										assign node179 = (inp[5]) ? node181 : 3'b110;
											assign node181 = (inp[1]) ? node183 : 3'b110;
												assign node183 = (inp[2]) ? 3'b001 : 3'b110;
					assign node186 = (inp[7]) ? 3'b000 : node187;
						assign node187 = (inp[11]) ? node189 : 3'b000;
							assign node189 = (inp[10]) ? node191 : 3'b000;
								assign node191 = (inp[8]) ? node199 : node192;
									assign node192 = (inp[0]) ? node194 : 3'b010;
										assign node194 = (inp[1]) ? node196 : 3'b010;
											assign node196 = (inp[5]) ? 3'b100 : 3'b010;
									assign node199 = (inp[2]) ? node201 : 3'b100;
										assign node201 = (inp[1]) ? node203 : 3'b100;
											assign node203 = (inp[5]) ? node205 : 3'b100;
												assign node205 = (inp[0]) ? 3'b000 : 3'b100;

endmodule