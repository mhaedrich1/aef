module dtc_split125_bm81 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node48;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node358;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node420;
	wire [3-1:0] node422;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;

	assign outp = (inp[9]) ? node166 : node1;
		assign node1 = (inp[3]) ? node123 : node2;
			assign node2 = (inp[6]) ? node82 : node3;
				assign node3 = (inp[4]) ? node31 : node4;
					assign node4 = (inp[7]) ? node10 : node5;
						assign node5 = (inp[10]) ? 3'b001 : node6;
							assign node6 = (inp[5]) ? 3'b000 : 3'b001;
						assign node10 = (inp[10]) ? node20 : node11;
							assign node11 = (inp[11]) ? node17 : node12;
								assign node12 = (inp[8]) ? 3'b100 : node13;
									assign node13 = (inp[5]) ? 3'b000 : 3'b100;
								assign node17 = (inp[0]) ? 3'b100 : 3'b101;
							assign node20 = (inp[1]) ? node26 : node21;
								assign node21 = (inp[0]) ? 3'b001 : node22;
									assign node22 = (inp[8]) ? 3'b101 : 3'b001;
								assign node26 = (inp[2]) ? 3'b101 : node27;
									assign node27 = (inp[5]) ? 3'b101 : 3'b001;
					assign node31 = (inp[10]) ? node55 : node32;
						assign node32 = (inp[7]) ? node48 : node33;
							assign node33 = (inp[0]) ? node41 : node34;
								assign node34 = (inp[1]) ? node36 : 3'b001;
									assign node36 = (inp[2]) ? node38 : 3'b010;
										assign node38 = (inp[5]) ? 3'b110 : 3'b100;
								assign node41 = (inp[2]) ? 3'b010 : node42;
									assign node42 = (inp[1]) ? 3'b110 : node43;
										assign node43 = (inp[8]) ? 3'b010 : 3'b110;
							assign node48 = (inp[11]) ? node50 : 3'b000;
								assign node50 = (inp[8]) ? 3'b100 : node51;
									assign node51 = (inp[1]) ? 3'b010 : 3'b100;
						assign node55 = (inp[7]) ? node71 : node56;
							assign node56 = (inp[2]) ? node68 : node57;
								assign node57 = (inp[0]) ? node61 : node58;
									assign node58 = (inp[8]) ? 3'b001 : 3'b011;
									assign node61 = (inp[11]) ? 3'b101 : node62;
										assign node62 = (inp[5]) ? 3'b001 : node63;
											assign node63 = (inp[8]) ? 3'b001 : 3'b101;
								assign node68 = (inp[0]) ? 3'b110 : 3'b001;
							assign node71 = (inp[2]) ? node79 : node72;
								assign node72 = (inp[0]) ? 3'b010 : node73;
									assign node73 = (inp[1]) ? 3'b110 : node74;
										assign node74 = (inp[5]) ? 3'b010 : 3'b110;
								assign node79 = (inp[0]) ? 3'b110 : 3'b001;
				assign node82 = (inp[4]) ? node112 : node83;
					assign node83 = (inp[10]) ? node95 : node84;
						assign node84 = (inp[7]) ? 3'b000 : node85;
							assign node85 = (inp[8]) ? node87 : 3'b100;
								assign node87 = (inp[11]) ? node89 : 3'b000;
									assign node89 = (inp[0]) ? node91 : 3'b100;
										assign node91 = (inp[5]) ? 3'b000 : 3'b100;
						assign node95 = (inp[7]) ? node103 : node96;
							assign node96 = (inp[1]) ? node100 : node97;
								assign node97 = (inp[11]) ? 3'b011 : 3'b010;
								assign node100 = (inp[8]) ? 3'b100 : 3'b110;
							assign node103 = (inp[5]) ? 3'b000 : node104;
								assign node104 = (inp[8]) ? node108 : node105;
									assign node105 = (inp[0]) ? 3'b100 : 3'b010;
									assign node108 = (inp[11]) ? 3'b100 : 3'b000;
					assign node112 = (inp[8]) ? 3'b000 : node113;
						assign node113 = (inp[7]) ? 3'b000 : node114;
							assign node114 = (inp[5]) ? node118 : node115;
								assign node115 = (inp[10]) ? 3'b010 : 3'b000;
								assign node118 = (inp[10]) ? 3'b100 : 3'b000;
			assign node123 = (inp[6]) ? 3'b000 : node124;
				assign node124 = (inp[4]) ? node152 : node125;
					assign node125 = (inp[10]) ? node139 : node126;
						assign node126 = (inp[7]) ? 3'b000 : node127;
							assign node127 = (inp[0]) ? 3'b100 : node128;
								assign node128 = (inp[8]) ? 3'b000 : node129;
									assign node129 = (inp[1]) ? 3'b100 : node130;
										assign node130 = (inp[11]) ? 3'b010 : node131;
											assign node131 = (inp[5]) ? 3'b000 : 3'b100;
						assign node139 = (inp[7]) ? node145 : node140;
							assign node140 = (inp[8]) ? 3'b010 : node141;
								assign node141 = (inp[0]) ? 3'b110 : 3'b010;
							assign node145 = (inp[2]) ? node149 : node146;
								assign node146 = (inp[8]) ? 3'b000 : 3'b100;
								assign node149 = (inp[0]) ? 3'b010 : 3'b100;
					assign node152 = (inp[7]) ? 3'b000 : node153;
						assign node153 = (inp[8]) ? node157 : node154;
							assign node154 = (inp[1]) ? 3'b000 : 3'b010;
							assign node157 = (inp[5]) ? 3'b000 : node158;
								assign node158 = (inp[10]) ? node160 : 3'b000;
									assign node160 = (inp[11]) ? 3'b100 : 3'b000;
		assign node166 = (inp[6]) ? node280 : node167;
			assign node167 = (inp[3]) ? node205 : node168;
				assign node168 = (inp[7]) ? node184 : node169;
					assign node169 = (inp[10]) ? 3'b111 : node170;
						assign node170 = (inp[4]) ? node172 : 3'b111;
							assign node172 = (inp[0]) ? node178 : node173;
								assign node173 = (inp[2]) ? 3'b011 : node174;
									assign node174 = (inp[11]) ? 3'b111 : 3'b011;
								assign node178 = (inp[5]) ? 3'b111 : node179;
									assign node179 = (inp[2]) ? 3'b001 : 3'b111;
					assign node184 = (inp[5]) ? node194 : node185;
						assign node185 = (inp[8]) ? node191 : node186;
							assign node186 = (inp[10]) ? 3'b111 : node187;
								assign node187 = (inp[1]) ? 3'b001 : 3'b101;
							assign node191 = (inp[4]) ? 3'b101 : 3'b111;
						assign node194 = (inp[4]) ? node202 : node195;
							assign node195 = (inp[8]) ? 3'b011 : node196;
								assign node196 = (inp[11]) ? node198 : 3'b111;
									assign node198 = (inp[2]) ? 3'b001 : 3'b111;
							assign node202 = (inp[10]) ? 3'b011 : 3'b001;
				assign node205 = (inp[11]) ? node237 : node206;
					assign node206 = (inp[7]) ? node222 : node207;
						assign node207 = (inp[8]) ? 3'b110 : node208;
							assign node208 = (inp[5]) ? node216 : node209;
								assign node209 = (inp[4]) ? node213 : node210;
									assign node210 = (inp[2]) ? 3'b101 : 3'b111;
									assign node213 = (inp[10]) ? 3'b101 : 3'b110;
								assign node216 = (inp[10]) ? 3'b001 : node217;
									assign node217 = (inp[4]) ? 3'b010 : 3'b001;
						assign node222 = (inp[10]) ? node230 : node223;
							assign node223 = (inp[4]) ? node225 : 3'b100;
								assign node225 = (inp[8]) ? 3'b000 : node226;
									assign node226 = (inp[5]) ? 3'b000 : 3'b100;
							assign node230 = (inp[0]) ? node232 : 3'b001;
								assign node232 = (inp[2]) ? 3'b010 : node233;
									assign node233 = (inp[4]) ? 3'b100 : 3'b110;
					assign node237 = (inp[4]) ? node259 : node238;
						assign node238 = (inp[5]) ? node250 : node239;
							assign node239 = (inp[0]) ? node245 : node240;
								assign node240 = (inp[10]) ? node242 : 3'b101;
									assign node242 = (inp[8]) ? 3'b011 : 3'b111;
								assign node245 = (inp[8]) ? node247 : 3'b011;
									assign node247 = (inp[7]) ? 3'b011 : 3'b111;
							assign node250 = (inp[8]) ? 3'b001 : node251;
								assign node251 = (inp[7]) ? node255 : node252;
									assign node252 = (inp[10]) ? 3'b111 : 3'b001;
									assign node255 = (inp[10]) ? 3'b101 : 3'b110;
						assign node259 = (inp[10]) ? node261 : 3'b110;
							assign node261 = (inp[0]) ? node269 : node262;
								assign node262 = (inp[8]) ? 3'b101 : node263;
									assign node263 = (inp[7]) ? node265 : 3'b011;
										assign node265 = (inp[5]) ? 3'b001 : 3'b101;
								assign node269 = (inp[7]) ? node271 : 3'b101;
									assign node271 = (inp[5]) ? node275 : node272;
										assign node272 = (inp[8]) ? 3'b110 : 3'b001;
										assign node275 = (inp[8]) ? node277 : 3'b110;
											assign node277 = (inp[2]) ? 3'b010 : 3'b110;
			assign node280 = (inp[3]) ? node378 : node281;
				assign node281 = (inp[10]) ? node331 : node282;
					assign node282 = (inp[8]) ? node308 : node283;
						assign node283 = (inp[2]) ? node295 : node284;
							assign node284 = (inp[7]) ? node288 : node285;
								assign node285 = (inp[11]) ? 3'b110 : 3'b010;
								assign node288 = (inp[0]) ? 3'b100 : node289;
									assign node289 = (inp[1]) ? node291 : 3'b010;
										assign node291 = (inp[11]) ? 3'b001 : 3'b000;
							assign node295 = (inp[0]) ? node303 : node296;
								assign node296 = (inp[1]) ? 3'b010 : node297;
									assign node297 = (inp[11]) ? node299 : 3'b110;
										assign node299 = (inp[4]) ? 3'b110 : 3'b101;
								assign node303 = (inp[11]) ? 3'b110 : node304;
									assign node304 = (inp[5]) ? 3'b010 : 3'b110;
						assign node308 = (inp[7]) ? node322 : node309;
							assign node309 = (inp[4]) ? node319 : node310;
								assign node310 = (inp[11]) ? node316 : node311;
									assign node311 = (inp[2]) ? node313 : 3'b001;
										assign node313 = (inp[0]) ? 3'b110 : 3'b011;
									assign node316 = (inp[0]) ? 3'b001 : 3'b000;
								assign node319 = (inp[0]) ? 3'b010 : 3'b100;
							assign node322 = (inp[11]) ? node326 : node323;
								assign node323 = (inp[4]) ? 3'b000 : 3'b100;
								assign node326 = (inp[1]) ? node328 : 3'b010;
									assign node328 = (inp[4]) ? 3'b100 : 3'b110;
					assign node331 = (inp[11]) ? node353 : node332;
						assign node332 = (inp[5]) ? node348 : node333;
							assign node333 = (inp[2]) ? node339 : node334;
								assign node334 = (inp[7]) ? 3'b110 : node335;
									assign node335 = (inp[0]) ? 3'b001 : 3'b011;
								assign node339 = (inp[7]) ? node343 : node340;
									assign node340 = (inp[0]) ? 3'b111 : 3'b101;
									assign node343 = (inp[4]) ? 3'b001 : node344;
										assign node344 = (inp[8]) ? 3'b001 : 3'b101;
							assign node348 = (inp[0]) ? 3'b001 : node349;
								assign node349 = (inp[1]) ? 3'b001 : 3'b110;
						assign node353 = (inp[5]) ? node367 : node354;
							assign node354 = (inp[8]) ? node362 : node355;
								assign node355 = (inp[4]) ? 3'b101 : node356;
									assign node356 = (inp[0]) ? node358 : 3'b111;
										assign node358 = (inp[7]) ? 3'b011 : 3'b111;
								assign node362 = (inp[4]) ? 3'b011 : node363;
									assign node363 = (inp[1]) ? 3'b111 : 3'b011;
							assign node367 = (inp[4]) ? node373 : node368;
								assign node368 = (inp[7]) ? node370 : 3'b111;
									assign node370 = (inp[1]) ? 3'b001 : 3'b101;
								assign node373 = (inp[7]) ? 3'b110 : node374;
									assign node374 = (inp[1]) ? 3'b001 : 3'b101;
				assign node378 = (inp[10]) ? node400 : node379;
					assign node379 = (inp[4]) ? 3'b000 : node380;
						assign node380 = (inp[7]) ? node390 : node381;
							assign node381 = (inp[1]) ? node385 : node382;
								assign node382 = (inp[11]) ? 3'b010 : 3'b100;
								assign node385 = (inp[11]) ? 3'b100 : node386;
									assign node386 = (inp[2]) ? 3'b000 : 3'b100;
							assign node390 = (inp[8]) ? 3'b000 : node391;
								assign node391 = (inp[5]) ? 3'b000 : node392;
									assign node392 = (inp[0]) ? 3'b000 : node393;
										assign node393 = (inp[11]) ? 3'b100 : 3'b000;
					assign node400 = (inp[7]) ? node418 : node401;
						assign node401 = (inp[8]) ? node415 : node402;
							assign node402 = (inp[5]) ? node408 : node403;
								assign node403 = (inp[11]) ? 3'b110 : node404;
									assign node404 = (inp[4]) ? 3'b010 : 3'b110;
								assign node408 = (inp[4]) ? 3'b100 : node409;
									assign node409 = (inp[11]) ? 3'b001 : node410;
										assign node410 = (inp[0]) ? 3'b010 : 3'b110;
							assign node415 = (inp[4]) ? 3'b100 : 3'b110;
						assign node418 = (inp[4]) ? node436 : node419;
							assign node419 = (inp[0]) ? node425 : node420;
								assign node420 = (inp[5]) ? node422 : 3'b010;
									assign node422 = (inp[2]) ? 3'b010 : 3'b100;
								assign node425 = (inp[11]) ? node431 : node426;
									assign node426 = (inp[5]) ? 3'b000 : node427;
										assign node427 = (inp[8]) ? 3'b000 : 3'b100;
									assign node431 = (inp[5]) ? 3'b100 : node432;
										assign node432 = (inp[1]) ? 3'b010 : 3'b110;
							assign node436 = (inp[0]) ? 3'b100 : node437;
								assign node437 = (inp[8]) ? 3'b000 : node438;
									assign node438 = (inp[11]) ? 3'b100 : 3'b000;

endmodule