module dtc_split66_bm37 (
	input  wire [8-1:0] inp,
	output wire [63-1:0] outp
);

	wire [63-1:0] node1;
	wire [63-1:0] node2;
	wire [63-1:0] node3;
	wire [63-1:0] node4;
	wire [63-1:0] node5;
	wire [63-1:0] node8;
	wire [63-1:0] node11;
	wire [63-1:0] node13;
	wire [63-1:0] node16;
	wire [63-1:0] node17;
	wire [63-1:0] node18;
	wire [63-1:0] node22;
	wire [63-1:0] node23;
	wire [63-1:0] node26;
	wire [63-1:0] node29;
	wire [63-1:0] node30;
	wire [63-1:0] node31;
	wire [63-1:0] node32;
	wire [63-1:0] node36;
	wire [63-1:0] node37;
	wire [63-1:0] node40;
	wire [63-1:0] node43;
	wire [63-1:0] node44;
	wire [63-1:0] node45;
	wire [63-1:0] node48;
	wire [63-1:0] node51;
	wire [63-1:0] node52;
	wire [63-1:0] node55;
	wire [63-1:0] node58;
	wire [63-1:0] node59;
	wire [63-1:0] node60;
	wire [63-1:0] node61;
	wire [63-1:0] node62;
	wire [63-1:0] node65;
	wire [63-1:0] node68;
	wire [63-1:0] node70;
	wire [63-1:0] node73;
	wire [63-1:0] node74;
	wire [63-1:0] node75;
	wire [63-1:0] node78;
	wire [63-1:0] node81;
	wire [63-1:0] node82;
	wire [63-1:0] node85;
	wire [63-1:0] node88;
	wire [63-1:0] node89;
	wire [63-1:0] node90;
	wire [63-1:0] node91;
	wire [63-1:0] node94;
	wire [63-1:0] node97;
	wire [63-1:0] node99;
	wire [63-1:0] node102;
	wire [63-1:0] node103;
	wire [63-1:0] node104;
	wire [63-1:0] node107;
	wire [63-1:0] node110;
	wire [63-1:0] node111;
	wire [63-1:0] node114;

	assign outp = (inp[7]) ? node58 : node1;
		assign node1 = (inp[6]) ? node29 : node2;
			assign node2 = (inp[1]) ? node16 : node3;
				assign node3 = (inp[3]) ? node11 : node4;
					assign node4 = (inp[2]) ? node8 : node5;
						assign node5 = (inp[4]) ? 63'b100111101001100000110001101110110010010101001100001101001010101 : 63'b100111101001100000110001101110110010010101001100001101001010101;
						assign node8 = (inp[0]) ? 63'b100111101001100000110001101110110010010101011100001101001010101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
					assign node11 = (inp[2]) ? node13 : 63'b100110101001100000110001101110110011010101001100000101001010101;
						assign node13 = (inp[4]) ? 63'b100110001001100000110001101110110011010101001100000101001000101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
				assign node16 = (inp[2]) ? node22 : node17;
					assign node17 = (inp[3]) ? 63'b100001101001100000010001101110010010010101001100101101000010101 : node18;
						assign node18 = (inp[4]) ? 63'b100111101001100000010001101110010010010101001100101101000000101 : 63'b100111101001100000010001101110010010010101001100101101000000101;
					assign node22 = (inp[3]) ? node26 : node23;
						assign node23 = (inp[4]) ? 63'b100111101001100000110001101110010010010101001100101101000000101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
						assign node26 = (inp[0]) ? 63'b100001101001100000110001101110010010010101011100101101000010101 : 63'b100001101001100000110001101110110011010101001100101101001010101;
			assign node29 = (inp[3]) ? node43 : node30;
				assign node30 = (inp[2]) ? node36 : node31;
					assign node31 = (inp[1]) ? 63'b100110101001100000110001101110110011010101000100001101001010001 : node32;
						assign node32 = (inp[5]) ? 63'b100110101001100000110001101110110001010101000101101101001010000 : 63'b100110101001100000110001101110110001010101000100101101001010000;
					assign node36 = (inp[0]) ? node40 : node37;
						assign node37 = (inp[5]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100111101001100000111001101110110011010001001100100101001010100;
						assign node40 = (inp[4]) ? 63'b100110101001100000110001101110110001010101010101101101001010000 : 63'b100111101001000000110001101110110011010100001100101101001010101;
				assign node43 = (inp[1]) ? node51 : node44;
					assign node44 = (inp[2]) ? node48 : node45;
						assign node45 = (inp[0]) ? 63'b100110101001100000110001101110110011010001001101001101001010101 : 63'b100110101001100000110001101110110011010001001100001101001010101;
						assign node48 = (inp[4]) ? 63'b100111101001100000110001101110110011010001001100101101001010101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
					assign node51 = (inp[2]) ? node55 : node52;
						assign node52 = (inp[5]) ? 63'b100110101001100000110001101110100011010101001100100101001010100 : 63'b100110101001100000110001101110100011010101001100100101001010100;
						assign node55 = (inp[0]) ? 63'b100110101001100000110001101110100011010101001100100101001010100 : 63'b100111101001100000110001101110110011010101001100001101001010101;
		assign node58 = (inp[2]) ? node88 : node59;
			assign node59 = (inp[3]) ? node73 : node60;
				assign node60 = (inp[1]) ? node68 : node61;
					assign node61 = (inp[6]) ? node65 : node62;
						assign node62 = (inp[5]) ? 63'b100111101001100000110001101110110011010101001000101101001000101 : 63'b100111101001100000110001101110110011010101001000101101001000101;
						assign node65 = (inp[4]) ? 63'b100111101001000000110001101000110111010101001100101100001010101 : 63'b100111101000000000110001100000110011010101001100101100001010101;
					assign node68 = (inp[6]) ? node70 : 63'b100111101001100000110001101110110011010101001100101101000010101;
						assign node70 = (inp[0]) ? 63'b100111101001100000110001001110110011010101001100101101000010101 : 63'b100111101001100000110001001110110011010101001100101101000010101;
				assign node73 = (inp[6]) ? node81 : node74;
					assign node74 = (inp[4]) ? node78 : node75;
						assign node75 = (inp[1]) ? 63'b100111101000000000110001100000110011010101001100101100001010101 : 63'b100001101000000000110001100000110011010101001100101100001010101;
						assign node78 = (inp[0]) ? 63'b000111101001001000110001101010110011000101001101101101001010101 : 63'b000111101001001000110001101010110011000101001100101101001010101;
					assign node81 = (inp[1]) ? node85 : node82;
						assign node82 = (inp[4]) ? 63'b100111101001100000100001101110110010010101001100101101000010101 : 63'b100111101011100000100001101110110010010101001100101101000010101;
						assign node85 = (inp[4]) ? 63'b100111101001000000110000100100110011010101101100101101001010101 : 63'b100111101000000000110000100100110011010101101100101101001010101;
			assign node88 = (inp[4]) ? node102 : node89;
				assign node89 = (inp[5]) ? node97 : node90;
					assign node90 = (inp[3]) ? node94 : node91;
						assign node91 = (inp[6]) ? 63'b100111101001100000010001101110110011010101001100000101001010101 : 63'b100111101001100000110001101110110011010101001100101101001010101;
						assign node94 = (inp[6]) ? 63'b100111101001100000110001101110110011010101001100101101001010101 : 63'b100001101001100000110001101110110011010101001100101101001010101;
					assign node97 = (inp[0]) ? node99 : 63'b100111101001100100110001101110110011010101001100101101001010101;
						assign node99 = (inp[1]) ? 63'b100111101001000000110001101110110011010100001100101101001110101 : 63'b100001101001000000110001101110110011000110001100101001001010101;
				assign node102 = (inp[0]) ? node110 : node103;
					assign node103 = (inp[5]) ? node107 : node104;
						assign node104 = (inp[6]) ? 63'b100111001001100000110001101110110001010101000100101101001000001 : 63'b100111100001000000110001101110110011000100001100101001001010101;
						assign node107 = (inp[1]) ? 63'b000111101001000000110001101000110011000101001100101100001010101 : 63'b100101101001110000110001101110110011010101001100101101001010101;
					assign node110 = (inp[6]) ? node114 : node111;
						assign node111 = (inp[3]) ? 63'b100111101000000000110001101001110011010101011101101100001010101 : 63'b100111101001100000110001101110110011010101011000101101000000101;
						assign node114 = (inp[1]) ? 63'b100111101001100000110001001110110011010101011100101101000010101 : 63'b100111101001100000100001101110110010010101011100101101000010101;

endmodule