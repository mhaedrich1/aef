module dtc_split33_bm80 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node389;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node401;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node415;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node423;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node472;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node549;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node557;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node563;
	wire [3-1:0] node566;
	wire [3-1:0] node567;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node583;
	wire [3-1:0] node585;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node608;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node635;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node672;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node720;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node749;
	wire [3-1:0] node752;
	wire [3-1:0] node753;
	wire [3-1:0] node756;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node767;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node773;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node781;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node788;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node803;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node807;
	wire [3-1:0] node810;
	wire [3-1:0] node813;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node825;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node833;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node850;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node857;
	wire [3-1:0] node860;
	wire [3-1:0] node864;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node879;
	wire [3-1:0] node881;
	wire [3-1:0] node884;
	wire [3-1:0] node886;
	wire [3-1:0] node887;
	wire [3-1:0] node890;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node905;
	wire [3-1:0] node907;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node916;
	wire [3-1:0] node917;
	wire [3-1:0] node918;
	wire [3-1:0] node923;
	wire [3-1:0] node925;
	wire [3-1:0] node928;
	wire [3-1:0] node930;
	wire [3-1:0] node932;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node951;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node968;
	wire [3-1:0] node971;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node977;
	wire [3-1:0] node981;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node997;
	wire [3-1:0] node999;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1013;
	wire [3-1:0] node1014;
	wire [3-1:0] node1015;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1027;
	wire [3-1:0] node1028;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1034;
	wire [3-1:0] node1037;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1045;
	wire [3-1:0] node1046;
	wire [3-1:0] node1049;
	wire [3-1:0] node1051;
	wire [3-1:0] node1054;
	wire [3-1:0] node1056;
	wire [3-1:0] node1058;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1066;
	wire [3-1:0] node1067;
	wire [3-1:0] node1071;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1083;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1090;
	wire [3-1:0] node1093;
	wire [3-1:0] node1094;
	wire [3-1:0] node1095;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1101;
	wire [3-1:0] node1103;
	wire [3-1:0] node1106;
	wire [3-1:0] node1108;
	wire [3-1:0] node1109;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1117;
	wire [3-1:0] node1121;
	wire [3-1:0] node1123;
	wire [3-1:0] node1124;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1134;
	wire [3-1:0] node1135;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1143;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1149;
	wire [3-1:0] node1150;
	wire [3-1:0] node1153;
	wire [3-1:0] node1158;
	wire [3-1:0] node1159;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1165;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1175;
	wire [3-1:0] node1178;
	wire [3-1:0] node1180;
	wire [3-1:0] node1183;
	wire [3-1:0] node1184;
	wire [3-1:0] node1185;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1190;
	wire [3-1:0] node1193;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1198;
	wire [3-1:0] node1200;
	wire [3-1:0] node1203;
	wire [3-1:0] node1205;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1214;
	wire [3-1:0] node1219;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1226;
	wire [3-1:0] node1229;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1234;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1238;
	wire [3-1:0] node1242;
	wire [3-1:0] node1244;
	wire [3-1:0] node1247;
	wire [3-1:0] node1249;
	wire [3-1:0] node1250;
	wire [3-1:0] node1253;
	wire [3-1:0] node1256;
	wire [3-1:0] node1258;
	wire [3-1:0] node1259;
	wire [3-1:0] node1262;
	wire [3-1:0] node1265;
	wire [3-1:0] node1266;
	wire [3-1:0] node1267;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1283;
	wire [3-1:0] node1284;
	wire [3-1:0] node1287;
	wire [3-1:0] node1290;
	wire [3-1:0] node1292;
	wire [3-1:0] node1293;
	wire [3-1:0] node1294;
	wire [3-1:0] node1298;
	wire [3-1:0] node1299;
	wire [3-1:0] node1300;
	wire [3-1:0] node1301;
	wire [3-1:0] node1304;
	wire [3-1:0] node1308;

	assign outp = (inp[6]) ? node526 : node1;
		assign node1 = (inp[3]) ? node393 : node2;
			assign node2 = (inp[9]) ? node240 : node3;
				assign node3 = (inp[4]) ? node121 : node4;
					assign node4 = (inp[7]) ? node62 : node5;
						assign node5 = (inp[0]) ? node33 : node6;
							assign node6 = (inp[2]) ? node12 : node7;
								assign node7 = (inp[8]) ? node9 : 3'b101;
									assign node9 = (inp[11]) ? 3'b001 : 3'b101;
								assign node12 = (inp[1]) ? node22 : node13;
									assign node13 = (inp[10]) ? node19 : node14;
										assign node14 = (inp[11]) ? 3'b101 : node15;
											assign node15 = (inp[5]) ? 3'b001 : 3'b011;
										assign node19 = (inp[8]) ? 3'b000 : 3'b001;
									assign node22 = (inp[5]) ? node26 : node23;
										assign node23 = (inp[8]) ? 3'b001 : 3'b110;
										assign node26 = (inp[11]) ? node30 : node27;
											assign node27 = (inp[8]) ? 3'b110 : 3'b001;
											assign node30 = (inp[10]) ? 3'b010 : 3'b110;
							assign node33 = (inp[2]) ? node49 : node34;
								assign node34 = (inp[11]) ? node46 : node35;
									assign node35 = (inp[8]) ? node41 : node36;
										assign node36 = (inp[5]) ? 3'b010 : node37;
											assign node37 = (inp[1]) ? 3'b010 : 3'b110;
										assign node41 = (inp[1]) ? 3'b110 : node42;
											assign node42 = (inp[5]) ? 3'b110 : 3'b010;
									assign node46 = (inp[10]) ? 3'b010 : 3'b000;
								assign node49 = (inp[1]) ? node59 : node50;
									assign node50 = (inp[8]) ? node56 : node51;
										assign node51 = (inp[5]) ? node53 : 3'b110;
											assign node53 = (inp[11]) ? 3'b010 : 3'b010;
										assign node56 = (inp[10]) ? 3'b110 : 3'b001;
									assign node59 = (inp[8]) ? 3'b110 : 3'b100;
						assign node62 = (inp[1]) ? node92 : node63;
							assign node63 = (inp[0]) ? node81 : node64;
								assign node64 = (inp[2]) ? node74 : node65;
									assign node65 = (inp[11]) ? 3'b001 : node66;
										assign node66 = (inp[5]) ? node70 : node67;
											assign node67 = (inp[10]) ? 3'b001 : 3'b000;
											assign node70 = (inp[8]) ? 3'b001 : 3'b000;
									assign node74 = (inp[8]) ? 3'b001 : node75;
										assign node75 = (inp[5]) ? node77 : 3'b001;
											assign node77 = (inp[10]) ? 3'b000 : 3'b001;
								assign node81 = (inp[5]) ? node85 : node82;
									assign node82 = (inp[8]) ? 3'b010 : 3'b001;
									assign node85 = (inp[8]) ? node89 : node86;
										assign node86 = (inp[10]) ? 3'b110 : 3'b001;
										assign node89 = (inp[10]) ? 3'b001 : 3'b101;
							assign node92 = (inp[2]) ? node106 : node93;
								assign node93 = (inp[10]) ? node99 : node94;
									assign node94 = (inp[11]) ? node96 : 3'b111;
										assign node96 = (inp[0]) ? 3'b101 : 3'b001;
									assign node99 = (inp[8]) ? 3'b001 : node100;
										assign node100 = (inp[0]) ? 3'b110 : node101;
											assign node101 = (inp[11]) ? 3'b001 : 3'b101;
								assign node106 = (inp[0]) ? node114 : node107;
									assign node107 = (inp[10]) ? 3'b001 : node108;
										assign node108 = (inp[5]) ? 3'b011 : node109;
											assign node109 = (inp[8]) ? 3'b111 : 3'b011;
									assign node114 = (inp[11]) ? 3'b001 : node115;
										assign node115 = (inp[10]) ? 3'b001 : node116;
											assign node116 = (inp[8]) ? 3'b101 : 3'b001;
					assign node121 = (inp[0]) ? node177 : node122;
						assign node122 = (inp[7]) ? node150 : node123;
							assign node123 = (inp[2]) ? node133 : node124;
								assign node124 = (inp[1]) ? 3'b110 : node125;
									assign node125 = (inp[8]) ? node129 : node126;
										assign node126 = (inp[11]) ? 3'b010 : 3'b100;
										assign node129 = (inp[10]) ? 3'b110 : 3'b100;
								assign node133 = (inp[1]) ? node139 : node134;
									assign node134 = (inp[11]) ? node136 : 3'b000;
										assign node136 = (inp[10]) ? 3'b110 : 3'b000;
									assign node139 = (inp[11]) ? node145 : node140;
										assign node140 = (inp[8]) ? node142 : 3'b010;
											assign node142 = (inp[10]) ? 3'b110 : 3'b000;
										assign node145 = (inp[8]) ? 3'b010 : node146;
											assign node146 = (inp[10]) ? 3'b000 : 3'b010;
							assign node150 = (inp[2]) ? node164 : node151;
								assign node151 = (inp[1]) ? node157 : node152;
									assign node152 = (inp[5]) ? node154 : 3'b111;
										assign node154 = (inp[8]) ? 3'b011 : 3'b001;
									assign node157 = (inp[5]) ? 3'b110 : node158;
										assign node158 = (inp[8]) ? 3'b001 : node159;
											assign node159 = (inp[10]) ? 3'b110 : 3'b101;
								assign node164 = (inp[10]) ? node170 : node165;
									assign node165 = (inp[1]) ? node167 : 3'b101;
										assign node167 = (inp[11]) ? 3'b101 : 3'b001;
									assign node170 = (inp[5]) ? node174 : node171;
										assign node171 = (inp[11]) ? 3'b001 : 3'b101;
										assign node174 = (inp[1]) ? 3'b110 : 3'b000;
						assign node177 = (inp[7]) ? node205 : node178;
							assign node178 = (inp[1]) ? node194 : node179;
								assign node179 = (inp[10]) ? node189 : node180;
									assign node180 = (inp[5]) ? node186 : node181;
										assign node181 = (inp[2]) ? 3'b010 : node182;
											assign node182 = (inp[8]) ? 3'b110 : 3'b010;
										assign node186 = (inp[8]) ? 3'b010 : 3'b100;
									assign node189 = (inp[8]) ? 3'b100 : node190;
										assign node190 = (inp[5]) ? 3'b000 : 3'b100;
								assign node194 = (inp[8]) ? node200 : node195;
									assign node195 = (inp[10]) ? 3'b000 : node196;
										assign node196 = (inp[5]) ? 3'b000 : 3'b100;
									assign node200 = (inp[10]) ? 3'b100 : node201;
										assign node201 = (inp[11]) ? 3'b100 : 3'b000;
							assign node205 = (inp[8]) ? node223 : node206;
								assign node206 = (inp[2]) ? node216 : node207;
									assign node207 = (inp[10]) ? node211 : node208;
										assign node208 = (inp[11]) ? 3'b100 : 3'b001;
										assign node211 = (inp[1]) ? 3'b010 : node212;
											assign node212 = (inp[11]) ? 3'b000 : 3'b010;
									assign node216 = (inp[11]) ? node220 : node217;
										assign node217 = (inp[1]) ? 3'b010 : 3'b110;
										assign node220 = (inp[1]) ? 3'b100 : 3'b110;
								assign node223 = (inp[2]) ? node229 : node224;
									assign node224 = (inp[1]) ? node226 : 3'b010;
										assign node226 = (inp[5]) ? 3'b100 : 3'b110;
									assign node229 = (inp[1]) ? node235 : node230;
										assign node230 = (inp[11]) ? node232 : 3'b110;
											assign node232 = (inp[5]) ? 3'b010 : 3'b110;
										assign node235 = (inp[10]) ? 3'b010 : node236;
											assign node236 = (inp[5]) ? 3'b010 : 3'b110;
				assign node240 = (inp[7]) ? node280 : node241;
					assign node241 = (inp[4]) ? node271 : node242;
						assign node242 = (inp[10]) ? node256 : node243;
							assign node243 = (inp[11]) ? node251 : node244;
								assign node244 = (inp[0]) ? node246 : 3'b010;
									assign node246 = (inp[1]) ? 3'b100 : node247;
										assign node247 = (inp[8]) ? 3'b010 : 3'b100;
								assign node251 = (inp[2]) ? node253 : 3'b000;
									assign node253 = (inp[8]) ? 3'b100 : 3'b000;
							assign node256 = (inp[0]) ? node266 : node257;
								assign node257 = (inp[8]) ? node263 : node258;
									assign node258 = (inp[5]) ? node260 : 3'b100;
										assign node260 = (inp[1]) ? 3'b100 : 3'b000;
									assign node263 = (inp[2]) ? 3'b100 : 3'b010;
								assign node266 = (inp[1]) ? 3'b000 : node267;
									assign node267 = (inp[2]) ? 3'b000 : 3'b100;
						assign node271 = (inp[0]) ? 3'b000 : node272;
							assign node272 = (inp[1]) ? 3'b000 : node273;
								assign node273 = (inp[5]) ? node275 : 3'b010;
									assign node275 = (inp[10]) ? 3'b000 : 3'b010;
					assign node280 = (inp[4]) ? node342 : node281;
						assign node281 = (inp[1]) ? node313 : node282;
							assign node282 = (inp[0]) ? node298 : node283;
								assign node283 = (inp[5]) ? node291 : node284;
									assign node284 = (inp[2]) ? 3'b101 : node285;
										assign node285 = (inp[10]) ? node287 : 3'b001;
											assign node287 = (inp[8]) ? 3'b001 : 3'b000;
									assign node291 = (inp[10]) ? 3'b100 : node292;
										assign node292 = (inp[8]) ? node294 : 3'b000;
											assign node294 = (inp[11]) ? 3'b000 : 3'b101;
								assign node298 = (inp[10]) ? node302 : node299;
									assign node299 = (inp[8]) ? 3'b000 : 3'b010;
									assign node302 = (inp[11]) ? node308 : node303;
										assign node303 = (inp[2]) ? 3'b010 : node304;
											assign node304 = (inp[8]) ? 3'b010 : 3'b000;
										assign node308 = (inp[2]) ? 3'b010 : node309;
											assign node309 = (inp[8]) ? 3'b110 : 3'b010;
							assign node313 = (inp[10]) ? node327 : node314;
								assign node314 = (inp[2]) ? node324 : node315;
									assign node315 = (inp[0]) ? node319 : node316;
										assign node316 = (inp[8]) ? 3'b101 : 3'b010;
										assign node319 = (inp[5]) ? node321 : 3'b110;
											assign node321 = (inp[8]) ? 3'b010 : 3'b100;
									assign node324 = (inp[0]) ? 3'b010 : 3'b110;
								assign node327 = (inp[0]) ? node335 : node328;
									assign node328 = (inp[5]) ? node330 : 3'b110;
										assign node330 = (inp[8]) ? 3'b110 : node331;
											assign node331 = (inp[11]) ? 3'b010 : 3'b001;
									assign node335 = (inp[11]) ? 3'b100 : node336;
										assign node336 = (inp[8]) ? 3'b010 : node337;
											assign node337 = (inp[2]) ? 3'b000 : 3'b100;
						assign node342 = (inp[10]) ? node370 : node343;
							assign node343 = (inp[11]) ? node361 : node344;
								assign node344 = (inp[1]) ? node352 : node345;
									assign node345 = (inp[5]) ? node349 : node346;
										assign node346 = (inp[8]) ? 3'b110 : 3'b010;
										assign node349 = (inp[8]) ? 3'b010 : 3'b100;
									assign node352 = (inp[0]) ? node358 : node353;
										assign node353 = (inp[5]) ? node355 : 3'b001;
											assign node355 = (inp[8]) ? 3'b110 : 3'b010;
										assign node358 = (inp[5]) ? 3'b000 : 3'b100;
								assign node361 = (inp[1]) ? node363 : 3'b100;
									assign node363 = (inp[0]) ? 3'b000 : node364;
										assign node364 = (inp[2]) ? 3'b100 : node365;
											assign node365 = (inp[5]) ? 3'b010 : 3'b110;
							assign node370 = (inp[0]) ? node384 : node371;
								assign node371 = (inp[1]) ? node379 : node372;
									assign node372 = (inp[8]) ? node374 : 3'b000;
										assign node374 = (inp[5]) ? node376 : 3'b100;
											assign node376 = (inp[11]) ? 3'b000 : 3'b100;
									assign node379 = (inp[8]) ? node381 : 3'b100;
										assign node381 = (inp[11]) ? 3'b100 : 3'b010;
								assign node384 = (inp[1]) ? 3'b000 : node385;
									assign node385 = (inp[8]) ? node389 : node386;
										assign node386 = (inp[5]) ? 3'b000 : 3'b100;
										assign node389 = (inp[5]) ? 3'b100 : 3'b000;
			assign node393 = (inp[9]) ? node507 : node394;
				assign node394 = (inp[4]) ? node472 : node395;
					assign node395 = (inp[7]) ? node427 : node396;
						assign node396 = (inp[11]) ? node420 : node397;
							assign node397 = (inp[10]) ? node411 : node398;
								assign node398 = (inp[1]) ? node404 : node399;
									assign node399 = (inp[5]) ? node401 : 3'b100;
										assign node401 = (inp[8]) ? 3'b100 : 3'b000;
									assign node404 = (inp[0]) ? 3'b000 : node405;
										assign node405 = (inp[8]) ? node407 : 3'b100;
											assign node407 = (inp[5]) ? 3'b010 : 3'b110;
								assign node411 = (inp[0]) ? 3'b000 : node412;
									assign node412 = (inp[2]) ? 3'b100 : node413;
										assign node413 = (inp[5]) ? node415 : 3'b000;
											assign node415 = (inp[8]) ? 3'b000 : 3'b000;
							assign node420 = (inp[0]) ? 3'b000 : node421;
								assign node421 = (inp[2]) ? node423 : 3'b000;
									assign node423 = (inp[8]) ? 3'b100 : 3'b000;
						assign node427 = (inp[0]) ? node453 : node428;
							assign node428 = (inp[5]) ? node434 : node429;
								assign node429 = (inp[8]) ? node431 : 3'b010;
									assign node431 = (inp[11]) ? 3'b000 : 3'b001;
								assign node434 = (inp[10]) ? node442 : node435;
									assign node435 = (inp[1]) ? node439 : node436;
										assign node436 = (inp[8]) ? 3'b000 : 3'b110;
										assign node439 = (inp[8]) ? 3'b110 : 3'b010;
									assign node442 = (inp[2]) ? node450 : node443;
										assign node443 = (inp[1]) ? node447 : node444;
											assign node444 = (inp[8]) ? 3'b110 : 3'b010;
											assign node447 = (inp[8]) ? 3'b010 : 3'b100;
										assign node450 = (inp[11]) ? 3'b100 : 3'b000;
							assign node453 = (inp[5]) ? node465 : node454;
								assign node454 = (inp[11]) ? node456 : 3'b010;
									assign node456 = (inp[1]) ? node462 : node457;
										assign node457 = (inp[10]) ? 3'b100 : node458;
											assign node458 = (inp[8]) ? 3'b010 : 3'b010;
										assign node462 = (inp[10]) ? 3'b000 : 3'b100;
								assign node465 = (inp[8]) ? 3'b100 : node466;
									assign node466 = (inp[1]) ? 3'b000 : node467;
										assign node467 = (inp[11]) ? 3'b000 : 3'b100;
					assign node472 = (inp[7]) ? node474 : 3'b000;
						assign node474 = (inp[10]) ? node498 : node475;
							assign node475 = (inp[5]) ? node487 : node476;
								assign node476 = (inp[11]) ? node480 : node477;
									assign node477 = (inp[1]) ? 3'b110 : 3'b100;
									assign node480 = (inp[2]) ? node482 : 3'b000;
										assign node482 = (inp[0]) ? node484 : 3'b100;
											assign node484 = (inp[8]) ? 3'b100 : 3'b000;
								assign node487 = (inp[1]) ? node489 : 3'b000;
									assign node489 = (inp[0]) ? 3'b000 : node490;
										assign node490 = (inp[8]) ? node494 : node491;
											assign node491 = (inp[11]) ? 3'b000 : 3'b100;
											assign node494 = (inp[11]) ? 3'b100 : 3'b010;
							assign node498 = (inp[5]) ? 3'b000 : node499;
								assign node499 = (inp[8]) ? 3'b000 : node500;
									assign node500 = (inp[11]) ? 3'b000 : node501;
										assign node501 = (inp[0]) ? 3'b000 : 3'b100;
				assign node507 = (inp[4]) ? 3'b000 : node508;
					assign node508 = (inp[7]) ? node510 : 3'b000;
						assign node510 = (inp[0]) ? 3'b000 : node511;
							assign node511 = (inp[1]) ? node517 : node512;
								assign node512 = (inp[5]) ? node514 : 3'b010;
									assign node514 = (inp[10]) ? 3'b000 : 3'b010;
								assign node517 = (inp[5]) ? 3'b000 : node518;
									assign node518 = (inp[10]) ? 3'b000 : node519;
										assign node519 = (inp[11]) ? 3'b100 : 3'b000;
		assign node526 = (inp[3]) ? node910 : node527;
			assign node527 = (inp[9]) ? node693 : node528;
				assign node528 = (inp[0]) ? node588 : node529;
					assign node529 = (inp[1]) ? node541 : node530;
						assign node530 = (inp[4]) ? node532 : 3'b111;
							assign node532 = (inp[7]) ? 3'b111 : node533;
								assign node533 = (inp[10]) ? node535 : 3'b111;
									assign node535 = (inp[2]) ? node537 : 3'b011;
										assign node537 = (inp[5]) ? 3'b111 : 3'b011;
						assign node541 = (inp[7]) ? node571 : node542;
							assign node542 = (inp[4]) ? node554 : node543;
								assign node543 = (inp[10]) ? node547 : node544;
									assign node544 = (inp[2]) ? 3'b111 : 3'b011;
									assign node547 = (inp[2]) ? 3'b011 : node548;
										assign node548 = (inp[8]) ? 3'b111 : node549;
											assign node549 = (inp[5]) ? 3'b010 : 3'b011;
								assign node554 = (inp[8]) ? node560 : node555;
									assign node555 = (inp[11]) ? node557 : 3'b101;
										assign node557 = (inp[10]) ? 3'b001 : 3'b101;
									assign node560 = (inp[11]) ? node566 : node561;
										assign node561 = (inp[5]) ? node563 : 3'b011;
											assign node563 = (inp[10]) ? 3'b101 : 3'b011;
										assign node566 = (inp[2]) ? 3'b101 : node567;
											assign node567 = (inp[10]) ? 3'b101 : 3'b011;
							assign node571 = (inp[4]) ? node573 : 3'b111;
								assign node573 = (inp[8]) ? node583 : node574;
									assign node574 = (inp[11]) ? node578 : node575;
										assign node575 = (inp[10]) ? 3'b011 : 3'b111;
										assign node578 = (inp[10]) ? 3'b101 : node579;
											assign node579 = (inp[5]) ? 3'b011 : 3'b101;
									assign node583 = (inp[10]) ? node585 : 3'b111;
										assign node585 = (inp[2]) ? 3'b111 : 3'b011;
					assign node588 = (inp[4]) ? node638 : node589;
						assign node589 = (inp[7]) ? node627 : node590;
							assign node590 = (inp[1]) ? node616 : node591;
								assign node591 = (inp[5]) ? node605 : node592;
									assign node592 = (inp[2]) ? node598 : node593;
										assign node593 = (inp[8]) ? 3'b111 : node594;
											assign node594 = (inp[10]) ? 3'b111 : 3'b011;
										assign node598 = (inp[10]) ? node602 : node599;
											assign node599 = (inp[8]) ? 3'b111 : 3'b011;
											assign node602 = (inp[8]) ? 3'b011 : 3'b111;
									assign node605 = (inp[11]) ? node611 : node606;
										assign node606 = (inp[8]) ? node608 : 3'b011;
											assign node608 = (inp[2]) ? 3'b011 : 3'b011;
										assign node611 = (inp[8]) ? 3'b011 : node612;
											assign node612 = (inp[10]) ? 3'b001 : 3'b101;
								assign node616 = (inp[8]) ? node622 : node617;
									assign node617 = (inp[5]) ? 3'b101 : node618;
										assign node618 = (inp[11]) ? 3'b001 : 3'b101;
									assign node622 = (inp[11]) ? 3'b001 : node623;
										assign node623 = (inp[2]) ? 3'b011 : 3'b111;
							assign node627 = (inp[11]) ? node633 : node628;
								assign node628 = (inp[1]) ? node630 : 3'b111;
									assign node630 = (inp[5]) ? 3'b101 : 3'b111;
								assign node633 = (inp[8]) ? node635 : 3'b011;
									assign node635 = (inp[2]) ? 3'b011 : 3'b111;
						assign node638 = (inp[1]) ? node668 : node639;
							assign node639 = (inp[5]) ? node655 : node640;
								assign node640 = (inp[2]) ? node648 : node641;
									assign node641 = (inp[8]) ? node645 : node642;
										assign node642 = (inp[11]) ? 3'b111 : 3'b011;
										assign node645 = (inp[11]) ? 3'b011 : 3'b111;
									assign node648 = (inp[11]) ? 3'b110 : node649;
										assign node649 = (inp[7]) ? 3'b111 : node650;
											assign node650 = (inp[8]) ? 3'b101 : 3'b001;
								assign node655 = (inp[11]) ? node661 : node656;
									assign node656 = (inp[2]) ? 3'b101 : node657;
										assign node657 = (inp[7]) ? 3'b011 : 3'b001;
									assign node661 = (inp[7]) ? 3'b101 : node662;
										assign node662 = (inp[10]) ? 3'b110 : node663;
											assign node663 = (inp[2]) ? 3'b001 : 3'b101;
							assign node668 = (inp[11]) ? node676 : node669;
								assign node669 = (inp[5]) ? 3'b001 : node670;
									assign node670 = (inp[10]) ? node672 : 3'b011;
										assign node672 = (inp[7]) ? 3'b101 : 3'b001;
								assign node676 = (inp[10]) ? node684 : node677;
									assign node677 = (inp[2]) ? 3'b001 : node678;
										assign node678 = (inp[8]) ? 3'b010 : node679;
											assign node679 = (inp[5]) ? 3'b000 : 3'b001;
									assign node684 = (inp[2]) ? node688 : node685;
										assign node685 = (inp[8]) ? 3'b001 : 3'b010;
										assign node688 = (inp[7]) ? 3'b110 : node689;
											assign node689 = (inp[8]) ? 3'b110 : 3'b010;
				assign node693 = (inp[0]) ? node781 : node694;
					assign node694 = (inp[4]) ? node730 : node695;
						assign node695 = (inp[7]) ? node717 : node696;
							assign node696 = (inp[1]) ? node706 : node697;
								assign node697 = (inp[8]) ? node699 : 3'b011;
									assign node699 = (inp[5]) ? node703 : node700;
										assign node700 = (inp[10]) ? 3'b011 : 3'b111;
										assign node703 = (inp[11]) ? 3'b101 : 3'b111;
								assign node706 = (inp[5]) ? node710 : node707;
									assign node707 = (inp[8]) ? 3'b011 : 3'b001;
									assign node710 = (inp[2]) ? node714 : node711;
										assign node711 = (inp[11]) ? 3'b101 : 3'b011;
										assign node714 = (inp[11]) ? 3'b001 : 3'b101;
							assign node717 = (inp[11]) ? node723 : node718;
								assign node718 = (inp[10]) ? node720 : 3'b111;
									assign node720 = (inp[8]) ? 3'b111 : 3'b101;
								assign node723 = (inp[8]) ? node725 : 3'b011;
									assign node725 = (inp[5]) ? 3'b111 : node726;
										assign node726 = (inp[1]) ? 3'b011 : 3'b111;
						assign node730 = (inp[7]) ? node744 : node731;
							assign node731 = (inp[1]) ? node739 : node732;
								assign node732 = (inp[11]) ? node736 : node733;
									assign node733 = (inp[10]) ? 3'b110 : 3'b001;
									assign node736 = (inp[10]) ? 3'b001 : 3'b101;
								assign node739 = (inp[2]) ? 3'b110 : node740;
									assign node740 = (inp[10]) ? 3'b110 : 3'b001;
							assign node744 = (inp[1]) ? node764 : node745;
								assign node745 = (inp[8]) ? node759 : node746;
									assign node746 = (inp[2]) ? node752 : node747;
										assign node747 = (inp[10]) ? node749 : 3'b011;
											assign node749 = (inp[11]) ? 3'b001 : 3'b101;
										assign node752 = (inp[5]) ? node756 : node753;
											assign node753 = (inp[10]) ? 3'b101 : 3'b011;
											assign node756 = (inp[10]) ? 3'b111 : 3'b101;
									assign node759 = (inp[10]) ? 3'b111 : node760;
										assign node760 = (inp[2]) ? 3'b011 : 3'b111;
								assign node764 = (inp[11]) ? node770 : node765;
									assign node765 = (inp[5]) ? node767 : 3'b101;
										assign node767 = (inp[2]) ? 3'b001 : 3'b101;
									assign node770 = (inp[2]) ? node776 : node771;
										assign node771 = (inp[8]) ? node773 : 3'b001;
											assign node773 = (inp[10]) ? 3'b001 : 3'b101;
										assign node776 = (inp[5]) ? 3'b110 : node777;
											assign node777 = (inp[8]) ? 3'b101 : 3'b001;
					assign node781 = (inp[4]) ? node841 : node782;
						assign node782 = (inp[1]) ? node820 : node783;
							assign node783 = (inp[7]) ? node803 : node784;
								assign node784 = (inp[8]) ? node792 : node785;
									assign node785 = (inp[10]) ? 3'b110 : node786;
										assign node786 = (inp[11]) ? node788 : 3'b001;
											assign node788 = (inp[5]) ? 3'b110 : 3'b001;
									assign node792 = (inp[11]) ? node798 : node793;
										assign node793 = (inp[2]) ? node795 : 3'b101;
											assign node795 = (inp[5]) ? 3'b001 : 3'b101;
										assign node798 = (inp[10]) ? 3'b001 : node799;
											assign node799 = (inp[5]) ? 3'b001 : 3'b101;
								assign node803 = (inp[10]) ? node813 : node804;
									assign node804 = (inp[5]) ? node810 : node805;
										assign node805 = (inp[2]) ? node807 : 3'b111;
											assign node807 = (inp[11]) ? 3'b011 : 3'b011;
										assign node810 = (inp[8]) ? 3'b011 : 3'b101;
									assign node813 = (inp[2]) ? node815 : 3'b011;
										assign node815 = (inp[11]) ? node817 : 3'b101;
											assign node817 = (inp[5]) ? 3'b001 : 3'b101;
							assign node820 = (inp[7]) ? node830 : node821;
								assign node821 = (inp[5]) ? 3'b010 : node822;
									assign node822 = (inp[2]) ? 3'b001 : node823;
										assign node823 = (inp[11]) ? node825 : 3'b001;
											assign node825 = (inp[8]) ? 3'b000 : 3'b010;
								assign node830 = (inp[2]) ? node836 : node831;
									assign node831 = (inp[10]) ? node833 : 3'b001;
										assign node833 = (inp[5]) ? 3'b001 : 3'b101;
									assign node836 = (inp[8]) ? 3'b001 : node837;
										assign node837 = (inp[5]) ? 3'b110 : 3'b001;
						assign node841 = (inp[10]) ? node871 : node842;
							assign node842 = (inp[7]) ? node854 : node843;
								assign node843 = (inp[8]) ? node847 : node844;
									assign node844 = (inp[5]) ? 3'b100 : 3'b010;
									assign node847 = (inp[1]) ? 3'b010 : node848;
										assign node848 = (inp[11]) ? node850 : 3'b110;
											assign node850 = (inp[2]) ? 3'b010 : 3'b110;
								assign node854 = (inp[1]) ? node864 : node855;
									assign node855 = (inp[2]) ? 3'b001 : node856;
										assign node856 = (inp[11]) ? node860 : node857;
											assign node857 = (inp[8]) ? 3'b101 : 3'b001;
											assign node860 = (inp[5]) ? 3'b001 : 3'b101;
									assign node864 = (inp[5]) ? node866 : 3'b001;
										assign node866 = (inp[2]) ? 3'b110 : node867;
											assign node867 = (inp[8]) ? 3'b010 : 3'b110;
							assign node871 = (inp[8]) ? node893 : node872;
								assign node872 = (inp[7]) ? node884 : node873;
									assign node873 = (inp[11]) ? node879 : node874;
										assign node874 = (inp[1]) ? 3'b100 : node875;
											assign node875 = (inp[5]) ? 3'b000 : 3'b010;
										assign node879 = (inp[5]) ? node881 : 3'b100;
											assign node881 = (inp[1]) ? 3'b000 : 3'b100;
									assign node884 = (inp[5]) ? node886 : 3'b110;
										assign node886 = (inp[11]) ? node890 : node887;
											assign node887 = (inp[1]) ? 3'b010 : 3'b110;
											assign node890 = (inp[2]) ? 3'b100 : 3'b000;
								assign node893 = (inp[2]) ? node903 : node894;
									assign node894 = (inp[7]) ? node900 : node895;
										assign node895 = (inp[1]) ? 3'b100 : node896;
											assign node896 = (inp[5]) ? 3'b010 : 3'b110;
										assign node900 = (inp[1]) ? 3'b010 : 3'b001;
									assign node903 = (inp[7]) ? node905 : 3'b010;
										assign node905 = (inp[1]) ? node907 : 3'b110;
											assign node907 = (inp[11]) ? 3'b010 : 3'b110;
			assign node910 = (inp[9]) ? node1128 : node911;
				assign node911 = (inp[7]) ? node1013 : node912;
					assign node912 = (inp[4]) ? node958 : node913;
						assign node913 = (inp[10]) ? node935 : node914;
							assign node914 = (inp[5]) ? node928 : node915;
								assign node915 = (inp[1]) ? node923 : node916;
									assign node916 = (inp[0]) ? 3'b001 : node917;
										assign node917 = (inp[11]) ? 3'b101 : node918;
											assign node918 = (inp[8]) ? 3'b111 : 3'b101;
									assign node923 = (inp[0]) ? node925 : 3'b001;
										assign node925 = (inp[2]) ? 3'b110 : 3'b111;
								assign node928 = (inp[2]) ? node930 : 3'b110;
									assign node930 = (inp[0]) ? node932 : 3'b001;
										assign node932 = (inp[8]) ? 3'b010 : 3'b100;
							assign node935 = (inp[8]) ? node945 : node936;
								assign node936 = (inp[5]) ? node940 : node937;
									assign node937 = (inp[0]) ? 3'b010 : 3'b110;
									assign node940 = (inp[1]) ? node942 : 3'b100;
										assign node942 = (inp[0]) ? 3'b100 : 3'b110;
								assign node945 = (inp[0]) ? node951 : node946;
									assign node946 = (inp[1]) ? 3'b001 : node947;
										assign node947 = (inp[2]) ? 3'b110 : 3'b100;
									assign node951 = (inp[1]) ? node955 : node952;
										assign node952 = (inp[11]) ? 3'b010 : 3'b110;
										assign node955 = (inp[2]) ? 3'b100 : 3'b110;
						assign node958 = (inp[0]) ? node990 : node959;
							assign node959 = (inp[1]) ? node971 : node960;
								assign node960 = (inp[5]) ? node968 : node961;
									assign node961 = (inp[8]) ? node963 : 3'b110;
										assign node963 = (inp[2]) ? 3'b000 : node964;
											assign node964 = (inp[10]) ? 3'b100 : 3'b000;
									assign node968 = (inp[8]) ? 3'b110 : 3'b000;
								assign node971 = (inp[5]) ? node981 : node972;
									assign node972 = (inp[11]) ? 3'b010 : node973;
										assign node973 = (inp[10]) ? node977 : node974;
											assign node974 = (inp[8]) ? 3'b001 : 3'b110;
											assign node977 = (inp[8]) ? 3'b110 : 3'b010;
									assign node981 = (inp[8]) ? node983 : 3'b100;
										assign node983 = (inp[10]) ? node987 : node984;
											assign node984 = (inp[2]) ? 3'b010 : 3'b110;
											assign node987 = (inp[2]) ? 3'b100 : 3'b010;
							assign node990 = (inp[1]) ? node1002 : node991;
								assign node991 = (inp[10]) ? node997 : node992;
									assign node992 = (inp[2]) ? 3'b010 : node993;
										assign node993 = (inp[8]) ? 3'b110 : 3'b010;
									assign node997 = (inp[8]) ? node999 : 3'b100;
										assign node999 = (inp[2]) ? 3'b010 : 3'b100;
								assign node1002 = (inp[11]) ? node1006 : node1003;
									assign node1003 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1006 = (inp[8]) ? 3'b100 : node1007;
										assign node1007 = (inp[10]) ? 3'b000 : node1008;
											assign node1008 = (inp[2]) ? 3'b100 : 3'b000;
					assign node1013 = (inp[0]) ? node1061 : node1014;
						assign node1014 = (inp[4]) ? node1040 : node1015;
							assign node1015 = (inp[10]) ? node1027 : node1016;
								assign node1016 = (inp[1]) ? node1022 : node1017;
									assign node1017 = (inp[8]) ? 3'b111 : node1018;
										assign node1018 = (inp[2]) ? 3'b011 : 3'b111;
									assign node1022 = (inp[11]) ? 3'b011 : node1023;
										assign node1023 = (inp[2]) ? 3'b011 : 3'b111;
								assign node1027 = (inp[1]) ? node1031 : node1028;
									assign node1028 = (inp[8]) ? 3'b011 : 3'b111;
									assign node1031 = (inp[11]) ? node1037 : node1032;
										assign node1032 = (inp[2]) ? node1034 : 3'b011;
											assign node1034 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1037 = (inp[8]) ? 3'b101 : 3'b001;
							assign node1040 = (inp[10]) ? node1054 : node1041;
								assign node1041 = (inp[11]) ? node1045 : node1042;
									assign node1042 = (inp[1]) ? 3'b001 : 3'b011;
									assign node1045 = (inp[5]) ? node1049 : node1046;
										assign node1046 = (inp[8]) ? 3'b101 : 3'b100;
										assign node1049 = (inp[8]) ? node1051 : 3'b001;
											assign node1051 = (inp[1]) ? 3'b001 : 3'b101;
								assign node1054 = (inp[8]) ? node1056 : 3'b110;
									assign node1056 = (inp[1]) ? node1058 : 3'b101;
										assign node1058 = (inp[2]) ? 3'b001 : 3'b101;
						assign node1061 = (inp[4]) ? node1093 : node1062;
							assign node1062 = (inp[1]) ? node1074 : node1063;
								assign node1063 = (inp[2]) ? node1071 : node1064;
									assign node1064 = (inp[11]) ? node1066 : 3'b001;
										assign node1066 = (inp[10]) ? 3'b101 : node1067;
											assign node1067 = (inp[5]) ? 3'b101 : 3'b011;
									assign node1071 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1074 = (inp[10]) ? node1080 : node1075;
									assign node1075 = (inp[8]) ? 3'b001 : node1076;
										assign node1076 = (inp[5]) ? 3'b110 : 3'b001;
									assign node1080 = (inp[11]) ? node1086 : node1081;
										assign node1081 = (inp[5]) ? node1083 : 3'b001;
											assign node1083 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1086 = (inp[8]) ? node1090 : node1087;
											assign node1087 = (inp[5]) ? 3'b010 : 3'b110;
											assign node1090 = (inp[2]) ? 3'b110 : 3'b010;
							assign node1093 = (inp[2]) ? node1113 : node1094;
								assign node1094 = (inp[11]) ? node1106 : node1095;
									assign node1095 = (inp[10]) ? node1101 : node1096;
										assign node1096 = (inp[5]) ? 3'b110 : node1097;
											assign node1097 = (inp[8]) ? 3'b101 : 3'b110;
										assign node1101 = (inp[5]) ? node1103 : 3'b010;
											assign node1103 = (inp[1]) ? 3'b100 : 3'b110;
									assign node1106 = (inp[8]) ? node1108 : 3'b010;
										assign node1108 = (inp[1]) ? 3'b100 : node1109;
											assign node1109 = (inp[10]) ? 3'b010 : 3'b110;
								assign node1113 = (inp[11]) ? node1121 : node1114;
									assign node1114 = (inp[5]) ? 3'b010 : node1115;
										assign node1115 = (inp[10]) ? node1117 : 3'b110;
											assign node1117 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1121 = (inp[10]) ? node1123 : 3'b010;
										assign node1123 = (inp[1]) ? 3'b100 : node1124;
											assign node1124 = (inp[8]) ? 3'b010 : 3'b000;
				assign node1128 = (inp[0]) ? node1232 : node1129;
					assign node1129 = (inp[4]) ? node1183 : node1130;
						assign node1130 = (inp[10]) ? node1158 : node1131;
							assign node1131 = (inp[11]) ? node1147 : node1132;
								assign node1132 = (inp[7]) ? node1140 : node1133;
									assign node1133 = (inp[5]) ? 3'b001 : node1134;
										assign node1134 = (inp[2]) ? 3'b100 : node1135;
											assign node1135 = (inp[8]) ? 3'b100 : 3'b001;
									assign node1140 = (inp[2]) ? 3'b001 : node1141;
										assign node1141 = (inp[1]) ? node1143 : 3'b001;
											assign node1143 = (inp[8]) ? 3'b001 : 3'b110;
								assign node1147 = (inp[5]) ? 3'b110 : node1148;
									assign node1148 = (inp[1]) ? 3'b100 : node1149;
										assign node1149 = (inp[8]) ? node1153 : node1150;
											assign node1150 = (inp[7]) ? 3'b101 : 3'b111;
											assign node1153 = (inp[7]) ? 3'b101 : 3'b001;
							assign node1158 = (inp[7]) ? node1168 : node1159;
								assign node1159 = (inp[5]) ? node1165 : node1160;
									assign node1160 = (inp[1]) ? 3'b010 : node1161;
										assign node1161 = (inp[11]) ? 3'b010 : 3'b110;
									assign node1165 = (inp[1]) ? 3'b100 : 3'b010;
								assign node1168 = (inp[5]) ? node1178 : node1169;
									assign node1169 = (inp[8]) ? node1171 : 3'b110;
										assign node1171 = (inp[2]) ? node1175 : node1172;
											assign node1172 = (inp[1]) ? 3'b001 : 3'b101;
											assign node1175 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1178 = (inp[1]) ? node1180 : 3'b110;
										assign node1180 = (inp[8]) ? 3'b110 : 3'b101;
						assign node1183 = (inp[1]) ? node1209 : node1184;
							assign node1184 = (inp[2]) ? node1196 : node1185;
								assign node1185 = (inp[10]) ? node1187 : 3'b110;
									assign node1187 = (inp[5]) ? node1193 : node1188;
										assign node1188 = (inp[7]) ? node1190 : 3'b010;
											assign node1190 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1193 = (inp[8]) ? 3'b100 : 3'b010;
								assign node1196 = (inp[11]) ? 3'b010 : node1197;
									assign node1197 = (inp[7]) ? node1203 : node1198;
										assign node1198 = (inp[5]) ? node1200 : 3'b110;
											assign node1200 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1203 = (inp[10]) ? node1205 : 3'b001;
											assign node1205 = (inp[5]) ? 3'b010 : 3'b110;
							assign node1209 = (inp[7]) ? node1219 : node1210;
								assign node1210 = (inp[10]) ? 3'b000 : node1211;
									assign node1211 = (inp[5]) ? 3'b000 : node1212;
										assign node1212 = (inp[11]) ? node1214 : 3'b100;
											assign node1214 = (inp[2]) ? 3'b100 : 3'b000;
								assign node1219 = (inp[8]) ? node1221 : 3'b100;
									assign node1221 = (inp[10]) ? node1229 : node1222;
										assign node1222 = (inp[5]) ? node1226 : node1223;
											assign node1223 = (inp[11]) ? 3'b110 : 3'b001;
											assign node1226 = (inp[2]) ? 3'b010 : 3'b010;
										assign node1229 = (inp[5]) ? 3'b100 : 3'b010;
					assign node1232 = (inp[4]) ? node1290 : node1233;
						assign node1233 = (inp[1]) ? node1265 : node1234;
							assign node1234 = (inp[2]) ? node1256 : node1235;
								assign node1235 = (inp[11]) ? node1247 : node1236;
									assign node1236 = (inp[5]) ? node1242 : node1237;
										assign node1237 = (inp[10]) ? 3'b110 : node1238;
											assign node1238 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1242 = (inp[7]) ? node1244 : 3'b100;
											assign node1244 = (inp[10]) ? 3'b000 : 3'b110;
									assign node1247 = (inp[8]) ? node1249 : 3'b101;
										assign node1249 = (inp[10]) ? node1253 : node1250;
											assign node1250 = (inp[5]) ? 3'b110 : 3'b000;
											assign node1253 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1256 = (inp[7]) ? node1258 : 3'b100;
									assign node1258 = (inp[11]) ? node1262 : node1259;
										assign node1259 = (inp[10]) ? 3'b010 : 3'b110;
										assign node1262 = (inp[10]) ? 3'b100 : 3'b110;
							assign node1265 = (inp[7]) ? node1271 : node1266;
								assign node1266 = (inp[11]) ? 3'b000 : node1267;
									assign node1267 = (inp[10]) ? 3'b000 : 3'b100;
								assign node1271 = (inp[10]) ? node1281 : node1272;
									assign node1272 = (inp[11]) ? node1274 : 3'b110;
										assign node1274 = (inp[8]) ? node1278 : node1275;
											assign node1275 = (inp[5]) ? 3'b100 : 3'b010;
											assign node1278 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1281 = (inp[11]) ? node1283 : 3'b010;
										assign node1283 = (inp[8]) ? node1287 : node1284;
											assign node1284 = (inp[5]) ? 3'b000 : 3'b100;
											assign node1287 = (inp[5]) ? 3'b100 : 3'b000;
						assign node1290 = (inp[7]) ? node1292 : 3'b000;
							assign node1292 = (inp[8]) ? node1298 : node1293;
								assign node1293 = (inp[10]) ? 3'b000 : node1294;
									assign node1294 = (inp[1]) ? 3'b000 : 3'b110;
								assign node1298 = (inp[11]) ? node1308 : node1299;
									assign node1299 = (inp[1]) ? 3'b100 : node1300;
										assign node1300 = (inp[5]) ? node1304 : node1301;
											assign node1301 = (inp[10]) ? 3'b010 : 3'b010;
											assign node1304 = (inp[10]) ? 3'b100 : 3'b010;
									assign node1308 = (inp[2]) ? 3'b100 : 3'b000;

endmodule