module dtc_split33_bm34 (
	input  wire [9-1:0] inp,
	output wire [5-1:0] outp
);

	wire [5-1:0] node1;
	wire [5-1:0] node2;
	wire [5-1:0] node3;
	wire [5-1:0] node4;
	wire [5-1:0] node5;
	wire [5-1:0] node6;
	wire [5-1:0] node8;
	wire [5-1:0] node11;
	wire [5-1:0] node12;
	wire [5-1:0] node15;
	wire [5-1:0] node18;
	wire [5-1:0] node19;
	wire [5-1:0] node20;
	wire [5-1:0] node24;
	wire [5-1:0] node25;
	wire [5-1:0] node29;
	wire [5-1:0] node30;
	wire [5-1:0] node31;
	wire [5-1:0] node32;
	wire [5-1:0] node36;
	wire [5-1:0] node39;
	wire [5-1:0] node40;
	wire [5-1:0] node43;
	wire [5-1:0] node45;
	wire [5-1:0] node48;
	wire [5-1:0] node49;
	wire [5-1:0] node50;
	wire [5-1:0] node51;
	wire [5-1:0] node53;
	wire [5-1:0] node57;
	wire [5-1:0] node58;
	wire [5-1:0] node62;
	wire [5-1:0] node63;
	wire [5-1:0] node64;
	wire [5-1:0] node65;
	wire [5-1:0] node69;
	wire [5-1:0] node72;
	wire [5-1:0] node73;
	wire [5-1:0] node76;
	wire [5-1:0] node79;
	wire [5-1:0] node80;
	wire [5-1:0] node81;
	wire [5-1:0] node82;
	wire [5-1:0] node83;
	wire [5-1:0] node86;
	wire [5-1:0] node89;
	wire [5-1:0] node90;
	wire [5-1:0] node91;
	wire [5-1:0] node95;
	wire [5-1:0] node98;
	wire [5-1:0] node100;
	wire [5-1:0] node101;
	wire [5-1:0] node103;
	wire [5-1:0] node106;
	wire [5-1:0] node108;
	wire [5-1:0] node111;
	wire [5-1:0] node112;
	wire [5-1:0] node113;
	wire [5-1:0] node114;
	wire [5-1:0] node117;
	wire [5-1:0] node120;
	wire [5-1:0] node121;
	wire [5-1:0] node122;
	wire [5-1:0] node127;
	wire [5-1:0] node128;
	wire [5-1:0] node130;
	wire [5-1:0] node132;
	wire [5-1:0] node135;
	wire [5-1:0] node136;
	wire [5-1:0] node137;
	wire [5-1:0] node140;
	wire [5-1:0] node143;
	wire [5-1:0] node145;
	wire [5-1:0] node148;
	wire [5-1:0] node149;
	wire [5-1:0] node150;
	wire [5-1:0] node151;
	wire [5-1:0] node153;
	wire [5-1:0] node155;
	wire [5-1:0] node156;
	wire [5-1:0] node160;
	wire [5-1:0] node162;
	wire [5-1:0] node164;
	wire [5-1:0] node166;
	wire [5-1:0] node169;
	wire [5-1:0] node170;
	wire [5-1:0] node171;
	wire [5-1:0] node174;
	wire [5-1:0] node176;
	wire [5-1:0] node179;
	wire [5-1:0] node180;
	wire [5-1:0] node182;
	wire [5-1:0] node184;
	wire [5-1:0] node187;
	wire [5-1:0] node188;
	wire [5-1:0] node191;
	wire [5-1:0] node193;
	wire [5-1:0] node196;
	wire [5-1:0] node197;
	wire [5-1:0] node198;
	wire [5-1:0] node199;
	wire [5-1:0] node200;
	wire [5-1:0] node202;
	wire [5-1:0] node205;
	wire [5-1:0] node208;
	wire [5-1:0] node209;
	wire [5-1:0] node210;
	wire [5-1:0] node214;
	wire [5-1:0] node217;
	wire [5-1:0] node218;
	wire [5-1:0] node219;
	wire [5-1:0] node221;
	wire [5-1:0] node224;
	wire [5-1:0] node227;
	wire [5-1:0] node228;
	wire [5-1:0] node231;
	wire [5-1:0] node232;
	wire [5-1:0] node236;
	wire [5-1:0] node237;
	wire [5-1:0] node238;
	wire [5-1:0] node239;
	wire [5-1:0] node241;
	wire [5-1:0] node246;
	wire [5-1:0] node247;
	wire [5-1:0] node249;
	wire [5-1:0] node250;
	wire [5-1:0] node253;
	wire [5-1:0] node256;
	wire [5-1:0] node258;
	wire [5-1:0] node259;
	wire [5-1:0] node262;

	assign outp = (inp[2]) ? node148 : node1;
		assign node1 = (inp[0]) ? node79 : node2;
			assign node2 = (inp[7]) ? node48 : node3;
				assign node3 = (inp[8]) ? node29 : node4;
					assign node4 = (inp[5]) ? node18 : node5;
						assign node5 = (inp[1]) ? node11 : node6;
							assign node6 = (inp[6]) ? node8 : 5'b00111;
								assign node8 = (inp[3]) ? 5'b10111 : 5'b10110;
							assign node11 = (inp[3]) ? node15 : node12;
								assign node12 = (inp[4]) ? 5'b01011 : 5'b00110;
								assign node15 = (inp[4]) ? 5'b00110 : 5'b00111;
						assign node18 = (inp[6]) ? node24 : node19;
							assign node19 = (inp[4]) ? 5'b00011 : node20;
								assign node20 = (inp[1]) ? 5'b11010 : 5'b01010;
							assign node24 = (inp[1]) ? 5'b01010 : node25;
								assign node25 = (inp[3]) ? 5'b11010 : 5'b11010;
					assign node29 = (inp[5]) ? node39 : node30;
						assign node30 = (inp[3]) ? node36 : node31;
							assign node31 = (inp[4]) ? 5'b10001 : node32;
								assign node32 = (inp[6]) ? 5'b11000 : 5'b01000;
							assign node36 = (inp[1]) ? 5'b00001 : 5'b10001;
						assign node39 = (inp[6]) ? node43 : node40;
							assign node40 = (inp[3]) ? 5'b00000 : 5'b10000;
							assign node43 = (inp[1]) ? node45 : 5'b11111;
								assign node45 = (inp[4]) ? 5'b01110 : 5'b01111;
				assign node48 = (inp[6]) ? node62 : node49;
					assign node49 = (inp[1]) ? node57 : node50;
						assign node50 = (inp[8]) ? 5'b00111 : node51;
							assign node51 = (inp[4]) ? node53 : 5'b00111;
								assign node53 = (inp[3]) ? 5'b00110 : 5'b00111;
						assign node57 = (inp[4]) ? 5'b10110 : node58;
							assign node58 = (inp[3]) ? 5'b10110 : 5'b11011;
					assign node62 = (inp[1]) ? node72 : node63;
						assign node63 = (inp[3]) ? node69 : node64;
							assign node64 = (inp[8]) ? 5'b10000 : node65;
								assign node65 = (inp[5]) ? 5'b10110 : 5'b11110;
							assign node69 = (inp[4]) ? 5'b11110 : 5'b11111;
						assign node72 = (inp[4]) ? node76 : node73;
							assign node73 = (inp[3]) ? 5'b01111 : 5'b00110;
							assign node76 = (inp[5]) ? 5'b01011 : 5'b01110;
			assign node79 = (inp[8]) ? node111 : node80;
				assign node80 = (inp[5]) ? node98 : node81;
					assign node81 = (inp[3]) ? node89 : node82;
						assign node82 = (inp[6]) ? node86 : node83;
							assign node83 = (inp[7]) ? 5'b10010 : 5'b00010;
							assign node86 = (inp[7]) ? 5'b10011 : 5'b10010;
						assign node89 = (inp[7]) ? node95 : node90;
							assign node90 = (inp[4]) ? 5'b00010 : node91;
								assign node91 = (inp[1]) ? 5'b00011 : 5'b10011;
							assign node95 = (inp[4]) ? 5'b01010 : 5'b01011;
					assign node98 = (inp[7]) ? node100 : 5'b00010;
						assign node100 = (inp[4]) ? node106 : node101;
							assign node101 = (inp[1]) ? node103 : 5'b10010;
								assign node103 = (inp[3]) ? 5'b10010 : 5'b00010;
							assign node106 = (inp[3]) ? node108 : 5'b00010;
								assign node108 = (inp[6]) ? 5'b10010 : 5'b00010;
				assign node111 = (inp[5]) ? node127 : node112;
					assign node112 = (inp[7]) ? node120 : node113;
						assign node113 = (inp[4]) ? node117 : node114;
							assign node114 = (inp[3]) ? 5'b10111 : 5'b11110;
							assign node117 = (inp[6]) ? 5'b00111 : 5'b10111;
						assign node120 = (inp[4]) ? 5'b01010 : node121;
							assign node121 = (inp[3]) ? 5'b00110 : node122;
								assign node122 = (inp[1]) ? 5'b00110 : 5'b10110;
					assign node127 = (inp[7]) ? node135 : node128;
						assign node128 = (inp[3]) ? node130 : 5'b11011;
							assign node130 = (inp[1]) ? node132 : 5'b11010;
								assign node132 = (inp[6]) ? 5'b01010 : 5'b11010;
						assign node135 = (inp[4]) ? node143 : node136;
							assign node136 = (inp[3]) ? node140 : node137;
								assign node137 = (inp[6]) ? 5'b11010 : 5'b01011;
								assign node140 = (inp[6]) ? 5'b00011 : 5'b10011;
							assign node143 = (inp[3]) ? node145 : 5'b10011;
								assign node145 = (inp[1]) ? 5'b00010 : 5'b10010;
		assign node148 = (inp[0]) ? node196 : node149;
			assign node149 = (inp[5]) ? node169 : node150;
				assign node150 = (inp[8]) ? node160 : node151;
					assign node151 = (inp[3]) ? node153 : 5'b01100;
						assign node153 = (inp[1]) ? node155 : 5'b11101;
							assign node155 = (inp[6]) ? 5'b00101 : node156;
								assign node156 = (inp[4]) ? 5'b10001 : 5'b10100;
					assign node160 = (inp[7]) ? node162 : 5'b11101;
						assign node162 = (inp[4]) ? node164 : 5'b11101;
							assign node164 = (inp[6]) ? node166 : 5'b11100;
								assign node166 = (inp[1]) ? 5'b01100 : 5'b11100;
				assign node169 = (inp[7]) ? node179 : node170;
					assign node170 = (inp[4]) ? node174 : node171;
						assign node171 = (inp[6]) ? 5'b11001 : 5'b11101;
						assign node174 = (inp[3]) ? node176 : 5'b01101;
							assign node176 = (inp[1]) ? 5'b01100 : 5'b11100;
					assign node179 = (inp[3]) ? node187 : node180;
						assign node180 = (inp[8]) ? node182 : 5'b01001;
							assign node182 = (inp[6]) ? node184 : 5'b01100;
								assign node184 = (inp[4]) ? 5'b00101 : 5'b01100;
						assign node187 = (inp[4]) ? node191 : node188;
							assign node188 = (inp[6]) ? 5'b00101 : 5'b10101;
							assign node191 = (inp[8]) ? node193 : 5'b10100;
								assign node193 = (inp[1]) ? 5'b00100 : 5'b00101;
			assign node196 = (inp[8]) ? node236 : node197;
				assign node197 = (inp[5]) ? node217 : node198;
					assign node198 = (inp[4]) ? node208 : node199;
						assign node199 = (inp[7]) ? node205 : node200;
							assign node200 = (inp[3]) ? node202 : 5'b00000;
								assign node202 = (inp[1]) ? 5'b00001 : 5'b10001;
							assign node205 = (inp[1]) ? 5'b01001 : 5'b11001;
						assign node208 = (inp[3]) ? node214 : node209;
							assign node209 = (inp[7]) ? 5'b00001 : node210;
								assign node210 = (inp[6]) ? 5'b11111 : 5'b11110;
							assign node214 = (inp[7]) ? 5'b11000 : 5'b10000;
					assign node217 = (inp[7]) ? node227 : node218;
						assign node218 = (inp[3]) ? node224 : node219;
							assign node219 = (inp[4]) ? node221 : 5'b01110;
								assign node221 = (inp[6]) ? 5'b10111 : 5'b00111;
							assign node224 = (inp[4]) ? 5'b01110 : 5'b01111;
						assign node227 = (inp[4]) ? node231 : node228;
							assign node228 = (inp[1]) ? 5'b00000 : 5'b10000;
							assign node231 = (inp[3]) ? 5'b00000 : node232;
								assign node232 = (inp[1]) ? 5'b01111 : 5'b11111;
				assign node236 = (inp[5]) ? node246 : node237;
					assign node237 = (inp[6]) ? 5'b01000 : node238;
						assign node238 = (inp[1]) ? 5'b10100 : node239;
							assign node239 = (inp[7]) ? node241 : 5'b01101;
								assign node241 = (inp[3]) ? 5'b00000 : 5'b00100;
					assign node246 = (inp[1]) ? node256 : node247;
						assign node247 = (inp[6]) ? node249 : 5'b01001;
							assign node249 = (inp[7]) ? node253 : node250;
								assign node250 = (inp[3]) ? 5'b11000 : 5'b11001;
								assign node253 = (inp[4]) ? 5'b10001 : 5'b11000;
						assign node256 = (inp[3]) ? node258 : 5'b00100;
							assign node258 = (inp[7]) ? node262 : node259;
								assign node259 = (inp[6]) ? 5'b01001 : 5'b11001;
								assign node262 = (inp[6]) ? 5'b00001 : 5'b10000;

endmodule