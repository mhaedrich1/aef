module dtc_split875_bm89 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node121;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node205;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node318;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node334;
	wire [3-1:0] node337;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node351;
	wire [3-1:0] node354;
	wire [3-1:0] node356;
	wire [3-1:0] node358;
	wire [3-1:0] node361;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node394;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node408;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node413;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node428;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node439;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node463;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node478;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node489;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node520;
	wire [3-1:0] node522;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node528;
	wire [3-1:0] node531;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node555;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node562;
	wire [3-1:0] node564;
	wire [3-1:0] node567;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node576;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node583;
	wire [3-1:0] node585;
	wire [3-1:0] node588;
	wire [3-1:0] node590;
	wire [3-1:0] node593;
	wire [3-1:0] node595;
	wire [3-1:0] node597;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node611;
	wire [3-1:0] node612;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node625;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node644;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node660;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node669;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node675;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node686;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node719;
	wire [3-1:0] node721;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node727;
	wire [3-1:0] node729;
	wire [3-1:0] node732;
	wire [3-1:0] node734;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node746;
	wire [3-1:0] node750;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node759;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node769;
	wire [3-1:0] node773;
	wire [3-1:0] node775;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node784;
	wire [3-1:0] node786;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node793;
	wire [3-1:0] node796;
	wire [3-1:0] node798;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node804;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node821;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node843;
	wire [3-1:0] node846;
	wire [3-1:0] node848;
	wire [3-1:0] node851;
	wire [3-1:0] node852;
	wire [3-1:0] node854;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node861;
	wire [3-1:0] node863;
	wire [3-1:0] node867;
	wire [3-1:0] node868;
	wire [3-1:0] node869;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node883;
	wire [3-1:0] node885;
	wire [3-1:0] node887;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node910;
	wire [3-1:0] node913;
	wire [3-1:0] node915;
	wire [3-1:0] node918;
	wire [3-1:0] node920;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node927;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node938;
	wire [3-1:0] node940;
	wire [3-1:0] node942;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node948;
	wire [3-1:0] node951;
	wire [3-1:0] node953;
	wire [3-1:0] node955;
	wire [3-1:0] node958;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node965;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node976;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node984;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node990;
	wire [3-1:0] node992;
	wire [3-1:0] node995;
	wire [3-1:0] node997;
	wire [3-1:0] node999;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1012;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1020;
	wire [3-1:0] node1023;
	wire [3-1:0] node1025;
	wire [3-1:0] node1027;
	wire [3-1:0] node1030;
	wire [3-1:0] node1032;
	wire [3-1:0] node1033;
	wire [3-1:0] node1038;
	wire [3-1:0] node1039;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;
	wire [3-1:0] node1049;
	wire [3-1:0] node1052;
	wire [3-1:0] node1055;
	wire [3-1:0] node1056;
	wire [3-1:0] node1059;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1066;
	wire [3-1:0] node1068;
	wire [3-1:0] node1070;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1078;
	wire [3-1:0] node1079;
	wire [3-1:0] node1082;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1091;
	wire [3-1:0] node1094;
	wire [3-1:0] node1096;
	wire [3-1:0] node1099;
	wire [3-1:0] node1101;
	wire [3-1:0] node1103;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1109;
	wire [3-1:0] node1111;
	wire [3-1:0] node1113;
	wire [3-1:0] node1116;
	wire [3-1:0] node1117;
	wire [3-1:0] node1120;
	wire [3-1:0] node1122;
	wire [3-1:0] node1125;
	wire [3-1:0] node1126;
	wire [3-1:0] node1127;
	wire [3-1:0] node1128;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1133;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1142;
	wire [3-1:0] node1144;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1151;
	wire [3-1:0] node1153;
	wire [3-1:0] node1156;
	wire [3-1:0] node1157;
	wire [3-1:0] node1158;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1162;
	wire [3-1:0] node1167;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1176;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1182;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1192;
	wire [3-1:0] node1196;
	wire [3-1:0] node1197;
	wire [3-1:0] node1199;
	wire [3-1:0] node1203;
	wire [3-1:0] node1205;
	wire [3-1:0] node1208;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1212;
	wire [3-1:0] node1214;
	wire [3-1:0] node1217;
	wire [3-1:0] node1218;
	wire [3-1:0] node1220;
	wire [3-1:0] node1224;
	wire [3-1:0] node1226;
	wire [3-1:0] node1229;
	wire [3-1:0] node1230;
	wire [3-1:0] node1231;
	wire [3-1:0] node1233;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1239;
	wire [3-1:0] node1240;
	wire [3-1:0] node1244;
	wire [3-1:0] node1246;
	wire [3-1:0] node1249;
	wire [3-1:0] node1250;
	wire [3-1:0] node1252;
	wire [3-1:0] node1254;
	wire [3-1:0] node1256;
	wire [3-1:0] node1259;
	wire [3-1:0] node1260;
	wire [3-1:0] node1262;
	wire [3-1:0] node1265;
	wire [3-1:0] node1267;
	wire [3-1:0] node1269;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1276;
	wire [3-1:0] node1277;
	wire [3-1:0] node1279;
	wire [3-1:0] node1283;
	wire [3-1:0] node1284;
	wire [3-1:0] node1285;
	wire [3-1:0] node1288;
	wire [3-1:0] node1290;
	wire [3-1:0] node1293;
	wire [3-1:0] node1294;
	wire [3-1:0] node1296;
	wire [3-1:0] node1298;
	wire [3-1:0] node1301;
	wire [3-1:0] node1303;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1312;
	wire [3-1:0] node1313;
	wire [3-1:0] node1314;
	wire [3-1:0] node1318;
	wire [3-1:0] node1319;
	wire [3-1:0] node1321;
	wire [3-1:0] node1324;
	wire [3-1:0] node1325;
	wire [3-1:0] node1328;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1335;
	wire [3-1:0] node1337;
	wire [3-1:0] node1339;
	wire [3-1:0] node1342;
	wire [3-1:0] node1343;
	wire [3-1:0] node1344;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1351;
	wire [3-1:0] node1353;
	wire [3-1:0] node1356;
	wire [3-1:0] node1357;
	wire [3-1:0] node1358;
	wire [3-1:0] node1360;
	wire [3-1:0] node1363;
	wire [3-1:0] node1365;
	wire [3-1:0] node1368;
	wire [3-1:0] node1370;
	wire [3-1:0] node1372;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1377;
	wire [3-1:0] node1379;
	wire [3-1:0] node1381;
	wire [3-1:0] node1385;
	wire [3-1:0] node1386;
	wire [3-1:0] node1387;
	wire [3-1:0] node1389;
	wire [3-1:0] node1392;
	wire [3-1:0] node1394;
	wire [3-1:0] node1396;
	wire [3-1:0] node1399;
	wire [3-1:0] node1400;
	wire [3-1:0] node1401;
	wire [3-1:0] node1403;
	wire [3-1:0] node1406;
	wire [3-1:0] node1408;
	wire [3-1:0] node1412;
	wire [3-1:0] node1413;
	wire [3-1:0] node1414;
	wire [3-1:0] node1415;
	wire [3-1:0] node1417;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1425;
	wire [3-1:0] node1426;
	wire [3-1:0] node1427;
	wire [3-1:0] node1428;
	wire [3-1:0] node1433;
	wire [3-1:0] node1434;
	wire [3-1:0] node1436;
	wire [3-1:0] node1439;
	wire [3-1:0] node1441;
	wire [3-1:0] node1444;
	wire [3-1:0] node1445;
	wire [3-1:0] node1446;
	wire [3-1:0] node1447;

	assign outp = (inp[6]) ? node824 : node1;
		assign node1 = (inp[9]) ? node417 : node2;
			assign node2 = (inp[3]) ? node270 : node3;
				assign node3 = (inp[4]) ? node135 : node4;
					assign node4 = (inp[7]) ? node36 : node5;
						assign node5 = (inp[10]) ? 3'b111 : node6;
							assign node6 = (inp[5]) ? node28 : node7;
								assign node7 = (inp[11]) ? node15 : node8;
									assign node8 = (inp[8]) ? node10 : 3'b101;
										assign node10 = (inp[1]) ? node12 : 3'b101;
											assign node12 = (inp[0]) ? 3'b011 : 3'b101;
									assign node15 = (inp[8]) ? node21 : node16;
										assign node16 = (inp[0]) ? node18 : 3'b101;
											assign node18 = (inp[2]) ? 3'b011 : 3'b101;
										assign node21 = (inp[2]) ? node23 : 3'b011;
											assign node23 = (inp[1]) ? node25 : 3'b011;
												assign node25 = (inp[0]) ? 3'b101 : 3'b011;
								assign node28 = (inp[11]) ? node30 : 3'b011;
									assign node30 = (inp[8]) ? 3'b101 : node31;
										assign node31 = (inp[2]) ? 3'b101 : 3'b011;
						assign node36 = (inp[10]) ? node82 : node37;
							assign node37 = (inp[11]) ? node59 : node38;
								assign node38 = (inp[8]) ? node48 : node39;
									assign node39 = (inp[5]) ? node43 : node40;
										assign node40 = (inp[0]) ? 3'b110 : 3'b010;
										assign node43 = (inp[1]) ? node45 : 3'b110;
											assign node45 = (inp[0]) ? 3'b010 : 3'b110;
									assign node48 = (inp[5]) ? node52 : node49;
										assign node49 = (inp[2]) ? 3'b010 : 3'b110;
										assign node52 = (inp[0]) ? node54 : 3'b000;
											assign node54 = (inp[2]) ? node56 : 3'b000;
												assign node56 = (inp[1]) ? 3'b100 : 3'b000;
								assign node59 = (inp[5]) ? node69 : node60;
									assign node60 = (inp[8]) ? node66 : node61;
										assign node61 = (inp[0]) ? node63 : 3'b111;
											assign node63 = (inp[2]) ? 3'b001 : 3'b011;
										assign node66 = (inp[2]) ? 3'b101 : 3'b001;
									assign node69 = (inp[8]) ? 3'b110 : node70;
										assign node70 = (inp[2]) ? node76 : node71;
											assign node71 = (inp[0]) ? node73 : 3'b001;
												assign node73 = (inp[1]) ? 3'b100 : 3'b001;
											assign node76 = (inp[1]) ? node78 : 3'b011;
												assign node78 = (inp[0]) ? 3'b110 : 3'b011;
							assign node82 = (inp[8]) ? node114 : node83;
								assign node83 = (inp[11]) ? node103 : node84;
									assign node84 = (inp[1]) ? node90 : node85;
										assign node85 = (inp[5]) ? 3'b101 : node86;
											assign node86 = (inp[0]) ? 3'b101 : 3'b001;
										assign node90 = (inp[2]) ? node96 : node91;
											assign node91 = (inp[5]) ? 3'b001 : node92;
												assign node92 = (inp[0]) ? 3'b101 : 3'b001;
											assign node96 = (inp[5]) ? node100 : node97;
												assign node97 = (inp[0]) ? 3'b101 : 3'b001;
												assign node100 = (inp[0]) ? 3'b001 : 3'b101;
									assign node103 = (inp[5]) ? node109 : node104;
										assign node104 = (inp[0]) ? node106 : 3'b101;
											assign node106 = (inp[1]) ? 3'b011 : 3'b001;
										assign node109 = (inp[2]) ? node111 : 3'b011;
											assign node111 = (inp[1]) ? 3'b101 : 3'b001;
								assign node114 = (inp[11]) ? node124 : node115;
									assign node115 = (inp[5]) ? node119 : node116;
										assign node116 = (inp[2]) ? 3'b001 : 3'b101;
										assign node119 = (inp[0]) ? node121 : 3'b010;
											assign node121 = (inp[2]) ? 3'b110 : 3'b010;
									assign node124 = (inp[5]) ? node130 : node125;
										assign node125 = (inp[2]) ? node127 : 3'b011;
											assign node127 = (inp[0]) ? 3'b101 : 3'b111;
										assign node130 = (inp[2]) ? node132 : 3'b101;
											assign node132 = (inp[1]) ? 3'b001 : 3'b101;
					assign node135 = (inp[10]) ? node191 : node136;
						assign node136 = (inp[7]) ? node156 : node137;
							assign node137 = (inp[8]) ? node147 : node138;
								assign node138 = (inp[11]) ? node140 : 3'b010;
									assign node140 = (inp[2]) ? 3'b110 : node141;
										assign node141 = (inp[0]) ? 3'b110 : node142;
											assign node142 = (inp[1]) ? 3'b110 : 3'b001;
								assign node147 = (inp[11]) ? node149 : 3'b100;
									assign node149 = (inp[1]) ? 3'b010 : node150;
										assign node150 = (inp[0]) ? 3'b110 : node151;
											assign node151 = (inp[2]) ? 3'b110 : 3'b101;
							assign node156 = (inp[5]) ? node174 : node157;
								assign node157 = (inp[11]) ? node165 : node158;
									assign node158 = (inp[8]) ? node160 : 3'b100;
										assign node160 = (inp[0]) ? node162 : 3'b100;
											assign node162 = (inp[1]) ? 3'b000 : 3'b100;
									assign node165 = (inp[8]) ? node169 : node166;
										assign node166 = (inp[2]) ? 3'b010 : 3'b100;
										assign node169 = (inp[2]) ? 3'b100 : node170;
											assign node170 = (inp[1]) ? 3'b100 : 3'b000;
								assign node174 = (inp[11]) ? node176 : 3'b000;
									assign node176 = (inp[8]) ? node182 : node177;
										assign node177 = (inp[2]) ? node179 : 3'b010;
											assign node179 = (inp[1]) ? 3'b100 : 3'b010;
										assign node182 = (inp[0]) ? 3'b000 : node183;
											assign node183 = (inp[2]) ? node187 : node184;
												assign node184 = (inp[1]) ? 3'b100 : 3'b000;
												assign node187 = (inp[1]) ? 3'b000 : 3'b100;
						assign node191 = (inp[7]) ? node235 : node192;
							assign node192 = (inp[8]) ? node214 : node193;
								assign node193 = (inp[11]) ? node209 : node194;
									assign node194 = (inp[1]) ? node202 : node195;
										assign node195 = (inp[5]) ? node197 : 3'b101;
											assign node197 = (inp[0]) ? node199 : 3'b101;
												assign node199 = (inp[2]) ? 3'b101 : 3'b001;
										assign node202 = (inp[2]) ? 3'b001 : node203;
											assign node203 = (inp[5]) ? node205 : 3'b101;
												assign node205 = (inp[0]) ? 3'b001 : 3'b101;
									assign node209 = (inp[0]) ? node211 : 3'b011;
										assign node211 = (inp[5]) ? 3'b101 : 3'b011;
								assign node214 = (inp[11]) ? node230 : node215;
									assign node215 = (inp[1]) ? node223 : node216;
										assign node216 = (inp[0]) ? node218 : 3'b001;
											assign node218 = (inp[5]) ? node220 : 3'b001;
												assign node220 = (inp[2]) ? 3'b001 : 3'b110;
										assign node223 = (inp[2]) ? 3'b110 : node224;
											assign node224 = (inp[5]) ? node226 : 3'b001;
												assign node226 = (inp[0]) ? 3'b110 : 3'b001;
									assign node230 = (inp[0]) ? node232 : 3'b101;
										assign node232 = (inp[5]) ? 3'b001 : 3'b101;
							assign node235 = (inp[11]) ? node247 : node236;
								assign node236 = (inp[8]) ? node242 : node237;
									assign node237 = (inp[5]) ? node239 : 3'b110;
										assign node239 = (inp[0]) ? 3'b010 : 3'b110;
									assign node242 = (inp[5]) ? node244 : 3'b010;
										assign node244 = (inp[0]) ? 3'b100 : 3'b010;
								assign node247 = (inp[8]) ? node257 : node248;
									assign node248 = (inp[0]) ? node250 : 3'b001;
										assign node250 = (inp[5]) ? node252 : 3'b001;
											assign node252 = (inp[1]) ? 3'b110 : node253;
												assign node253 = (inp[2]) ? 3'b110 : 3'b001;
									assign node257 = (inp[5]) ? node265 : node258;
										assign node258 = (inp[2]) ? node262 : node259;
											assign node259 = (inp[0]) ? 3'b101 : 3'b001;
											assign node262 = (inp[0]) ? 3'b110 : 3'b010;
										assign node265 = (inp[1]) ? node267 : 3'b110;
											assign node267 = (inp[0]) ? 3'b010 : 3'b110;
				assign node270 = (inp[4]) ? node406 : node271;
					assign node271 = (inp[7]) ? node361 : node272;
						assign node272 = (inp[10]) ? node310 : node273;
							assign node273 = (inp[11]) ? node283 : node274;
								assign node274 = (inp[8]) ? 3'b000 : node275;
									assign node275 = (inp[1]) ? node277 : 3'b100;
										assign node277 = (inp[5]) ? node279 : 3'b100;
											assign node279 = (inp[0]) ? 3'b000 : 3'b100;
								assign node283 = (inp[5]) ? node297 : node284;
									assign node284 = (inp[2]) ? node290 : node285;
										assign node285 = (inp[0]) ? 3'b010 : node286;
											assign node286 = (inp[8]) ? 3'b010 : 3'b110;
										assign node290 = (inp[8]) ? node294 : node291;
											assign node291 = (inp[0]) ? 3'b010 : 3'b110;
											assign node294 = (inp[1]) ? 3'b100 : 3'b110;
									assign node297 = (inp[8]) ? node303 : node298;
										assign node298 = (inp[0]) ? node300 : 3'b010;
											assign node300 = (inp[1]) ? 3'b100 : 3'b010;
										assign node303 = (inp[0]) ? node305 : 3'b100;
											assign node305 = (inp[2]) ? node307 : 3'b100;
												assign node307 = (inp[1]) ? 3'b000 : 3'b100;
							assign node310 = (inp[11]) ? node330 : node311;
								assign node311 = (inp[8]) ? node321 : node312;
									assign node312 = (inp[5]) ? node316 : node313;
										assign node313 = (inp[0]) ? 3'b110 : 3'b010;
										assign node316 = (inp[1]) ? node318 : 3'b110;
											assign node318 = (inp[0]) ? 3'b010 : 3'b110;
									assign node321 = (inp[5]) ? node325 : node322;
										assign node322 = (inp[2]) ? 3'b010 : 3'b110;
										assign node325 = (inp[2]) ? node327 : 3'b000;
											assign node327 = (inp[1]) ? 3'b100 : 3'b000;
								assign node330 = (inp[5]) ? node342 : node331;
									assign node331 = (inp[8]) ? node337 : node332;
										assign node332 = (inp[0]) ? node334 : 3'b111;
											assign node334 = (inp[2]) ? 3'b001 : 3'b011;
										assign node337 = (inp[2]) ? node339 : 3'b001;
											assign node339 = (inp[0]) ? 3'b110 : 3'b101;
									assign node342 = (inp[8]) ? node354 : node343;
										assign node343 = (inp[2]) ? node349 : node344;
											assign node344 = (inp[1]) ? node346 : 3'b001;
												assign node346 = (inp[0]) ? 3'b100 : 3'b001;
											assign node349 = (inp[0]) ? node351 : 3'b011;
												assign node351 = (inp[1]) ? 3'b110 : 3'b011;
										assign node354 = (inp[2]) ? node356 : 3'b110;
											assign node356 = (inp[0]) ? node358 : 3'b110;
												assign node358 = (inp[1]) ? 3'b010 : 3'b110;
						assign node361 = (inp[10]) ? node363 : 3'b000;
							assign node363 = (inp[8]) ? node391 : node364;
								assign node364 = (inp[11]) ? node370 : node365;
									assign node365 = (inp[0]) ? node367 : 3'b100;
										assign node367 = (inp[5]) ? 3'b000 : 3'b100;
									assign node370 = (inp[0]) ? node380 : node371;
										assign node371 = (inp[5]) ? node373 : 3'b010;
											assign node373 = (inp[1]) ? node377 : node374;
												assign node374 = (inp[2]) ? 3'b010 : 3'b000;
												assign node377 = (inp[2]) ? 3'b000 : 3'b010;
										assign node380 = (inp[5]) ? node384 : node381;
											assign node381 = (inp[2]) ? 3'b010 : 3'b000;
											assign node384 = (inp[1]) ? node388 : node385;
												assign node385 = (inp[2]) ? 3'b110 : 3'b000;
												assign node388 = (inp[2]) ? 3'b100 : 3'b110;
								assign node391 = (inp[11]) ? node397 : node392;
									assign node392 = (inp[5]) ? node394 : 3'b000;
										assign node394 = (inp[0]) ? 3'b100 : 3'b000;
									assign node397 = (inp[5]) ? node401 : node398;
										assign node398 = (inp[0]) ? 3'b100 : 3'b000;
										assign node401 = (inp[0]) ? node403 : 3'b100;
											assign node403 = (inp[1]) ? 3'b000 : 3'b100;
					assign node406 = (inp[10]) ? node408 : 3'b000;
						assign node408 = (inp[11]) ? node410 : 3'b000;
							assign node410 = (inp[7]) ? 3'b000 : node411;
								assign node411 = (inp[8]) ? node413 : 3'b100;
									assign node413 = (inp[5]) ? 3'b000 : 3'b100;
			assign node417 = (inp[7]) ? node513 : node418;
				assign node418 = (inp[3]) ? node420 : 3'b111;
					assign node420 = (inp[4]) ? node452 : node421;
						assign node421 = (inp[10]) ? 3'b111 : node422;
							assign node422 = (inp[5]) ? node444 : node423;
								assign node423 = (inp[8]) ? node431 : node424;
									assign node424 = (inp[2]) ? node426 : 3'b101;
										assign node426 = (inp[11]) ? node428 : 3'b101;
											assign node428 = (inp[0]) ? 3'b011 : 3'b101;
									assign node431 = (inp[11]) ? node437 : node432;
										assign node432 = (inp[0]) ? node434 : 3'b101;
											assign node434 = (inp[1]) ? 3'b011 : 3'b101;
										assign node437 = (inp[1]) ? node439 : 3'b011;
											assign node439 = (inp[2]) ? node441 : 3'b011;
												assign node441 = (inp[0]) ? 3'b101 : 3'b011;
								assign node444 = (inp[11]) ? node446 : 3'b011;
									assign node446 = (inp[8]) ? 3'b101 : node447;
										assign node447 = (inp[2]) ? 3'b101 : 3'b011;
						assign node452 = (inp[10]) ? node472 : node453;
							assign node453 = (inp[8]) ? node463 : node454;
								assign node454 = (inp[11]) ? node456 : 3'b010;
									assign node456 = (inp[2]) ? 3'b110 : node457;
										assign node457 = (inp[0]) ? 3'b110 : node458;
											assign node458 = (inp[1]) ? 3'b110 : 3'b001;
								assign node463 = (inp[11]) ? node465 : 3'b100;
									assign node465 = (inp[1]) ? 3'b010 : node466;
										assign node466 = (inp[2]) ? 3'b110 : node467;
											assign node467 = (inp[0]) ? 3'b110 : 3'b101;
							assign node472 = (inp[8]) ? node494 : node473;
								assign node473 = (inp[11]) ? node489 : node474;
									assign node474 = (inp[1]) ? node482 : node475;
										assign node475 = (inp[2]) ? 3'b101 : node476;
											assign node476 = (inp[5]) ? node478 : 3'b101;
												assign node478 = (inp[0]) ? 3'b001 : 3'b101;
										assign node482 = (inp[2]) ? 3'b001 : node483;
											assign node483 = (inp[5]) ? node485 : 3'b101;
												assign node485 = (inp[0]) ? 3'b001 : 3'b101;
									assign node489 = (inp[0]) ? node491 : 3'b011;
										assign node491 = (inp[5]) ? 3'b101 : 3'b011;
								assign node494 = (inp[11]) ? node508 : node495;
									assign node495 = (inp[1]) ? node503 : node496;
										assign node496 = (inp[5]) ? node498 : 3'b001;
											assign node498 = (inp[0]) ? node500 : 3'b001;
												assign node500 = (inp[2]) ? 3'b001 : 3'b110;
										assign node503 = (inp[5]) ? 3'b110 : node504;
											assign node504 = (inp[2]) ? 3'b110 : 3'b001;
									assign node508 = (inp[5]) ? node510 : 3'b101;
										assign node510 = (inp[0]) ? 3'b001 : 3'b101;
				assign node513 = (inp[10]) ? node683 : node514;
					assign node514 = (inp[4]) ? node600 : node515;
						assign node515 = (inp[3]) ? node543 : node516;
							assign node516 = (inp[5]) ? node536 : node517;
								assign node517 = (inp[8]) ? node525 : node518;
									assign node518 = (inp[0]) ? node520 : 3'b110;
										assign node520 = (inp[2]) ? node522 : 3'b110;
											assign node522 = (inp[11]) ? 3'b000 : 3'b110;
									assign node525 = (inp[11]) ? node531 : node526;
										assign node526 = (inp[0]) ? node528 : 3'b110;
											assign node528 = (inp[1]) ? 3'b000 : 3'b110;
										assign node531 = (inp[2]) ? node533 : 3'b000;
											assign node533 = (inp[0]) ? 3'b110 : 3'b000;
								assign node536 = (inp[11]) ? node538 : 3'b000;
									assign node538 = (inp[2]) ? 3'b110 : node539;
										assign node539 = (inp[8]) ? 3'b110 : 3'b000;
							assign node543 = (inp[11]) ? node567 : node544;
								assign node544 = (inp[8]) ? node558 : node545;
									assign node545 = (inp[1]) ? node551 : node546;
										assign node546 = (inp[5]) ? 3'b110 : node547;
											assign node547 = (inp[0]) ? 3'b110 : 3'b010;
										assign node551 = (inp[0]) ? node555 : node552;
											assign node552 = (inp[5]) ? 3'b110 : 3'b010;
											assign node555 = (inp[5]) ? 3'b010 : 3'b110;
									assign node558 = (inp[5]) ? node562 : node559;
										assign node559 = (inp[2]) ? 3'b010 : 3'b110;
										assign node562 = (inp[0]) ? node564 : 3'b000;
											assign node564 = (inp[1]) ? 3'b100 : 3'b000;
								assign node567 = (inp[5]) ? node581 : node568;
									assign node568 = (inp[8]) ? node574 : node569;
										assign node569 = (inp[0]) ? node571 : 3'b111;
											assign node571 = (inp[2]) ? 3'b001 : 3'b011;
										assign node574 = (inp[2]) ? node576 : 3'b001;
											assign node576 = (inp[0]) ? node578 : 3'b101;
												assign node578 = (inp[1]) ? 3'b110 : 3'b101;
									assign node581 = (inp[8]) ? node593 : node582;
										assign node582 = (inp[2]) ? node588 : node583;
											assign node583 = (inp[1]) ? node585 : 3'b001;
												assign node585 = (inp[0]) ? 3'b100 : 3'b001;
											assign node588 = (inp[1]) ? node590 : 3'b011;
												assign node590 = (inp[0]) ? 3'b110 : 3'b011;
										assign node593 = (inp[0]) ? node595 : 3'b110;
											assign node595 = (inp[2]) ? node597 : 3'b110;
												assign node597 = (inp[1]) ? 3'b010 : 3'b110;
						assign node600 = (inp[3]) ? node640 : node601;
							assign node601 = (inp[8]) ? node621 : node602;
								assign node602 = (inp[11]) ? node604 : 3'b001;
									assign node604 = (inp[2]) ? node616 : node605;
										assign node605 = (inp[5]) ? node611 : node606;
											assign node606 = (inp[0]) ? 3'b101 : node607;
												assign node607 = (inp[1]) ? 3'b101 : 3'b011;
											assign node611 = (inp[0]) ? 3'b100 : node612;
												assign node612 = (inp[1]) ? 3'b100 : 3'b010;
										assign node616 = (inp[5]) ? 3'b101 : node617;
											assign node617 = (inp[0]) ? 3'b100 : 3'b101;
								assign node621 = (inp[11]) ? node625 : node622;
									assign node622 = (inp[5]) ? 3'b110 : 3'b111;
									assign node625 = (inp[1]) ? node637 : node626;
										assign node626 = (inp[5]) ? node632 : node627;
											assign node627 = (inp[0]) ? 3'b100 : node628;
												assign node628 = (inp[2]) ? 3'b100 : 3'b110;
											assign node632 = (inp[2]) ? 3'b101 : node633;
												assign node633 = (inp[0]) ? 3'b101 : 3'b111;
										assign node637 = (inp[5]) ? 3'b001 : 3'b000;
							assign node640 = (inp[5]) ? node660 : node641;
								assign node641 = (inp[11]) ? node649 : node642;
									assign node642 = (inp[1]) ? node644 : 3'b100;
										assign node644 = (inp[8]) ? node646 : 3'b100;
											assign node646 = (inp[0]) ? 3'b000 : 3'b100;
									assign node649 = (inp[8]) ? node655 : node650;
										assign node650 = (inp[1]) ? 3'b010 : node651;
											assign node651 = (inp[2]) ? 3'b010 : 3'b100;
										assign node655 = (inp[2]) ? 3'b100 : node656;
											assign node656 = (inp[1]) ? 3'b100 : 3'b000;
								assign node660 = (inp[11]) ? node662 : 3'b000;
									assign node662 = (inp[8]) ? node672 : node663;
										assign node663 = (inp[0]) ? node665 : 3'b010;
											assign node665 = (inp[1]) ? node669 : node666;
												assign node666 = (inp[2]) ? 3'b010 : 3'b100;
												assign node669 = (inp[2]) ? 3'b100 : 3'b010;
										assign node672 = (inp[0]) ? node678 : node673;
											assign node673 = (inp[1]) ? node675 : 3'b100;
												assign node675 = (inp[2]) ? 3'b000 : 3'b100;
											assign node678 = (inp[1]) ? 3'b100 : node679;
												assign node679 = (inp[2]) ? 3'b100 : 3'b000;
					assign node683 = (inp[4]) ? node739 : node684;
						assign node684 = (inp[3]) ? node686 : 3'b100;
							assign node686 = (inp[8]) ? node712 : node687;
								assign node687 = (inp[11]) ? node697 : node688;
									assign node688 = (inp[1]) ? node690 : 3'b101;
										assign node690 = (inp[0]) ? node694 : node691;
											assign node691 = (inp[5]) ? 3'b101 : 3'b001;
											assign node694 = (inp[5]) ? 3'b001 : 3'b101;
									assign node697 = (inp[0]) ? node703 : node698;
										assign node698 = (inp[5]) ? node700 : 3'b101;
											assign node700 = (inp[2]) ? 3'b001 : 3'b011;
										assign node703 = (inp[5]) ? node707 : node704;
											assign node704 = (inp[2]) ? 3'b011 : 3'b001;
											assign node707 = (inp[2]) ? 3'b001 : node708;
												assign node708 = (inp[1]) ? 3'b111 : 3'b011;
								assign node712 = (inp[11]) ? node724 : node713;
									assign node713 = (inp[5]) ? node717 : node714;
										assign node714 = (inp[2]) ? 3'b001 : 3'b101;
										assign node717 = (inp[2]) ? node719 : 3'b010;
											assign node719 = (inp[1]) ? node721 : 3'b010;
												assign node721 = (inp[0]) ? 3'b110 : 3'b010;
									assign node724 = (inp[5]) ? node732 : node725;
										assign node725 = (inp[2]) ? node727 : 3'b011;
											assign node727 = (inp[1]) ? node729 : 3'b111;
												assign node729 = (inp[0]) ? 3'b101 : 3'b111;
										assign node732 = (inp[0]) ? node734 : 3'b101;
											assign node734 = (inp[1]) ? node736 : 3'b101;
												assign node736 = (inp[2]) ? 3'b001 : 3'b101;
						assign node739 = (inp[3]) ? node789 : node740;
							assign node740 = (inp[1]) ? node764 : node741;
								assign node741 = (inp[8]) ? node753 : node742;
									assign node742 = (inp[11]) ? node750 : node743;
										assign node743 = (inp[2]) ? 3'b111 : node744;
											assign node744 = (inp[5]) ? node746 : 3'b111;
												assign node746 = (inp[0]) ? 3'b011 : 3'b111;
										assign node750 = (inp[0]) ? 3'b111 : 3'b001;
									assign node753 = (inp[11]) ? node759 : node754;
										assign node754 = (inp[2]) ? 3'b011 : node755;
											assign node755 = (inp[5]) ? 3'b101 : 3'b011;
										assign node759 = (inp[0]) ? node761 : 3'b111;
											assign node761 = (inp[5]) ? 3'b011 : 3'b111;
								assign node764 = (inp[8]) ? node778 : node765;
									assign node765 = (inp[11]) ? node773 : node766;
										assign node766 = (inp[2]) ? 3'b011 : node767;
											assign node767 = (inp[0]) ? node769 : 3'b111;
												assign node769 = (inp[5]) ? 3'b011 : 3'b111;
										assign node773 = (inp[5]) ? node775 : 3'b001;
											assign node775 = (inp[0]) ? 3'b111 : 3'b001;
									assign node778 = (inp[11]) ? node784 : node779;
										assign node779 = (inp[2]) ? 3'b101 : node780;
											assign node780 = (inp[5]) ? 3'b101 : 3'b011;
										assign node784 = (inp[5]) ? node786 : 3'b111;
											assign node786 = (inp[0]) ? 3'b011 : 3'b111;
							assign node789 = (inp[11]) ? node801 : node790;
								assign node790 = (inp[8]) ? node796 : node791;
									assign node791 = (inp[0]) ? node793 : 3'b110;
										assign node793 = (inp[5]) ? 3'b010 : 3'b110;
									assign node796 = (inp[0]) ? node798 : 3'b010;
										assign node798 = (inp[5]) ? 3'b100 : 3'b010;
								assign node801 = (inp[8]) ? node811 : node802;
									assign node802 = (inp[5]) ? node804 : 3'b001;
										assign node804 = (inp[0]) ? node806 : 3'b001;
											assign node806 = (inp[2]) ? 3'b110 : node807;
												assign node807 = (inp[1]) ? 3'b110 : 3'b001;
									assign node811 = (inp[5]) ? node819 : node812;
										assign node812 = (inp[2]) ? node816 : node813;
											assign node813 = (inp[0]) ? 3'b101 : 3'b001;
											assign node816 = (inp[0]) ? 3'b110 : 3'b010;
										assign node819 = (inp[1]) ? node821 : 3'b110;
											assign node821 = (inp[0]) ? 3'b010 : 3'b110;
		assign node824 = (inp[9]) ? node1004 : node825;
			assign node825 = (inp[3]) ? 3'b000 : node826;
				assign node826 = (inp[7]) ? node958 : node827;
					assign node827 = (inp[10]) ? node867 : node828;
						assign node828 = (inp[4]) ? 3'b000 : node829;
							assign node829 = (inp[11]) ? node841 : node830;
								assign node830 = (inp[8]) ? 3'b000 : node831;
									assign node831 = (inp[5]) ? node833 : 3'b100;
										assign node833 = (inp[0]) ? node835 : 3'b100;
											assign node835 = (inp[1]) ? 3'b000 : node836;
												assign node836 = (inp[2]) ? 3'b000 : 3'b100;
								assign node841 = (inp[8]) ? node851 : node842;
									assign node842 = (inp[0]) ? node846 : node843;
										assign node843 = (inp[5]) ? 3'b010 : 3'b110;
										assign node846 = (inp[1]) ? node848 : 3'b010;
											assign node848 = (inp[5]) ? 3'b100 : 3'b010;
									assign node851 = (inp[5]) ? node859 : node852;
										assign node852 = (inp[2]) ? node854 : 3'b010;
											assign node854 = (inp[0]) ? node856 : 3'b110;
												assign node856 = (inp[1]) ? 3'b100 : 3'b110;
										assign node859 = (inp[1]) ? node861 : 3'b100;
											assign node861 = (inp[2]) ? node863 : 3'b100;
												assign node863 = (inp[0]) ? 3'b000 : 3'b100;
						assign node867 = (inp[4]) ? node923 : node868;
							assign node868 = (inp[11]) ? node890 : node869;
								assign node869 = (inp[8]) ? node879 : node870;
									assign node870 = (inp[0]) ? node874 : node871;
										assign node871 = (inp[5]) ? 3'b110 : 3'b010;
										assign node874 = (inp[5]) ? node876 : 3'b110;
											assign node876 = (inp[1]) ? 3'b010 : 3'b110;
									assign node879 = (inp[5]) ? node883 : node880;
										assign node880 = (inp[2]) ? 3'b010 : 3'b110;
										assign node883 = (inp[1]) ? node885 : 3'b000;
											assign node885 = (inp[2]) ? node887 : 3'b000;
												assign node887 = (inp[0]) ? 3'b100 : 3'b000;
								assign node890 = (inp[5]) ? node906 : node891;
									assign node891 = (inp[2]) ? node897 : node892;
										assign node892 = (inp[8]) ? 3'b001 : node893;
											assign node893 = (inp[0]) ? 3'b011 : 3'b111;
										assign node897 = (inp[1]) ? node903 : node898;
											assign node898 = (inp[0]) ? node900 : 3'b111;
												assign node900 = (inp[8]) ? 3'b101 : 3'b001;
											assign node903 = (inp[0]) ? 3'b110 : 3'b101;
									assign node906 = (inp[8]) ? node918 : node907;
										assign node907 = (inp[2]) ? node913 : node908;
											assign node908 = (inp[1]) ? node910 : 3'b001;
												assign node910 = (inp[0]) ? 3'b100 : 3'b001;
											assign node913 = (inp[1]) ? node915 : 3'b011;
												assign node915 = (inp[0]) ? 3'b110 : 3'b011;
										assign node918 = (inp[2]) ? node920 : 3'b110;
											assign node920 = (inp[0]) ? 3'b010 : 3'b110;
							assign node923 = (inp[11]) ? node931 : node924;
								assign node924 = (inp[8]) ? 3'b000 : node925;
									assign node925 = (inp[5]) ? node927 : 3'b100;
										assign node927 = (inp[0]) ? 3'b000 : 3'b100;
								assign node931 = (inp[5]) ? node945 : node932;
									assign node932 = (inp[0]) ? node938 : node933;
										assign node933 = (inp[2]) ? 3'b110 : node934;
											assign node934 = (inp[8]) ? 3'b010 : 3'b110;
										assign node938 = (inp[2]) ? node940 : 3'b010;
											assign node940 = (inp[8]) ? node942 : 3'b010;
												assign node942 = (inp[1]) ? 3'b100 : 3'b110;
									assign node945 = (inp[8]) ? node951 : node946;
										assign node946 = (inp[0]) ? node948 : 3'b010;
											assign node948 = (inp[1]) ? 3'b100 : 3'b010;
										assign node951 = (inp[0]) ? node953 : 3'b100;
											assign node953 = (inp[1]) ? node955 : 3'b100;
												assign node955 = (inp[2]) ? 3'b000 : 3'b100;
					assign node958 = (inp[10]) ? node960 : 3'b000;
						assign node960 = (inp[4]) ? 3'b000 : node961;
							assign node961 = (inp[11]) ? node973 : node962;
								assign node962 = (inp[8]) ? 3'b000 : node963;
									assign node963 = (inp[0]) ? node965 : 3'b100;
										assign node965 = (inp[5]) ? node967 : 3'b100;
											assign node967 = (inp[1]) ? 3'b000 : node968;
												assign node968 = (inp[2]) ? 3'b000 : 3'b100;
								assign node973 = (inp[8]) ? node987 : node974;
									assign node974 = (inp[1]) ? node980 : node975;
										assign node975 = (inp[5]) ? 3'b010 : node976;
											assign node976 = (inp[0]) ? 3'b010 : 3'b110;
										assign node980 = (inp[0]) ? node984 : node981;
											assign node981 = (inp[5]) ? 3'b010 : 3'b110;
											assign node984 = (inp[5]) ? 3'b100 : 3'b010;
									assign node987 = (inp[5]) ? node995 : node988;
										assign node988 = (inp[2]) ? node990 : 3'b010;
											assign node990 = (inp[0]) ? node992 : 3'b110;
												assign node992 = (inp[1]) ? 3'b100 : 3'b110;
										assign node995 = (inp[1]) ? node997 : 3'b100;
											assign node997 = (inp[2]) ? node999 : 3'b100;
												assign node999 = (inp[0]) ? 3'b000 : 3'b100;
			assign node1004 = (inp[3]) ? node1272 : node1005;
				assign node1005 = (inp[4]) ? node1125 : node1006;
					assign node1006 = (inp[7]) ? node1038 : node1007;
						assign node1007 = (inp[10]) ? 3'b011 : node1008;
							assign node1008 = (inp[5]) ? node1030 : node1009;
								assign node1009 = (inp[8]) ? node1017 : node1010;
									assign node1010 = (inp[2]) ? node1012 : 3'b001;
										assign node1012 = (inp[11]) ? node1014 : 3'b001;
											assign node1014 = (inp[0]) ? 3'b011 : 3'b001;
									assign node1017 = (inp[11]) ? node1023 : node1018;
										assign node1018 = (inp[1]) ? node1020 : 3'b001;
											assign node1020 = (inp[0]) ? 3'b011 : 3'b001;
										assign node1023 = (inp[2]) ? node1025 : 3'b011;
											assign node1025 = (inp[1]) ? node1027 : 3'b011;
												assign node1027 = (inp[0]) ? 3'b001 : 3'b011;
								assign node1030 = (inp[11]) ? node1032 : 3'b011;
									assign node1032 = (inp[2]) ? 3'b001 : node1033;
										assign node1033 = (inp[8]) ? 3'b001 : 3'b011;
						assign node1038 = (inp[10]) ? node1106 : node1039;
							assign node1039 = (inp[11]) ? node1073 : node1040;
								assign node1040 = (inp[8]) ? node1062 : node1041;
									assign node1041 = (inp[1]) ? node1047 : node1042;
										assign node1042 = (inp[0]) ? 3'b110 : node1043;
											assign node1043 = (inp[5]) ? 3'b110 : 3'b010;
										assign node1047 = (inp[2]) ? node1055 : node1048;
											assign node1048 = (inp[5]) ? node1052 : node1049;
												assign node1049 = (inp[0]) ? 3'b110 : 3'b010;
												assign node1052 = (inp[0]) ? 3'b010 : 3'b110;
											assign node1055 = (inp[0]) ? node1059 : node1056;
												assign node1056 = (inp[5]) ? 3'b110 : 3'b010;
												assign node1059 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1062 = (inp[5]) ? node1066 : node1063;
										assign node1063 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1066 = (inp[2]) ? node1068 : 3'b000;
											assign node1068 = (inp[1]) ? node1070 : 3'b000;
												assign node1070 = (inp[0]) ? 3'b100 : 3'b000;
								assign node1073 = (inp[5]) ? node1087 : node1074;
									assign node1074 = (inp[0]) ? node1078 : node1075;
										assign node1075 = (inp[8]) ? 3'b101 : 3'b111;
										assign node1078 = (inp[2]) ? node1082 : node1079;
											assign node1079 = (inp[8]) ? 3'b001 : 3'b011;
											assign node1082 = (inp[8]) ? node1084 : 3'b001;
												assign node1084 = (inp[1]) ? 3'b110 : 3'b101;
									assign node1087 = (inp[8]) ? node1099 : node1088;
										assign node1088 = (inp[2]) ? node1094 : node1089;
											assign node1089 = (inp[0]) ? node1091 : 3'b001;
												assign node1091 = (inp[1]) ? 3'b100 : 3'b001;
											assign node1094 = (inp[0]) ? node1096 : 3'b011;
												assign node1096 = (inp[1]) ? 3'b110 : 3'b011;
										assign node1099 = (inp[2]) ? node1101 : 3'b110;
											assign node1101 = (inp[1]) ? node1103 : 3'b110;
												assign node1103 = (inp[0]) ? 3'b010 : 3'b110;
							assign node1106 = (inp[5]) ? node1116 : node1107;
								assign node1107 = (inp[11]) ? node1109 : 3'b001;
									assign node1109 = (inp[1]) ? node1111 : 3'b011;
										assign node1111 = (inp[8]) ? node1113 : 3'b011;
											assign node1113 = (inp[0]) ? 3'b101 : 3'b111;
								assign node1116 = (inp[11]) ? node1120 : node1117;
									assign node1117 = (inp[8]) ? 3'b110 : 3'b111;
									assign node1120 = (inp[1]) ? node1122 : 3'b101;
										assign node1122 = (inp[8]) ? 3'b001 : 3'b101;
					assign node1125 = (inp[10]) ? node1185 : node1126;
						assign node1126 = (inp[5]) ? node1156 : node1127;
							assign node1127 = (inp[8]) ? node1139 : node1128;
								assign node1128 = (inp[11]) ? node1130 : 3'b010;
									assign node1130 = (inp[7]) ? 3'b010 : node1131;
										assign node1131 = (inp[0]) ? 3'b110 : node1132;
											assign node1132 = (inp[2]) ? 3'b110 : node1133;
												assign node1133 = (inp[1]) ? 3'b110 : 3'b001;
								assign node1139 = (inp[11]) ? node1147 : node1140;
									assign node1140 = (inp[7]) ? node1142 : 3'b100;
										assign node1142 = (inp[1]) ? node1144 : 3'b010;
											assign node1144 = (inp[0]) ? 3'b000 : 3'b010;
									assign node1147 = (inp[7]) ? node1151 : node1148;
										assign node1148 = (inp[1]) ? 3'b010 : 3'b110;
										assign node1151 = (inp[1]) ? node1153 : 3'b110;
											assign node1153 = (inp[0]) ? 3'b100 : 3'b110;
							assign node1156 = (inp[7]) ? node1176 : node1157;
								assign node1157 = (inp[8]) ? node1167 : node1158;
									assign node1158 = (inp[11]) ? node1160 : 3'b010;
										assign node1160 = (inp[2]) ? 3'b110 : node1161;
											assign node1161 = (inp[0]) ? 3'b110 : node1162;
												assign node1162 = (inp[1]) ? 3'b110 : 3'b001;
									assign node1167 = (inp[11]) ? node1169 : 3'b100;
										assign node1169 = (inp[1]) ? 3'b010 : node1170;
											assign node1170 = (inp[2]) ? 3'b110 : node1171;
												assign node1171 = (inp[0]) ? 3'b110 : 3'b101;
								assign node1176 = (inp[11]) ? node1178 : 3'b000;
									assign node1178 = (inp[8]) ? node1182 : node1179;
										assign node1179 = (inp[0]) ? 3'b100 : 3'b000;
										assign node1182 = (inp[0]) ? 3'b000 : 3'b100;
						assign node1185 = (inp[7]) ? node1229 : node1186;
							assign node1186 = (inp[8]) ? node1208 : node1187;
								assign node1187 = (inp[11]) ? node1203 : node1188;
									assign node1188 = (inp[1]) ? node1196 : node1189;
										assign node1189 = (inp[2]) ? 3'b101 : node1190;
											assign node1190 = (inp[0]) ? node1192 : 3'b101;
												assign node1192 = (inp[5]) ? 3'b001 : 3'b101;
										assign node1196 = (inp[2]) ? 3'b001 : node1197;
											assign node1197 = (inp[0]) ? node1199 : 3'b101;
												assign node1199 = (inp[5]) ? 3'b001 : 3'b101;
									assign node1203 = (inp[0]) ? node1205 : 3'b011;
										assign node1205 = (inp[5]) ? 3'b101 : 3'b011;
								assign node1208 = (inp[11]) ? node1224 : node1209;
									assign node1209 = (inp[1]) ? node1217 : node1210;
										assign node1210 = (inp[0]) ? node1212 : 3'b001;
											assign node1212 = (inp[5]) ? node1214 : 3'b001;
												assign node1214 = (inp[2]) ? 3'b001 : 3'b110;
										assign node1217 = (inp[2]) ? 3'b110 : node1218;
											assign node1218 = (inp[5]) ? node1220 : 3'b001;
												assign node1220 = (inp[0]) ? 3'b110 : 3'b001;
									assign node1224 = (inp[0]) ? node1226 : 3'b101;
										assign node1226 = (inp[5]) ? 3'b001 : 3'b101;
							assign node1229 = (inp[11]) ? node1249 : node1230;
								assign node1230 = (inp[0]) ? node1236 : node1231;
									assign node1231 = (inp[5]) ? node1233 : 3'b110;
										assign node1233 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1236 = (inp[8]) ? node1244 : node1237;
										assign node1237 = (inp[5]) ? node1239 : 3'b110;
											assign node1239 = (inp[1]) ? 3'b010 : node1240;
												assign node1240 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1244 = (inp[1]) ? node1246 : 3'b010;
											assign node1246 = (inp[5]) ? 3'b100 : 3'b010;
								assign node1249 = (inp[5]) ? node1259 : node1250;
									assign node1250 = (inp[0]) ? node1252 : 3'b001;
										assign node1252 = (inp[2]) ? node1254 : 3'b001;
											assign node1254 = (inp[1]) ? node1256 : 3'b001;
												assign node1256 = (inp[8]) ? 3'b110 : 3'b001;
									assign node1259 = (inp[8]) ? node1265 : node1260;
										assign node1260 = (inp[1]) ? node1262 : 3'b101;
											assign node1262 = (inp[0]) ? 3'b110 : 3'b101;
										assign node1265 = (inp[2]) ? node1267 : 3'b110;
											assign node1267 = (inp[0]) ? node1269 : 3'b110;
												assign node1269 = (inp[1]) ? 3'b010 : 3'b110;
				assign node1272 = (inp[10]) ? node1308 : node1273;
					assign node1273 = (inp[4]) ? 3'b000 : node1274;
						assign node1274 = (inp[7]) ? 3'b000 : node1275;
							assign node1275 = (inp[11]) ? node1283 : node1276;
								assign node1276 = (inp[8]) ? 3'b000 : node1277;
									assign node1277 = (inp[5]) ? node1279 : 3'b100;
										assign node1279 = (inp[0]) ? 3'b000 : 3'b100;
								assign node1283 = (inp[8]) ? node1293 : node1284;
									assign node1284 = (inp[0]) ? node1288 : node1285;
										assign node1285 = (inp[5]) ? 3'b010 : 3'b110;
										assign node1288 = (inp[5]) ? node1290 : 3'b010;
											assign node1290 = (inp[1]) ? 3'b100 : 3'b010;
									assign node1293 = (inp[5]) ? node1301 : node1294;
										assign node1294 = (inp[2]) ? node1296 : 3'b010;
											assign node1296 = (inp[0]) ? node1298 : 3'b110;
												assign node1298 = (inp[1]) ? 3'b100 : 3'b110;
										assign node1301 = (inp[1]) ? node1303 : 3'b100;
											assign node1303 = (inp[0]) ? 3'b000 : 3'b100;
					assign node1308 = (inp[4]) ? node1412 : node1309;
						assign node1309 = (inp[7]) ? node1375 : node1310;
							assign node1310 = (inp[11]) ? node1342 : node1311;
								assign node1311 = (inp[8]) ? node1331 : node1312;
									assign node1312 = (inp[1]) ? node1318 : node1313;
										assign node1313 = (inp[5]) ? 3'b110 : node1314;
											assign node1314 = (inp[0]) ? 3'b110 : 3'b010;
										assign node1318 = (inp[2]) ? node1324 : node1319;
											assign node1319 = (inp[5]) ? node1321 : 3'b010;
												assign node1321 = (inp[0]) ? 3'b010 : 3'b110;
											assign node1324 = (inp[0]) ? node1328 : node1325;
												assign node1325 = (inp[5]) ? 3'b110 : 3'b010;
												assign node1328 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1331 = (inp[5]) ? node1335 : node1332;
										assign node1332 = (inp[2]) ? 3'b010 : 3'b110;
										assign node1335 = (inp[2]) ? node1337 : 3'b000;
											assign node1337 = (inp[1]) ? node1339 : 3'b000;
												assign node1339 = (inp[0]) ? 3'b100 : 3'b000;
								assign node1342 = (inp[5]) ? node1356 : node1343;
									assign node1343 = (inp[8]) ? node1349 : node1344;
										assign node1344 = (inp[0]) ? node1346 : 3'b111;
											assign node1346 = (inp[2]) ? 3'b001 : 3'b011;
										assign node1349 = (inp[2]) ? node1351 : 3'b001;
											assign node1351 = (inp[0]) ? node1353 : 3'b101;
												assign node1353 = (inp[1]) ? 3'b110 : 3'b101;
									assign node1356 = (inp[8]) ? node1368 : node1357;
										assign node1357 = (inp[2]) ? node1363 : node1358;
											assign node1358 = (inp[0]) ? node1360 : 3'b001;
												assign node1360 = (inp[1]) ? 3'b100 : 3'b001;
											assign node1363 = (inp[1]) ? node1365 : 3'b011;
												assign node1365 = (inp[0]) ? 3'b110 : 3'b011;
										assign node1368 = (inp[1]) ? node1370 : 3'b110;
											assign node1370 = (inp[2]) ? node1372 : 3'b110;
												assign node1372 = (inp[0]) ? 3'b010 : 3'b110;
							assign node1375 = (inp[11]) ? node1385 : node1376;
								assign node1376 = (inp[5]) ? 3'b000 : node1377;
									assign node1377 = (inp[1]) ? node1379 : 3'b100;
										assign node1379 = (inp[8]) ? node1381 : 3'b100;
											assign node1381 = (inp[0]) ? 3'b000 : 3'b100;
								assign node1385 = (inp[5]) ? node1399 : node1386;
									assign node1386 = (inp[8]) ? node1392 : node1387;
										assign node1387 = (inp[2]) ? node1389 : 3'b110;
											assign node1389 = (inp[0]) ? 3'b010 : 3'b110;
										assign node1392 = (inp[0]) ? node1394 : 3'b010;
											assign node1394 = (inp[1]) ? node1396 : 3'b010;
												assign node1396 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1399 = (inp[8]) ? 3'b100 : node1400;
										assign node1400 = (inp[2]) ? node1406 : node1401;
											assign node1401 = (inp[0]) ? node1403 : 3'b010;
												assign node1403 = (inp[1]) ? 3'b000 : 3'b010;
											assign node1406 = (inp[1]) ? node1408 : 3'b110;
												assign node1408 = (inp[0]) ? 3'b100 : 3'b110;
						assign node1412 = (inp[7]) ? node1444 : node1413;
							assign node1413 = (inp[11]) ? node1425 : node1414;
								assign node1414 = (inp[8]) ? 3'b000 : node1415;
									assign node1415 = (inp[5]) ? node1417 : 3'b100;
										assign node1417 = (inp[0]) ? node1419 : 3'b100;
											assign node1419 = (inp[1]) ? 3'b000 : node1420;
												assign node1420 = (inp[2]) ? 3'b000 : 3'b100;
								assign node1425 = (inp[5]) ? node1433 : node1426;
									assign node1426 = (inp[0]) ? 3'b010 : node1427;
										assign node1427 = (inp[2]) ? 3'b110 : node1428;
											assign node1428 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1433 = (inp[8]) ? node1439 : node1434;
										assign node1434 = (inp[1]) ? node1436 : 3'b010;
											assign node1436 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1439 = (inp[1]) ? node1441 : 3'b100;
											assign node1441 = (inp[2]) ? 3'b000 : 3'b100;
							assign node1444 = (inp[8]) ? 3'b000 : node1445;
								assign node1445 = (inp[5]) ? 3'b000 : node1446;
									assign node1446 = (inp[2]) ? 3'b000 : node1447;
										assign node1447 = (inp[11]) ? 3'b100 : 3'b000;

endmodule