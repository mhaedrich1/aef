module dtc_split5_bm98 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node290;
	wire [3-1:0] node294;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node316;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node323;
	wire [3-1:0] node327;
	wire [3-1:0] node329;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node359;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node378;
	wire [3-1:0] node380;
	wire [3-1:0] node384;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node397;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node405;
	wire [3-1:0] node407;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node425;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node448;
	wire [3-1:0] node450;
	wire [3-1:0] node452;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node468;
	wire [3-1:0] node470;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node481;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node488;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node504;
	wire [3-1:0] node506;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node513;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node520;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node538;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node581;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node624;

	assign outp = (inp[0]) ? node226 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b111;
			assign node3 = (inp[3]) ? node153 : node4;
				assign node4 = (inp[9]) ? node44 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b100;
						assign node7 = (inp[7]) ? node11 : node8;
							assign node8 = (inp[1]) ? 3'b000 : 3'b100;
							assign node11 = (inp[1]) ? node25 : node12;
								assign node12 = (inp[2]) ? node18 : node13;
									assign node13 = (inp[10]) ? node15 : 3'b000;
										assign node15 = (inp[5]) ? 3'b000 : 3'b100;
									assign node18 = (inp[10]) ? node20 : 3'b100;
										assign node20 = (inp[11]) ? node22 : 3'b100;
											assign node22 = (inp[5]) ? 3'b100 : 3'b000;
								assign node25 = (inp[8]) ? node37 : node26;
									assign node26 = (inp[10]) ? node32 : node27;
										assign node27 = (inp[2]) ? 3'b100 : node28;
											assign node28 = (inp[5]) ? 3'b100 : 3'b101;
										assign node32 = (inp[2]) ? 3'b101 : node33;
											assign node33 = (inp[5]) ? 3'b100 : 3'b100;
									assign node37 = (inp[11]) ? node39 : 3'b100;
										assign node39 = (inp[5]) ? node41 : 3'b100;
											assign node41 = (inp[2]) ? 3'b100 : 3'b100;
					assign node44 = (inp[1]) ? node92 : node45;
						assign node45 = (inp[4]) ? node61 : node46;
							assign node46 = (inp[2]) ? node56 : node47;
								assign node47 = (inp[7]) ? 3'b001 : node48;
									assign node48 = (inp[8]) ? node50 : 3'b101;
										assign node50 = (inp[10]) ? 3'b001 : node51;
											assign node51 = (inp[5]) ? 3'b101 : 3'b001;
								assign node56 = (inp[5]) ? 3'b101 : node57;
									assign node57 = (inp[11]) ? 3'b101 : 3'b001;
							assign node61 = (inp[7]) ? node77 : node62;
								assign node62 = (inp[8]) ? node72 : node63;
									assign node63 = (inp[10]) ? node67 : node64;
										assign node64 = (inp[2]) ? 3'b001 : 3'b111;
										assign node67 = (inp[11]) ? node69 : 3'b101;
											assign node69 = (inp[2]) ? 3'b111 : 3'b101;
									assign node72 = (inp[2]) ? node74 : 3'b101;
										assign node74 = (inp[5]) ? 3'b101 : 3'b111;
								assign node77 = (inp[2]) ? node85 : node78;
									assign node78 = (inp[11]) ? node82 : node79;
										assign node79 = (inp[5]) ? 3'b111 : 3'b011;
										assign node82 = (inp[5]) ? 3'b011 : 3'b111;
									assign node85 = (inp[11]) ? node89 : node86;
										assign node86 = (inp[8]) ? 3'b101 : 3'b001;
										assign node89 = (inp[8]) ? 3'b001 : 3'b101;
						assign node92 = (inp[4]) ? node112 : node93;
							assign node93 = (inp[2]) ? node105 : node94;
								assign node94 = (inp[7]) ? 3'b001 : node95;
									assign node95 = (inp[8]) ? node97 : 3'b100;
										assign node97 = (inp[5]) ? node101 : node98;
											assign node98 = (inp[11]) ? 3'b100 : 3'b001;
											assign node101 = (inp[11]) ? 3'b001 : 3'b100;
								assign node105 = (inp[5]) ? node107 : 3'b100;
									assign node107 = (inp[11]) ? node109 : 3'b100;
										assign node109 = (inp[7]) ? 3'b100 : 3'b001;
							assign node112 = (inp[7]) ? node134 : node113;
								assign node113 = (inp[2]) ? node125 : node114;
									assign node114 = (inp[11]) ? node120 : node115;
										assign node115 = (inp[8]) ? node117 : 3'b110;
											assign node117 = (inp[10]) ? 3'b110 : 3'b100;
										assign node120 = (inp[5]) ? node122 : 3'b100;
											assign node122 = (inp[8]) ? 3'b110 : 3'b100;
									assign node125 = (inp[11]) ? node127 : 3'b100;
										assign node127 = (inp[5]) ? node131 : node128;
											assign node128 = (inp[10]) ? 3'b001 : 3'b010;
											assign node131 = (inp[10]) ? 3'b110 : 3'b100;
								assign node134 = (inp[8]) ? node144 : node135;
									assign node135 = (inp[11]) ? node141 : node136;
										assign node136 = (inp[2]) ? 3'b001 : node137;
											assign node137 = (inp[5]) ? 3'b110 : 3'b001;
										assign node141 = (inp[2]) ? 3'b110 : 3'b001;
									assign node144 = (inp[11]) ? node150 : node145;
										assign node145 = (inp[2]) ? 3'b110 : node146;
											assign node146 = (inp[5]) ? 3'b110 : 3'b001;
										assign node150 = (inp[5]) ? 3'b001 : 3'b110;
				assign node153 = (inp[9]) ? node173 : node154;
					assign node154 = (inp[4]) ? node156 : 3'b010;
						assign node156 = (inp[1]) ? node158 : 3'b010;
							assign node158 = (inp[7]) ? node160 : 3'b010;
								assign node160 = (inp[2]) ? node166 : node161;
									assign node161 = (inp[5]) ? node163 : 3'b110;
										assign node163 = (inp[8]) ? 3'b010 : 3'b110;
									assign node166 = (inp[10]) ? node168 : 3'b010;
										assign node168 = (inp[8]) ? node170 : 3'b110;
											assign node170 = (inp[5]) ? 3'b010 : 3'b010;
					assign node173 = (inp[1]) ? node175 : 3'b111;
						assign node175 = (inp[7]) ? node197 : node176;
							assign node176 = (inp[4]) ? node190 : node177;
								assign node177 = (inp[2]) ? node185 : node178;
									assign node178 = (inp[11]) ? node182 : node179;
										assign node179 = (inp[8]) ? 3'b111 : 3'b011;
										assign node182 = (inp[5]) ? 3'b111 : 3'b011;
									assign node185 = (inp[5]) ? 3'b011 : node186;
										assign node186 = (inp[11]) ? 3'b011 : 3'b111;
								assign node190 = (inp[2]) ? node192 : 3'b001;
									assign node192 = (inp[8]) ? node194 : 3'b001;
										assign node194 = (inp[10]) ? 3'b111 : 3'b011;
							assign node197 = (inp[2]) ? node213 : node198;
								assign node198 = (inp[4]) ? node200 : 3'b101;
									assign node200 = (inp[10]) ? node206 : node201;
										assign node201 = (inp[5]) ? node203 : 3'b011;
											assign node203 = (inp[11]) ? 3'b111 : 3'b011;
										assign node206 = (inp[5]) ? node210 : node207;
											assign node207 = (inp[11]) ? 3'b011 : 3'b111;
											assign node210 = (inp[11]) ? 3'b111 : 3'b011;
								assign node213 = (inp[4]) ? node215 : 3'b001;
									assign node215 = (inp[11]) ? node221 : node216;
										assign node216 = (inp[8]) ? node218 : 3'b101;
											assign node218 = (inp[10]) ? 3'b001 : 3'b001;
										assign node221 = (inp[5]) ? 3'b011 : node222;
											assign node222 = (inp[10]) ? 3'b101 : 3'b001;
		assign node226 = (inp[3]) ? node366 : node227;
			assign node227 = (inp[6]) ? node327 : node228;
				assign node228 = (inp[9]) ? node252 : node229;
					assign node229 = (inp[4]) ? node231 : 3'b010;
						assign node231 = (inp[7]) ? node235 : node232;
							assign node232 = (inp[1]) ? 3'b000 : 3'b010;
							assign node235 = (inp[1]) ? 3'b010 : node236;
								assign node236 = (inp[2]) ? node244 : node237;
									assign node237 = (inp[10]) ? node239 : 3'b000;
										assign node239 = (inp[8]) ? node241 : 3'b010;
											assign node241 = (inp[5]) ? 3'b010 : 3'b000;
									assign node244 = (inp[5]) ? node246 : 3'b010;
										assign node246 = (inp[8]) ? 3'b010 : node247;
											assign node247 = (inp[10]) ? 3'b000 : 3'b000;
					assign node252 = (inp[2]) ? node284 : node253;
						assign node253 = (inp[4]) ? node263 : node254;
							assign node254 = (inp[7]) ? 3'b000 : node255;
								assign node255 = (inp[11]) ? node259 : node256;
									assign node256 = (inp[5]) ? 3'b010 : 3'b000;
									assign node259 = (inp[5]) ? 3'b000 : 3'b010;
							assign node263 = (inp[7]) ? node265 : 3'b010;
								assign node265 = (inp[1]) ? node275 : node266;
									assign node266 = (inp[8]) ? 3'b010 : node267;
										assign node267 = (inp[5]) ? node271 : node268;
											assign node268 = (inp[11]) ? 3'b010 : 3'b000;
											assign node271 = (inp[10]) ? 3'b000 : 3'b010;
									assign node275 = (inp[10]) ? node277 : 3'b000;
										assign node277 = (inp[11]) ? node281 : node278;
											assign node278 = (inp[5]) ? 3'b010 : 3'b000;
											assign node281 = (inp[5]) ? 3'b000 : 3'b010;
						assign node284 = (inp[7]) ? node310 : node285;
							assign node285 = (inp[5]) ? node299 : node286;
								assign node286 = (inp[11]) ? node294 : node287;
									assign node287 = (inp[10]) ? 3'b000 : node288;
										assign node288 = (inp[4]) ? node290 : 3'b000;
											assign node290 = (inp[8]) ? 3'b010 : 3'b000;
									assign node294 = (inp[4]) ? node296 : 3'b010;
										assign node296 = (inp[1]) ? 3'b010 : 3'b000;
								assign node299 = (inp[11]) ? node307 : node300;
									assign node300 = (inp[4]) ? node302 : 3'b010;
										assign node302 = (inp[10]) ? 3'b010 : node303;
											assign node303 = (inp[8]) ? 3'b010 : 3'b000;
									assign node307 = (inp[4]) ? 3'b010 : 3'b000;
							assign node310 = (inp[4]) ? node312 : 3'b010;
								assign node312 = (inp[1]) ? node320 : node313;
									assign node313 = (inp[10]) ? 3'b010 : node314;
										assign node314 = (inp[5]) ? node316 : 3'b000;
											assign node316 = (inp[11]) ? 3'b000 : 3'b010;
									assign node320 = (inp[11]) ? 3'b110 : node321;
										assign node321 = (inp[8]) ? node323 : 3'b100;
											assign node323 = (inp[5]) ? 3'b100 : 3'b010;
				assign node327 = (inp[4]) ? node329 : 3'b000;
					assign node329 = (inp[9]) ? node331 : 3'b000;
						assign node331 = (inp[1]) ? node363 : node332;
							assign node332 = (inp[11]) ? node348 : node333;
								assign node333 = (inp[10]) ? node343 : node334;
									assign node334 = (inp[5]) ? node338 : node335;
										assign node335 = (inp[2]) ? 3'b110 : 3'b010;
										assign node338 = (inp[8]) ? 3'b110 : node339;
											assign node339 = (inp[2]) ? 3'b010 : 3'b110;
									assign node343 = (inp[2]) ? 3'b010 : node344;
										assign node344 = (inp[5]) ? 3'b100 : 3'b010;
								assign node348 = (inp[2]) ? node356 : node349;
									assign node349 = (inp[5]) ? node353 : node350;
										assign node350 = (inp[10]) ? 3'b100 : 3'b110;
										assign node353 = (inp[10]) ? 3'b010 : 3'b000;
									assign node356 = (inp[7]) ? 3'b100 : node357;
										assign node357 = (inp[8]) ? node359 : 3'b100;
											assign node359 = (inp[5]) ? 3'b100 : 3'b000;
							assign node363 = (inp[7]) ? 3'b000 : 3'b100;
			assign node366 = (inp[9]) ? node456 : node367;
				assign node367 = (inp[4]) ? node373 : node368;
					assign node368 = (inp[6]) ? 3'b000 : node369;
						assign node369 = (inp[1]) ? 3'b000 : 3'b001;
					assign node373 = (inp[7]) ? node411 : node374;
						assign node374 = (inp[1]) ? node392 : node375;
							assign node375 = (inp[6]) ? 3'b001 : node376;
								assign node376 = (inp[2]) ? node384 : node377;
									assign node377 = (inp[11]) ? 3'b011 : node378;
										assign node378 = (inp[8]) ? node380 : 3'b111;
											assign node380 = (inp[10]) ? 3'b111 : 3'b011;
									assign node384 = (inp[5]) ? node386 : 3'b101;
										assign node386 = (inp[10]) ? 3'b011 : node387;
											assign node387 = (inp[8]) ? 3'b101 : 3'b001;
							assign node392 = (inp[6]) ? 3'b100 : node393;
								assign node393 = (inp[11]) ? node401 : node394;
									assign node394 = (inp[2]) ? 3'b001 : node395;
										assign node395 = (inp[8]) ? node397 : 3'b101;
											assign node397 = (inp[10]) ? 3'b101 : 3'b001;
									assign node401 = (inp[2]) ? node405 : node402;
										assign node402 = (inp[8]) ? 3'b101 : 3'b001;
										assign node405 = (inp[8]) ? node407 : 3'b110;
											assign node407 = (inp[10]) ? 3'b001 : 3'b110;
						assign node411 = (inp[1]) ? node433 : node412;
							assign node412 = (inp[6]) ? node416 : node413;
								assign node413 = (inp[2]) ? 3'b001 : 3'b101;
								assign node416 = (inp[10]) ? node428 : node417;
									assign node417 = (inp[2]) ? node423 : node418;
										assign node418 = (inp[11]) ? node420 : 3'b100;
											assign node420 = (inp[5]) ? 3'b010 : 3'b100;
										assign node423 = (inp[11]) ? node425 : 3'b000;
											assign node425 = (inp[5]) ? 3'b110 : 3'b010;
									assign node428 = (inp[5]) ? 3'b010 : node429;
										assign node429 = (inp[2]) ? 3'b110 : 3'b010;
							assign node433 = (inp[6]) ? 3'b000 : node434;
								assign node434 = (inp[2]) ? node448 : node435;
									assign node435 = (inp[10]) ? node443 : node436;
										assign node436 = (inp[5]) ? node440 : node437;
											assign node437 = (inp[11]) ? 3'b110 : 3'b010;
											assign node440 = (inp[11]) ? 3'b010 : 3'b110;
										assign node443 = (inp[8]) ? 3'b010 : node444;
											assign node444 = (inp[5]) ? 3'b010 : 3'b010;
									assign node448 = (inp[11]) ? node450 : 3'b010;
										assign node450 = (inp[8]) ? node452 : 3'b100;
											assign node452 = (inp[10]) ? 3'b000 : 3'b000;
				assign node456 = (inp[6]) ? node524 : node457;
					assign node457 = (inp[1]) ? node459 : 3'b111;
						assign node459 = (inp[4]) ? node497 : node460;
							assign node460 = (inp[11]) ? node484 : node461;
								assign node461 = (inp[8]) ? node473 : node462;
									assign node462 = (inp[7]) ? node468 : node463;
										assign node463 = (inp[10]) ? 3'b010 : node464;
											assign node464 = (inp[2]) ? 3'b110 : 3'b010;
										assign node468 = (inp[5]) ? node470 : 3'b110;
											assign node470 = (inp[2]) ? 3'b110 : 3'b010;
									assign node473 = (inp[5]) ? node479 : node474;
										assign node474 = (inp[10]) ? node476 : 3'b001;
											assign node476 = (inp[2]) ? 3'b001 : 3'b001;
										assign node479 = (inp[10]) ? node481 : 3'b001;
											assign node481 = (inp[7]) ? 3'b010 : 3'b110;
								assign node484 = (inp[8]) ? node492 : node485;
									assign node485 = (inp[5]) ? 3'b001 : node486;
										assign node486 = (inp[2]) ? node488 : 3'b001;
											assign node488 = (inp[10]) ? 3'b001 : 3'b101;
									assign node492 = (inp[10]) ? node494 : 3'b001;
										assign node494 = (inp[5]) ? 3'b001 : 3'b010;
							assign node497 = (inp[7]) ? node509 : node498;
								assign node498 = (inp[5]) ? node504 : node499;
									assign node499 = (inp[11]) ? 3'b111 : node500;
										assign node500 = (inp[8]) ? 3'b111 : 3'b011;
									assign node504 = (inp[11]) ? node506 : 3'b011;
										assign node506 = (inp[10]) ? 3'b111 : 3'b011;
								assign node509 = (inp[2]) ? node517 : node510;
									assign node510 = (inp[8]) ? 3'b001 : node511;
										assign node511 = (inp[11]) ? node513 : 3'b001;
											assign node513 = (inp[5]) ? 3'b011 : 3'b001;
									assign node517 = (inp[8]) ? 3'b101 : node518;
										assign node518 = (inp[10]) ? node520 : 3'b101;
											assign node520 = (inp[11]) ? 3'b011 : 3'b001;
					assign node524 = (inp[1]) ? node586 : node525;
						assign node525 = (inp[7]) ? node559 : node526;
							assign node526 = (inp[4]) ? node550 : node527;
								assign node527 = (inp[2]) ? node541 : node528;
									assign node528 = (inp[8]) ? node534 : node529;
										assign node529 = (inp[5]) ? 3'b001 : node530;
											assign node530 = (inp[11]) ? 3'b001 : 3'b101;
										assign node534 = (inp[5]) ? node538 : node535;
											assign node535 = (inp[11]) ? 3'b001 : 3'b101;
											assign node538 = (inp[11]) ? 3'b101 : 3'b001;
									assign node541 = (inp[10]) ? 3'b101 : node542;
										assign node542 = (inp[8]) ? node546 : node543;
											assign node543 = (inp[11]) ? 3'b101 : 3'b001;
											assign node546 = (inp[5]) ? 3'b101 : 3'b001;
								assign node550 = (inp[2]) ? node552 : 3'b010;
									assign node552 = (inp[8]) ? node556 : node553;
										assign node553 = (inp[10]) ? 3'b010 : 3'b101;
										assign node556 = (inp[10]) ? 3'b101 : 3'b001;
							assign node559 = (inp[4]) ? node563 : node560;
								assign node560 = (inp[2]) ? 3'b010 : 3'b110;
								assign node563 = (inp[2]) ? node575 : node564;
									assign node564 = (inp[8]) ? node570 : node565;
										assign node565 = (inp[10]) ? 3'b001 : node566;
											assign node566 = (inp[5]) ? 3'b001 : 3'b101;
										assign node570 = (inp[11]) ? 3'b101 : node571;
											assign node571 = (inp[10]) ? 3'b101 : 3'b001;
									assign node575 = (inp[11]) ? node581 : node576;
										assign node576 = (inp[10]) ? 3'b110 : node577;
											assign node577 = (inp[8]) ? 3'b010 : 3'b110;
										assign node581 = (inp[8]) ? node583 : 3'b001;
											assign node583 = (inp[5]) ? 3'b000 : 3'b110;
						assign node586 = (inp[7]) ? node608 : node587;
							assign node587 = (inp[4]) ? node595 : node588;
								assign node588 = (inp[5]) ? node592 : node589;
									assign node589 = (inp[11]) ? 3'b010 : 3'b110;
									assign node592 = (inp[11]) ? 3'b110 : 3'b010;
								assign node595 = (inp[2]) ? node601 : node596;
									assign node596 = (inp[10]) ? node598 : 3'b000;
										assign node598 = (inp[8]) ? 3'b000 : 3'b001;
									assign node601 = (inp[8]) ? node605 : node602;
										assign node602 = (inp[10]) ? 3'b001 : 3'b110;
										assign node605 = (inp[10]) ? 3'b110 : 3'b010;
							assign node608 = (inp[2]) ? node616 : node609;
								assign node609 = (inp[4]) ? node611 : 3'b100;
									assign node611 = (inp[5]) ? node613 : 3'b110;
										assign node613 = (inp[11]) ? 3'b110 : 3'b010;
								assign node616 = (inp[4]) ? node618 : 3'b000;
									assign node618 = (inp[11]) ? node622 : node619;
										assign node619 = (inp[8]) ? 3'b000 : 3'b100;
										assign node622 = (inp[8]) ? node624 : 3'b010;
											assign node624 = (inp[5]) ? 3'b100 : 3'b000;

endmodule