module dtc_split875_bm51 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node5;
	wire [2-1:0] node7;
	wire [2-1:0] node9;
	wire [2-1:0] node12;
	wire [2-1:0] node13;
	wire [2-1:0] node15;
	wire [2-1:0] node18;
	wire [2-1:0] node20;
	wire [2-1:0] node23;
	wire [2-1:0] node24;
	wire [2-1:0] node25;
	wire [2-1:0] node29;
	wire [2-1:0] node30;
	wire [2-1:0] node33;
	wire [2-1:0] node34;
	wire [2-1:0] node38;
	wire [2-1:0] node39;
	wire [2-1:0] node40;
	wire [2-1:0] node43;
	wire [2-1:0] node46;
	wire [2-1:0] node47;
	wire [2-1:0] node50;
	wire [2-1:0] node53;
	wire [2-1:0] node54;
	wire [2-1:0] node55;
	wire [2-1:0] node56;
	wire [2-1:0] node59;
	wire [2-1:0] node62;
	wire [2-1:0] node63;
	wire [2-1:0] node66;
	wire [2-1:0] node69;
	wire [2-1:0] node70;
	wire [2-1:0] node71;
	wire [2-1:0] node75;
	wire [2-1:0] node76;
	wire [2-1:0] node80;
	wire [2-1:0] node81;
	wire [2-1:0] node82;
	wire [2-1:0] node83;
	wire [2-1:0] node84;
	wire [2-1:0] node86;
	wire [2-1:0] node89;
	wire [2-1:0] node90;
	wire [2-1:0] node93;
	wire [2-1:0] node96;
	wire [2-1:0] node97;
	wire [2-1:0] node98;
	wire [2-1:0] node99;
	wire [2-1:0] node104;
	wire [2-1:0] node107;
	wire [2-1:0] node108;
	wire [2-1:0] node109;
	wire [2-1:0] node113;
	wire [2-1:0] node114;
	wire [2-1:0] node118;
	wire [2-1:0] node119;
	wire [2-1:0] node120;
	wire [2-1:0] node121;
	wire [2-1:0] node122;
	wire [2-1:0] node123;
	wire [2-1:0] node127;
	wire [2-1:0] node128;
	wire [2-1:0] node133;
	wire [2-1:0] node134;
	wire [2-1:0] node135;
	wire [2-1:0] node136;
	wire [2-1:0] node140;
	wire [2-1:0] node141;
	wire [2-1:0] node146;
	wire [2-1:0] node147;

	assign outp = (inp[6]) ? node80 : node1;
		assign node1 = (inp[2]) ? node53 : node2;
			assign node2 = (inp[0]) ? node38 : node3;
				assign node3 = (inp[7]) ? node23 : node4;
					assign node4 = (inp[4]) ? node12 : node5;
						assign node5 = (inp[5]) ? node7 : 2'b00;
							assign node7 = (inp[3]) ? node9 : 2'b01;
								assign node9 = (inp[1]) ? 2'b00 : 2'b01;
						assign node12 = (inp[5]) ? node18 : node13;
							assign node13 = (inp[3]) ? node15 : 2'b01;
								assign node15 = (inp[1]) ? 2'b00 : 2'b01;
							assign node18 = (inp[1]) ? node20 : 2'b00;
								assign node20 = (inp[3]) ? 2'b01 : 2'b00;
					assign node23 = (inp[5]) ? node29 : node24;
						assign node24 = (inp[4]) ? 2'b11 : node25;
							assign node25 = (inp[3]) ? 2'b10 : 2'b11;
						assign node29 = (inp[4]) ? node33 : node30;
							assign node30 = (inp[3]) ? 2'b11 : 2'b10;
							assign node33 = (inp[3]) ? 2'b10 : node34;
								assign node34 = (inp[1]) ? 2'b11 : 2'b10;
				assign node38 = (inp[1]) ? node46 : node39;
					assign node39 = (inp[5]) ? node43 : node40;
						assign node40 = (inp[3]) ? 2'b11 : 2'b10;
						assign node43 = (inp[3]) ? 2'b10 : 2'b11;
					assign node46 = (inp[3]) ? node50 : node47;
						assign node47 = (inp[5]) ? 2'b11 : 2'b10;
						assign node50 = (inp[5]) ? 2'b10 : 2'b11;
			assign node53 = (inp[0]) ? node69 : node54;
				assign node54 = (inp[7]) ? node62 : node55;
					assign node55 = (inp[1]) ? node59 : node56;
						assign node56 = (inp[4]) ? 2'b11 : 2'b10;
						assign node59 = (inp[4]) ? 2'b10 : 2'b11;
					assign node62 = (inp[3]) ? node66 : node63;
						assign node63 = (inp[4]) ? 2'b01 : 2'b00;
						assign node66 = (inp[4]) ? 2'b00 : 2'b01;
				assign node69 = (inp[3]) ? node75 : node70;
					assign node70 = (inp[1]) ? 2'b01 : node71;
						assign node71 = (inp[7]) ? 2'b01 : 2'b00;
					assign node75 = (inp[7]) ? 2'b00 : node76;
						assign node76 = (inp[1]) ? 2'b00 : 2'b01;
		assign node80 = (inp[7]) ? node118 : node81;
			assign node81 = (inp[0]) ? node107 : node82;
				assign node82 = (inp[5]) ? node96 : node83;
					assign node83 = (inp[4]) ? node89 : node84;
						assign node84 = (inp[1]) ? node86 : 2'b10;
							assign node86 = (inp[2]) ? 2'b11 : 2'b10;
						assign node89 = (inp[1]) ? node93 : node90;
							assign node90 = (inp[2]) ? 2'b11 : 2'b10;
							assign node93 = (inp[2]) ? 2'b10 : 2'b11;
					assign node96 = (inp[4]) ? node104 : node97;
						assign node97 = (inp[1]) ? 2'b11 : node98;
							assign node98 = (inp[2]) ? 2'b10 : node99;
								assign node99 = (inp[3]) ? 2'b10 : 2'b11;
						assign node104 = (inp[1]) ? 2'b10 : 2'b11;
				assign node107 = (inp[1]) ? node113 : node108;
					assign node108 = (inp[2]) ? 2'b01 : node109;
						assign node109 = (inp[5]) ? 2'b01 : 2'b00;
					assign node113 = (inp[5]) ? 2'b00 : node114;
						assign node114 = (inp[2]) ? 2'b00 : 2'b01;
			assign node118 = (inp[2]) ? node146 : node119;
				assign node119 = (inp[5]) ? node133 : node120;
					assign node120 = (inp[0]) ? 2'b01 : node121;
						assign node121 = (inp[4]) ? node127 : node122;
							assign node122 = (inp[3]) ? 2'b00 : node123;
								assign node123 = (inp[1]) ? 2'b00 : 2'b01;
							assign node127 = (inp[1]) ? 2'b01 : node128;
								assign node128 = (inp[3]) ? 2'b01 : 2'b00;
					assign node133 = (inp[0]) ? 2'b00 : node134;
						assign node134 = (inp[4]) ? node140 : node135;
							assign node135 = (inp[3]) ? 2'b01 : node136;
								assign node136 = (inp[1]) ? 2'b01 : 2'b00;
							assign node140 = (inp[1]) ? 2'b00 : node141;
								assign node141 = (inp[3]) ? 2'b00 : 2'b01;
				assign node146 = (inp[4]) ? 2'b00 : node147;
					assign node147 = (inp[0]) ? 2'b00 : 2'b01;

endmodule