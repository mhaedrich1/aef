module dtc_split66_bm77 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node262;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node275;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node332;
	wire [3-1:0] node333;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node384;
	wire [3-1:0] node387;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node410;
	wire [3-1:0] node411;
	wire [3-1:0] node412;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node460;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node465;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node471;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node495;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node502;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node512;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node519;
	wire [3-1:0] node522;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node532;
	wire [3-1:0] node534;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node541;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node613;
	wire [3-1:0] node615;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node626;
	wire [3-1:0] node628;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node637;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node644;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node658;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node664;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node671;
	wire [3-1:0] node673;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node680;
	wire [3-1:0] node681;
	wire [3-1:0] node682;
	wire [3-1:0] node684;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node714;
	wire [3-1:0] node717;
	wire [3-1:0] node718;
	wire [3-1:0] node719;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node758;
	wire [3-1:0] node761;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node809;
	wire [3-1:0] node811;
	wire [3-1:0] node813;
	wire [3-1:0] node815;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node825;
	wire [3-1:0] node826;
	wire [3-1:0] node828;
	wire [3-1:0] node832;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node837;
	wire [3-1:0] node840;

	assign outp = (inp[3]) ? node108 : node1;
		assign node1 = (inp[4]) ? node3 : 3'b000;
			assign node3 = (inp[6]) ? 3'b000 : node4;
				assign node4 = (inp[0]) ? node6 : 3'b000;
					assign node6 = (inp[7]) ? node90 : node7;
						assign node7 = (inp[5]) ? node45 : node8;
							assign node8 = (inp[9]) ? node22 : node9;
								assign node9 = (inp[8]) ? node17 : node10;
									assign node10 = (inp[11]) ? node14 : node11;
										assign node11 = (inp[10]) ? 3'b000 : 3'b100;
										assign node14 = (inp[10]) ? 3'b100 : 3'b000;
									assign node17 = (inp[11]) ? node19 : 3'b100;
										assign node19 = (inp[10]) ? 3'b000 : 3'b100;
								assign node22 = (inp[1]) ? node24 : 3'b000;
									assign node24 = (inp[2]) ? node34 : node25;
										assign node25 = (inp[10]) ? 3'b100 : node26;
											assign node26 = (inp[11]) ? node30 : node27;
												assign node27 = (inp[8]) ? 3'b100 : 3'b000;
												assign node30 = (inp[8]) ? 3'b000 : 3'b100;
										assign node34 = (inp[11]) ? node42 : node35;
											assign node35 = (inp[10]) ? node39 : node36;
												assign node36 = (inp[8]) ? 3'b000 : 3'b100;
												assign node39 = (inp[8]) ? 3'b100 : 3'b010;
											assign node42 = (inp[8]) ? 3'b010 : 3'b110;
							assign node45 = (inp[1]) ? node65 : node46;
								assign node46 = (inp[10]) ? node54 : node47;
									assign node47 = (inp[8]) ? 3'b000 : node48;
										assign node48 = (inp[2]) ? 3'b100 : node49;
											assign node49 = (inp[11]) ? 3'b000 : 3'b100;
									assign node54 = (inp[8]) ? node60 : node55;
										assign node55 = (inp[9]) ? node57 : 3'b010;
											assign node57 = (inp[11]) ? 3'b010 : 3'b000;
										assign node60 = (inp[11]) ? 3'b100 : node61;
											assign node61 = (inp[9]) ? 3'b000 : 3'b100;
								assign node65 = (inp[10]) ? node77 : node66;
									assign node66 = (inp[9]) ? node70 : node67;
										assign node67 = (inp[8]) ? 3'b000 : 3'b100;
										assign node70 = (inp[2]) ? node74 : node71;
											assign node71 = (inp[8]) ? 3'b100 : 3'b010;
											assign node74 = (inp[8]) ? 3'b010 : 3'b110;
									assign node77 = (inp[2]) ? node83 : node78;
										assign node78 = (inp[9]) ? node80 : 3'b010;
											assign node80 = (inp[8]) ? 3'b010 : 3'b110;
										assign node83 = (inp[8]) ? node87 : node84;
											assign node84 = (inp[9]) ? 3'b001 : 3'b010;
											assign node87 = (inp[11]) ? 3'b100 : 3'b110;
						assign node90 = (inp[1]) ? node92 : 3'b000;
							assign node92 = (inp[9]) ? node94 : 3'b000;
								assign node94 = (inp[2]) ? node96 : 3'b000;
									assign node96 = (inp[11]) ? node100 : node97;
										assign node97 = (inp[8]) ? 3'b000 : 3'b010;
										assign node100 = (inp[5]) ? node102 : 3'b000;
											assign node102 = (inp[8]) ? 3'b100 : node103;
												assign node103 = (inp[10]) ? 3'b010 : 3'b100;
		assign node108 = (inp[0]) ? node284 : node109;
			assign node109 = (inp[6]) ? node267 : node110;
				assign node110 = (inp[4]) ? node142 : node111;
					assign node111 = (inp[7]) ? 3'b000 : node112;
						assign node112 = (inp[5]) ? node114 : 3'b000;
							assign node114 = (inp[9]) ? node116 : 3'b000;
								assign node116 = (inp[1]) ? node124 : node117;
									assign node117 = (inp[10]) ? node119 : 3'b000;
										assign node119 = (inp[8]) ? 3'b000 : node120;
											assign node120 = (inp[2]) ? 3'b100 : 3'b000;
									assign node124 = (inp[10]) ? node134 : node125;
										assign node125 = (inp[8]) ? node131 : node126;
											assign node126 = (inp[2]) ? node128 : 3'b100;
												assign node128 = (inp[11]) ? 3'b010 : 3'b100;
											assign node131 = (inp[11]) ? 3'b100 : 3'b000;
										assign node134 = (inp[8]) ? node136 : 3'b010;
											assign node136 = (inp[11]) ? 3'b010 : node137;
												assign node137 = (inp[2]) ? 3'b100 : 3'b000;
					assign node142 = (inp[1]) ? node192 : node143;
						assign node143 = (inp[7]) ? node181 : node144;
							assign node144 = (inp[9]) ? node154 : node145;
								assign node145 = (inp[2]) ? node147 : 3'b000;
									assign node147 = (inp[10]) ? node149 : 3'b000;
										assign node149 = (inp[8]) ? 3'b000 : node150;
											assign node150 = (inp[5]) ? 3'b100 : 3'b000;
								assign node154 = (inp[2]) ? node170 : node155;
									assign node155 = (inp[10]) ? node161 : node156;
										assign node156 = (inp[8]) ? 3'b000 : node157;
											assign node157 = (inp[5]) ? 3'b100 : 3'b000;
										assign node161 = (inp[5]) ? node167 : node162;
											assign node162 = (inp[8]) ? 3'b000 : node163;
												assign node163 = (inp[11]) ? 3'b100 : 3'b000;
											assign node167 = (inp[8]) ? 3'b100 : 3'b010;
									assign node170 = (inp[5]) ? node176 : node171;
										assign node171 = (inp[10]) ? node173 : 3'b000;
											assign node173 = (inp[8]) ? 3'b000 : 3'b010;
										assign node176 = (inp[11]) ? 3'b010 : node177;
											assign node177 = (inp[8]) ? 3'b010 : 3'b110;
							assign node181 = (inp[10]) ? node183 : 3'b000;
								assign node183 = (inp[9]) ? node185 : 3'b000;
									assign node185 = (inp[8]) ? 3'b000 : node186;
										assign node186 = (inp[2]) ? node188 : 3'b000;
											assign node188 = (inp[5]) ? 3'b100 : 3'b000;
						assign node192 = (inp[7]) ? node236 : node193;
							assign node193 = (inp[9]) ? node203 : node194;
								assign node194 = (inp[10]) ? node196 : 3'b100;
									assign node196 = (inp[8]) ? 3'b100 : node197;
										assign node197 = (inp[2]) ? 3'b110 : node198;
											assign node198 = (inp[5]) ? 3'b110 : 3'b100;
								assign node203 = (inp[5]) ? node221 : node204;
									assign node204 = (inp[11]) ? node216 : node205;
										assign node205 = (inp[10]) ? node213 : node206;
											assign node206 = (inp[8]) ? node210 : node207;
												assign node207 = (inp[2]) ? 3'b110 : 3'b010;
												assign node210 = (inp[2]) ? 3'b010 : 3'b000;
											assign node213 = (inp[2]) ? 3'b001 : 3'b100;
										assign node216 = (inp[10]) ? node218 : 3'b010;
											assign node218 = (inp[2]) ? 3'b110 : 3'b010;
									assign node221 = (inp[2]) ? node229 : node222;
										assign node222 = (inp[11]) ? node226 : node223;
											assign node223 = (inp[8]) ? 3'b010 : 3'b110;
											assign node226 = (inp[10]) ? 3'b110 : 3'b001;
										assign node229 = (inp[11]) ? node231 : 3'b001;
											assign node231 = (inp[10]) ? node233 : 3'b101;
												assign node233 = (inp[8]) ? 3'b101 : 3'b011;
							assign node236 = (inp[9]) ? node238 : 3'b000;
								assign node238 = (inp[5]) ? node254 : node239;
									assign node239 = (inp[2]) ? node241 : 3'b000;
										assign node241 = (inp[8]) ? node249 : node242;
											assign node242 = (inp[11]) ? node246 : node243;
												assign node243 = (inp[10]) ? 3'b100 : 3'b000;
												assign node246 = (inp[10]) ? 3'b010 : 3'b100;
											assign node249 = (inp[11]) ? node251 : 3'b000;
												assign node251 = (inp[10]) ? 3'b100 : 3'b000;
									assign node254 = (inp[10]) ? node262 : node255;
										assign node255 = (inp[11]) ? 3'b100 : node256;
											assign node256 = (inp[8]) ? node258 : 3'b010;
												assign node258 = (inp[2]) ? 3'b100 : 3'b000;
										assign node262 = (inp[11]) ? node264 : 3'b010;
											assign node264 = (inp[2]) ? 3'b110 : 3'b010;
				assign node267 = (inp[1]) ? node269 : 3'b000;
					assign node269 = (inp[5]) ? node271 : 3'b000;
						assign node271 = (inp[10]) ? node273 : 3'b000;
							assign node273 = (inp[4]) ? node275 : 3'b000;
								assign node275 = (inp[9]) ? node277 : 3'b000;
									assign node277 = (inp[8]) ? 3'b000 : node278;
										assign node278 = (inp[2]) ? node280 : 3'b000;
											assign node280 = (inp[7]) ? 3'b000 : 3'b100;
			assign node284 = (inp[6]) ? node676 : node285;
				assign node285 = (inp[7]) ? node507 : node286;
					assign node286 = (inp[4]) ? node390 : node287;
						assign node287 = (inp[11]) ? node339 : node288;
							assign node288 = (inp[9]) ? node304 : node289;
								assign node289 = (inp[5]) ? node297 : node290;
									assign node290 = (inp[8]) ? node294 : node291;
										assign node291 = (inp[10]) ? 3'b110 : 3'b001;
										assign node294 = (inp[10]) ? 3'b001 : 3'b010;
									assign node297 = (inp[10]) ? node301 : node298;
										assign node298 = (inp[8]) ? 3'b101 : 3'b010;
										assign node301 = (inp[8]) ? 3'b010 : 3'b101;
								assign node304 = (inp[1]) ? node316 : node305;
									assign node305 = (inp[8]) ? node313 : node306;
										assign node306 = (inp[2]) ? node308 : 3'b010;
											assign node308 = (inp[5]) ? 3'b110 : node309;
												assign node309 = (inp[10]) ? 3'b110 : 3'b010;
										assign node313 = (inp[2]) ? 3'b010 : 3'b100;
									assign node316 = (inp[10]) ? node324 : node317;
										assign node317 = (inp[5]) ? 3'b101 : node318;
											assign node318 = (inp[2]) ? 3'b110 : node319;
												assign node319 = (inp[8]) ? 3'b010 : 3'b110;
										assign node324 = (inp[5]) ? node332 : node325;
											assign node325 = (inp[8]) ? node329 : node326;
												assign node326 = (inp[2]) ? 3'b101 : 3'b001;
												assign node329 = (inp[2]) ? 3'b001 : 3'b110;
											assign node332 = (inp[2]) ? node336 : node333;
												assign node333 = (inp[8]) ? 3'b101 : 3'b011;
												assign node336 = (inp[8]) ? 3'b011 : 3'b111;
							assign node339 = (inp[8]) ? node365 : node340;
								assign node340 = (inp[5]) ? node352 : node341;
									assign node341 = (inp[10]) ? node349 : node342;
										assign node342 = (inp[9]) ? node344 : 3'b101;
											assign node344 = (inp[1]) ? node346 : 3'b100;
												assign node346 = (inp[2]) ? 3'b101 : 3'b001;
										assign node349 = (inp[9]) ? 3'b101 : 3'b001;
									assign node352 = (inp[10]) ? node358 : node353;
										assign node353 = (inp[9]) ? node355 : 3'b001;
											assign node355 = (inp[1]) ? 3'b011 : 3'b001;
										assign node358 = (inp[9]) ? node360 : 3'b101;
											assign node360 = (inp[1]) ? 3'b011 : node361;
												assign node361 = (inp[2]) ? 3'b101 : 3'b001;
								assign node365 = (inp[1]) ? node379 : node366;
									assign node366 = (inp[10]) ? node372 : node367;
										assign node367 = (inp[5]) ? 3'b110 : node368;
											assign node368 = (inp[9]) ? 3'b000 : 3'b010;
										assign node372 = (inp[9]) ? node376 : node373;
											assign node373 = (inp[5]) ? 3'b001 : 3'b101;
											assign node376 = (inp[2]) ? 3'b010 : 3'b110;
									assign node379 = (inp[5]) ? node381 : 3'b101;
										assign node381 = (inp[10]) ? node387 : node382;
											assign node382 = (inp[9]) ? node384 : 3'b110;
												assign node384 = (inp[2]) ? 3'b101 : 3'b001;
											assign node387 = (inp[9]) ? 3'b101 : 3'b001;
						assign node390 = (inp[1]) ? node460 : node391;
							assign node391 = (inp[9]) ? node421 : node392;
								assign node392 = (inp[11]) ? node406 : node393;
									assign node393 = (inp[2]) ? 3'b101 : node394;
										assign node394 = (inp[10]) ? node400 : node395;
											assign node395 = (inp[8]) ? 3'b101 : node396;
												assign node396 = (inp[5]) ? 3'b111 : 3'b101;
											assign node400 = (inp[8]) ? 3'b111 : node401;
												assign node401 = (inp[5]) ? 3'b101 : 3'b111;
									assign node406 = (inp[8]) ? node410 : node407;
										assign node407 = (inp[10]) ? 3'b101 : 3'b111;
										assign node410 = (inp[10]) ? node416 : node411;
											assign node411 = (inp[2]) ? 3'b101 : node412;
												assign node412 = (inp[5]) ? 3'b101 : 3'b111;
											assign node416 = (inp[5]) ? 3'b111 : node417;
												assign node417 = (inp[2]) ? 3'b111 : 3'b101;
								assign node421 = (inp[5]) ? node437 : node422;
									assign node422 = (inp[10]) ? node430 : node423;
										assign node423 = (inp[8]) ? node427 : node424;
											assign node424 = (inp[2]) ? 3'b011 : 3'b001;
											assign node427 = (inp[2]) ? 3'b001 : 3'b110;
										assign node430 = (inp[8]) ? node434 : node431;
											assign node431 = (inp[2]) ? 3'b011 : 3'b101;
											assign node434 = (inp[2]) ? 3'b101 : 3'b001;
									assign node437 = (inp[10]) ? node449 : node438;
										assign node438 = (inp[8]) ? node444 : node439;
											assign node439 = (inp[11]) ? node441 : 3'b101;
												assign node441 = (inp[2]) ? 3'b111 : 3'b011;
											assign node444 = (inp[11]) ? 3'b101 : node445;
												assign node445 = (inp[2]) ? 3'b101 : 3'b001;
										assign node449 = (inp[8]) ? node455 : node450;
											assign node450 = (inp[11]) ? 3'b111 : node451;
												assign node451 = (inp[2]) ? 3'b111 : 3'b011;
											assign node455 = (inp[11]) ? 3'b011 : node456;
												assign node456 = (inp[2]) ? 3'b011 : 3'b101;
							assign node460 = (inp[2]) ? node492 : node461;
								assign node461 = (inp[9]) ? node475 : node462;
									assign node462 = (inp[5]) ? node468 : node463;
										assign node463 = (inp[10]) ? node465 : 3'b011;
											assign node465 = (inp[11]) ? 3'b001 : 3'b011;
										assign node468 = (inp[11]) ? 3'b011 : node469;
											assign node469 = (inp[8]) ? node471 : 3'b001;
												assign node471 = (inp[10]) ? 3'b011 : 3'b001;
									assign node475 = (inp[11]) ? node487 : node476;
										assign node476 = (inp[8]) ? node482 : node477;
											assign node477 = (inp[10]) ? 3'b111 : node478;
												assign node478 = (inp[5]) ? 3'b111 : 3'b011;
											assign node482 = (inp[10]) ? node484 : 3'b011;
												assign node484 = (inp[5]) ? 3'b111 : 3'b011;
										assign node487 = (inp[8]) ? node489 : 3'b111;
											assign node489 = (inp[5]) ? 3'b111 : 3'b011;
								assign node492 = (inp[9]) ? node498 : node493;
									assign node493 = (inp[8]) ? node495 : 3'b111;
										assign node495 = (inp[5]) ? 3'b111 : 3'b101;
									assign node498 = (inp[10]) ? 3'b111 : node499;
										assign node499 = (inp[5]) ? 3'b111 : node500;
											assign node500 = (inp[8]) ? node502 : 3'b111;
												assign node502 = (inp[11]) ? 3'b111 : 3'b011;
					assign node507 = (inp[4]) ? node585 : node508;
						assign node508 = (inp[9]) ? node522 : node509;
							assign node509 = (inp[11]) ? node515 : node510;
								assign node510 = (inp[10]) ? node512 : 3'b110;
									assign node512 = (inp[8]) ? 3'b110 : 3'b010;
								assign node515 = (inp[8]) ? node519 : node516;
									assign node516 = (inp[10]) ? 3'b110 : 3'b010;
									assign node519 = (inp[10]) ? 3'b010 : 3'b110;
							assign node522 = (inp[10]) ? node552 : node523;
								assign node523 = (inp[1]) ? node537 : node524;
									assign node524 = (inp[2]) ? node532 : node525;
										assign node525 = (inp[5]) ? node527 : 3'b000;
											assign node527 = (inp[8]) ? 3'b100 : node528;
												assign node528 = (inp[11]) ? 3'b100 : 3'b000;
										assign node532 = (inp[11]) ? node534 : 3'b100;
											assign node534 = (inp[8]) ? 3'b110 : 3'b010;
									assign node537 = (inp[5]) ? node545 : node538;
										assign node538 = (inp[11]) ? 3'b100 : node539;
											assign node539 = (inp[8]) ? node541 : 3'b100;
												assign node541 = (inp[2]) ? 3'b100 : 3'b110;
										assign node545 = (inp[2]) ? node549 : node546;
											assign node546 = (inp[8]) ? 3'b100 : 3'b110;
											assign node549 = (inp[8]) ? 3'b110 : 3'b001;
								assign node552 = (inp[1]) ? node568 : node553;
									assign node553 = (inp[5]) ? node559 : node554;
										assign node554 = (inp[8]) ? node556 : 3'b000;
											assign node556 = (inp[2]) ? 3'b100 : 3'b000;
										assign node559 = (inp[8]) ? node561 : 3'b010;
											assign node561 = (inp[11]) ? node565 : node562;
												assign node562 = (inp[2]) ? 3'b100 : 3'b000;
												assign node565 = (inp[2]) ? 3'b010 : 3'b000;
									assign node568 = (inp[11]) ? node580 : node569;
										assign node569 = (inp[2]) ? node575 : node570;
											assign node570 = (inp[5]) ? 3'b010 : node571;
												assign node571 = (inp[8]) ? 3'b100 : 3'b010;
											assign node575 = (inp[5]) ? 3'b110 : node576;
												assign node576 = (inp[8]) ? 3'b010 : 3'b110;
										assign node580 = (inp[8]) ? 3'b010 : node581;
											assign node581 = (inp[5]) ? 3'b001 : 3'b010;
						assign node585 = (inp[5]) ? node631 : node586;
							assign node586 = (inp[9]) ? node602 : node587;
								assign node587 = (inp[10]) ? node595 : node588;
									assign node588 = (inp[11]) ? node592 : node589;
										assign node589 = (inp[8]) ? 3'b000 : 3'b010;
										assign node592 = (inp[8]) ? 3'b010 : 3'b110;
									assign node595 = (inp[8]) ? node599 : node596;
										assign node596 = (inp[11]) ? 3'b001 : 3'b100;
										assign node599 = (inp[11]) ? 3'b110 : 3'b010;
								assign node602 = (inp[1]) ? node618 : node603;
									assign node603 = (inp[2]) ? node609 : node604;
										assign node604 = (inp[8]) ? 3'b100 : node605;
											assign node605 = (inp[10]) ? 3'b110 : 3'b010;
										assign node609 = (inp[8]) ? node613 : node610;
											assign node610 = (inp[10]) ? 3'b001 : 3'b110;
											assign node613 = (inp[11]) ? node615 : 3'b100;
												assign node615 = (inp[10]) ? 3'b110 : 3'b010;
									assign node618 = (inp[2]) ? node626 : node619;
										assign node619 = (inp[8]) ? node621 : 3'b001;
											assign node621 = (inp[10]) ? 3'b001 : node622;
												assign node622 = (inp[11]) ? 3'b111 : 3'b110;
										assign node626 = (inp[8]) ? node628 : 3'b101;
											assign node628 = (inp[10]) ? 3'b101 : 3'b001;
							assign node631 = (inp[10]) ? node653 : node632;
								assign node632 = (inp[8]) ? node644 : node633;
									assign node633 = (inp[9]) ? node637 : node634;
										assign node634 = (inp[11]) ? 3'b101 : 3'b001;
										assign node637 = (inp[1]) ? node639 : 3'b101;
											assign node639 = (inp[11]) ? 3'b011 : node640;
												assign node640 = (inp[2]) ? 3'b011 : 3'b101;
									assign node644 = (inp[9]) ? node646 : 3'b010;
										assign node646 = (inp[1]) ? node650 : node647;
											assign node647 = (inp[11]) ? 3'b001 : 3'b000;
											assign node650 = (inp[2]) ? 3'b101 : 3'b001;
								assign node653 = (inp[9]) ? node661 : node654;
									assign node654 = (inp[11]) ? node658 : node655;
										assign node655 = (inp[8]) ? 3'b001 : 3'b101;
										assign node658 = (inp[8]) ? 3'b101 : 3'b011;
									assign node661 = (inp[2]) ? node667 : node662;
										assign node662 = (inp[1]) ? node664 : 3'b110;
											assign node664 = (inp[11]) ? 3'b011 : 3'b101;
										assign node667 = (inp[1]) ? node671 : node668;
											assign node668 = (inp[11]) ? 3'b011 : 3'b101;
											assign node671 = (inp[8]) ? node673 : 3'b111;
												assign node673 = (inp[11]) ? 3'b111 : 3'b011;
				assign node676 = (inp[4]) ? node698 : node677;
					assign node677 = (inp[8]) ? 3'b000 : node678;
						assign node678 = (inp[9]) ? node680 : 3'b000;
							assign node680 = (inp[7]) ? 3'b000 : node681;
								assign node681 = (inp[10]) ? node687 : node682;
									assign node682 = (inp[1]) ? node684 : 3'b000;
										assign node684 = (inp[2]) ? 3'b010 : 3'b000;
									assign node687 = (inp[2]) ? node693 : node688;
										assign node688 = (inp[5]) ? node690 : 3'b000;
											assign node690 = (inp[11]) ? 3'b100 : 3'b000;
										assign node693 = (inp[5]) ? 3'b110 : 3'b100;
					assign node698 = (inp[7]) ? node806 : node699;
						assign node699 = (inp[8]) ? node747 : node700;
							assign node700 = (inp[10]) ? node726 : node701;
								assign node701 = (inp[5]) ? node711 : node702;
									assign node702 = (inp[9]) ? node704 : 3'b100;
										assign node704 = (inp[1]) ? node708 : node705;
											assign node705 = (inp[11]) ? 3'b100 : 3'b000;
											assign node708 = (inp[2]) ? 3'b110 : 3'b010;
									assign node711 = (inp[2]) ? node717 : node712;
										assign node712 = (inp[11]) ? node714 : 3'b110;
											assign node714 = (inp[9]) ? 3'b100 : 3'b110;
										assign node717 = (inp[1]) ? node723 : node718;
											assign node718 = (inp[9]) ? 3'b010 : node719;
												assign node719 = (inp[11]) ? 3'b110 : 3'b010;
											assign node723 = (inp[9]) ? 3'b001 : 3'b010;
								assign node726 = (inp[5]) ? node736 : node727;
									assign node727 = (inp[9]) ? node729 : 3'b010;
										assign node729 = (inp[2]) ? node733 : node730;
											assign node730 = (inp[1]) ? 3'b010 : 3'b000;
											assign node733 = (inp[1]) ? 3'b001 : 3'b100;
									assign node736 = (inp[11]) ? node742 : node737;
										assign node737 = (inp[1]) ? node739 : 3'b010;
											assign node739 = (inp[9]) ? 3'b101 : 3'b110;
										assign node742 = (inp[9]) ? node744 : 3'b001;
											assign node744 = (inp[1]) ? 3'b101 : 3'b110;
							assign node747 = (inp[1]) ? node773 : node748;
								assign node748 = (inp[10]) ? node764 : node749;
									assign node749 = (inp[9]) ? node755 : node750;
										assign node750 = (inp[5]) ? 3'b100 : node751;
											assign node751 = (inp[11]) ? 3'b000 : 3'b110;
										assign node755 = (inp[2]) ? node761 : node756;
											assign node756 = (inp[11]) ? node758 : 3'b000;
												assign node758 = (inp[5]) ? 3'b000 : 3'b100;
											assign node761 = (inp[5]) ? 3'b100 : 3'b000;
									assign node764 = (inp[5]) ? node768 : node765;
										assign node765 = (inp[11]) ? 3'b100 : 3'b000;
										assign node768 = (inp[9]) ? node770 : 3'b010;
											assign node770 = (inp[2]) ? 3'b010 : 3'b100;
								assign node773 = (inp[9]) ? node783 : node774;
									assign node774 = (inp[5]) ? 3'b100 : node775;
										assign node775 = (inp[11]) ? node779 : node776;
											assign node776 = (inp[10]) ? 3'b000 : 3'b110;
											assign node779 = (inp[10]) ? 3'b100 : 3'b000;
									assign node783 = (inp[11]) ? node791 : node784;
										assign node784 = (inp[5]) ? node786 : 3'b100;
											assign node786 = (inp[2]) ? 3'b110 : node787;
												assign node787 = (inp[10]) ? 3'b110 : 3'b010;
										assign node791 = (inp[2]) ? node799 : node792;
											assign node792 = (inp[10]) ? node796 : node793;
												assign node793 = (inp[5]) ? 3'b010 : 3'b110;
												assign node796 = (inp[5]) ? 3'b110 : 3'b010;
											assign node799 = (inp[10]) ? node803 : node800;
												assign node800 = (inp[5]) ? 3'b110 : 3'b010;
												assign node803 = (inp[5]) ? 3'b001 : 3'b110;
						assign node806 = (inp[5]) ? node820 : node807;
							assign node807 = (inp[2]) ? node809 : 3'b000;
								assign node809 = (inp[9]) ? node811 : 3'b000;
									assign node811 = (inp[11]) ? node813 : 3'b000;
										assign node813 = (inp[8]) ? node815 : 3'b100;
											assign node815 = (inp[1]) ? node817 : 3'b000;
												assign node817 = (inp[10]) ? 3'b100 : 3'b000;
							assign node820 = (inp[8]) ? node832 : node821;
								assign node821 = (inp[9]) ? node825 : node822;
									assign node822 = (inp[10]) ? 3'b100 : 3'b000;
									assign node825 = (inp[1]) ? 3'b010 : node826;
										assign node826 = (inp[2]) ? node828 : 3'b000;
											assign node828 = (inp[10]) ? 3'b100 : 3'b000;
								assign node832 = (inp[9]) ? node834 : 3'b000;
									assign node834 = (inp[10]) ? node840 : node835;
										assign node835 = (inp[1]) ? node837 : 3'b000;
											assign node837 = (inp[2]) ? 3'b100 : 3'b000;
										assign node840 = (inp[11]) ? 3'b010 : 3'b000;

endmodule