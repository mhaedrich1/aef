module dtc_split75_bm63 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node13;
	wire [4-1:0] node15;
	wire [4-1:0] node16;
	wire [4-1:0] node19;
	wire [4-1:0] node22;
	wire [4-1:0] node23;
	wire [4-1:0] node26;
	wire [4-1:0] node29;
	wire [4-1:0] node30;
	wire [4-1:0] node32;
	wire [4-1:0] node35;
	wire [4-1:0] node36;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node42;
	wire [4-1:0] node43;
	wire [4-1:0] node46;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node51;
	wire [4-1:0] node54;
	wire [4-1:0] node57;
	wire [4-1:0] node59;
	wire [4-1:0] node62;
	wire [4-1:0] node63;
	wire [4-1:0] node64;
	wire [4-1:0] node67;
	wire [4-1:0] node70;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node76;
	wire [4-1:0] node80;
	wire [4-1:0] node81;
	wire [4-1:0] node82;
	wire [4-1:0] node84;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node92;
	wire [4-1:0] node93;
	wire [4-1:0] node94;
	wire [4-1:0] node98;
	wire [4-1:0] node99;
	wire [4-1:0] node102;
	wire [4-1:0] node105;
	wire [4-1:0] node106;
	wire [4-1:0] node107;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node113;
	wire [4-1:0] node116;
	wire [4-1:0] node117;
	wire [4-1:0] node120;
	wire [4-1:0] node123;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node129;
	wire [4-1:0] node133;
	wire [4-1:0] node135;
	wire [4-1:0] node136;
	wire [4-1:0] node139;
	wire [4-1:0] node142;
	wire [4-1:0] node143;
	wire [4-1:0] node144;
	wire [4-1:0] node145;
	wire [4-1:0] node146;
	wire [4-1:0] node147;
	wire [4-1:0] node149;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node157;
	wire [4-1:0] node158;
	wire [4-1:0] node160;
	wire [4-1:0] node163;
	wire [4-1:0] node165;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node170;
	wire [4-1:0] node172;
	wire [4-1:0] node175;
	wire [4-1:0] node176;
	wire [4-1:0] node180;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node186;
	wire [4-1:0] node189;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node192;
	wire [4-1:0] node194;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node202;
	wire [4-1:0] node204;
	wire [4-1:0] node207;
	wire [4-1:0] node208;
	wire [4-1:0] node209;
	wire [4-1:0] node212;
	wire [4-1:0] node215;
	wire [4-1:0] node217;
	wire [4-1:0] node218;
	wire [4-1:0] node221;
	wire [4-1:0] node224;
	wire [4-1:0] node225;
	wire [4-1:0] node226;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node230;
	wire [4-1:0] node233;
	wire [4-1:0] node235;
	wire [4-1:0] node238;
	wire [4-1:0] node239;
	wire [4-1:0] node242;
	wire [4-1:0] node245;
	wire [4-1:0] node246;
	wire [4-1:0] node247;
	wire [4-1:0] node249;
	wire [4-1:0] node252;
	wire [4-1:0] node254;
	wire [4-1:0] node257;
	wire [4-1:0] node258;
	wire [4-1:0] node260;
	wire [4-1:0] node263;
	wire [4-1:0] node266;
	wire [4-1:0] node267;
	wire [4-1:0] node268;
	wire [4-1:0] node269;
	wire [4-1:0] node273;
	wire [4-1:0] node274;
	wire [4-1:0] node276;
	wire [4-1:0] node279;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node287;
	wire [4-1:0] node289;
	wire [4-1:0] node292;
	wire [4-1:0] node293;
	wire [4-1:0] node295;
	wire [4-1:0] node298;
	wire [4-1:0] node300;
	wire [4-1:0] node303;
	wire [4-1:0] node304;
	wire [4-1:0] node305;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node310;
	wire [4-1:0] node313;
	wire [4-1:0] node315;
	wire [4-1:0] node318;
	wire [4-1:0] node319;
	wire [4-1:0] node321;
	wire [4-1:0] node324;
	wire [4-1:0] node326;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node331;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node337;
	wire [4-1:0] node340;
	wire [4-1:0] node341;
	wire [4-1:0] node344;
	wire [4-1:0] node347;
	wire [4-1:0] node348;
	wire [4-1:0] node349;
	wire [4-1:0] node350;
	wire [4-1:0] node353;
	wire [4-1:0] node356;
	wire [4-1:0] node357;
	wire [4-1:0] node360;
	wire [4-1:0] node363;
	wire [4-1:0] node364;
	wire [4-1:0] node365;
	wire [4-1:0] node369;
	wire [4-1:0] node371;
	wire [4-1:0] node374;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node377;
	wire [4-1:0] node379;
	wire [4-1:0] node380;
	wire [4-1:0] node384;
	wire [4-1:0] node385;
	wire [4-1:0] node387;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node395;
	wire [4-1:0] node398;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node416;
	wire [4-1:0] node419;
	wire [4-1:0] node421;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node427;
	wire [4-1:0] node430;
	wire [4-1:0] node431;
	wire [4-1:0] node432;
	wire [4-1:0] node435;
	wire [4-1:0] node439;
	wire [4-1:0] node440;
	wire [4-1:0] node441;
	wire [4-1:0] node442;
	wire [4-1:0] node443;
	wire [4-1:0] node445;
	wire [4-1:0] node448;
	wire [4-1:0] node450;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node456;
	wire [4-1:0] node457;
	wire [4-1:0] node460;
	wire [4-1:0] node463;
	wire [4-1:0] node464;
	wire [4-1:0] node465;
	wire [4-1:0] node468;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node475;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node483;
	wire [4-1:0] node487;
	wire [4-1:0] node489;
	wire [4-1:0] node492;
	wire [4-1:0] node493;
	wire [4-1:0] node494;
	wire [4-1:0] node497;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node503;
	wire [4-1:0] node506;
	wire [4-1:0] node507;
	wire [4-1:0] node510;
	wire [4-1:0] node513;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node522;
	wire [4-1:0] node524;
	wire [4-1:0] node527;
	wire [4-1:0] node528;
	wire [4-1:0] node529;
	wire [4-1:0] node533;
	wire [4-1:0] node536;
	wire [4-1:0] node537;
	wire [4-1:0] node538;
	wire [4-1:0] node539;
	wire [4-1:0] node544;
	wire [4-1:0] node545;
	wire [4-1:0] node549;
	wire [4-1:0] node550;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node556;
	wire [4-1:0] node559;
	wire [4-1:0] node560;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node569;
	wire [4-1:0] node570;
	wire [4-1:0] node571;
	wire [4-1:0] node573;
	wire [4-1:0] node576;
	wire [4-1:0] node579;
	wire [4-1:0] node581;
	wire [4-1:0] node584;
	wire [4-1:0] node585;
	wire [4-1:0] node586;
	wire [4-1:0] node587;
	wire [4-1:0] node588;
	wire [4-1:0] node589;
	wire [4-1:0] node590;
	wire [4-1:0] node593;
	wire [4-1:0] node595;
	wire [4-1:0] node598;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node604;
	wire [4-1:0] node607;
	wire [4-1:0] node608;
	wire [4-1:0] node612;
	wire [4-1:0] node614;
	wire [4-1:0] node617;
	wire [4-1:0] node618;
	wire [4-1:0] node619;
	wire [4-1:0] node621;
	wire [4-1:0] node622;
	wire [4-1:0] node625;
	wire [4-1:0] node628;
	wire [4-1:0] node630;
	wire [4-1:0] node631;
	wire [4-1:0] node635;
	wire [4-1:0] node636;
	wire [4-1:0] node638;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node645;
	wire [4-1:0] node648;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node653;
	wire [4-1:0] node655;
	wire [4-1:0] node658;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node665;
	wire [4-1:0] node666;
	wire [4-1:0] node668;
	wire [4-1:0] node671;
	wire [4-1:0] node672;
	wire [4-1:0] node673;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node683;
	wire [4-1:0] node684;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node690;
	wire [4-1:0] node693;
	wire [4-1:0] node694;
	wire [4-1:0] node698;
	wire [4-1:0] node699;
	wire [4-1:0] node700;
	wire [4-1:0] node704;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node714;
	wire [4-1:0] node717;
	wire [4-1:0] node718;
	wire [4-1:0] node721;
	wire [4-1:0] node724;
	wire [4-1:0] node725;
	wire [4-1:0] node726;
	wire [4-1:0] node729;
	wire [4-1:0] node732;
	wire [4-1:0] node733;
	wire [4-1:0] node736;
	wire [4-1:0] node739;
	wire [4-1:0] node740;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node745;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node755;
	wire [4-1:0] node758;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node765;
	wire [4-1:0] node768;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node774;
	wire [4-1:0] node775;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node784;
	wire [4-1:0] node787;
	wire [4-1:0] node788;
	wire [4-1:0] node792;
	wire [4-1:0] node793;
	wire [4-1:0] node794;
	wire [4-1:0] node795;
	wire [4-1:0] node798;
	wire [4-1:0] node801;
	wire [4-1:0] node804;
	wire [4-1:0] node805;
	wire [4-1:0] node806;
	wire [4-1:0] node809;
	wire [4-1:0] node812;
	wire [4-1:0] node813;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node824;
	wire [4-1:0] node826;
	wire [4-1:0] node829;
	wire [4-1:0] node831;
	wire [4-1:0] node832;
	wire [4-1:0] node835;
	wire [4-1:0] node838;
	wire [4-1:0] node839;
	wire [4-1:0] node841;
	wire [4-1:0] node844;
	wire [4-1:0] node845;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node851;
	wire [4-1:0] node852;
	wire [4-1:0] node853;
	wire [4-1:0] node856;
	wire [4-1:0] node859;
	wire [4-1:0] node861;
	wire [4-1:0] node864;
	wire [4-1:0] node865;
	wire [4-1:0] node866;
	wire [4-1:0] node869;
	wire [4-1:0] node872;
	wire [4-1:0] node874;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node879;
	wire [4-1:0] node880;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node887;
	wire [4-1:0] node891;
	wire [4-1:0] node892;
	wire [4-1:0] node895;
	wire [4-1:0] node898;
	wire [4-1:0] node899;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node904;
	wire [4-1:0] node906;
	wire [4-1:0] node910;
	wire [4-1:0] node911;
	wire [4-1:0] node912;
	wire [4-1:0] node915;
	wire [4-1:0] node918;
	wire [4-1:0] node919;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node925;
	wire [4-1:0] node926;
	wire [4-1:0] node929;
	wire [4-1:0] node932;
	wire [4-1:0] node934;
	wire [4-1:0] node937;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node947;
	wire [4-1:0] node951;
	wire [4-1:0] node953;
	wire [4-1:0] node954;
	wire [4-1:0] node957;
	wire [4-1:0] node960;
	wire [4-1:0] node961;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node966;
	wire [4-1:0] node969;
	wire [4-1:0] node972;
	wire [4-1:0] node973;
	wire [4-1:0] node974;
	wire [4-1:0] node977;
	wire [4-1:0] node980;
	wire [4-1:0] node981;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node989;
	wire [4-1:0] node992;
	wire [4-1:0] node994;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node1001;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1006;
	wire [4-1:0] node1007;
	wire [4-1:0] node1010;
	wire [4-1:0] node1013;
	wire [4-1:0] node1016;
	wire [4-1:0] node1018;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1025;
	wire [4-1:0] node1028;
	wire [4-1:0] node1029;
	wire [4-1:0] node1030;
	wire [4-1:0] node1033;
	wire [4-1:0] node1036;
	wire [4-1:0] node1037;
	wire [4-1:0] node1040;
	wire [4-1:0] node1043;
	wire [4-1:0] node1044;
	wire [4-1:0] node1045;
	wire [4-1:0] node1046;
	wire [4-1:0] node1049;
	wire [4-1:0] node1052;
	wire [4-1:0] node1054;
	wire [4-1:0] node1057;
	wire [4-1:0] node1059;
	wire [4-1:0] node1060;
	wire [4-1:0] node1064;
	wire [4-1:0] node1065;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1074;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1081;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1086;
	wire [4-1:0] node1089;
	wire [4-1:0] node1092;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1097;
	wire [4-1:0] node1100;
	wire [4-1:0] node1101;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1112;
	wire [4-1:0] node1116;
	wire [4-1:0] node1117;
	wire [4-1:0] node1119;
	wire [4-1:0] node1123;
	wire [4-1:0] node1124;
	wire [4-1:0] node1126;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1132;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1139;
	wire [4-1:0] node1140;
	wire [4-1:0] node1142;
	wire [4-1:0] node1145;
	wire [4-1:0] node1147;
	wire [4-1:0] node1150;
	wire [4-1:0] node1152;
	wire [4-1:0] node1153;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1169;
	wire [4-1:0] node1170;
	wire [4-1:0] node1171;
	wire [4-1:0] node1176;
	wire [4-1:0] node1177;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1182;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1188;
	wire [4-1:0] node1191;
	wire [4-1:0] node1193;
	wire [4-1:0] node1196;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1203;
	wire [4-1:0] node1206;
	wire [4-1:0] node1207;
	wire [4-1:0] node1208;
	wire [4-1:0] node1212;
	wire [4-1:0] node1213;
	wire [4-1:0] node1217;
	wire [4-1:0] node1218;
	wire [4-1:0] node1219;
	wire [4-1:0] node1220;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1224;
	wire [4-1:0] node1225;
	wire [4-1:0] node1228;
	wire [4-1:0] node1230;
	wire [4-1:0] node1233;
	wire [4-1:0] node1235;
	wire [4-1:0] node1237;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1243;
	wire [4-1:0] node1246;
	wire [4-1:0] node1247;
	wire [4-1:0] node1249;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1256;
	wire [4-1:0] node1259;
	wire [4-1:0] node1260;
	wire [4-1:0] node1263;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1269;
	wire [4-1:0] node1271;
	wire [4-1:0] node1274;
	wire [4-1:0] node1275;
	wire [4-1:0] node1276;
	wire [4-1:0] node1277;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1284;
	wire [4-1:0] node1287;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1293;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1300;
	wire [4-1:0] node1301;
	wire [4-1:0] node1302;
	wire [4-1:0] node1303;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1312;
	wire [4-1:0] node1313;
	wire [4-1:0] node1314;
	wire [4-1:0] node1315;
	wire [4-1:0] node1320;
	wire [4-1:0] node1322;
	wire [4-1:0] node1324;
	wire [4-1:0] node1327;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1332;
	wire [4-1:0] node1335;
	wire [4-1:0] node1336;
	wire [4-1:0] node1337;
	wire [4-1:0] node1341;
	wire [4-1:0] node1342;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1350;
	wire [4-1:0] node1352;
	wire [4-1:0] node1355;
	wire [4-1:0] node1357;
	wire [4-1:0] node1360;
	wire [4-1:0] node1361;
	wire [4-1:0] node1363;
	wire [4-1:0] node1366;
	wire [4-1:0] node1367;
	wire [4-1:0] node1371;
	wire [4-1:0] node1372;
	wire [4-1:0] node1373;
	wire [4-1:0] node1375;
	wire [4-1:0] node1376;
	wire [4-1:0] node1380;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1386;
	wire [4-1:0] node1389;
	wire [4-1:0] node1390;
	wire [4-1:0] node1391;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1396;
	wire [4-1:0] node1400;
	wire [4-1:0] node1401;
	wire [4-1:0] node1404;
	wire [4-1:0] node1406;
	wire [4-1:0] node1409;
	wire [4-1:0] node1410;
	wire [4-1:0] node1411;
	wire [4-1:0] node1415;
	wire [4-1:0] node1416;
	wire [4-1:0] node1417;
	wire [4-1:0] node1421;
	wire [4-1:0] node1423;
	wire [4-1:0] node1426;
	wire [4-1:0] node1427;
	wire [4-1:0] node1428;
	wire [4-1:0] node1429;
	wire [4-1:0] node1430;
	wire [4-1:0] node1432;
	wire [4-1:0] node1435;
	wire [4-1:0] node1436;
	wire [4-1:0] node1438;
	wire [4-1:0] node1439;
	wire [4-1:0] node1443;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1450;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1453;
	wire [4-1:0] node1455;
	wire [4-1:0] node1458;
	wire [4-1:0] node1460;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1472;
	wire [4-1:0] node1474;
	wire [4-1:0] node1475;
	wire [4-1:0] node1476;
	wire [4-1:0] node1480;
	wire [4-1:0] node1483;
	wire [4-1:0] node1484;
	wire [4-1:0] node1485;
	wire [4-1:0] node1487;
	wire [4-1:0] node1488;
	wire [4-1:0] node1491;
	wire [4-1:0] node1492;
	wire [4-1:0] node1496;
	wire [4-1:0] node1497;
	wire [4-1:0] node1498;
	wire [4-1:0] node1500;
	wire [4-1:0] node1503;
	wire [4-1:0] node1506;
	wire [4-1:0] node1507;
	wire [4-1:0] node1509;
	wire [4-1:0] node1513;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1520;
	wire [4-1:0] node1521;
	wire [4-1:0] node1525;
	wire [4-1:0] node1526;
	wire [4-1:0] node1528;
	wire [4-1:0] node1530;
	wire [4-1:0] node1533;
	wire [4-1:0] node1536;
	wire [4-1:0] node1537;
	wire [4-1:0] node1538;
	wire [4-1:0] node1539;
	wire [4-1:0] node1540;
	wire [4-1:0] node1542;
	wire [4-1:0] node1545;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1550;
	wire [4-1:0] node1553;
	wire [4-1:0] node1555;
	wire [4-1:0] node1558;
	wire [4-1:0] node1560;
	wire [4-1:0] node1563;
	wire [4-1:0] node1564;
	wire [4-1:0] node1566;
	wire [4-1:0] node1569;
	wire [4-1:0] node1570;
	wire [4-1:0] node1572;
	wire [4-1:0] node1573;
	wire [4-1:0] node1577;
	wire [4-1:0] node1578;
	wire [4-1:0] node1582;
	wire [4-1:0] node1583;
	wire [4-1:0] node1584;
	wire [4-1:0] node1585;
	wire [4-1:0] node1586;
	wire [4-1:0] node1589;
	wire [4-1:0] node1592;
	wire [4-1:0] node1593;
	wire [4-1:0] node1595;
	wire [4-1:0] node1599;
	wire [4-1:0] node1600;
	wire [4-1:0] node1601;
	wire [4-1:0] node1604;
	wire [4-1:0] node1606;
	wire [4-1:0] node1609;
	wire [4-1:0] node1611;
	wire [4-1:0] node1613;
	wire [4-1:0] node1616;
	wire [4-1:0] node1617;
	wire [4-1:0] node1618;
	wire [4-1:0] node1620;
	wire [4-1:0] node1622;
	wire [4-1:0] node1625;
	wire [4-1:0] node1626;
	wire [4-1:0] node1630;
	wire [4-1:0] node1631;
	wire [4-1:0] node1632;
	wire [4-1:0] node1636;
	wire [4-1:0] node1637;
	wire [4-1:0] node1639;
	wire [4-1:0] node1643;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1646;
	wire [4-1:0] node1647;
	wire [4-1:0] node1648;
	wire [4-1:0] node1649;
	wire [4-1:0] node1651;
	wire [4-1:0] node1652;
	wire [4-1:0] node1656;
	wire [4-1:0] node1657;
	wire [4-1:0] node1660;
	wire [4-1:0] node1663;
	wire [4-1:0] node1664;
	wire [4-1:0] node1665;
	wire [4-1:0] node1666;
	wire [4-1:0] node1671;
	wire [4-1:0] node1672;
	wire [4-1:0] node1675;
	wire [4-1:0] node1677;
	wire [4-1:0] node1680;
	wire [4-1:0] node1681;
	wire [4-1:0] node1682;
	wire [4-1:0] node1683;
	wire [4-1:0] node1687;
	wire [4-1:0] node1688;
	wire [4-1:0] node1691;
	wire [4-1:0] node1694;
	wire [4-1:0] node1695;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1702;
	wire [4-1:0] node1703;
	wire [4-1:0] node1705;
	wire [4-1:0] node1709;
	wire [4-1:0] node1710;
	wire [4-1:0] node1711;
	wire [4-1:0] node1712;
	wire [4-1:0] node1713;
	wire [4-1:0] node1715;
	wire [4-1:0] node1719;
	wire [4-1:0] node1720;
	wire [4-1:0] node1723;
	wire [4-1:0] node1726;
	wire [4-1:0] node1727;
	wire [4-1:0] node1728;
	wire [4-1:0] node1729;
	wire [4-1:0] node1733;
	wire [4-1:0] node1735;
	wire [4-1:0] node1738;
	wire [4-1:0] node1739;
	wire [4-1:0] node1742;
	wire [4-1:0] node1744;
	wire [4-1:0] node1747;
	wire [4-1:0] node1748;
	wire [4-1:0] node1749;
	wire [4-1:0] node1752;
	wire [4-1:0] node1753;
	wire [4-1:0] node1756;
	wire [4-1:0] node1758;
	wire [4-1:0] node1761;
	wire [4-1:0] node1762;
	wire [4-1:0] node1763;
	wire [4-1:0] node1766;
	wire [4-1:0] node1769;
	wire [4-1:0] node1770;
	wire [4-1:0] node1774;
	wire [4-1:0] node1775;
	wire [4-1:0] node1776;
	wire [4-1:0] node1777;
	wire [4-1:0] node1778;
	wire [4-1:0] node1779;
	wire [4-1:0] node1782;
	wire [4-1:0] node1785;
	wire [4-1:0] node1787;
	wire [4-1:0] node1788;
	wire [4-1:0] node1792;
	wire [4-1:0] node1793;
	wire [4-1:0] node1796;
	wire [4-1:0] node1797;
	wire [4-1:0] node1800;
	wire [4-1:0] node1802;
	wire [4-1:0] node1805;
	wire [4-1:0] node1806;
	wire [4-1:0] node1807;
	wire [4-1:0] node1808;
	wire [4-1:0] node1809;
	wire [4-1:0] node1813;
	wire [4-1:0] node1816;
	wire [4-1:0] node1818;
	wire [4-1:0] node1819;
	wire [4-1:0] node1823;
	wire [4-1:0] node1824;
	wire [4-1:0] node1826;
	wire [4-1:0] node1829;
	wire [4-1:0] node1830;
	wire [4-1:0] node1833;
	wire [4-1:0] node1835;
	wire [4-1:0] node1838;
	wire [4-1:0] node1839;
	wire [4-1:0] node1840;
	wire [4-1:0] node1841;
	wire [4-1:0] node1843;
	wire [4-1:0] node1846;
	wire [4-1:0] node1848;
	wire [4-1:0] node1851;
	wire [4-1:0] node1852;
	wire [4-1:0] node1855;
	wire [4-1:0] node1856;
	wire [4-1:0] node1858;
	wire [4-1:0] node1861;
	wire [4-1:0] node1863;
	wire [4-1:0] node1866;
	wire [4-1:0] node1867;
	wire [4-1:0] node1868;
	wire [4-1:0] node1869;
	wire [4-1:0] node1870;
	wire [4-1:0] node1873;
	wire [4-1:0] node1876;
	wire [4-1:0] node1878;
	wire [4-1:0] node1881;
	wire [4-1:0] node1882;
	wire [4-1:0] node1886;
	wire [4-1:0] node1887;
	wire [4-1:0] node1889;
	wire [4-1:0] node1891;
	wire [4-1:0] node1894;
	wire [4-1:0] node1895;
	wire [4-1:0] node1896;
	wire [4-1:0] node1899;
	wire [4-1:0] node1903;
	wire [4-1:0] node1904;
	wire [4-1:0] node1905;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1908;
	wire [4-1:0] node1909;
	wire [4-1:0] node1912;
	wire [4-1:0] node1913;
	wire [4-1:0] node1917;
	wire [4-1:0] node1918;
	wire [4-1:0] node1919;
	wire [4-1:0] node1924;
	wire [4-1:0] node1925;
	wire [4-1:0] node1926;
	wire [4-1:0] node1928;
	wire [4-1:0] node1931;
	wire [4-1:0] node1933;
	wire [4-1:0] node1936;
	wire [4-1:0] node1937;
	wire [4-1:0] node1939;
	wire [4-1:0] node1942;
	wire [4-1:0] node1945;
	wire [4-1:0] node1946;
	wire [4-1:0] node1947;
	wire [4-1:0] node1949;
	wire [4-1:0] node1950;
	wire [4-1:0] node1953;
	wire [4-1:0] node1956;
	wire [4-1:0] node1957;
	wire [4-1:0] node1958;
	wire [4-1:0] node1961;
	wire [4-1:0] node1965;
	wire [4-1:0] node1966;
	wire [4-1:0] node1967;
	wire [4-1:0] node1968;
	wire [4-1:0] node1972;
	wire [4-1:0] node1973;
	wire [4-1:0] node1976;
	wire [4-1:0] node1979;
	wire [4-1:0] node1980;
	wire [4-1:0] node1981;
	wire [4-1:0] node1986;
	wire [4-1:0] node1987;
	wire [4-1:0] node1988;
	wire [4-1:0] node1989;
	wire [4-1:0] node1990;
	wire [4-1:0] node1994;
	wire [4-1:0] node1995;
	wire [4-1:0] node1996;
	wire [4-1:0] node2000;
	wire [4-1:0] node2002;
	wire [4-1:0] node2005;
	wire [4-1:0] node2006;
	wire [4-1:0] node2007;
	wire [4-1:0] node2010;
	wire [4-1:0] node2012;
	wire [4-1:0] node2015;
	wire [4-1:0] node2017;
	wire [4-1:0] node2020;
	wire [4-1:0] node2021;
	wire [4-1:0] node2022;
	wire [4-1:0] node2023;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2030;
	wire [4-1:0] node2033;
	wire [4-1:0] node2035;
	wire [4-1:0] node2038;
	wire [4-1:0] node2039;
	wire [4-1:0] node2040;
	wire [4-1:0] node2041;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2050;
	wire [4-1:0] node2052;
	wire [4-1:0] node2053;
	wire [4-1:0] node2057;
	wire [4-1:0] node2058;
	wire [4-1:0] node2059;
	wire [4-1:0] node2060;
	wire [4-1:0] node2061;
	wire [4-1:0] node2064;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2070;
	wire [4-1:0] node2071;
	wire [4-1:0] node2075;
	wire [4-1:0] node2076;
	wire [4-1:0] node2077;
	wire [4-1:0] node2080;
	wire [4-1:0] node2083;
	wire [4-1:0] node2084;
	wire [4-1:0] node2085;
	wire [4-1:0] node2088;
	wire [4-1:0] node2091;
	wire [4-1:0] node2092;
	wire [4-1:0] node2095;
	wire [4-1:0] node2098;
	wire [4-1:0] node2099;
	wire [4-1:0] node2100;
	wire [4-1:0] node2101;
	wire [4-1:0] node2103;
	wire [4-1:0] node2106;
	wire [4-1:0] node2109;
	wire [4-1:0] node2110;
	wire [4-1:0] node2114;
	wire [4-1:0] node2115;
	wire [4-1:0] node2116;
	wire [4-1:0] node2117;
	wire [4-1:0] node2120;
	wire [4-1:0] node2124;
	wire [4-1:0] node2125;
	wire [4-1:0] node2126;
	wire [4-1:0] node2129;
	wire [4-1:0] node2133;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2136;
	wire [4-1:0] node2137;
	wire [4-1:0] node2138;
	wire [4-1:0] node2142;
	wire [4-1:0] node2145;
	wire [4-1:0] node2146;
	wire [4-1:0] node2149;
	wire [4-1:0] node2151;
	wire [4-1:0] node2154;
	wire [4-1:0] node2155;
	wire [4-1:0] node2157;
	wire [4-1:0] node2159;
	wire [4-1:0] node2162;
	wire [4-1:0] node2164;
	wire [4-1:0] node2166;
	wire [4-1:0] node2169;
	wire [4-1:0] node2170;
	wire [4-1:0] node2171;
	wire [4-1:0] node2172;
	wire [4-1:0] node2173;
	wire [4-1:0] node2176;
	wire [4-1:0] node2180;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2186;
	wire [4-1:0] node2189;
	wire [4-1:0] node2190;
	wire [4-1:0] node2191;
	wire [4-1:0] node2193;
	wire [4-1:0] node2196;
	wire [4-1:0] node2198;
	wire [4-1:0] node2201;
	wire [4-1:0] node2204;
	wire [4-1:0] node2205;
	wire [4-1:0] node2206;
	wire [4-1:0] node2207;
	wire [4-1:0] node2208;
	wire [4-1:0] node2209;
	wire [4-1:0] node2210;
	wire [4-1:0] node2211;
	wire [4-1:0] node2212;
	wire [4-1:0] node2215;
	wire [4-1:0] node2217;
	wire [4-1:0] node2220;
	wire [4-1:0] node2221;
	wire [4-1:0] node2222;
	wire [4-1:0] node2225;
	wire [4-1:0] node2228;
	wire [4-1:0] node2230;
	wire [4-1:0] node2233;
	wire [4-1:0] node2234;
	wire [4-1:0] node2235;
	wire [4-1:0] node2236;
	wire [4-1:0] node2237;
	wire [4-1:0] node2240;
	wire [4-1:0] node2243;
	wire [4-1:0] node2245;
	wire [4-1:0] node2248;
	wire [4-1:0] node2249;
	wire [4-1:0] node2250;
	wire [4-1:0] node2253;
	wire [4-1:0] node2257;
	wire [4-1:0] node2258;
	wire [4-1:0] node2259;
	wire [4-1:0] node2260;
	wire [4-1:0] node2263;
	wire [4-1:0] node2267;
	wire [4-1:0] node2268;
	wire [4-1:0] node2271;
	wire [4-1:0] node2274;
	wire [4-1:0] node2275;
	wire [4-1:0] node2276;
	wire [4-1:0] node2277;
	wire [4-1:0] node2280;
	wire [4-1:0] node2282;
	wire [4-1:0] node2285;
	wire [4-1:0] node2286;
	wire [4-1:0] node2287;
	wire [4-1:0] node2291;
	wire [4-1:0] node2293;
	wire [4-1:0] node2294;
	wire [4-1:0] node2297;
	wire [4-1:0] node2300;
	wire [4-1:0] node2301;
	wire [4-1:0] node2302;
	wire [4-1:0] node2303;
	wire [4-1:0] node2304;
	wire [4-1:0] node2307;
	wire [4-1:0] node2310;
	wire [4-1:0] node2311;
	wire [4-1:0] node2314;
	wire [4-1:0] node2317;
	wire [4-1:0] node2318;
	wire [4-1:0] node2319;
	wire [4-1:0] node2322;
	wire [4-1:0] node2325;
	wire [4-1:0] node2326;
	wire [4-1:0] node2329;
	wire [4-1:0] node2332;
	wire [4-1:0] node2333;
	wire [4-1:0] node2334;
	wire [4-1:0] node2335;
	wire [4-1:0] node2338;
	wire [4-1:0] node2341;
	wire [4-1:0] node2342;
	wire [4-1:0] node2345;
	wire [4-1:0] node2348;
	wire [4-1:0] node2350;
	wire [4-1:0] node2351;
	wire [4-1:0] node2354;
	wire [4-1:0] node2357;
	wire [4-1:0] node2358;
	wire [4-1:0] node2359;
	wire [4-1:0] node2360;
	wire [4-1:0] node2361;
	wire [4-1:0] node2362;
	wire [4-1:0] node2365;
	wire [4-1:0] node2368;
	wire [4-1:0] node2369;
	wire [4-1:0] node2372;
	wire [4-1:0] node2375;
	wire [4-1:0] node2376;
	wire [4-1:0] node2377;
	wire [4-1:0] node2379;
	wire [4-1:0] node2383;
	wire [4-1:0] node2384;
	wire [4-1:0] node2386;
	wire [4-1:0] node2389;
	wire [4-1:0] node2391;
	wire [4-1:0] node2394;
	wire [4-1:0] node2395;
	wire [4-1:0] node2396;
	wire [4-1:0] node2397;
	wire [4-1:0] node2400;
	wire [4-1:0] node2403;
	wire [4-1:0] node2404;
	wire [4-1:0] node2407;
	wire [4-1:0] node2410;
	wire [4-1:0] node2411;
	wire [4-1:0] node2412;
	wire [4-1:0] node2413;
	wire [4-1:0] node2418;
	wire [4-1:0] node2419;
	wire [4-1:0] node2421;
	wire [4-1:0] node2424;
	wire [4-1:0] node2425;
	wire [4-1:0] node2428;
	wire [4-1:0] node2431;
	wire [4-1:0] node2432;
	wire [4-1:0] node2433;
	wire [4-1:0] node2434;
	wire [4-1:0] node2435;
	wire [4-1:0] node2439;
	wire [4-1:0] node2440;
	wire [4-1:0] node2443;
	wire [4-1:0] node2445;
	wire [4-1:0] node2448;
	wire [4-1:0] node2449;
	wire [4-1:0] node2450;
	wire [4-1:0] node2451;
	wire [4-1:0] node2454;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2461;
	wire [4-1:0] node2464;
	wire [4-1:0] node2465;
	wire [4-1:0] node2466;
	wire [4-1:0] node2470;
	wire [4-1:0] node2471;
	wire [4-1:0] node2474;
	wire [4-1:0] node2477;
	wire [4-1:0] node2478;
	wire [4-1:0] node2479;
	wire [4-1:0] node2480;
	wire [4-1:0] node2483;
	wire [4-1:0] node2486;
	wire [4-1:0] node2487;
	wire [4-1:0] node2489;
	wire [4-1:0] node2492;
	wire [4-1:0] node2495;
	wire [4-1:0] node2496;
	wire [4-1:0] node2497;
	wire [4-1:0] node2498;
	wire [4-1:0] node2501;
	wire [4-1:0] node2504;
	wire [4-1:0] node2505;
	wire [4-1:0] node2508;
	wire [4-1:0] node2511;
	wire [4-1:0] node2512;
	wire [4-1:0] node2515;
	wire [4-1:0] node2518;
	wire [4-1:0] node2519;
	wire [4-1:0] node2520;
	wire [4-1:0] node2521;
	wire [4-1:0] node2522;
	wire [4-1:0] node2523;
	wire [4-1:0] node2524;
	wire [4-1:0] node2527;
	wire [4-1:0] node2530;
	wire [4-1:0] node2531;
	wire [4-1:0] node2532;
	wire [4-1:0] node2535;
	wire [4-1:0] node2539;
	wire [4-1:0] node2540;
	wire [4-1:0] node2542;
	wire [4-1:0] node2545;
	wire [4-1:0] node2546;
	wire [4-1:0] node2547;
	wire [4-1:0] node2550;
	wire [4-1:0] node2553;
	wire [4-1:0] node2555;
	wire [4-1:0] node2558;
	wire [4-1:0] node2559;
	wire [4-1:0] node2560;
	wire [4-1:0] node2561;
	wire [4-1:0] node2564;
	wire [4-1:0] node2567;
	wire [4-1:0] node2568;
	wire [4-1:0] node2569;
	wire [4-1:0] node2572;
	wire [4-1:0] node2575;
	wire [4-1:0] node2577;
	wire [4-1:0] node2580;
	wire [4-1:0] node2581;
	wire [4-1:0] node2582;
	wire [4-1:0] node2583;
	wire [4-1:0] node2587;
	wire [4-1:0] node2590;
	wire [4-1:0] node2591;
	wire [4-1:0] node2594;
	wire [4-1:0] node2596;
	wire [4-1:0] node2599;
	wire [4-1:0] node2600;
	wire [4-1:0] node2601;
	wire [4-1:0] node2602;
	wire [4-1:0] node2603;
	wire [4-1:0] node2606;
	wire [4-1:0] node2607;
	wire [4-1:0] node2610;
	wire [4-1:0] node2613;
	wire [4-1:0] node2615;
	wire [4-1:0] node2617;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2622;
	wire [4-1:0] node2623;
	wire [4-1:0] node2626;
	wire [4-1:0] node2629;
	wire [4-1:0] node2630;
	wire [4-1:0] node2633;
	wire [4-1:0] node2636;
	wire [4-1:0] node2638;
	wire [4-1:0] node2640;
	wire [4-1:0] node2643;
	wire [4-1:0] node2644;
	wire [4-1:0] node2645;
	wire [4-1:0] node2646;
	wire [4-1:0] node2647;
	wire [4-1:0] node2651;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2656;
	wire [4-1:0] node2659;
	wire [4-1:0] node2662;
	wire [4-1:0] node2663;
	wire [4-1:0] node2667;
	wire [4-1:0] node2668;
	wire [4-1:0] node2669;
	wire [4-1:0] node2672;
	wire [4-1:0] node2673;
	wire [4-1:0] node2677;
	wire [4-1:0] node2678;
	wire [4-1:0] node2681;
	wire [4-1:0] node2682;
	wire [4-1:0] node2685;
	wire [4-1:0] node2688;
	wire [4-1:0] node2689;
	wire [4-1:0] node2690;
	wire [4-1:0] node2691;
	wire [4-1:0] node2692;
	wire [4-1:0] node2693;
	wire [4-1:0] node2695;
	wire [4-1:0] node2699;
	wire [4-1:0] node2700;
	wire [4-1:0] node2701;
	wire [4-1:0] node2704;
	wire [4-1:0] node2707;
	wire [4-1:0] node2708;
	wire [4-1:0] node2711;
	wire [4-1:0] node2714;
	wire [4-1:0] node2715;
	wire [4-1:0] node2716;
	wire [4-1:0] node2718;
	wire [4-1:0] node2722;
	wire [4-1:0] node2723;
	wire [4-1:0] node2724;
	wire [4-1:0] node2727;
	wire [4-1:0] node2730;
	wire [4-1:0] node2732;
	wire [4-1:0] node2735;
	wire [4-1:0] node2736;
	wire [4-1:0] node2737;
	wire [4-1:0] node2738;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2745;
	wire [4-1:0] node2748;
	wire [4-1:0] node2749;
	wire [4-1:0] node2750;
	wire [4-1:0] node2754;
	wire [4-1:0] node2757;
	wire [4-1:0] node2758;
	wire [4-1:0] node2761;
	wire [4-1:0] node2762;
	wire [4-1:0] node2765;
	wire [4-1:0] node2766;
	wire [4-1:0] node2769;
	wire [4-1:0] node2772;
	wire [4-1:0] node2773;
	wire [4-1:0] node2774;
	wire [4-1:0] node2775;
	wire [4-1:0] node2776;
	wire [4-1:0] node2777;
	wire [4-1:0] node2781;
	wire [4-1:0] node2784;
	wire [4-1:0] node2785;
	wire [4-1:0] node2788;
	wire [4-1:0] node2791;
	wire [4-1:0] node2792;
	wire [4-1:0] node2793;
	wire [4-1:0] node2794;
	wire [4-1:0] node2797;
	wire [4-1:0] node2800;
	wire [4-1:0] node2801;
	wire [4-1:0] node2804;
	wire [4-1:0] node2807;
	wire [4-1:0] node2808;
	wire [4-1:0] node2809;
	wire [4-1:0] node2812;
	wire [4-1:0] node2815;
	wire [4-1:0] node2817;
	wire [4-1:0] node2820;
	wire [4-1:0] node2821;
	wire [4-1:0] node2822;
	wire [4-1:0] node2823;
	wire [4-1:0] node2824;
	wire [4-1:0] node2827;
	wire [4-1:0] node2830;
	wire [4-1:0] node2831;
	wire [4-1:0] node2835;
	wire [4-1:0] node2836;
	wire [4-1:0] node2838;
	wire [4-1:0] node2841;
	wire [4-1:0] node2842;
	wire [4-1:0] node2845;
	wire [4-1:0] node2848;
	wire [4-1:0] node2849;
	wire [4-1:0] node2850;
	wire [4-1:0] node2854;
	wire [4-1:0] node2855;
	wire [4-1:0] node2858;
	wire [4-1:0] node2860;
	wire [4-1:0] node2863;
	wire [4-1:0] node2864;
	wire [4-1:0] node2865;
	wire [4-1:0] node2866;
	wire [4-1:0] node2867;
	wire [4-1:0] node2868;
	wire [4-1:0] node2869;
	wire [4-1:0] node2870;
	wire [4-1:0] node2872;
	wire [4-1:0] node2875;
	wire [4-1:0] node2878;
	wire [4-1:0] node2880;
	wire [4-1:0] node2883;
	wire [4-1:0] node2884;
	wire [4-1:0] node2885;
	wire [4-1:0] node2888;
	wire [4-1:0] node2891;
	wire [4-1:0] node2892;
	wire [4-1:0] node2893;
	wire [4-1:0] node2897;
	wire [4-1:0] node2898;
	wire [4-1:0] node2901;
	wire [4-1:0] node2904;
	wire [4-1:0] node2905;
	wire [4-1:0] node2906;
	wire [4-1:0] node2907;
	wire [4-1:0] node2908;
	wire [4-1:0] node2912;
	wire [4-1:0] node2915;
	wire [4-1:0] node2916;
	wire [4-1:0] node2917;
	wire [4-1:0] node2920;
	wire [4-1:0] node2924;
	wire [4-1:0] node2926;
	wire [4-1:0] node2927;
	wire [4-1:0] node2928;
	wire [4-1:0] node2932;
	wire [4-1:0] node2933;
	wire [4-1:0] node2936;
	wire [4-1:0] node2939;
	wire [4-1:0] node2940;
	wire [4-1:0] node2941;
	wire [4-1:0] node2942;
	wire [4-1:0] node2943;
	wire [4-1:0] node2944;
	wire [4-1:0] node2947;
	wire [4-1:0] node2950;
	wire [4-1:0] node2951;
	wire [4-1:0] node2954;
	wire [4-1:0] node2957;
	wire [4-1:0] node2958;
	wire [4-1:0] node2959;
	wire [4-1:0] node2963;
	wire [4-1:0] node2964;
	wire [4-1:0] node2967;
	wire [4-1:0] node2970;
	wire [4-1:0] node2971;
	wire [4-1:0] node2972;
	wire [4-1:0] node2974;
	wire [4-1:0] node2977;
	wire [4-1:0] node2979;
	wire [4-1:0] node2982;
	wire [4-1:0] node2983;
	wire [4-1:0] node2986;
	wire [4-1:0] node2989;
	wire [4-1:0] node2990;
	wire [4-1:0] node2992;
	wire [4-1:0] node2994;
	wire [4-1:0] node2995;
	wire [4-1:0] node2998;
	wire [4-1:0] node3001;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3006;
	wire [4-1:0] node3007;
	wire [4-1:0] node3011;
	wire [4-1:0] node3013;
	wire [4-1:0] node3014;
	wire [4-1:0] node3018;
	wire [4-1:0] node3019;
	wire [4-1:0] node3020;
	wire [4-1:0] node3021;
	wire [4-1:0] node3022;
	wire [4-1:0] node3023;
	wire [4-1:0] node3026;
	wire [4-1:0] node3027;
	wire [4-1:0] node3031;
	wire [4-1:0] node3033;
	wire [4-1:0] node3036;
	wire [4-1:0] node3037;
	wire [4-1:0] node3040;
	wire [4-1:0] node3042;
	wire [4-1:0] node3043;
	wire [4-1:0] node3047;
	wire [4-1:0] node3048;
	wire [4-1:0] node3049;
	wire [4-1:0] node3051;
	wire [4-1:0] node3052;
	wire [4-1:0] node3056;
	wire [4-1:0] node3057;
	wire [4-1:0] node3059;
	wire [4-1:0] node3062;
	wire [4-1:0] node3064;
	wire [4-1:0] node3067;
	wire [4-1:0] node3068;
	wire [4-1:0] node3071;
	wire [4-1:0] node3072;
	wire [4-1:0] node3075;
	wire [4-1:0] node3077;
	wire [4-1:0] node3080;
	wire [4-1:0] node3081;
	wire [4-1:0] node3082;
	wire [4-1:0] node3083;
	wire [4-1:0] node3085;
	wire [4-1:0] node3088;
	wire [4-1:0] node3089;
	wire [4-1:0] node3090;
	wire [4-1:0] node3094;
	wire [4-1:0] node3095;
	wire [4-1:0] node3098;
	wire [4-1:0] node3101;
	wire [4-1:0] node3102;
	wire [4-1:0] node3103;
	wire [4-1:0] node3104;
	wire [4-1:0] node3108;
	wire [4-1:0] node3109;
	wire [4-1:0] node3113;
	wire [4-1:0] node3115;
	wire [4-1:0] node3116;
	wire [4-1:0] node3119;
	wire [4-1:0] node3122;
	wire [4-1:0] node3123;
	wire [4-1:0] node3124;
	wire [4-1:0] node3125;
	wire [4-1:0] node3128;
	wire [4-1:0] node3131;
	wire [4-1:0] node3132;
	wire [4-1:0] node3134;
	wire [4-1:0] node3137;
	wire [4-1:0] node3139;
	wire [4-1:0] node3142;
	wire [4-1:0] node3143;
	wire [4-1:0] node3144;
	wire [4-1:0] node3147;
	wire [4-1:0] node3148;
	wire [4-1:0] node3152;
	wire [4-1:0] node3153;
	wire [4-1:0] node3156;
	wire [4-1:0] node3158;
	wire [4-1:0] node3161;
	wire [4-1:0] node3162;
	wire [4-1:0] node3163;
	wire [4-1:0] node3164;
	wire [4-1:0] node3165;
	wire [4-1:0] node3166;
	wire [4-1:0] node3167;
	wire [4-1:0] node3168;
	wire [4-1:0] node3172;
	wire [4-1:0] node3175;
	wire [4-1:0] node3176;
	wire [4-1:0] node3177;
	wire [4-1:0] node3181;
	wire [4-1:0] node3182;
	wire [4-1:0] node3186;
	wire [4-1:0] node3187;
	wire [4-1:0] node3189;
	wire [4-1:0] node3192;
	wire [4-1:0] node3194;
	wire [4-1:0] node3195;
	wire [4-1:0] node3199;
	wire [4-1:0] node3200;
	wire [4-1:0] node3201;
	wire [4-1:0] node3202;
	wire [4-1:0] node3203;
	wire [4-1:0] node3208;
	wire [4-1:0] node3211;
	wire [4-1:0] node3212;
	wire [4-1:0] node3213;
	wire [4-1:0] node3214;
	wire [4-1:0] node3218;
	wire [4-1:0] node3220;
	wire [4-1:0] node3223;
	wire [4-1:0] node3225;
	wire [4-1:0] node3228;
	wire [4-1:0] node3229;
	wire [4-1:0] node3230;
	wire [4-1:0] node3231;
	wire [4-1:0] node3232;
	wire [4-1:0] node3235;
	wire [4-1:0] node3238;
	wire [4-1:0] node3240;
	wire [4-1:0] node3243;
	wire [4-1:0] node3244;
	wire [4-1:0] node3245;
	wire [4-1:0] node3246;
	wire [4-1:0] node3249;
	wire [4-1:0] node3252;
	wire [4-1:0] node3253;
	wire [4-1:0] node3256;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3263;
	wire [4-1:0] node3265;
	wire [4-1:0] node3268;
	wire [4-1:0] node3269;
	wire [4-1:0] node3270;
	wire [4-1:0] node3271;
	wire [4-1:0] node3273;
	wire [4-1:0] node3276;
	wire [4-1:0] node3279;
	wire [4-1:0] node3280;
	wire [4-1:0] node3283;
	wire [4-1:0] node3286;
	wire [4-1:0] node3287;
	wire [4-1:0] node3288;
	wire [4-1:0] node3291;
	wire [4-1:0] node3294;
	wire [4-1:0] node3295;
	wire [4-1:0] node3296;
	wire [4-1:0] node3299;
	wire [4-1:0] node3302;
	wire [4-1:0] node3303;
	wire [4-1:0] node3307;
	wire [4-1:0] node3308;
	wire [4-1:0] node3309;
	wire [4-1:0] node3310;
	wire [4-1:0] node3311;
	wire [4-1:0] node3312;
	wire [4-1:0] node3315;
	wire [4-1:0] node3318;
	wire [4-1:0] node3319;
	wire [4-1:0] node3322;
	wire [4-1:0] node3323;
	wire [4-1:0] node3326;
	wire [4-1:0] node3329;
	wire [4-1:0] node3330;
	wire [4-1:0] node3331;
	wire [4-1:0] node3332;
	wire [4-1:0] node3335;
	wire [4-1:0] node3338;
	wire [4-1:0] node3339;
	wire [4-1:0] node3342;
	wire [4-1:0] node3345;
	wire [4-1:0] node3346;
	wire [4-1:0] node3349;
	wire [4-1:0] node3350;
	wire [4-1:0] node3353;
	wire [4-1:0] node3356;
	wire [4-1:0] node3357;
	wire [4-1:0] node3358;
	wire [4-1:0] node3359;
	wire [4-1:0] node3362;
	wire [4-1:0] node3364;
	wire [4-1:0] node3367;
	wire [4-1:0] node3368;
	wire [4-1:0] node3371;
	wire [4-1:0] node3373;
	wire [4-1:0] node3376;
	wire [4-1:0] node3377;
	wire [4-1:0] node3380;
	wire [4-1:0] node3381;
	wire [4-1:0] node3384;
	wire [4-1:0] node3386;
	wire [4-1:0] node3389;
	wire [4-1:0] node3390;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3393;
	wire [4-1:0] node3395;
	wire [4-1:0] node3398;
	wire [4-1:0] node3401;
	wire [4-1:0] node3402;
	wire [4-1:0] node3405;
	wire [4-1:0] node3406;
	wire [4-1:0] node3410;
	wire [4-1:0] node3411;
	wire [4-1:0] node3412;
	wire [4-1:0] node3415;
	wire [4-1:0] node3416;
	wire [4-1:0] node3420;
	wire [4-1:0] node3422;
	wire [4-1:0] node3425;
	wire [4-1:0] node3426;
	wire [4-1:0] node3427;
	wire [4-1:0] node3428;
	wire [4-1:0] node3430;
	wire [4-1:0] node3433;
	wire [4-1:0] node3435;
	wire [4-1:0] node3438;
	wire [4-1:0] node3439;
	wire [4-1:0] node3442;
	wire [4-1:0] node3443;
	wire [4-1:0] node3446;
	wire [4-1:0] node3449;
	wire [4-1:0] node3450;
	wire [4-1:0] node3451;
	wire [4-1:0] node3455;
	wire [4-1:0] node3456;
	wire [4-1:0] node3459;
	wire [4-1:0] node3461;
	wire [4-1:0] node3464;
	wire [4-1:0] node3465;
	wire [4-1:0] node3466;
	wire [4-1:0] node3467;
	wire [4-1:0] node3468;
	wire [4-1:0] node3469;
	wire [4-1:0] node3470;
	wire [4-1:0] node3471;
	wire [4-1:0] node3472;
	wire [4-1:0] node3473;
	wire [4-1:0] node3477;
	wire [4-1:0] node3478;
	wire [4-1:0] node3482;
	wire [4-1:0] node3485;
	wire [4-1:0] node3486;
	wire [4-1:0] node3487;
	wire [4-1:0] node3489;
	wire [4-1:0] node3492;
	wire [4-1:0] node3494;
	wire [4-1:0] node3497;
	wire [4-1:0] node3499;
	wire [4-1:0] node3502;
	wire [4-1:0] node3503;
	wire [4-1:0] node3504;
	wire [4-1:0] node3506;
	wire [4-1:0] node3507;
	wire [4-1:0] node3511;
	wire [4-1:0] node3512;
	wire [4-1:0] node3514;
	wire [4-1:0] node3517;
	wire [4-1:0] node3520;
	wire [4-1:0] node3521;
	wire [4-1:0] node3522;
	wire [4-1:0] node3524;
	wire [4-1:0] node3527;
	wire [4-1:0] node3529;
	wire [4-1:0] node3532;
	wire [4-1:0] node3533;
	wire [4-1:0] node3535;
	wire [4-1:0] node3538;
	wire [4-1:0] node3540;
	wire [4-1:0] node3543;
	wire [4-1:0] node3544;
	wire [4-1:0] node3545;
	wire [4-1:0] node3546;
	wire [4-1:0] node3547;
	wire [4-1:0] node3551;
	wire [4-1:0] node3552;
	wire [4-1:0] node3556;
	wire [4-1:0] node3557;
	wire [4-1:0] node3558;
	wire [4-1:0] node3560;
	wire [4-1:0] node3564;
	wire [4-1:0] node3565;
	wire [4-1:0] node3567;
	wire [4-1:0] node3570;
	wire [4-1:0] node3573;
	wire [4-1:0] node3574;
	wire [4-1:0] node3575;
	wire [4-1:0] node3576;
	wire [4-1:0] node3578;
	wire [4-1:0] node3581;
	wire [4-1:0] node3583;
	wire [4-1:0] node3586;
	wire [4-1:0] node3588;
	wire [4-1:0] node3591;
	wire [4-1:0] node3592;
	wire [4-1:0] node3593;
	wire [4-1:0] node3594;
	wire [4-1:0] node3598;
	wire [4-1:0] node3599;
	wire [4-1:0] node3602;
	wire [4-1:0] node3605;
	wire [4-1:0] node3606;
	wire [4-1:0] node3607;
	wire [4-1:0] node3610;
	wire [4-1:0] node3613;
	wire [4-1:0] node3614;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3620;
	wire [4-1:0] node3621;
	wire [4-1:0] node3622;
	wire [4-1:0] node3623;
	wire [4-1:0] node3626;
	wire [4-1:0] node3629;
	wire [4-1:0] node3630;
	wire [4-1:0] node3633;
	wire [4-1:0] node3635;
	wire [4-1:0] node3638;
	wire [4-1:0] node3639;
	wire [4-1:0] node3640;
	wire [4-1:0] node3642;
	wire [4-1:0] node3646;
	wire [4-1:0] node3648;
	wire [4-1:0] node3649;
	wire [4-1:0] node3653;
	wire [4-1:0] node3654;
	wire [4-1:0] node3655;
	wire [4-1:0] node3656;
	wire [4-1:0] node3659;
	wire [4-1:0] node3661;
	wire [4-1:0] node3664;
	wire [4-1:0] node3665;
	wire [4-1:0] node3669;
	wire [4-1:0] node3670;
	wire [4-1:0] node3671;
	wire [4-1:0] node3673;
	wire [4-1:0] node3677;
	wire [4-1:0] node3678;
	wire [4-1:0] node3679;
	wire [4-1:0] node3682;
	wire [4-1:0] node3686;
	wire [4-1:0] node3687;
	wire [4-1:0] node3688;
	wire [4-1:0] node3689;
	wire [4-1:0] node3691;
	wire [4-1:0] node3692;
	wire [4-1:0] node3696;
	wire [4-1:0] node3698;
	wire [4-1:0] node3699;
	wire [4-1:0] node3702;
	wire [4-1:0] node3705;
	wire [4-1:0] node3706;
	wire [4-1:0] node3707;
	wire [4-1:0] node3709;
	wire [4-1:0] node3712;
	wire [4-1:0] node3713;
	wire [4-1:0] node3716;
	wire [4-1:0] node3719;
	wire [4-1:0] node3720;
	wire [4-1:0] node3721;
	wire [4-1:0] node3725;
	wire [4-1:0] node3726;
	wire [4-1:0] node3729;
	wire [4-1:0] node3732;
	wire [4-1:0] node3733;
	wire [4-1:0] node3734;
	wire [4-1:0] node3735;
	wire [4-1:0] node3736;
	wire [4-1:0] node3740;
	wire [4-1:0] node3741;
	wire [4-1:0] node3744;
	wire [4-1:0] node3747;
	wire [4-1:0] node3748;
	wire [4-1:0] node3750;
	wire [4-1:0] node3753;
	wire [4-1:0] node3754;
	wire [4-1:0] node3757;
	wire [4-1:0] node3760;
	wire [4-1:0] node3761;
	wire [4-1:0] node3762;
	wire [4-1:0] node3763;
	wire [4-1:0] node3767;
	wire [4-1:0] node3768;
	wire [4-1:0] node3771;
	wire [4-1:0] node3774;
	wire [4-1:0] node3775;
	wire [4-1:0] node3776;
	wire [4-1:0] node3781;
	wire [4-1:0] node3782;
	wire [4-1:0] node3783;
	wire [4-1:0] node3784;
	wire [4-1:0] node3785;
	wire [4-1:0] node3786;
	wire [4-1:0] node3787;
	wire [4-1:0] node3788;
	wire [4-1:0] node3791;
	wire [4-1:0] node3794;
	wire [4-1:0] node3795;
	wire [4-1:0] node3798;
	wire [4-1:0] node3801;
	wire [4-1:0] node3802;
	wire [4-1:0] node3803;
	wire [4-1:0] node3806;
	wire [4-1:0] node3809;
	wire [4-1:0] node3810;
	wire [4-1:0] node3813;
	wire [4-1:0] node3816;
	wire [4-1:0] node3817;
	wire [4-1:0] node3819;
	wire [4-1:0] node3820;
	wire [4-1:0] node3824;
	wire [4-1:0] node3825;
	wire [4-1:0] node3826;
	wire [4-1:0] node3830;
	wire [4-1:0] node3832;
	wire [4-1:0] node3835;
	wire [4-1:0] node3836;
	wire [4-1:0] node3837;
	wire [4-1:0] node3838;
	wire [4-1:0] node3839;
	wire [4-1:0] node3843;
	wire [4-1:0] node3846;
	wire [4-1:0] node3847;
	wire [4-1:0] node3850;
	wire [4-1:0] node3853;
	wire [4-1:0] node3854;
	wire [4-1:0] node3855;
	wire [4-1:0] node3856;
	wire [4-1:0] node3860;
	wire [4-1:0] node3863;
	wire [4-1:0] node3864;
	wire [4-1:0] node3866;
	wire [4-1:0] node3869;
	wire [4-1:0] node3870;
	wire [4-1:0] node3874;
	wire [4-1:0] node3875;
	wire [4-1:0] node3876;
	wire [4-1:0] node3877;
	wire [4-1:0] node3878;
	wire [4-1:0] node3880;
	wire [4-1:0] node3884;
	wire [4-1:0] node3885;
	wire [4-1:0] node3888;
	wire [4-1:0] node3889;
	wire [4-1:0] node3892;
	wire [4-1:0] node3895;
	wire [4-1:0] node3896;
	wire [4-1:0] node3897;
	wire [4-1:0] node3900;
	wire [4-1:0] node3901;
	wire [4-1:0] node3904;
	wire [4-1:0] node3907;
	wire [4-1:0] node3910;
	wire [4-1:0] node3911;
	wire [4-1:0] node3912;
	wire [4-1:0] node3913;
	wire [4-1:0] node3915;
	wire [4-1:0] node3918;
	wire [4-1:0] node3920;
	wire [4-1:0] node3923;
	wire [4-1:0] node3924;
	wire [4-1:0] node3925;
	wire [4-1:0] node3929;
	wire [4-1:0] node3930;
	wire [4-1:0] node3933;
	wire [4-1:0] node3936;
	wire [4-1:0] node3937;
	wire [4-1:0] node3938;
	wire [4-1:0] node3941;
	wire [4-1:0] node3944;
	wire [4-1:0] node3945;
	wire [4-1:0] node3946;
	wire [4-1:0] node3949;
	wire [4-1:0] node3952;
	wire [4-1:0] node3955;
	wire [4-1:0] node3956;
	wire [4-1:0] node3957;
	wire [4-1:0] node3958;
	wire [4-1:0] node3959;
	wire [4-1:0] node3960;
	wire [4-1:0] node3963;
	wire [4-1:0] node3966;
	wire [4-1:0] node3967;
	wire [4-1:0] node3968;
	wire [4-1:0] node3972;
	wire [4-1:0] node3974;
	wire [4-1:0] node3977;
	wire [4-1:0] node3978;
	wire [4-1:0] node3979;
	wire [4-1:0] node3982;
	wire [4-1:0] node3984;
	wire [4-1:0] node3987;
	wire [4-1:0] node3988;
	wire [4-1:0] node3989;
	wire [4-1:0] node3992;
	wire [4-1:0] node3996;
	wire [4-1:0] node3997;
	wire [4-1:0] node3998;
	wire [4-1:0] node3999;
	wire [4-1:0] node4002;
	wire [4-1:0] node4005;
	wire [4-1:0] node4006;
	wire [4-1:0] node4008;
	wire [4-1:0] node4012;
	wire [4-1:0] node4013;
	wire [4-1:0] node4014;
	wire [4-1:0] node4015;
	wire [4-1:0] node4018;
	wire [4-1:0] node4021;
	wire [4-1:0] node4022;
	wire [4-1:0] node4025;
	wire [4-1:0] node4028;
	wire [4-1:0] node4029;
	wire [4-1:0] node4030;
	wire [4-1:0] node4033;
	wire [4-1:0] node4036;
	wire [4-1:0] node4037;
	wire [4-1:0] node4040;
	wire [4-1:0] node4043;
	wire [4-1:0] node4044;
	wire [4-1:0] node4045;
	wire [4-1:0] node4046;
	wire [4-1:0] node4047;
	wire [4-1:0] node4050;
	wire [4-1:0] node4051;
	wire [4-1:0] node4054;
	wire [4-1:0] node4057;
	wire [4-1:0] node4058;
	wire [4-1:0] node4059;
	wire [4-1:0] node4062;
	wire [4-1:0] node4066;
	wire [4-1:0] node4067;
	wire [4-1:0] node4069;
	wire [4-1:0] node4071;
	wire [4-1:0] node4074;
	wire [4-1:0] node4075;
	wire [4-1:0] node4078;
	wire [4-1:0] node4079;
	wire [4-1:0] node4083;
	wire [4-1:0] node4084;
	wire [4-1:0] node4085;
	wire [4-1:0] node4086;
	wire [4-1:0] node4087;
	wire [4-1:0] node4090;
	wire [4-1:0] node4094;
	wire [4-1:0] node4095;
	wire [4-1:0] node4098;
	wire [4-1:0] node4099;
	wire [4-1:0] node4102;
	wire [4-1:0] node4105;
	wire [4-1:0] node4106;
	wire [4-1:0] node4107;
	wire [4-1:0] node4111;
	wire [4-1:0] node4113;
	wire [4-1:0] node4116;
	wire [4-1:0] node4117;
	wire [4-1:0] node4118;
	wire [4-1:0] node4119;
	wire [4-1:0] node4120;
	wire [4-1:0] node4121;
	wire [4-1:0] node4122;
	wire [4-1:0] node4124;
	wire [4-1:0] node4125;
	wire [4-1:0] node4130;
	wire [4-1:0] node4131;
	wire [4-1:0] node4133;
	wire [4-1:0] node4135;
	wire [4-1:0] node4138;
	wire [4-1:0] node4139;
	wire [4-1:0] node4142;
	wire [4-1:0] node4144;
	wire [4-1:0] node4147;
	wire [4-1:0] node4148;
	wire [4-1:0] node4149;
	wire [4-1:0] node4150;
	wire [4-1:0] node4153;
	wire [4-1:0] node4155;
	wire [4-1:0] node4158;
	wire [4-1:0] node4159;
	wire [4-1:0] node4162;
	wire [4-1:0] node4165;
	wire [4-1:0] node4166;
	wire [4-1:0] node4167;
	wire [4-1:0] node4169;
	wire [4-1:0] node4172;
	wire [4-1:0] node4173;
	wire [4-1:0] node4177;
	wire [4-1:0] node4178;
	wire [4-1:0] node4179;
	wire [4-1:0] node4182;
	wire [4-1:0] node4185;
	wire [4-1:0] node4186;
	wire [4-1:0] node4190;
	wire [4-1:0] node4191;
	wire [4-1:0] node4192;
	wire [4-1:0] node4193;
	wire [4-1:0] node4194;
	wire [4-1:0] node4195;
	wire [4-1:0] node4198;
	wire [4-1:0] node4201;
	wire [4-1:0] node4203;
	wire [4-1:0] node4206;
	wire [4-1:0] node4207;
	wire [4-1:0] node4210;
	wire [4-1:0] node4211;
	wire [4-1:0] node4214;
	wire [4-1:0] node4217;
	wire [4-1:0] node4218;
	wire [4-1:0] node4219;
	wire [4-1:0] node4220;
	wire [4-1:0] node4224;
	wire [4-1:0] node4226;
	wire [4-1:0] node4229;
	wire [4-1:0] node4230;
	wire [4-1:0] node4232;
	wire [4-1:0] node4235;
	wire [4-1:0] node4238;
	wire [4-1:0] node4239;
	wire [4-1:0] node4240;
	wire [4-1:0] node4242;
	wire [4-1:0] node4244;
	wire [4-1:0] node4247;
	wire [4-1:0] node4248;
	wire [4-1:0] node4249;
	wire [4-1:0] node4252;
	wire [4-1:0] node4255;
	wire [4-1:0] node4256;
	wire [4-1:0] node4260;
	wire [4-1:0] node4261;
	wire [4-1:0] node4262;
	wire [4-1:0] node4263;
	wire [4-1:0] node4266;
	wire [4-1:0] node4269;
	wire [4-1:0] node4270;
	wire [4-1:0] node4273;
	wire [4-1:0] node4276;
	wire [4-1:0] node4277;
	wire [4-1:0] node4278;
	wire [4-1:0] node4282;
	wire [4-1:0] node4285;
	wire [4-1:0] node4286;
	wire [4-1:0] node4287;
	wire [4-1:0] node4288;
	wire [4-1:0] node4289;
	wire [4-1:0] node4290;
	wire [4-1:0] node4291;
	wire [4-1:0] node4294;
	wire [4-1:0] node4298;
	wire [4-1:0] node4299;
	wire [4-1:0] node4301;
	wire [4-1:0] node4305;
	wire [4-1:0] node4307;
	wire [4-1:0] node4308;
	wire [4-1:0] node4309;
	wire [4-1:0] node4313;
	wire [4-1:0] node4314;
	wire [4-1:0] node4318;
	wire [4-1:0] node4319;
	wire [4-1:0] node4320;
	wire [4-1:0] node4321;
	wire [4-1:0] node4325;
	wire [4-1:0] node4326;
	wire [4-1:0] node4327;
	wire [4-1:0] node4332;
	wire [4-1:0] node4333;
	wire [4-1:0] node4335;
	wire [4-1:0] node4338;
	wire [4-1:0] node4339;
	wire [4-1:0] node4340;
	wire [4-1:0] node4344;
	wire [4-1:0] node4347;
	wire [4-1:0] node4348;
	wire [4-1:0] node4349;
	wire [4-1:0] node4350;
	wire [4-1:0] node4351;
	wire [4-1:0] node4353;
	wire [4-1:0] node4356;
	wire [4-1:0] node4358;
	wire [4-1:0] node4361;
	wire [4-1:0] node4362;
	wire [4-1:0] node4366;
	wire [4-1:0] node4367;
	wire [4-1:0] node4368;
	wire [4-1:0] node4369;
	wire [4-1:0] node4373;
	wire [4-1:0] node4375;
	wire [4-1:0] node4378;
	wire [4-1:0] node4379;
	wire [4-1:0] node4383;
	wire [4-1:0] node4384;
	wire [4-1:0] node4385;
	wire [4-1:0] node4387;
	wire [4-1:0] node4389;
	wire [4-1:0] node4392;
	wire [4-1:0] node4393;
	wire [4-1:0] node4395;
	wire [4-1:0] node4398;
	wire [4-1:0] node4400;
	wire [4-1:0] node4403;
	wire [4-1:0] node4404;
	wire [4-1:0] node4405;
	wire [4-1:0] node4406;
	wire [4-1:0] node4410;
	wire [4-1:0] node4411;
	wire [4-1:0] node4415;
	wire [4-1:0] node4417;
	wire [4-1:0] node4420;
	wire [4-1:0] node4421;
	wire [4-1:0] node4422;
	wire [4-1:0] node4423;
	wire [4-1:0] node4424;
	wire [4-1:0] node4425;
	wire [4-1:0] node4428;
	wire [4-1:0] node4429;
	wire [4-1:0] node4433;
	wire [4-1:0] node4434;
	wire [4-1:0] node4435;
	wire [4-1:0] node4438;
	wire [4-1:0] node4439;
	wire [4-1:0] node4442;
	wire [4-1:0] node4445;
	wire [4-1:0] node4446;
	wire [4-1:0] node4448;
	wire [4-1:0] node4451;
	wire [4-1:0] node4452;
	wire [4-1:0] node4456;
	wire [4-1:0] node4457;
	wire [4-1:0] node4458;
	wire [4-1:0] node4459;
	wire [4-1:0] node4460;
	wire [4-1:0] node4464;
	wire [4-1:0] node4466;
	wire [4-1:0] node4469;
	wire [4-1:0] node4470;
	wire [4-1:0] node4471;
	wire [4-1:0] node4475;
	wire [4-1:0] node4478;
	wire [4-1:0] node4479;
	wire [4-1:0] node4482;
	wire [4-1:0] node4483;
	wire [4-1:0] node4485;
	wire [4-1:0] node4488;
	wire [4-1:0] node4491;
	wire [4-1:0] node4492;
	wire [4-1:0] node4493;
	wire [4-1:0] node4494;
	wire [4-1:0] node4495;
	wire [4-1:0] node4496;
	wire [4-1:0] node4501;
	wire [4-1:0] node4502;
	wire [4-1:0] node4504;
	wire [4-1:0] node4507;
	wire [4-1:0] node4508;
	wire [4-1:0] node4511;
	wire [4-1:0] node4514;
	wire [4-1:0] node4515;
	wire [4-1:0] node4517;
	wire [4-1:0] node4519;
	wire [4-1:0] node4522;
	wire [4-1:0] node4523;
	wire [4-1:0] node4524;
	wire [4-1:0] node4527;
	wire [4-1:0] node4530;
	wire [4-1:0] node4532;
	wire [4-1:0] node4535;
	wire [4-1:0] node4536;
	wire [4-1:0] node4537;
	wire [4-1:0] node4538;
	wire [4-1:0] node4540;
	wire [4-1:0] node4543;
	wire [4-1:0] node4546;
	wire [4-1:0] node4547;
	wire [4-1:0] node4548;
	wire [4-1:0] node4553;
	wire [4-1:0] node4554;
	wire [4-1:0] node4555;
	wire [4-1:0] node4557;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4565;
	wire [4-1:0] node4567;
	wire [4-1:0] node4568;
	wire [4-1:0] node4571;
	wire [4-1:0] node4574;
	wire [4-1:0] node4575;
	wire [4-1:0] node4576;
	wire [4-1:0] node4577;
	wire [4-1:0] node4578;
	wire [4-1:0] node4579;
	wire [4-1:0] node4582;
	wire [4-1:0] node4585;
	wire [4-1:0] node4587;
	wire [4-1:0] node4588;
	wire [4-1:0] node4591;
	wire [4-1:0] node4594;
	wire [4-1:0] node4595;
	wire [4-1:0] node4596;
	wire [4-1:0] node4598;
	wire [4-1:0] node4601;
	wire [4-1:0] node4603;
	wire [4-1:0] node4606;
	wire [4-1:0] node4607;
	wire [4-1:0] node4609;
	wire [4-1:0] node4612;
	wire [4-1:0] node4615;
	wire [4-1:0] node4616;
	wire [4-1:0] node4617;
	wire [4-1:0] node4619;
	wire [4-1:0] node4621;
	wire [4-1:0] node4624;
	wire [4-1:0] node4625;
	wire [4-1:0] node4626;
	wire [4-1:0] node4630;
	wire [4-1:0] node4632;
	wire [4-1:0] node4635;
	wire [4-1:0] node4636;
	wire [4-1:0] node4637;
	wire [4-1:0] node4640;
	wire [4-1:0] node4643;
	wire [4-1:0] node4644;
	wire [4-1:0] node4646;
	wire [4-1:0] node4649;
	wire [4-1:0] node4650;
	wire [4-1:0] node4653;
	wire [4-1:0] node4656;
	wire [4-1:0] node4657;
	wire [4-1:0] node4658;
	wire [4-1:0] node4659;
	wire [4-1:0] node4660;
	wire [4-1:0] node4661;
	wire [4-1:0] node4665;
	wire [4-1:0] node4668;
	wire [4-1:0] node4669;
	wire [4-1:0] node4671;
	wire [4-1:0] node4674;
	wire [4-1:0] node4677;
	wire [4-1:0] node4678;
	wire [4-1:0] node4679;
	wire [4-1:0] node4681;
	wire [4-1:0] node4684;
	wire [4-1:0] node4687;
	wire [4-1:0] node4688;
	wire [4-1:0] node4691;
	wire [4-1:0] node4693;
	wire [4-1:0] node4696;
	wire [4-1:0] node4697;
	wire [4-1:0] node4698;
	wire [4-1:0] node4699;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4707;
	wire [4-1:0] node4709;
	wire [4-1:0] node4710;
	wire [4-1:0] node4714;
	wire [4-1:0] node4715;
	wire [4-1:0] node4716;
	wire [4-1:0] node4717;
	wire [4-1:0] node4721;
	wire [4-1:0] node4722;
	wire [4-1:0] node4725;
	wire [4-1:0] node4728;
	wire [4-1:0] node4729;
	wire [4-1:0] node4730;
	wire [4-1:0] node4734;
	wire [4-1:0] node4736;
	wire [4-1:0] node4739;
	wire [4-1:0] node4740;
	wire [4-1:0] node4741;
	wire [4-1:0] node4742;
	wire [4-1:0] node4743;
	wire [4-1:0] node4744;
	wire [4-1:0] node4745;
	wire [4-1:0] node4746;
	wire [4-1:0] node4747;
	wire [4-1:0] node4748;
	wire [4-1:0] node4751;
	wire [4-1:0] node4753;
	wire [4-1:0] node4756;
	wire [4-1:0] node4757;
	wire [4-1:0] node4758;
	wire [4-1:0] node4762;
	wire [4-1:0] node4765;
	wire [4-1:0] node4766;
	wire [4-1:0] node4767;
	wire [4-1:0] node4768;
	wire [4-1:0] node4769;
	wire [4-1:0] node4772;
	wire [4-1:0] node4775;
	wire [4-1:0] node4776;
	wire [4-1:0] node4779;
	wire [4-1:0] node4782;
	wire [4-1:0] node4784;
	wire [4-1:0] node4787;
	wire [4-1:0] node4788;
	wire [4-1:0] node4789;
	wire [4-1:0] node4791;
	wire [4-1:0] node4794;
	wire [4-1:0] node4797;
	wire [4-1:0] node4798;
	wire [4-1:0] node4799;
	wire [4-1:0] node4803;
	wire [4-1:0] node4806;
	wire [4-1:0] node4807;
	wire [4-1:0] node4808;
	wire [4-1:0] node4809;
	wire [4-1:0] node4811;
	wire [4-1:0] node4812;
	wire [4-1:0] node4815;
	wire [4-1:0] node4818;
	wire [4-1:0] node4820;
	wire [4-1:0] node4822;
	wire [4-1:0] node4825;
	wire [4-1:0] node4826;
	wire [4-1:0] node4827;
	wire [4-1:0] node4828;
	wire [4-1:0] node4831;
	wire [4-1:0] node4835;
	wire [4-1:0] node4836;
	wire [4-1:0] node4839;
	wire [4-1:0] node4840;
	wire [4-1:0] node4844;
	wire [4-1:0] node4845;
	wire [4-1:0] node4846;
	wire [4-1:0] node4847;
	wire [4-1:0] node4849;
	wire [4-1:0] node4852;
	wire [4-1:0] node4854;
	wire [4-1:0] node4857;
	wire [4-1:0] node4858;
	wire [4-1:0] node4861;
	wire [4-1:0] node4862;
	wire [4-1:0] node4865;
	wire [4-1:0] node4868;
	wire [4-1:0] node4869;
	wire [4-1:0] node4870;
	wire [4-1:0] node4872;
	wire [4-1:0] node4876;
	wire [4-1:0] node4877;
	wire [4-1:0] node4878;
	wire [4-1:0] node4881;
	wire [4-1:0] node4884;
	wire [4-1:0] node4886;
	wire [4-1:0] node4889;
	wire [4-1:0] node4890;
	wire [4-1:0] node4891;
	wire [4-1:0] node4892;
	wire [4-1:0] node4893;
	wire [4-1:0] node4894;
	wire [4-1:0] node4897;
	wire [4-1:0] node4898;
	wire [4-1:0] node4902;
	wire [4-1:0] node4903;
	wire [4-1:0] node4906;
	wire [4-1:0] node4909;
	wire [4-1:0] node4910;
	wire [4-1:0] node4911;
	wire [4-1:0] node4912;
	wire [4-1:0] node4916;
	wire [4-1:0] node4917;
	wire [4-1:0] node4920;
	wire [4-1:0] node4923;
	wire [4-1:0] node4924;
	wire [4-1:0] node4927;
	wire [4-1:0] node4930;
	wire [4-1:0] node4931;
	wire [4-1:0] node4932;
	wire [4-1:0] node4933;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4941;
	wire [4-1:0] node4942;
	wire [4-1:0] node4943;
	wire [4-1:0] node4946;
	wire [4-1:0] node4949;
	wire [4-1:0] node4950;
	wire [4-1:0] node4953;
	wire [4-1:0] node4956;
	wire [4-1:0] node4957;
	wire [4-1:0] node4959;
	wire [4-1:0] node4962;
	wire [4-1:0] node4964;
	wire [4-1:0] node4965;
	wire [4-1:0] node4968;
	wire [4-1:0] node4971;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4974;
	wire [4-1:0] node4975;
	wire [4-1:0] node4977;
	wire [4-1:0] node4981;
	wire [4-1:0] node4982;
	wire [4-1:0] node4985;
	wire [4-1:0] node4986;
	wire [4-1:0] node4990;
	wire [4-1:0] node4991;
	wire [4-1:0] node4992;
	wire [4-1:0] node4995;
	wire [4-1:0] node4996;
	wire [4-1:0] node5000;
	wire [4-1:0] node5002;
	wire [4-1:0] node5003;
	wire [4-1:0] node5006;
	wire [4-1:0] node5009;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5015;
	wire [4-1:0] node5016;
	wire [4-1:0] node5019;
	wire [4-1:0] node5022;
	wire [4-1:0] node5023;
	wire [4-1:0] node5024;
	wire [4-1:0] node5027;
	wire [4-1:0] node5030;
	wire [4-1:0] node5033;
	wire [4-1:0] node5034;
	wire [4-1:0] node5035;
	wire [4-1:0] node5036;
	wire [4-1:0] node5040;
	wire [4-1:0] node5041;
	wire [4-1:0] node5046;
	wire [4-1:0] node5047;
	wire [4-1:0] node5048;
	wire [4-1:0] node5049;
	wire [4-1:0] node5050;
	wire [4-1:0] node5051;
	wire [4-1:0] node5053;
	wire [4-1:0] node5054;
	wire [4-1:0] node5058;
	wire [4-1:0] node5059;
	wire [4-1:0] node5063;
	wire [4-1:0] node5064;
	wire [4-1:0] node5065;
	wire [4-1:0] node5066;
	wire [4-1:0] node5070;
	wire [4-1:0] node5071;
	wire [4-1:0] node5074;
	wire [4-1:0] node5077;
	wire [4-1:0] node5078;
	wire [4-1:0] node5082;
	wire [4-1:0] node5083;
	wire [4-1:0] node5084;
	wire [4-1:0] node5085;
	wire [4-1:0] node5086;
	wire [4-1:0] node5090;
	wire [4-1:0] node5093;
	wire [4-1:0] node5095;
	wire [4-1:0] node5098;
	wire [4-1:0] node5099;
	wire [4-1:0] node5100;
	wire [4-1:0] node5101;
	wire [4-1:0] node5105;
	wire [4-1:0] node5108;
	wire [4-1:0] node5111;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5114;
	wire [4-1:0] node5115;
	wire [4-1:0] node5116;
	wire [4-1:0] node5120;
	wire [4-1:0] node5122;
	wire [4-1:0] node5125;
	wire [4-1:0] node5127;
	wire [4-1:0] node5128;
	wire [4-1:0] node5131;
	wire [4-1:0] node5134;
	wire [4-1:0] node5135;
	wire [4-1:0] node5136;
	wire [4-1:0] node5139;
	wire [4-1:0] node5142;
	wire [4-1:0] node5143;
	wire [4-1:0] node5146;
	wire [4-1:0] node5149;
	wire [4-1:0] node5150;
	wire [4-1:0] node5151;
	wire [4-1:0] node5153;
	wire [4-1:0] node5154;
	wire [4-1:0] node5158;
	wire [4-1:0] node5159;
	wire [4-1:0] node5160;
	wire [4-1:0] node5163;
	wire [4-1:0] node5166;
	wire [4-1:0] node5168;
	wire [4-1:0] node5171;
	wire [4-1:0] node5172;
	wire [4-1:0] node5174;
	wire [4-1:0] node5177;
	wire [4-1:0] node5179;
	wire [4-1:0] node5182;
	wire [4-1:0] node5183;
	wire [4-1:0] node5184;
	wire [4-1:0] node5185;
	wire [4-1:0] node5186;
	wire [4-1:0] node5188;
	wire [4-1:0] node5191;
	wire [4-1:0] node5192;
	wire [4-1:0] node5195;
	wire [4-1:0] node5198;
	wire [4-1:0] node5199;
	wire [4-1:0] node5200;
	wire [4-1:0] node5204;
	wire [4-1:0] node5205;
	wire [4-1:0] node5206;
	wire [4-1:0] node5210;
	wire [4-1:0] node5211;
	wire [4-1:0] node5215;
	wire [4-1:0] node5216;
	wire [4-1:0] node5217;
	wire [4-1:0] node5220;
	wire [4-1:0] node5221;
	wire [4-1:0] node5223;
	wire [4-1:0] node5227;
	wire [4-1:0] node5230;
	wire [4-1:0] node5231;
	wire [4-1:0] node5232;
	wire [4-1:0] node5233;
	wire [4-1:0] node5234;
	wire [4-1:0] node5236;
	wire [4-1:0] node5239;
	wire [4-1:0] node5240;
	wire [4-1:0] node5243;
	wire [4-1:0] node5246;
	wire [4-1:0] node5247;
	wire [4-1:0] node5251;
	wire [4-1:0] node5252;
	wire [4-1:0] node5253;
	wire [4-1:0] node5254;
	wire [4-1:0] node5258;
	wire [4-1:0] node5259;
	wire [4-1:0] node5263;
	wire [4-1:0] node5264;
	wire [4-1:0] node5267;
	wire [4-1:0] node5268;
	wire [4-1:0] node5272;
	wire [4-1:0] node5273;
	wire [4-1:0] node5274;
	wire [4-1:0] node5275;
	wire [4-1:0] node5279;
	wire [4-1:0] node5280;
	wire [4-1:0] node5283;
	wire [4-1:0] node5286;
	wire [4-1:0] node5289;
	wire [4-1:0] node5290;
	wire [4-1:0] node5291;
	wire [4-1:0] node5292;
	wire [4-1:0] node5293;
	wire [4-1:0] node5294;
	wire [4-1:0] node5295;
	wire [4-1:0] node5296;
	wire [4-1:0] node5299;
	wire [4-1:0] node5300;
	wire [4-1:0] node5303;
	wire [4-1:0] node5306;
	wire [4-1:0] node5307;
	wire [4-1:0] node5311;
	wire [4-1:0] node5312;
	wire [4-1:0] node5313;
	wire [4-1:0] node5314;
	wire [4-1:0] node5318;
	wire [4-1:0] node5319;
	wire [4-1:0] node5322;
	wire [4-1:0] node5325;
	wire [4-1:0] node5326;
	wire [4-1:0] node5329;
	wire [4-1:0] node5330;
	wire [4-1:0] node5334;
	wire [4-1:0] node5335;
	wire [4-1:0] node5336;
	wire [4-1:0] node5338;
	wire [4-1:0] node5339;
	wire [4-1:0] node5342;
	wire [4-1:0] node5345;
	wire [4-1:0] node5346;
	wire [4-1:0] node5347;
	wire [4-1:0] node5351;
	wire [4-1:0] node5352;
	wire [4-1:0] node5355;
	wire [4-1:0] node5358;
	wire [4-1:0] node5359;
	wire [4-1:0] node5361;
	wire [4-1:0] node5364;
	wire [4-1:0] node5365;
	wire [4-1:0] node5366;
	wire [4-1:0] node5370;
	wire [4-1:0] node5373;
	wire [4-1:0] node5374;
	wire [4-1:0] node5375;
	wire [4-1:0] node5376;
	wire [4-1:0] node5377;
	wire [4-1:0] node5378;
	wire [4-1:0] node5382;
	wire [4-1:0] node5385;
	wire [4-1:0] node5386;
	wire [4-1:0] node5389;
	wire [4-1:0] node5392;
	wire [4-1:0] node5393;
	wire [4-1:0] node5394;
	wire [4-1:0] node5396;
	wire [4-1:0] node5399;
	wire [4-1:0] node5401;
	wire [4-1:0] node5404;
	wire [4-1:0] node5405;
	wire [4-1:0] node5407;
	wire [4-1:0] node5410;
	wire [4-1:0] node5413;
	wire [4-1:0] node5414;
	wire [4-1:0] node5415;
	wire [4-1:0] node5417;
	wire [4-1:0] node5418;
	wire [4-1:0] node5422;
	wire [4-1:0] node5423;
	wire [4-1:0] node5425;
	wire [4-1:0] node5429;
	wire [4-1:0] node5430;
	wire [4-1:0] node5432;
	wire [4-1:0] node5435;
	wire [4-1:0] node5436;
	wire [4-1:0] node5439;
	wire [4-1:0] node5440;
	wire [4-1:0] node5444;
	wire [4-1:0] node5445;
	wire [4-1:0] node5446;
	wire [4-1:0] node5447;
	wire [4-1:0] node5448;
	wire [4-1:0] node5449;
	wire [4-1:0] node5452;
	wire [4-1:0] node5453;
	wire [4-1:0] node5456;
	wire [4-1:0] node5459;
	wire [4-1:0] node5460;
	wire [4-1:0] node5463;
	wire [4-1:0] node5466;
	wire [4-1:0] node5467;
	wire [4-1:0] node5468;
	wire [4-1:0] node5470;
	wire [4-1:0] node5473;
	wire [4-1:0] node5476;
	wire [4-1:0] node5477;
	wire [4-1:0] node5479;
	wire [4-1:0] node5482;
	wire [4-1:0] node5484;
	wire [4-1:0] node5487;
	wire [4-1:0] node5488;
	wire [4-1:0] node5489;
	wire [4-1:0] node5490;
	wire [4-1:0] node5494;
	wire [4-1:0] node5496;
	wire [4-1:0] node5499;
	wire [4-1:0] node5500;
	wire [4-1:0] node5501;
	wire [4-1:0] node5503;
	wire [4-1:0] node5506;
	wire [4-1:0] node5507;
	wire [4-1:0] node5511;
	wire [4-1:0] node5512;
	wire [4-1:0] node5513;
	wire [4-1:0] node5517;
	wire [4-1:0] node5520;
	wire [4-1:0] node5521;
	wire [4-1:0] node5522;
	wire [4-1:0] node5523;
	wire [4-1:0] node5524;
	wire [4-1:0] node5526;
	wire [4-1:0] node5529;
	wire [4-1:0] node5531;
	wire [4-1:0] node5534;
	wire [4-1:0] node5535;
	wire [4-1:0] node5538;
	wire [4-1:0] node5541;
	wire [4-1:0] node5542;
	wire [4-1:0] node5543;
	wire [4-1:0] node5546;
	wire [4-1:0] node5548;
	wire [4-1:0] node5551;
	wire [4-1:0] node5552;
	wire [4-1:0] node5554;
	wire [4-1:0] node5557;
	wire [4-1:0] node5558;
	wire [4-1:0] node5561;
	wire [4-1:0] node5564;
	wire [4-1:0] node5565;
	wire [4-1:0] node5566;
	wire [4-1:0] node5567;
	wire [4-1:0] node5569;
	wire [4-1:0] node5572;
	wire [4-1:0] node5574;
	wire [4-1:0] node5577;
	wire [4-1:0] node5578;
	wire [4-1:0] node5579;
	wire [4-1:0] node5582;
	wire [4-1:0] node5585;
	wire [4-1:0] node5587;
	wire [4-1:0] node5590;
	wire [4-1:0] node5591;
	wire [4-1:0] node5592;
	wire [4-1:0] node5595;
	wire [4-1:0] node5597;
	wire [4-1:0] node5600;
	wire [4-1:0] node5603;
	wire [4-1:0] node5604;
	wire [4-1:0] node5605;
	wire [4-1:0] node5606;
	wire [4-1:0] node5607;
	wire [4-1:0] node5608;
	wire [4-1:0] node5609;
	wire [4-1:0] node5611;
	wire [4-1:0] node5614;
	wire [4-1:0] node5617;
	wire [4-1:0] node5619;
	wire [4-1:0] node5620;
	wire [4-1:0] node5624;
	wire [4-1:0] node5625;
	wire [4-1:0] node5627;
	wire [4-1:0] node5629;
	wire [4-1:0] node5632;
	wire [4-1:0] node5633;
	wire [4-1:0] node5636;
	wire [4-1:0] node5639;
	wire [4-1:0] node5640;
	wire [4-1:0] node5641;
	wire [4-1:0] node5642;
	wire [4-1:0] node5645;
	wire [4-1:0] node5647;
	wire [4-1:0] node5650;
	wire [4-1:0] node5651;
	wire [4-1:0] node5652;
	wire [4-1:0] node5656;
	wire [4-1:0] node5659;
	wire [4-1:0] node5660;
	wire [4-1:0] node5661;
	wire [4-1:0] node5664;
	wire [4-1:0] node5667;
	wire [4-1:0] node5668;
	wire [4-1:0] node5669;
	wire [4-1:0] node5674;
	wire [4-1:0] node5675;
	wire [4-1:0] node5676;
	wire [4-1:0] node5677;
	wire [4-1:0] node5680;
	wire [4-1:0] node5681;
	wire [4-1:0] node5684;
	wire [4-1:0] node5687;
	wire [4-1:0] node5688;
	wire [4-1:0] node5689;
	wire [4-1:0] node5691;
	wire [4-1:0] node5694;
	wire [4-1:0] node5696;
	wire [4-1:0] node5699;
	wire [4-1:0] node5700;
	wire [4-1:0] node5701;
	wire [4-1:0] node5705;
	wire [4-1:0] node5708;
	wire [4-1:0] node5709;
	wire [4-1:0] node5710;
	wire [4-1:0] node5711;
	wire [4-1:0] node5712;
	wire [4-1:0] node5715;
	wire [4-1:0] node5718;
	wire [4-1:0] node5720;
	wire [4-1:0] node5723;
	wire [4-1:0] node5724;
	wire [4-1:0] node5725;
	wire [4-1:0] node5729;
	wire [4-1:0] node5732;
	wire [4-1:0] node5733;
	wire [4-1:0] node5734;
	wire [4-1:0] node5737;
	wire [4-1:0] node5740;
	wire [4-1:0] node5741;
	wire [4-1:0] node5742;
	wire [4-1:0] node5746;
	wire [4-1:0] node5747;
	wire [4-1:0] node5751;
	wire [4-1:0] node5752;
	wire [4-1:0] node5753;
	wire [4-1:0] node5754;
	wire [4-1:0] node5755;
	wire [4-1:0] node5756;
	wire [4-1:0] node5758;
	wire [4-1:0] node5761;
	wire [4-1:0] node5762;
	wire [4-1:0] node5766;
	wire [4-1:0] node5767;
	wire [4-1:0] node5768;
	wire [4-1:0] node5771;
	wire [4-1:0] node5774;
	wire [4-1:0] node5775;
	wire [4-1:0] node5779;
	wire [4-1:0] node5780;
	wire [4-1:0] node5781;
	wire [4-1:0] node5784;
	wire [4-1:0] node5787;
	wire [4-1:0] node5788;
	wire [4-1:0] node5789;
	wire [4-1:0] node5793;
	wire [4-1:0] node5796;
	wire [4-1:0] node5797;
	wire [4-1:0] node5798;
	wire [4-1:0] node5799;
	wire [4-1:0] node5802;
	wire [4-1:0] node5803;
	wire [4-1:0] node5806;
	wire [4-1:0] node5809;
	wire [4-1:0] node5810;
	wire [4-1:0] node5813;
	wire [4-1:0] node5816;
	wire [4-1:0] node5817;
	wire [4-1:0] node5818;
	wire [4-1:0] node5819;
	wire [4-1:0] node5823;
	wire [4-1:0] node5824;
	wire [4-1:0] node5828;
	wire [4-1:0] node5829;
	wire [4-1:0] node5831;
	wire [4-1:0] node5834;
	wire [4-1:0] node5837;
	wire [4-1:0] node5838;
	wire [4-1:0] node5839;
	wire [4-1:0] node5840;
	wire [4-1:0] node5841;
	wire [4-1:0] node5844;
	wire [4-1:0] node5846;
	wire [4-1:0] node5849;
	wire [4-1:0] node5850;
	wire [4-1:0] node5852;
	wire [4-1:0] node5855;
	wire [4-1:0] node5858;
	wire [4-1:0] node5859;
	wire [4-1:0] node5860;
	wire [4-1:0] node5861;
	wire [4-1:0] node5864;
	wire [4-1:0] node5867;
	wire [4-1:0] node5868;
	wire [4-1:0] node5872;
	wire [4-1:0] node5873;
	wire [4-1:0] node5874;
	wire [4-1:0] node5878;
	wire [4-1:0] node5881;
	wire [4-1:0] node5882;
	wire [4-1:0] node5883;
	wire [4-1:0] node5884;
	wire [4-1:0] node5888;
	wire [4-1:0] node5889;
	wire [4-1:0] node5890;
	wire [4-1:0] node5894;
	wire [4-1:0] node5897;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5902;
	wire [4-1:0] node5903;
	wire [4-1:0] node5906;
	wire [4-1:0] node5909;
	wire [4-1:0] node5912;
	wire [4-1:0] node5913;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5916;
	wire [4-1:0] node5917;
	wire [4-1:0] node5918;
	wire [4-1:0] node5920;
	wire [4-1:0] node5923;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5928;
	wire [4-1:0] node5930;
	wire [4-1:0] node5933;
	wire [4-1:0] node5935;
	wire [4-1:0] node5938;
	wire [4-1:0] node5939;
	wire [4-1:0] node5941;
	wire [4-1:0] node5942;
	wire [4-1:0] node5945;
	wire [4-1:0] node5946;
	wire [4-1:0] node5950;
	wire [4-1:0] node5951;
	wire [4-1:0] node5952;
	wire [4-1:0] node5954;
	wire [4-1:0] node5957;
	wire [4-1:0] node5960;
	wire [4-1:0] node5961;
	wire [4-1:0] node5963;
	wire [4-1:0] node5966;
	wire [4-1:0] node5969;
	wire [4-1:0] node5970;
	wire [4-1:0] node5971;
	wire [4-1:0] node5974;
	wire [4-1:0] node5975;
	wire [4-1:0] node5976;
	wire [4-1:0] node5980;
	wire [4-1:0] node5981;
	wire [4-1:0] node5982;
	wire [4-1:0] node5986;
	wire [4-1:0] node5989;
	wire [4-1:0] node5990;
	wire [4-1:0] node5991;
	wire [4-1:0] node5992;
	wire [4-1:0] node5995;
	wire [4-1:0] node5996;
	wire [4-1:0] node6000;
	wire [4-1:0] node6001;
	wire [4-1:0] node6003;
	wire [4-1:0] node6006;
	wire [4-1:0] node6007;
	wire [4-1:0] node6010;
	wire [4-1:0] node6013;
	wire [4-1:0] node6014;
	wire [4-1:0] node6015;
	wire [4-1:0] node6018;
	wire [4-1:0] node6020;
	wire [4-1:0] node6023;
	wire [4-1:0] node6024;
	wire [4-1:0] node6025;
	wire [4-1:0] node6030;
	wire [4-1:0] node6031;
	wire [4-1:0] node6032;
	wire [4-1:0] node6033;
	wire [4-1:0] node6034;
	wire [4-1:0] node6035;
	wire [4-1:0] node6038;
	wire [4-1:0] node6039;
	wire [4-1:0] node6043;
	wire [4-1:0] node6045;
	wire [4-1:0] node6047;
	wire [4-1:0] node6050;
	wire [4-1:0] node6051;
	wire [4-1:0] node6052;
	wire [4-1:0] node6053;
	wire [4-1:0] node6057;
	wire [4-1:0] node6058;
	wire [4-1:0] node6062;
	wire [4-1:0] node6063;
	wire [4-1:0] node6066;
	wire [4-1:0] node6069;
	wire [4-1:0] node6070;
	wire [4-1:0] node6071;
	wire [4-1:0] node6072;
	wire [4-1:0] node6073;
	wire [4-1:0] node6077;
	wire [4-1:0] node6079;
	wire [4-1:0] node6082;
	wire [4-1:0] node6083;
	wire [4-1:0] node6085;
	wire [4-1:0] node6088;
	wire [4-1:0] node6091;
	wire [4-1:0] node6092;
	wire [4-1:0] node6093;
	wire [4-1:0] node6094;
	wire [4-1:0] node6097;
	wire [4-1:0] node6100;
	wire [4-1:0] node6103;
	wire [4-1:0] node6104;
	wire [4-1:0] node6107;
	wire [4-1:0] node6108;
	wire [4-1:0] node6112;
	wire [4-1:0] node6113;
	wire [4-1:0] node6114;
	wire [4-1:0] node6115;
	wire [4-1:0] node6117;
	wire [4-1:0] node6119;
	wire [4-1:0] node6122;
	wire [4-1:0] node6124;
	wire [4-1:0] node6126;
	wire [4-1:0] node6129;
	wire [4-1:0] node6130;
	wire [4-1:0] node6131;
	wire [4-1:0] node6134;
	wire [4-1:0] node6136;
	wire [4-1:0] node6139;
	wire [4-1:0] node6140;
	wire [4-1:0] node6141;
	wire [4-1:0] node6144;
	wire [4-1:0] node6147;
	wire [4-1:0] node6148;
	wire [4-1:0] node6151;
	wire [4-1:0] node6154;
	wire [4-1:0] node6155;
	wire [4-1:0] node6156;
	wire [4-1:0] node6158;
	wire [4-1:0] node6161;
	wire [4-1:0] node6162;
	wire [4-1:0] node6164;
	wire [4-1:0] node6167;
	wire [4-1:0] node6169;
	wire [4-1:0] node6172;
	wire [4-1:0] node6174;
	wire [4-1:0] node6175;
	wire [4-1:0] node6177;
	wire [4-1:0] node6181;
	wire [4-1:0] node6182;
	wire [4-1:0] node6183;
	wire [4-1:0] node6184;
	wire [4-1:0] node6185;
	wire [4-1:0] node6186;
	wire [4-1:0] node6187;
	wire [4-1:0] node6189;
	wire [4-1:0] node6192;
	wire [4-1:0] node6193;
	wire [4-1:0] node6196;
	wire [4-1:0] node6199;
	wire [4-1:0] node6200;
	wire [4-1:0] node6201;
	wire [4-1:0] node6204;
	wire [4-1:0] node6207;
	wire [4-1:0] node6209;
	wire [4-1:0] node6212;
	wire [4-1:0] node6213;
	wire [4-1:0] node6214;
	wire [4-1:0] node6215;
	wire [4-1:0] node6218;
	wire [4-1:0] node6221;
	wire [4-1:0] node6222;
	wire [4-1:0] node6226;
	wire [4-1:0] node6227;
	wire [4-1:0] node6228;
	wire [4-1:0] node6231;
	wire [4-1:0] node6234;
	wire [4-1:0] node6235;
	wire [4-1:0] node6238;
	wire [4-1:0] node6241;
	wire [4-1:0] node6242;
	wire [4-1:0] node6243;
	wire [4-1:0] node6244;
	wire [4-1:0] node6246;
	wire [4-1:0] node6250;
	wire [4-1:0] node6251;
	wire [4-1:0] node6252;
	wire [4-1:0] node6255;
	wire [4-1:0] node6258;
	wire [4-1:0] node6261;
	wire [4-1:0] node6262;
	wire [4-1:0] node6263;
	wire [4-1:0] node6264;
	wire [4-1:0] node6268;
	wire [4-1:0] node6271;
	wire [4-1:0] node6272;
	wire [4-1:0] node6275;
	wire [4-1:0] node6277;
	wire [4-1:0] node6280;
	wire [4-1:0] node6281;
	wire [4-1:0] node6282;
	wire [4-1:0] node6283;
	wire [4-1:0] node6284;
	wire [4-1:0] node6286;
	wire [4-1:0] node6289;
	wire [4-1:0] node6292;
	wire [4-1:0] node6293;
	wire [4-1:0] node6294;
	wire [4-1:0] node6298;
	wire [4-1:0] node6299;
	wire [4-1:0] node6302;
	wire [4-1:0] node6305;
	wire [4-1:0] node6306;
	wire [4-1:0] node6307;
	wire [4-1:0] node6308;
	wire [4-1:0] node6312;
	wire [4-1:0] node6315;
	wire [4-1:0] node6316;
	wire [4-1:0] node6319;
	wire [4-1:0] node6321;
	wire [4-1:0] node6324;
	wire [4-1:0] node6325;
	wire [4-1:0] node6326;
	wire [4-1:0] node6327;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6335;
	wire [4-1:0] node6336;
	wire [4-1:0] node6337;
	wire [4-1:0] node6341;
	wire [4-1:0] node6342;
	wire [4-1:0] node6345;
	wire [4-1:0] node6348;
	wire [4-1:0] node6349;
	wire [4-1:0] node6350;
	wire [4-1:0] node6352;
	wire [4-1:0] node6355;
	wire [4-1:0] node6358;
	wire [4-1:0] node6359;
	wire [4-1:0] node6361;
	wire [4-1:0] node6364;
	wire [4-1:0] node6367;
	wire [4-1:0] node6368;
	wire [4-1:0] node6369;
	wire [4-1:0] node6370;
	wire [4-1:0] node6371;
	wire [4-1:0] node6372;
	wire [4-1:0] node6373;
	wire [4-1:0] node6378;
	wire [4-1:0] node6379;
	wire [4-1:0] node6381;
	wire [4-1:0] node6384;
	wire [4-1:0] node6385;
	wire [4-1:0] node6389;
	wire [4-1:0] node6391;
	wire [4-1:0] node6392;
	wire [4-1:0] node6394;
	wire [4-1:0] node6397;
	wire [4-1:0] node6398;
	wire [4-1:0] node6402;
	wire [4-1:0] node6403;
	wire [4-1:0] node6404;
	wire [4-1:0] node6405;
	wire [4-1:0] node6407;
	wire [4-1:0] node6410;
	wire [4-1:0] node6411;
	wire [4-1:0] node6415;
	wire [4-1:0] node6416;
	wire [4-1:0] node6417;
	wire [4-1:0] node6421;
	wire [4-1:0] node6424;
	wire [4-1:0] node6425;
	wire [4-1:0] node6426;
	wire [4-1:0] node6427;
	wire [4-1:0] node6431;
	wire [4-1:0] node6433;
	wire [4-1:0] node6436;
	wire [4-1:0] node6438;
	wire [4-1:0] node6439;
	wire [4-1:0] node6443;
	wire [4-1:0] node6444;
	wire [4-1:0] node6445;
	wire [4-1:0] node6446;
	wire [4-1:0] node6447;
	wire [4-1:0] node6448;
	wire [4-1:0] node6451;
	wire [4-1:0] node6454;
	wire [4-1:0] node6456;
	wire [4-1:0] node6459;
	wire [4-1:0] node6460;
	wire [4-1:0] node6461;
	wire [4-1:0] node6464;
	wire [4-1:0] node6467;
	wire [4-1:0] node6468;
	wire [4-1:0] node6471;
	wire [4-1:0] node6474;
	wire [4-1:0] node6475;
	wire [4-1:0] node6476;
	wire [4-1:0] node6478;
	wire [4-1:0] node6481;
	wire [4-1:0] node6482;
	wire [4-1:0] node6485;
	wire [4-1:0] node6488;
	wire [4-1:0] node6489;
	wire [4-1:0] node6491;
	wire [4-1:0] node6494;
	wire [4-1:0] node6496;
	wire [4-1:0] node6499;
	wire [4-1:0] node6500;
	wire [4-1:0] node6501;
	wire [4-1:0] node6502;
	wire [4-1:0] node6505;
	wire [4-1:0] node6506;
	wire [4-1:0] node6510;
	wire [4-1:0] node6511;
	wire [4-1:0] node6514;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6519;
	wire [4-1:0] node6522;
	wire [4-1:0] node6524;
	wire [4-1:0] node6527;
	wire [4-1:0] node6528;
	wire [4-1:0] node6530;
	wire [4-1:0] node6533;
	wire [4-1:0] node6536;
	wire [4-1:0] node6537;
	wire [4-1:0] node6538;
	wire [4-1:0] node6539;
	wire [4-1:0] node6540;
	wire [4-1:0] node6541;
	wire [4-1:0] node6542;
	wire [4-1:0] node6544;
	wire [4-1:0] node6545;
	wire [4-1:0] node6549;
	wire [4-1:0] node6550;
	wire [4-1:0] node6553;
	wire [4-1:0] node6555;
	wire [4-1:0] node6558;
	wire [4-1:0] node6559;
	wire [4-1:0] node6560;
	wire [4-1:0] node6563;
	wire [4-1:0] node6566;
	wire [4-1:0] node6567;
	wire [4-1:0] node6568;
	wire [4-1:0] node6572;
	wire [4-1:0] node6574;
	wire [4-1:0] node6577;
	wire [4-1:0] node6578;
	wire [4-1:0] node6579;
	wire [4-1:0] node6580;
	wire [4-1:0] node6583;
	wire [4-1:0] node6584;
	wire [4-1:0] node6588;
	wire [4-1:0] node6589;
	wire [4-1:0] node6590;
	wire [4-1:0] node6594;
	wire [4-1:0] node6595;
	wire [4-1:0] node6598;
	wire [4-1:0] node6601;
	wire [4-1:0] node6602;
	wire [4-1:0] node6603;
	wire [4-1:0] node6604;
	wire [4-1:0] node6608;
	wire [4-1:0] node6611;
	wire [4-1:0] node6613;
	wire [4-1:0] node6616;
	wire [4-1:0] node6617;
	wire [4-1:0] node6618;
	wire [4-1:0] node6619;
	wire [4-1:0] node6621;
	wire [4-1:0] node6624;
	wire [4-1:0] node6625;
	wire [4-1:0] node6628;
	wire [4-1:0] node6629;
	wire [4-1:0] node6632;
	wire [4-1:0] node6635;
	wire [4-1:0] node6636;
	wire [4-1:0] node6637;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6645;
	wire [4-1:0] node6646;
	wire [4-1:0] node6647;
	wire [4-1:0] node6652;
	wire [4-1:0] node6653;
	wire [4-1:0] node6654;
	wire [4-1:0] node6655;
	wire [4-1:0] node6656;
	wire [4-1:0] node6660;
	wire [4-1:0] node6661;
	wire [4-1:0] node6664;
	wire [4-1:0] node6667;
	wire [4-1:0] node6668;
	wire [4-1:0] node6671;
	wire [4-1:0] node6672;
	wire [4-1:0] node6676;
	wire [4-1:0] node6677;
	wire [4-1:0] node6679;
	wire [4-1:0] node6682;
	wire [4-1:0] node6684;
	wire [4-1:0] node6686;
	wire [4-1:0] node6689;
	wire [4-1:0] node6690;
	wire [4-1:0] node6691;
	wire [4-1:0] node6692;
	wire [4-1:0] node6693;
	wire [4-1:0] node6696;
	wire [4-1:0] node6697;
	wire [4-1:0] node6698;
	wire [4-1:0] node6701;
	wire [4-1:0] node6704;
	wire [4-1:0] node6705;
	wire [4-1:0] node6709;
	wire [4-1:0] node6710;
	wire [4-1:0] node6711;
	wire [4-1:0] node6714;
	wire [4-1:0] node6715;
	wire [4-1:0] node6719;
	wire [4-1:0] node6720;
	wire [4-1:0] node6721;
	wire [4-1:0] node6725;
	wire [4-1:0] node6728;
	wire [4-1:0] node6729;
	wire [4-1:0] node6730;
	wire [4-1:0] node6731;
	wire [4-1:0] node6735;
	wire [4-1:0] node6736;
	wire [4-1:0] node6737;
	wire [4-1:0] node6740;
	wire [4-1:0] node6743;
	wire [4-1:0] node6746;
	wire [4-1:0] node6747;
	wire [4-1:0] node6748;
	wire [4-1:0] node6751;
	wire [4-1:0] node6754;
	wire [4-1:0] node6755;
	wire [4-1:0] node6756;
	wire [4-1:0] node6759;
	wire [4-1:0] node6763;
	wire [4-1:0] node6764;
	wire [4-1:0] node6765;
	wire [4-1:0] node6766;
	wire [4-1:0] node6767;
	wire [4-1:0] node6769;
	wire [4-1:0] node6773;
	wire [4-1:0] node6774;
	wire [4-1:0] node6776;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6783;
	wire [4-1:0] node6786;
	wire [4-1:0] node6787;
	wire [4-1:0] node6788;
	wire [4-1:0] node6789;
	wire [4-1:0] node6792;
	wire [4-1:0] node6795;
	wire [4-1:0] node6798;
	wire [4-1:0] node6799;
	wire [4-1:0] node6802;
	wire [4-1:0] node6803;
	wire [4-1:0] node6806;
	wire [4-1:0] node6809;
	wire [4-1:0] node6810;
	wire [4-1:0] node6811;
	wire [4-1:0] node6812;
	wire [4-1:0] node6813;
	wire [4-1:0] node6817;
	wire [4-1:0] node6819;
	wire [4-1:0] node6822;
	wire [4-1:0] node6824;
	wire [4-1:0] node6827;
	wire [4-1:0] node6828;
	wire [4-1:0] node6829;
	wire [4-1:0] node6830;
	wire [4-1:0] node6834;
	wire [4-1:0] node6837;
	wire [4-1:0] node6838;
	wire [4-1:0] node6840;
	wire [4-1:0] node6844;
	wire [4-1:0] node6845;
	wire [4-1:0] node6846;
	wire [4-1:0] node6847;
	wire [4-1:0] node6848;
	wire [4-1:0] node6849;
	wire [4-1:0] node6851;
	wire [4-1:0] node6854;
	wire [4-1:0] node6856;
	wire [4-1:0] node6859;
	wire [4-1:0] node6860;
	wire [4-1:0] node6861;
	wire [4-1:0] node6864;
	wire [4-1:0] node6865;
	wire [4-1:0] node6869;
	wire [4-1:0] node6870;
	wire [4-1:0] node6871;
	wire [4-1:0] node6874;
	wire [4-1:0] node6877;
	wire [4-1:0] node6879;
	wire [4-1:0] node6882;
	wire [4-1:0] node6883;
	wire [4-1:0] node6884;
	wire [4-1:0] node6885;
	wire [4-1:0] node6886;
	wire [4-1:0] node6890;
	wire [4-1:0] node6891;
	wire [4-1:0] node6894;
	wire [4-1:0] node6897;
	wire [4-1:0] node6898;
	wire [4-1:0] node6901;
	wire [4-1:0] node6904;
	wire [4-1:0] node6905;
	wire [4-1:0] node6906;
	wire [4-1:0] node6907;
	wire [4-1:0] node6910;
	wire [4-1:0] node6913;
	wire [4-1:0] node6914;
	wire [4-1:0] node6918;
	wire [4-1:0] node6919;
	wire [4-1:0] node6920;
	wire [4-1:0] node6923;
	wire [4-1:0] node6926;
	wire [4-1:0] node6927;
	wire [4-1:0] node6931;
	wire [4-1:0] node6932;
	wire [4-1:0] node6933;
	wire [4-1:0] node6934;
	wire [4-1:0] node6937;
	wire [4-1:0] node6938;
	wire [4-1:0] node6939;
	wire [4-1:0] node6943;
	wire [4-1:0] node6946;
	wire [4-1:0] node6947;
	wire [4-1:0] node6949;
	wire [4-1:0] node6951;
	wire [4-1:0] node6954;
	wire [4-1:0] node6955;
	wire [4-1:0] node6956;
	wire [4-1:0] node6959;
	wire [4-1:0] node6962;
	wire [4-1:0] node6965;
	wire [4-1:0] node6966;
	wire [4-1:0] node6967;
	wire [4-1:0] node6968;
	wire [4-1:0] node6969;
	wire [4-1:0] node6972;
	wire [4-1:0] node6976;
	wire [4-1:0] node6978;
	wire [4-1:0] node6980;
	wire [4-1:0] node6983;
	wire [4-1:0] node6984;
	wire [4-1:0] node6985;
	wire [4-1:0] node6986;
	wire [4-1:0] node6989;
	wire [4-1:0] node6993;
	wire [4-1:0] node6994;
	wire [4-1:0] node6995;
	wire [4-1:0] node7000;
	wire [4-1:0] node7001;
	wire [4-1:0] node7002;
	wire [4-1:0] node7003;
	wire [4-1:0] node7004;
	wire [4-1:0] node7005;
	wire [4-1:0] node7008;
	wire [4-1:0] node7011;
	wire [4-1:0] node7013;
	wire [4-1:0] node7014;
	wire [4-1:0] node7017;
	wire [4-1:0] node7020;
	wire [4-1:0] node7021;
	wire [4-1:0] node7022;
	wire [4-1:0] node7023;
	wire [4-1:0] node7026;
	wire [4-1:0] node7029;
	wire [4-1:0] node7030;
	wire [4-1:0] node7033;
	wire [4-1:0] node7036;
	wire [4-1:0] node7037;
	wire [4-1:0] node7040;
	wire [4-1:0] node7043;
	wire [4-1:0] node7044;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7048;
	wire [4-1:0] node7051;
	wire [4-1:0] node7053;
	wire [4-1:0] node7056;
	wire [4-1:0] node7057;
	wire [4-1:0] node7060;
	wire [4-1:0] node7061;
	wire [4-1:0] node7064;
	wire [4-1:0] node7067;
	wire [4-1:0] node7068;
	wire [4-1:0] node7069;
	wire [4-1:0] node7070;
	wire [4-1:0] node7074;
	wire [4-1:0] node7075;
	wire [4-1:0] node7079;
	wire [4-1:0] node7080;
	wire [4-1:0] node7083;
	wire [4-1:0] node7086;
	wire [4-1:0] node7087;
	wire [4-1:0] node7088;
	wire [4-1:0] node7089;
	wire [4-1:0] node7090;
	wire [4-1:0] node7093;
	wire [4-1:0] node7096;
	wire [4-1:0] node7097;
	wire [4-1:0] node7098;
	wire [4-1:0] node7102;
	wire [4-1:0] node7104;
	wire [4-1:0] node7107;
	wire [4-1:0] node7108;
	wire [4-1:0] node7109;
	wire [4-1:0] node7110;
	wire [4-1:0] node7113;
	wire [4-1:0] node7116;
	wire [4-1:0] node7117;
	wire [4-1:0] node7121;
	wire [4-1:0] node7122;
	wire [4-1:0] node7125;
	wire [4-1:0] node7127;
	wire [4-1:0] node7130;
	wire [4-1:0] node7131;
	wire [4-1:0] node7132;
	wire [4-1:0] node7133;
	wire [4-1:0] node7134;
	wire [4-1:0] node7137;
	wire [4-1:0] node7140;
	wire [4-1:0] node7143;
	wire [4-1:0] node7144;
	wire [4-1:0] node7147;
	wire [4-1:0] node7150;
	wire [4-1:0] node7151;
	wire [4-1:0] node7152;
	wire [4-1:0] node7153;
	wire [4-1:0] node7156;
	wire [4-1:0] node7159;
	wire [4-1:0] node7160;
	wire [4-1:0] node7163;
	wire [4-1:0] node7166;
	wire [4-1:0] node7168;
	wire [4-1:0] node7171;
	wire [4-1:0] node7172;
	wire [4-1:0] node7173;
	wire [4-1:0] node7174;
	wire [4-1:0] node7175;
	wire [4-1:0] node7176;
	wire [4-1:0] node7177;
	wire [4-1:0] node7178;
	wire [4-1:0] node7181;
	wire [4-1:0] node7182;
	wire [4-1:0] node7183;
	wire [4-1:0] node7186;
	wire [4-1:0] node7189;
	wire [4-1:0] node7190;
	wire [4-1:0] node7191;
	wire [4-1:0] node7196;
	wire [4-1:0] node7197;
	wire [4-1:0] node7200;
	wire [4-1:0] node7201;
	wire [4-1:0] node7202;
	wire [4-1:0] node7203;
	wire [4-1:0] node7206;
	wire [4-1:0] node7209;
	wire [4-1:0] node7210;
	wire [4-1:0] node7213;
	wire [4-1:0] node7216;
	wire [4-1:0] node7217;
	wire [4-1:0] node7220;
	wire [4-1:0] node7223;
	wire [4-1:0] node7224;
	wire [4-1:0] node7225;
	wire [4-1:0] node7226;
	wire [4-1:0] node7227;
	wire [4-1:0] node7228;
	wire [4-1:0] node7232;
	wire [4-1:0] node7234;
	wire [4-1:0] node7237;
	wire [4-1:0] node7238;
	wire [4-1:0] node7241;
	wire [4-1:0] node7244;
	wire [4-1:0] node7245;
	wire [4-1:0] node7246;
	wire [4-1:0] node7249;
	wire [4-1:0] node7252;
	wire [4-1:0] node7253;
	wire [4-1:0] node7256;
	wire [4-1:0] node7258;
	wire [4-1:0] node7261;
	wire [4-1:0] node7262;
	wire [4-1:0] node7263;
	wire [4-1:0] node7266;
	wire [4-1:0] node7267;
	wire [4-1:0] node7270;
	wire [4-1:0] node7271;
	wire [4-1:0] node7275;
	wire [4-1:0] node7276;
	wire [4-1:0] node7279;
	wire [4-1:0] node7280;
	wire [4-1:0] node7282;
	wire [4-1:0] node7285;
	wire [4-1:0] node7288;
	wire [4-1:0] node7289;
	wire [4-1:0] node7290;
	wire [4-1:0] node7291;
	wire [4-1:0] node7292;
	wire [4-1:0] node7293;
	wire [4-1:0] node7294;
	wire [4-1:0] node7297;
	wire [4-1:0] node7300;
	wire [4-1:0] node7301;
	wire [4-1:0] node7304;
	wire [4-1:0] node7307;
	wire [4-1:0] node7308;
	wire [4-1:0] node7309;
	wire [4-1:0] node7312;
	wire [4-1:0] node7315;
	wire [4-1:0] node7316;
	wire [4-1:0] node7320;
	wire [4-1:0] node7321;
	wire [4-1:0] node7323;
	wire [4-1:0] node7324;
	wire [4-1:0] node7327;
	wire [4-1:0] node7330;
	wire [4-1:0] node7332;
	wire [4-1:0] node7334;
	wire [4-1:0] node7337;
	wire [4-1:0] node7338;
	wire [4-1:0] node7339;
	wire [4-1:0] node7341;
	wire [4-1:0] node7344;
	wire [4-1:0] node7345;
	wire [4-1:0] node7346;
	wire [4-1:0] node7350;
	wire [4-1:0] node7351;
	wire [4-1:0] node7355;
	wire [4-1:0] node7356;
	wire [4-1:0] node7357;
	wire [4-1:0] node7358;
	wire [4-1:0] node7362;
	wire [4-1:0] node7363;
	wire [4-1:0] node7367;
	wire [4-1:0] node7368;
	wire [4-1:0] node7369;
	wire [4-1:0] node7372;
	wire [4-1:0] node7375;
	wire [4-1:0] node7377;
	wire [4-1:0] node7380;
	wire [4-1:0] node7381;
	wire [4-1:0] node7382;
	wire [4-1:0] node7383;
	wire [4-1:0] node7384;
	wire [4-1:0] node7385;
	wire [4-1:0] node7388;
	wire [4-1:0] node7391;
	wire [4-1:0] node7392;
	wire [4-1:0] node7395;
	wire [4-1:0] node7398;
	wire [4-1:0] node7399;
	wire [4-1:0] node7400;
	wire [4-1:0] node7403;
	wire [4-1:0] node7406;
	wire [4-1:0] node7407;
	wire [4-1:0] node7410;
	wire [4-1:0] node7413;
	wire [4-1:0] node7414;
	wire [4-1:0] node7415;
	wire [4-1:0] node7417;
	wire [4-1:0] node7420;
	wire [4-1:0] node7422;
	wire [4-1:0] node7425;
	wire [4-1:0] node7427;
	wire [4-1:0] node7429;
	wire [4-1:0] node7432;
	wire [4-1:0] node7433;
	wire [4-1:0] node7434;
	wire [4-1:0] node7435;
	wire [4-1:0] node7436;
	wire [4-1:0] node7439;
	wire [4-1:0] node7443;
	wire [4-1:0] node7445;
	wire [4-1:0] node7447;
	wire [4-1:0] node7450;
	wire [4-1:0] node7451;
	wire [4-1:0] node7452;
	wire [4-1:0] node7453;
	wire [4-1:0] node7456;
	wire [4-1:0] node7459;
	wire [4-1:0] node7460;
	wire [4-1:0] node7463;
	wire [4-1:0] node7466;
	wire [4-1:0] node7467;
	wire [4-1:0] node7469;
	wire [4-1:0] node7472;
	wire [4-1:0] node7473;
	wire [4-1:0] node7476;
	wire [4-1:0] node7479;
	wire [4-1:0] node7480;
	wire [4-1:0] node7481;
	wire [4-1:0] node7482;
	wire [4-1:0] node7483;
	wire [4-1:0] node7484;
	wire [4-1:0] node7485;
	wire [4-1:0] node7488;
	wire [4-1:0] node7489;
	wire [4-1:0] node7492;
	wire [4-1:0] node7495;
	wire [4-1:0] node7496;
	wire [4-1:0] node7499;
	wire [4-1:0] node7500;
	wire [4-1:0] node7503;
	wire [4-1:0] node7506;
	wire [4-1:0] node7507;
	wire [4-1:0] node7508;
	wire [4-1:0] node7510;
	wire [4-1:0] node7514;
	wire [4-1:0] node7515;
	wire [4-1:0] node7516;
	wire [4-1:0] node7521;
	wire [4-1:0] node7522;
	wire [4-1:0] node7523;
	wire [4-1:0] node7524;
	wire [4-1:0] node7525;
	wire [4-1:0] node7528;
	wire [4-1:0] node7531;
	wire [4-1:0] node7534;
	wire [4-1:0] node7535;
	wire [4-1:0] node7536;
	wire [4-1:0] node7539;
	wire [4-1:0] node7542;
	wire [4-1:0] node7544;
	wire [4-1:0] node7547;
	wire [4-1:0] node7548;
	wire [4-1:0] node7549;
	wire [4-1:0] node7550;
	wire [4-1:0] node7554;
	wire [4-1:0] node7557;
	wire [4-1:0] node7560;
	wire [4-1:0] node7561;
	wire [4-1:0] node7562;
	wire [4-1:0] node7563;
	wire [4-1:0] node7564;
	wire [4-1:0] node7565;
	wire [4-1:0] node7569;
	wire [4-1:0] node7570;
	wire [4-1:0] node7574;
	wire [4-1:0] node7575;
	wire [4-1:0] node7576;
	wire [4-1:0] node7580;
	wire [4-1:0] node7581;
	wire [4-1:0] node7585;
	wire [4-1:0] node7586;
	wire [4-1:0] node7587;
	wire [4-1:0] node7590;
	wire [4-1:0] node7591;
	wire [4-1:0] node7595;
	wire [4-1:0] node7596;
	wire [4-1:0] node7597;
	wire [4-1:0] node7600;
	wire [4-1:0] node7603;
	wire [4-1:0] node7606;
	wire [4-1:0] node7607;
	wire [4-1:0] node7608;
	wire [4-1:0] node7609;
	wire [4-1:0] node7610;
	wire [4-1:0] node7613;
	wire [4-1:0] node7616;
	wire [4-1:0] node7617;
	wire [4-1:0] node7621;
	wire [4-1:0] node7622;
	wire [4-1:0] node7624;
	wire [4-1:0] node7628;
	wire [4-1:0] node7629;
	wire [4-1:0] node7630;
	wire [4-1:0] node7633;
	wire [4-1:0] node7634;
	wire [4-1:0] node7638;
	wire [4-1:0] node7639;
	wire [4-1:0] node7640;
	wire [4-1:0] node7644;
	wire [4-1:0] node7646;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7651;
	wire [4-1:0] node7652;
	wire [4-1:0] node7653;
	wire [4-1:0] node7654;
	wire [4-1:0] node7657;
	wire [4-1:0] node7660;
	wire [4-1:0] node7661;
	wire [4-1:0] node7662;
	wire [4-1:0] node7665;
	wire [4-1:0] node7668;
	wire [4-1:0] node7670;
	wire [4-1:0] node7673;
	wire [4-1:0] node7674;
	wire [4-1:0] node7675;
	wire [4-1:0] node7676;
	wire [4-1:0] node7679;
	wire [4-1:0] node7682;
	wire [4-1:0] node7684;
	wire [4-1:0] node7687;
	wire [4-1:0] node7689;
	wire [4-1:0] node7690;
	wire [4-1:0] node7693;
	wire [4-1:0] node7696;
	wire [4-1:0] node7697;
	wire [4-1:0] node7698;
	wire [4-1:0] node7699;
	wire [4-1:0] node7700;
	wire [4-1:0] node7704;
	wire [4-1:0] node7705;
	wire [4-1:0] node7709;
	wire [4-1:0] node7710;
	wire [4-1:0] node7713;
	wire [4-1:0] node7715;
	wire [4-1:0] node7718;
	wire [4-1:0] node7719;
	wire [4-1:0] node7720;
	wire [4-1:0] node7721;
	wire [4-1:0] node7724;
	wire [4-1:0] node7727;
	wire [4-1:0] node7729;
	wire [4-1:0] node7732;
	wire [4-1:0] node7733;
	wire [4-1:0] node7736;
	wire [4-1:0] node7739;
	wire [4-1:0] node7740;
	wire [4-1:0] node7741;
	wire [4-1:0] node7742;
	wire [4-1:0] node7743;
	wire [4-1:0] node7746;
	wire [4-1:0] node7749;
	wire [4-1:0] node7750;
	wire [4-1:0] node7752;
	wire [4-1:0] node7756;
	wire [4-1:0] node7757;
	wire [4-1:0] node7758;
	wire [4-1:0] node7759;
	wire [4-1:0] node7763;
	wire [4-1:0] node7766;
	wire [4-1:0] node7767;
	wire [4-1:0] node7768;
	wire [4-1:0] node7773;
	wire [4-1:0] node7774;
	wire [4-1:0] node7775;
	wire [4-1:0] node7776;
	wire [4-1:0] node7779;
	wire [4-1:0] node7780;
	wire [4-1:0] node7783;
	wire [4-1:0] node7786;
	wire [4-1:0] node7787;
	wire [4-1:0] node7790;
	wire [4-1:0] node7793;
	wire [4-1:0] node7794;
	wire [4-1:0] node7797;
	wire [4-1:0] node7800;
	wire [4-1:0] node7801;
	wire [4-1:0] node7802;
	wire [4-1:0] node7803;
	wire [4-1:0] node7804;
	wire [4-1:0] node7805;
	wire [4-1:0] node7806;
	wire [4-1:0] node7809;
	wire [4-1:0] node7811;
	wire [4-1:0] node7813;
	wire [4-1:0] node7816;
	wire [4-1:0] node7817;
	wire [4-1:0] node7819;
	wire [4-1:0] node7822;
	wire [4-1:0] node7823;
	wire [4-1:0] node7826;
	wire [4-1:0] node7828;
	wire [4-1:0] node7831;
	wire [4-1:0] node7832;
	wire [4-1:0] node7833;
	wire [4-1:0] node7834;
	wire [4-1:0] node7835;
	wire [4-1:0] node7839;
	wire [4-1:0] node7840;
	wire [4-1:0] node7843;
	wire [4-1:0] node7846;
	wire [4-1:0] node7847;
	wire [4-1:0] node7850;
	wire [4-1:0] node7851;
	wire [4-1:0] node7854;
	wire [4-1:0] node7857;
	wire [4-1:0] node7858;
	wire [4-1:0] node7859;
	wire [4-1:0] node7861;
	wire [4-1:0] node7864;
	wire [4-1:0] node7866;
	wire [4-1:0] node7869;
	wire [4-1:0] node7870;
	wire [4-1:0] node7871;
	wire [4-1:0] node7874;
	wire [4-1:0] node7878;
	wire [4-1:0] node7879;
	wire [4-1:0] node7880;
	wire [4-1:0] node7881;
	wire [4-1:0] node7883;
	wire [4-1:0] node7884;
	wire [4-1:0] node7888;
	wire [4-1:0] node7889;
	wire [4-1:0] node7892;
	wire [4-1:0] node7894;
	wire [4-1:0] node7897;
	wire [4-1:0] node7898;
	wire [4-1:0] node7900;
	wire [4-1:0] node7901;
	wire [4-1:0] node7905;
	wire [4-1:0] node7906;
	wire [4-1:0] node7907;
	wire [4-1:0] node7910;
	wire [4-1:0] node7913;
	wire [4-1:0] node7914;
	wire [4-1:0] node7918;
	wire [4-1:0] node7919;
	wire [4-1:0] node7921;
	wire [4-1:0] node7924;
	wire [4-1:0] node7925;
	wire [4-1:0] node7926;
	wire [4-1:0] node7929;
	wire [4-1:0] node7932;
	wire [4-1:0] node7933;
	wire [4-1:0] node7935;
	wire [4-1:0] node7939;
	wire [4-1:0] node7940;
	wire [4-1:0] node7941;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7945;
	wire [4-1:0] node7948;
	wire [4-1:0] node7949;
	wire [4-1:0] node7950;
	wire [4-1:0] node7953;
	wire [4-1:0] node7956;
	wire [4-1:0] node7958;
	wire [4-1:0] node7961;
	wire [4-1:0] node7962;
	wire [4-1:0] node7963;
	wire [4-1:0] node7966;
	wire [4-1:0] node7969;
	wire [4-1:0] node7972;
	wire [4-1:0] node7973;
	wire [4-1:0] node7974;
	wire [4-1:0] node7975;
	wire [4-1:0] node7978;
	wire [4-1:0] node7979;
	wire [4-1:0] node7983;
	wire [4-1:0] node7984;
	wire [4-1:0] node7987;
	wire [4-1:0] node7990;
	wire [4-1:0] node7991;
	wire [4-1:0] node7992;
	wire [4-1:0] node7994;
	wire [4-1:0] node7997;
	wire [4-1:0] node7998;
	wire [4-1:0] node8002;
	wire [4-1:0] node8003;
	wire [4-1:0] node8006;
	wire [4-1:0] node8009;
	wire [4-1:0] node8010;
	wire [4-1:0] node8011;
	wire [4-1:0] node8012;
	wire [4-1:0] node8013;
	wire [4-1:0] node8014;
	wire [4-1:0] node8019;
	wire [4-1:0] node8020;
	wire [4-1:0] node8021;
	wire [4-1:0] node8024;
	wire [4-1:0] node8027;
	wire [4-1:0] node8030;
	wire [4-1:0] node8031;
	wire [4-1:0] node8033;
	wire [4-1:0] node8034;
	wire [4-1:0] node8037;
	wire [4-1:0] node8040;
	wire [4-1:0] node8041;
	wire [4-1:0] node8044;
	wire [4-1:0] node8045;
	wire [4-1:0] node8048;
	wire [4-1:0] node8051;
	wire [4-1:0] node8052;
	wire [4-1:0] node8053;
	wire [4-1:0] node8054;
	wire [4-1:0] node8055;
	wire [4-1:0] node8058;
	wire [4-1:0] node8062;
	wire [4-1:0] node8063;
	wire [4-1:0] node8064;
	wire [4-1:0] node8068;
	wire [4-1:0] node8071;
	wire [4-1:0] node8072;
	wire [4-1:0] node8073;
	wire [4-1:0] node8074;
	wire [4-1:0] node8077;
	wire [4-1:0] node8080;
	wire [4-1:0] node8082;
	wire [4-1:0] node8085;
	wire [4-1:0] node8088;
	wire [4-1:0] node8089;
	wire [4-1:0] node8090;
	wire [4-1:0] node8091;
	wire [4-1:0] node8092;
	wire [4-1:0] node8093;
	wire [4-1:0] node8094;
	wire [4-1:0] node8097;
	wire [4-1:0] node8098;
	wire [4-1:0] node8101;
	wire [4-1:0] node8104;
	wire [4-1:0] node8106;
	wire [4-1:0] node8108;
	wire [4-1:0] node8111;
	wire [4-1:0] node8112;
	wire [4-1:0] node8113;
	wire [4-1:0] node8115;
	wire [4-1:0] node8119;
	wire [4-1:0] node8120;
	wire [4-1:0] node8122;
	wire [4-1:0] node8125;
	wire [4-1:0] node8128;
	wire [4-1:0] node8129;
	wire [4-1:0] node8130;
	wire [4-1:0] node8131;
	wire [4-1:0] node8133;
	wire [4-1:0] node8136;
	wire [4-1:0] node8139;
	wire [4-1:0] node8140;
	wire [4-1:0] node8143;
	wire [4-1:0] node8144;
	wire [4-1:0] node8148;
	wire [4-1:0] node8149;
	wire [4-1:0] node8150;
	wire [4-1:0] node8152;
	wire [4-1:0] node8155;
	wire [4-1:0] node8158;
	wire [4-1:0] node8160;
	wire [4-1:0] node8163;
	wire [4-1:0] node8164;
	wire [4-1:0] node8165;
	wire [4-1:0] node8166;
	wire [4-1:0] node8167;
	wire [4-1:0] node8170;
	wire [4-1:0] node8173;
	wire [4-1:0] node8175;
	wire [4-1:0] node8176;
	wire [4-1:0] node8179;
	wire [4-1:0] node8182;
	wire [4-1:0] node8183;
	wire [4-1:0] node8186;
	wire [4-1:0] node8187;
	wire [4-1:0] node8190;
	wire [4-1:0] node8191;
	wire [4-1:0] node8195;
	wire [4-1:0] node8196;
	wire [4-1:0] node8197;
	wire [4-1:0] node8198;
	wire [4-1:0] node8199;
	wire [4-1:0] node8203;
	wire [4-1:0] node8205;
	wire [4-1:0] node8208;
	wire [4-1:0] node8209;
	wire [4-1:0] node8210;
	wire [4-1:0] node8214;
	wire [4-1:0] node8216;
	wire [4-1:0] node8219;
	wire [4-1:0] node8220;
	wire [4-1:0] node8221;
	wire [4-1:0] node8223;
	wire [4-1:0] node8227;
	wire [4-1:0] node8228;
	wire [4-1:0] node8230;
	wire [4-1:0] node8233;
	wire [4-1:0] node8234;
	wire [4-1:0] node8237;
	wire [4-1:0] node8240;
	wire [4-1:0] node8241;
	wire [4-1:0] node8242;
	wire [4-1:0] node8243;
	wire [4-1:0] node8244;
	wire [4-1:0] node8247;
	wire [4-1:0] node8248;
	wire [4-1:0] node8249;
	wire [4-1:0] node8252;
	wire [4-1:0] node8255;
	wire [4-1:0] node8256;
	wire [4-1:0] node8259;
	wire [4-1:0] node8262;
	wire [4-1:0] node8263;
	wire [4-1:0] node8264;
	wire [4-1:0] node8266;
	wire [4-1:0] node8269;
	wire [4-1:0] node8270;
	wire [4-1:0] node8273;
	wire [4-1:0] node8276;
	wire [4-1:0] node8278;
	wire [4-1:0] node8279;
	wire [4-1:0] node8282;
	wire [4-1:0] node8285;
	wire [4-1:0] node8286;
	wire [4-1:0] node8287;
	wire [4-1:0] node8288;
	wire [4-1:0] node8291;
	wire [4-1:0] node8292;
	wire [4-1:0] node8295;
	wire [4-1:0] node8298;
	wire [4-1:0] node8299;
	wire [4-1:0] node8302;
	wire [4-1:0] node8303;
	wire [4-1:0] node8306;
	wire [4-1:0] node8309;
	wire [4-1:0] node8310;
	wire [4-1:0] node8311;
	wire [4-1:0] node8312;
	wire [4-1:0] node8315;
	wire [4-1:0] node8318;
	wire [4-1:0] node8319;
	wire [4-1:0] node8323;
	wire [4-1:0] node8324;
	wire [4-1:0] node8327;
	wire [4-1:0] node8330;
	wire [4-1:0] node8331;
	wire [4-1:0] node8332;
	wire [4-1:0] node8333;
	wire [4-1:0] node8334;
	wire [4-1:0] node8336;
	wire [4-1:0] node8339;
	wire [4-1:0] node8340;
	wire [4-1:0] node8343;
	wire [4-1:0] node8346;
	wire [4-1:0] node8347;
	wire [4-1:0] node8348;
	wire [4-1:0] node8351;
	wire [4-1:0] node8354;
	wire [4-1:0] node8355;
	wire [4-1:0] node8359;
	wire [4-1:0] node8360;
	wire [4-1:0] node8361;
	wire [4-1:0] node8363;
	wire [4-1:0] node8366;
	wire [4-1:0] node8369;
	wire [4-1:0] node8371;
	wire [4-1:0] node8374;
	wire [4-1:0] node8375;
	wire [4-1:0] node8376;
	wire [4-1:0] node8377;
	wire [4-1:0] node8378;
	wire [4-1:0] node8382;
	wire [4-1:0] node8383;
	wire [4-1:0] node8387;
	wire [4-1:0] node8388;
	wire [4-1:0] node8389;
	wire [4-1:0] node8393;
	wire [4-1:0] node8395;
	wire [4-1:0] node8398;
	wire [4-1:0] node8399;
	wire [4-1:0] node8400;
	wire [4-1:0] node8401;
	wire [4-1:0] node8406;
	wire [4-1:0] node8407;
	wire [4-1:0] node8411;
	wire [4-1:0] node8412;
	wire [4-1:0] node8413;
	wire [4-1:0] node8414;
	wire [4-1:0] node8415;
	wire [4-1:0] node8416;
	wire [4-1:0] node8417;
	wire [4-1:0] node8418;
	wire [4-1:0] node8420;
	wire [4-1:0] node8423;
	wire [4-1:0] node8425;
	wire [4-1:0] node8426;
	wire [4-1:0] node8429;
	wire [4-1:0] node8432;
	wire [4-1:0] node8434;
	wire [4-1:0] node8436;
	wire [4-1:0] node8439;
	wire [4-1:0] node8440;
	wire [4-1:0] node8441;
	wire [4-1:0] node8442;
	wire [4-1:0] node8445;
	wire [4-1:0] node8447;
	wire [4-1:0] node8450;
	wire [4-1:0] node8451;
	wire [4-1:0] node8453;
	wire [4-1:0] node8456;
	wire [4-1:0] node8458;
	wire [4-1:0] node8461;
	wire [4-1:0] node8462;
	wire [4-1:0] node8463;
	wire [4-1:0] node8464;
	wire [4-1:0] node8467;
	wire [4-1:0] node8471;
	wire [4-1:0] node8472;
	wire [4-1:0] node8475;
	wire [4-1:0] node8477;
	wire [4-1:0] node8480;
	wire [4-1:0] node8481;
	wire [4-1:0] node8482;
	wire [4-1:0] node8483;
	wire [4-1:0] node8484;
	wire [4-1:0] node8488;
	wire [4-1:0] node8489;
	wire [4-1:0] node8490;
	wire [4-1:0] node8494;
	wire [4-1:0] node8497;
	wire [4-1:0] node8498;
	wire [4-1:0] node8499;
	wire [4-1:0] node8502;
	wire [4-1:0] node8505;
	wire [4-1:0] node8506;
	wire [4-1:0] node8507;
	wire [4-1:0] node8510;
	wire [4-1:0] node8513;
	wire [4-1:0] node8514;
	wire [4-1:0] node8518;
	wire [4-1:0] node8519;
	wire [4-1:0] node8520;
	wire [4-1:0] node8522;
	wire [4-1:0] node8525;
	wire [4-1:0] node8526;
	wire [4-1:0] node8528;
	wire [4-1:0] node8531;
	wire [4-1:0] node8533;
	wire [4-1:0] node8536;
	wire [4-1:0] node8537;
	wire [4-1:0] node8539;
	wire [4-1:0] node8541;
	wire [4-1:0] node8544;
	wire [4-1:0] node8545;
	wire [4-1:0] node8548;
	wire [4-1:0] node8549;
	wire [4-1:0] node8553;
	wire [4-1:0] node8554;
	wire [4-1:0] node8555;
	wire [4-1:0] node8556;
	wire [4-1:0] node8557;
	wire [4-1:0] node8558;
	wire [4-1:0] node8560;
	wire [4-1:0] node8563;
	wire [4-1:0] node8566;
	wire [4-1:0] node8567;
	wire [4-1:0] node8568;
	wire [4-1:0] node8572;
	wire [4-1:0] node8573;
	wire [4-1:0] node8576;
	wire [4-1:0] node8579;
	wire [4-1:0] node8580;
	wire [4-1:0] node8581;
	wire [4-1:0] node8582;
	wire [4-1:0] node8585;
	wire [4-1:0] node8588;
	wire [4-1:0] node8589;
	wire [4-1:0] node8592;
	wire [4-1:0] node8595;
	wire [4-1:0] node8596;
	wire [4-1:0] node8597;
	wire [4-1:0] node8601;
	wire [4-1:0] node8603;
	wire [4-1:0] node8606;
	wire [4-1:0] node8607;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8610;
	wire [4-1:0] node8613;
	wire [4-1:0] node8616;
	wire [4-1:0] node8618;
	wire [4-1:0] node8621;
	wire [4-1:0] node8622;
	wire [4-1:0] node8625;
	wire [4-1:0] node8628;
	wire [4-1:0] node8629;
	wire [4-1:0] node8630;
	wire [4-1:0] node8631;
	wire [4-1:0] node8635;
	wire [4-1:0] node8636;
	wire [4-1:0] node8639;
	wire [4-1:0] node8642;
	wire [4-1:0] node8643;
	wire [4-1:0] node8644;
	wire [4-1:0] node8647;
	wire [4-1:0] node8650;
	wire [4-1:0] node8653;
	wire [4-1:0] node8654;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8657;
	wire [4-1:0] node8658;
	wire [4-1:0] node8663;
	wire [4-1:0] node8665;
	wire [4-1:0] node8668;
	wire [4-1:0] node8669;
	wire [4-1:0] node8670;
	wire [4-1:0] node8671;
	wire [4-1:0] node8675;
	wire [4-1:0] node8678;
	wire [4-1:0] node8679;
	wire [4-1:0] node8682;
	wire [4-1:0] node8685;
	wire [4-1:0] node8686;
	wire [4-1:0] node8687;
	wire [4-1:0] node8688;
	wire [4-1:0] node8690;
	wire [4-1:0] node8694;
	wire [4-1:0] node8695;
	wire [4-1:0] node8699;
	wire [4-1:0] node8700;
	wire [4-1:0] node8701;
	wire [4-1:0] node8703;
	wire [4-1:0] node8707;
	wire [4-1:0] node8708;
	wire [4-1:0] node8709;
	wire [4-1:0] node8713;
	wire [4-1:0] node8715;
	wire [4-1:0] node8718;
	wire [4-1:0] node8719;
	wire [4-1:0] node8720;
	wire [4-1:0] node8721;
	wire [4-1:0] node8722;
	wire [4-1:0] node8723;
	wire [4-1:0] node8725;
	wire [4-1:0] node8728;
	wire [4-1:0] node8729;
	wire [4-1:0] node8731;
	wire [4-1:0] node8734;
	wire [4-1:0] node8735;
	wire [4-1:0] node8739;
	wire [4-1:0] node8740;
	wire [4-1:0] node8742;
	wire [4-1:0] node8743;
	wire [4-1:0] node8747;
	wire [4-1:0] node8748;
	wire [4-1:0] node8751;
	wire [4-1:0] node8754;
	wire [4-1:0] node8755;
	wire [4-1:0] node8756;
	wire [4-1:0] node8757;
	wire [4-1:0] node8760;
	wire [4-1:0] node8762;
	wire [4-1:0] node8765;
	wire [4-1:0] node8767;
	wire [4-1:0] node8770;
	wire [4-1:0] node8771;
	wire [4-1:0] node8772;
	wire [4-1:0] node8774;
	wire [4-1:0] node8777;
	wire [4-1:0] node8780;
	wire [4-1:0] node8781;
	wire [4-1:0] node8784;
	wire [4-1:0] node8787;
	wire [4-1:0] node8788;
	wire [4-1:0] node8789;
	wire [4-1:0] node8790;
	wire [4-1:0] node8791;
	wire [4-1:0] node8792;
	wire [4-1:0] node8796;
	wire [4-1:0] node8797;
	wire [4-1:0] node8800;
	wire [4-1:0] node8803;
	wire [4-1:0] node8804;
	wire [4-1:0] node8806;
	wire [4-1:0] node8809;
	wire [4-1:0] node8810;
	wire [4-1:0] node8813;
	wire [4-1:0] node8816;
	wire [4-1:0] node8817;
	wire [4-1:0] node8818;
	wire [4-1:0] node8821;
	wire [4-1:0] node8824;
	wire [4-1:0] node8825;
	wire [4-1:0] node8829;
	wire [4-1:0] node8830;
	wire [4-1:0] node8831;
	wire [4-1:0] node8832;
	wire [4-1:0] node8833;
	wire [4-1:0] node8837;
	wire [4-1:0] node8838;
	wire [4-1:0] node8842;
	wire [4-1:0] node8843;
	wire [4-1:0] node8846;
	wire [4-1:0] node8849;
	wire [4-1:0] node8851;
	wire [4-1:0] node8852;
	wire [4-1:0] node8855;
	wire [4-1:0] node8856;
	wire [4-1:0] node8860;
	wire [4-1:0] node8861;
	wire [4-1:0] node8862;
	wire [4-1:0] node8863;
	wire [4-1:0] node8864;
	wire [4-1:0] node8865;
	wire [4-1:0] node8866;
	wire [4-1:0] node8869;
	wire [4-1:0] node8872;
	wire [4-1:0] node8875;
	wire [4-1:0] node8876;
	wire [4-1:0] node8878;
	wire [4-1:0] node8881;
	wire [4-1:0] node8884;
	wire [4-1:0] node8885;
	wire [4-1:0] node8886;
	wire [4-1:0] node8888;
	wire [4-1:0] node8891;
	wire [4-1:0] node8892;
	wire [4-1:0] node8895;
	wire [4-1:0] node8898;
	wire [4-1:0] node8901;
	wire [4-1:0] node8902;
	wire [4-1:0] node8903;
	wire [4-1:0] node8904;
	wire [4-1:0] node8907;
	wire [4-1:0] node8910;
	wire [4-1:0] node8911;
	wire [4-1:0] node8912;
	wire [4-1:0] node8915;
	wire [4-1:0] node8918;
	wire [4-1:0] node8921;
	wire [4-1:0] node8924;
	wire [4-1:0] node8925;
	wire [4-1:0] node8926;
	wire [4-1:0] node8927;
	wire [4-1:0] node8929;
	wire [4-1:0] node8930;
	wire [4-1:0] node8933;
	wire [4-1:0] node8936;
	wire [4-1:0] node8937;
	wire [4-1:0] node8938;
	wire [4-1:0] node8941;
	wire [4-1:0] node8945;
	wire [4-1:0] node8946;
	wire [4-1:0] node8947;
	wire [4-1:0] node8950;
	wire [4-1:0] node8952;
	wire [4-1:0] node8955;
	wire [4-1:0] node8956;
	wire [4-1:0] node8958;
	wire [4-1:0] node8961;
	wire [4-1:0] node8964;
	wire [4-1:0] node8965;
	wire [4-1:0] node8966;
	wire [4-1:0] node8967;
	wire [4-1:0] node8971;
	wire [4-1:0] node8973;
	wire [4-1:0] node8976;
	wire [4-1:0] node8979;
	wire [4-1:0] node8980;
	wire [4-1:0] node8981;
	wire [4-1:0] node8982;
	wire [4-1:0] node8983;
	wire [4-1:0] node8984;
	wire [4-1:0] node8985;
	wire [4-1:0] node8986;
	wire [4-1:0] node8989;
	wire [4-1:0] node8990;
	wire [4-1:0] node8994;
	wire [4-1:0] node8995;
	wire [4-1:0] node8997;
	wire [4-1:0] node9000;
	wire [4-1:0] node9003;
	wire [4-1:0] node9004;
	wire [4-1:0] node9005;
	wire [4-1:0] node9009;
	wire [4-1:0] node9010;
	wire [4-1:0] node9012;
	wire [4-1:0] node9015;
	wire [4-1:0] node9016;
	wire [4-1:0] node9020;
	wire [4-1:0] node9021;
	wire [4-1:0] node9022;
	wire [4-1:0] node9023;
	wire [4-1:0] node9025;
	wire [4-1:0] node9028;
	wire [4-1:0] node9030;
	wire [4-1:0] node9033;
	wire [4-1:0] node9034;
	wire [4-1:0] node9035;
	wire [4-1:0] node9039;
	wire [4-1:0] node9040;
	wire [4-1:0] node9043;
	wire [4-1:0] node9046;
	wire [4-1:0] node9047;
	wire [4-1:0] node9048;
	wire [4-1:0] node9049;
	wire [4-1:0] node9052;
	wire [4-1:0] node9055;
	wire [4-1:0] node9057;
	wire [4-1:0] node9060;
	wire [4-1:0] node9061;
	wire [4-1:0] node9063;
	wire [4-1:0] node9066;
	wire [4-1:0] node9068;
	wire [4-1:0] node9071;
	wire [4-1:0] node9072;
	wire [4-1:0] node9073;
	wire [4-1:0] node9074;
	wire [4-1:0] node9075;
	wire [4-1:0] node9077;
	wire [4-1:0] node9080;
	wire [4-1:0] node9081;
	wire [4-1:0] node9084;
	wire [4-1:0] node9087;
	wire [4-1:0] node9088;
	wire [4-1:0] node9089;
	wire [4-1:0] node9094;
	wire [4-1:0] node9095;
	wire [4-1:0] node9096;
	wire [4-1:0] node9097;
	wire [4-1:0] node9101;
	wire [4-1:0] node9103;
	wire [4-1:0] node9106;
	wire [4-1:0] node9107;
	wire [4-1:0] node9110;
	wire [4-1:0] node9111;
	wire [4-1:0] node9115;
	wire [4-1:0] node9116;
	wire [4-1:0] node9117;
	wire [4-1:0] node9118;
	wire [4-1:0] node9122;
	wire [4-1:0] node9123;
	wire [4-1:0] node9124;
	wire [4-1:0] node9128;
	wire [4-1:0] node9131;
	wire [4-1:0] node9132;
	wire [4-1:0] node9133;
	wire [4-1:0] node9135;
	wire [4-1:0] node9140;
	wire [4-1:0] node9141;
	wire [4-1:0] node9142;
	wire [4-1:0] node9143;
	wire [4-1:0] node9144;
	wire [4-1:0] node9145;
	wire [4-1:0] node9148;
	wire [4-1:0] node9151;
	wire [4-1:0] node9152;
	wire [4-1:0] node9155;
	wire [4-1:0] node9157;
	wire [4-1:0] node9160;
	wire [4-1:0] node9161;
	wire [4-1:0] node9162;
	wire [4-1:0] node9166;
	wire [4-1:0] node9167;
	wire [4-1:0] node9168;
	wire [4-1:0] node9171;
	wire [4-1:0] node9174;
	wire [4-1:0] node9177;
	wire [4-1:0] node9178;
	wire [4-1:0] node9179;
	wire [4-1:0] node9180;
	wire [4-1:0] node9181;
	wire [4-1:0] node9184;
	wire [4-1:0] node9187;
	wire [4-1:0] node9188;
	wire [4-1:0] node9191;
	wire [4-1:0] node9194;
	wire [4-1:0] node9195;
	wire [4-1:0] node9198;
	wire [4-1:0] node9201;
	wire [4-1:0] node9203;
	wire [4-1:0] node9204;
	wire [4-1:0] node9205;
	wire [4-1:0] node9208;
	wire [4-1:0] node9211;
	wire [4-1:0] node9213;
	wire [4-1:0] node9216;
	wire [4-1:0] node9217;
	wire [4-1:0] node9218;
	wire [4-1:0] node9219;
	wire [4-1:0] node9220;
	wire [4-1:0] node9222;
	wire [4-1:0] node9225;
	wire [4-1:0] node9226;
	wire [4-1:0] node9229;
	wire [4-1:0] node9232;
	wire [4-1:0] node9233;
	wire [4-1:0] node9236;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9243;
	wire [4-1:0] node9246;
	wire [4-1:0] node9249;
	wire [4-1:0] node9250;
	wire [4-1:0] node9251;
	wire [4-1:0] node9255;
	wire [4-1:0] node9257;
	wire [4-1:0] node9260;
	wire [4-1:0] node9261;
	wire [4-1:0] node9262;
	wire [4-1:0] node9264;
	wire [4-1:0] node9267;
	wire [4-1:0] node9268;
	wire [4-1:0] node9269;
	wire [4-1:0] node9272;
	wire [4-1:0] node9275;
	wire [4-1:0] node9276;
	wire [4-1:0] node9280;
	wire [4-1:0] node9281;
	wire [4-1:0] node9282;
	wire [4-1:0] node9286;
	wire [4-1:0] node9289;
	wire [4-1:0] node9290;
	wire [4-1:0] node9291;
	wire [4-1:0] node9292;
	wire [4-1:0] node9293;
	wire [4-1:0] node9294;
	wire [4-1:0] node9295;
	wire [4-1:0] node9297;
	wire [4-1:0] node9301;
	wire [4-1:0] node9302;
	wire [4-1:0] node9304;
	wire [4-1:0] node9307;
	wire [4-1:0] node9308;
	wire [4-1:0] node9312;
	wire [4-1:0] node9313;
	wire [4-1:0] node9314;
	wire [4-1:0] node9317;
	wire [4-1:0] node9318;
	wire [4-1:0] node9321;
	wire [4-1:0] node9324;
	wire [4-1:0] node9325;
	wire [4-1:0] node9326;
	wire [4-1:0] node9330;
	wire [4-1:0] node9331;
	wire [4-1:0] node9334;
	wire [4-1:0] node9337;
	wire [4-1:0] node9338;
	wire [4-1:0] node9339;
	wire [4-1:0] node9340;
	wire [4-1:0] node9343;
	wire [4-1:0] node9346;
	wire [4-1:0] node9347;
	wire [4-1:0] node9350;
	wire [4-1:0] node9352;
	wire [4-1:0] node9355;
	wire [4-1:0] node9356;
	wire [4-1:0] node9357;
	wire [4-1:0] node9358;
	wire [4-1:0] node9361;
	wire [4-1:0] node9364;
	wire [4-1:0] node9366;
	wire [4-1:0] node9369;
	wire [4-1:0] node9370;
	wire [4-1:0] node9371;
	wire [4-1:0] node9374;
	wire [4-1:0] node9378;
	wire [4-1:0] node9379;
	wire [4-1:0] node9380;
	wire [4-1:0] node9381;
	wire [4-1:0] node9382;
	wire [4-1:0] node9384;
	wire [4-1:0] node9387;
	wire [4-1:0] node9389;
	wire [4-1:0] node9392;
	wire [4-1:0] node9393;
	wire [4-1:0] node9395;
	wire [4-1:0] node9398;
	wire [4-1:0] node9400;
	wire [4-1:0] node9403;
	wire [4-1:0] node9404;
	wire [4-1:0] node9405;
	wire [4-1:0] node9406;
	wire [4-1:0] node9409;
	wire [4-1:0] node9412;
	wire [4-1:0] node9413;
	wire [4-1:0] node9416;
	wire [4-1:0] node9419;
	wire [4-1:0] node9420;
	wire [4-1:0] node9421;
	wire [4-1:0] node9425;
	wire [4-1:0] node9427;
	wire [4-1:0] node9430;
	wire [4-1:0] node9431;
	wire [4-1:0] node9432;
	wire [4-1:0] node9434;
	wire [4-1:0] node9435;
	wire [4-1:0] node9438;
	wire [4-1:0] node9441;
	wire [4-1:0] node9442;
	wire [4-1:0] node9444;
	wire [4-1:0] node9447;
	wire [4-1:0] node9448;
	wire [4-1:0] node9452;
	wire [4-1:0] node9453;
	wire [4-1:0] node9454;
	wire [4-1:0] node9455;
	wire [4-1:0] node9460;
	wire [4-1:0] node9462;
	wire [4-1:0] node9463;
	wire [4-1:0] node9467;
	wire [4-1:0] node9468;
	wire [4-1:0] node9469;
	wire [4-1:0] node9470;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9475;
	wire [4-1:0] node9478;
	wire [4-1:0] node9479;
	wire [4-1:0] node9481;
	wire [4-1:0] node9484;
	wire [4-1:0] node9487;
	wire [4-1:0] node9488;
	wire [4-1:0] node9490;
	wire [4-1:0] node9493;
	wire [4-1:0] node9495;
	wire [4-1:0] node9498;
	wire [4-1:0] node9499;
	wire [4-1:0] node9500;
	wire [4-1:0] node9501;
	wire [4-1:0] node9503;
	wire [4-1:0] node9506;
	wire [4-1:0] node9507;
	wire [4-1:0] node9510;
	wire [4-1:0] node9513;
	wire [4-1:0] node9514;
	wire [4-1:0] node9515;
	wire [4-1:0] node9518;
	wire [4-1:0] node9521;
	wire [4-1:0] node9524;
	wire [4-1:0] node9525;
	wire [4-1:0] node9526;
	wire [4-1:0] node9528;
	wire [4-1:0] node9531;
	wire [4-1:0] node9534;
	wire [4-1:0] node9535;
	wire [4-1:0] node9536;
	wire [4-1:0] node9540;
	wire [4-1:0] node9541;
	wire [4-1:0] node9544;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9549;
	wire [4-1:0] node9550;
	wire [4-1:0] node9551;
	wire [4-1:0] node9554;
	wire [4-1:0] node9555;
	wire [4-1:0] node9558;
	wire [4-1:0] node9561;
	wire [4-1:0] node9562;
	wire [4-1:0] node9564;
	wire [4-1:0] node9567;
	wire [4-1:0] node9570;
	wire [4-1:0] node9571;
	wire [4-1:0] node9572;
	wire [4-1:0] node9573;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9583;
	wire [4-1:0] node9584;
	wire [4-1:0] node9585;
	wire [4-1:0] node9586;
	wire [4-1:0] node9589;
	wire [4-1:0] node9590;
	wire [4-1:0] node9593;
	wire [4-1:0] node9596;
	wire [4-1:0] node9597;
	wire [4-1:0] node9598;
	wire [4-1:0] node9601;
	wire [4-1:0] node9604;
	wire [4-1:0] node9607;
	wire [4-1:0] node9608;
	wire [4-1:0] node9609;
	wire [4-1:0] node9610;
	wire [4-1:0] node9613;
	wire [4-1:0] node9616;
	wire [4-1:0] node9617;
	wire [4-1:0] node9621;
	wire [4-1:0] node9624;
	wire [4-1:0] node9625;
	wire [4-1:0] node9626;
	wire [4-1:0] node9627;
	wire [4-1:0] node9628;
	wire [4-1:0] node9629;
	wire [4-1:0] node9630;
	wire [4-1:0] node9631;
	wire [4-1:0] node9632;
	wire [4-1:0] node9634;
	wire [4-1:0] node9636;
	wire [4-1:0] node9638;
	wire [4-1:0] node9641;
	wire [4-1:0] node9643;
	wire [4-1:0] node9644;
	wire [4-1:0] node9645;
	wire [4-1:0] node9648;
	wire [4-1:0] node9652;
	wire [4-1:0] node9653;
	wire [4-1:0] node9654;
	wire [4-1:0] node9656;
	wire [4-1:0] node9657;
	wire [4-1:0] node9660;
	wire [4-1:0] node9663;
	wire [4-1:0] node9664;
	wire [4-1:0] node9666;
	wire [4-1:0] node9669;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9674;
	wire [4-1:0] node9677;
	wire [4-1:0] node9680;
	wire [4-1:0] node9682;
	wire [4-1:0] node9683;
	wire [4-1:0] node9687;
	wire [4-1:0] node9688;
	wire [4-1:0] node9689;
	wire [4-1:0] node9691;
	wire [4-1:0] node9692;
	wire [4-1:0] node9694;
	wire [4-1:0] node9697;
	wire [4-1:0] node9698;
	wire [4-1:0] node9702;
	wire [4-1:0] node9704;
	wire [4-1:0] node9705;
	wire [4-1:0] node9706;
	wire [4-1:0] node9710;
	wire [4-1:0] node9711;
	wire [4-1:0] node9715;
	wire [4-1:0] node9716;
	wire [4-1:0] node9717;
	wire [4-1:0] node9719;
	wire [4-1:0] node9721;
	wire [4-1:0] node9724;
	wire [4-1:0] node9725;
	wire [4-1:0] node9726;
	wire [4-1:0] node9730;
	wire [4-1:0] node9733;
	wire [4-1:0] node9734;
	wire [4-1:0] node9735;
	wire [4-1:0] node9737;
	wire [4-1:0] node9740;
	wire [4-1:0] node9742;
	wire [4-1:0] node9743;
	wire [4-1:0] node9746;
	wire [4-1:0] node9749;
	wire [4-1:0] node9750;
	wire [4-1:0] node9752;
	wire [4-1:0] node9755;
	wire [4-1:0] node9756;
	wire [4-1:0] node9760;
	wire [4-1:0] node9761;
	wire [4-1:0] node9762;
	wire [4-1:0] node9763;
	wire [4-1:0] node9764;
	wire [4-1:0] node9766;
	wire [4-1:0] node9767;
	wire [4-1:0] node9771;
	wire [4-1:0] node9773;
	wire [4-1:0] node9774;
	wire [4-1:0] node9778;
	wire [4-1:0] node9779;
	wire [4-1:0] node9780;
	wire [4-1:0] node9782;
	wire [4-1:0] node9785;
	wire [4-1:0] node9787;
	wire [4-1:0] node9790;
	wire [4-1:0] node9792;
	wire [4-1:0] node9794;
	wire [4-1:0] node9797;
	wire [4-1:0] node9798;
	wire [4-1:0] node9799;
	wire [4-1:0] node9800;
	wire [4-1:0] node9802;
	wire [4-1:0] node9805;
	wire [4-1:0] node9807;
	wire [4-1:0] node9810;
	wire [4-1:0] node9811;
	wire [4-1:0] node9814;
	wire [4-1:0] node9817;
	wire [4-1:0] node9818;
	wire [4-1:0] node9819;
	wire [4-1:0] node9820;
	wire [4-1:0] node9824;
	wire [4-1:0] node9827;
	wire [4-1:0] node9828;
	wire [4-1:0] node9831;
	wire [4-1:0] node9833;
	wire [4-1:0] node9834;
	wire [4-1:0] node9837;
	wire [4-1:0] node9840;
	wire [4-1:0] node9841;
	wire [4-1:0] node9842;
	wire [4-1:0] node9843;
	wire [4-1:0] node9844;
	wire [4-1:0] node9847;
	wire [4-1:0] node9848;
	wire [4-1:0] node9852;
	wire [4-1:0] node9853;
	wire [4-1:0] node9855;
	wire [4-1:0] node9859;
	wire [4-1:0] node9860;
	wire [4-1:0] node9861;
	wire [4-1:0] node9862;
	wire [4-1:0] node9865;
	wire [4-1:0] node9868;
	wire [4-1:0] node9870;
	wire [4-1:0] node9871;
	wire [4-1:0] node9875;
	wire [4-1:0] node9877;
	wire [4-1:0] node9879;
	wire [4-1:0] node9882;
	wire [4-1:0] node9883;
	wire [4-1:0] node9884;
	wire [4-1:0] node9885;
	wire [4-1:0] node9886;
	wire [4-1:0] node9889;
	wire [4-1:0] node9892;
	wire [4-1:0] node9895;
	wire [4-1:0] node9896;
	wire [4-1:0] node9899;
	wire [4-1:0] node9900;
	wire [4-1:0] node9904;
	wire [4-1:0] node9905;
	wire [4-1:0] node9906;
	wire [4-1:0] node9907;
	wire [4-1:0] node9908;
	wire [4-1:0] node9911;
	wire [4-1:0] node9914;
	wire [4-1:0] node9915;
	wire [4-1:0] node9919;
	wire [4-1:0] node9920;
	wire [4-1:0] node9923;
	wire [4-1:0] node9926;
	wire [4-1:0] node9927;
	wire [4-1:0] node9928;
	wire [4-1:0] node9931;
	wire [4-1:0] node9934;
	wire [4-1:0] node9936;
	wire [4-1:0] node9939;
	wire [4-1:0] node9940;
	wire [4-1:0] node9941;
	wire [4-1:0] node9942;
	wire [4-1:0] node9943;
	wire [4-1:0] node9944;
	wire [4-1:0] node9945;
	wire [4-1:0] node9948;
	wire [4-1:0] node9951;
	wire [4-1:0] node9952;
	wire [4-1:0] node9954;
	wire [4-1:0] node9957;
	wire [4-1:0] node9958;
	wire [4-1:0] node9962;
	wire [4-1:0] node9963;
	wire [4-1:0] node9964;
	wire [4-1:0] node9967;
	wire [4-1:0] node9969;
	wire [4-1:0] node9972;
	wire [4-1:0] node9973;
	wire [4-1:0] node9977;
	wire [4-1:0] node9978;
	wire [4-1:0] node9979;
	wire [4-1:0] node9980;
	wire [4-1:0] node9981;
	wire [4-1:0] node9983;
	wire [4-1:0] node9986;
	wire [4-1:0] node9987;
	wire [4-1:0] node9990;
	wire [4-1:0] node9993;
	wire [4-1:0] node9994;
	wire [4-1:0] node9998;
	wire [4-1:0] node9999;
	wire [4-1:0] node10002;
	wire [4-1:0] node10003;
	wire [4-1:0] node10007;
	wire [4-1:0] node10008;
	wire [4-1:0] node10010;
	wire [4-1:0] node10013;
	wire [4-1:0] node10014;
	wire [4-1:0] node10017;
	wire [4-1:0] node10018;
	wire [4-1:0] node10022;
	wire [4-1:0] node10023;
	wire [4-1:0] node10024;
	wire [4-1:0] node10025;
	wire [4-1:0] node10026;
	wire [4-1:0] node10027;
	wire [4-1:0] node10031;
	wire [4-1:0] node10032;
	wire [4-1:0] node10036;
	wire [4-1:0] node10037;
	wire [4-1:0] node10038;
	wire [4-1:0] node10041;
	wire [4-1:0] node10044;
	wire [4-1:0] node10045;
	wire [4-1:0] node10046;
	wire [4-1:0] node10051;
	wire [4-1:0] node10052;
	wire [4-1:0] node10053;
	wire [4-1:0] node10056;
	wire [4-1:0] node10059;
	wire [4-1:0] node10060;
	wire [4-1:0] node10064;
	wire [4-1:0] node10065;
	wire [4-1:0] node10066;
	wire [4-1:0] node10067;
	wire [4-1:0] node10068;
	wire [4-1:0] node10071;
	wire [4-1:0] node10074;
	wire [4-1:0] node10077;
	wire [4-1:0] node10078;
	wire [4-1:0] node10081;
	wire [4-1:0] node10082;
	wire [4-1:0] node10086;
	wire [4-1:0] node10087;
	wire [4-1:0] node10088;
	wire [4-1:0] node10090;
	wire [4-1:0] node10094;
	wire [4-1:0] node10095;
	wire [4-1:0] node10098;
	wire [4-1:0] node10099;
	wire [4-1:0] node10103;
	wire [4-1:0] node10104;
	wire [4-1:0] node10105;
	wire [4-1:0] node10106;
	wire [4-1:0] node10107;
	wire [4-1:0] node10108;
	wire [4-1:0] node10110;
	wire [4-1:0] node10114;
	wire [4-1:0] node10115;
	wire [4-1:0] node10117;
	wire [4-1:0] node10120;
	wire [4-1:0] node10123;
	wire [4-1:0] node10124;
	wire [4-1:0] node10125;
	wire [4-1:0] node10128;
	wire [4-1:0] node10131;
	wire [4-1:0] node10132;
	wire [4-1:0] node10133;
	wire [4-1:0] node10136;
	wire [4-1:0] node10138;
	wire [4-1:0] node10142;
	wire [4-1:0] node10143;
	wire [4-1:0] node10144;
	wire [4-1:0] node10145;
	wire [4-1:0] node10146;
	wire [4-1:0] node10147;
	wire [4-1:0] node10151;
	wire [4-1:0] node10152;
	wire [4-1:0] node10155;
	wire [4-1:0] node10158;
	wire [4-1:0] node10160;
	wire [4-1:0] node10163;
	wire [4-1:0] node10164;
	wire [4-1:0] node10165;
	wire [4-1:0] node10168;
	wire [4-1:0] node10171;
	wire [4-1:0] node10173;
	wire [4-1:0] node10176;
	wire [4-1:0] node10177;
	wire [4-1:0] node10178;
	wire [4-1:0] node10180;
	wire [4-1:0] node10183;
	wire [4-1:0] node10185;
	wire [4-1:0] node10188;
	wire [4-1:0] node10189;
	wire [4-1:0] node10191;
	wire [4-1:0] node10194;
	wire [4-1:0] node10196;
	wire [4-1:0] node10199;
	wire [4-1:0] node10200;
	wire [4-1:0] node10201;
	wire [4-1:0] node10202;
	wire [4-1:0] node10203;
	wire [4-1:0] node10204;
	wire [4-1:0] node10208;
	wire [4-1:0] node10209;
	wire [4-1:0] node10212;
	wire [4-1:0] node10215;
	wire [4-1:0] node10216;
	wire [4-1:0] node10217;
	wire [4-1:0] node10220;
	wire [4-1:0] node10223;
	wire [4-1:0] node10224;
	wire [4-1:0] node10228;
	wire [4-1:0] node10229;
	wire [4-1:0] node10230;
	wire [4-1:0] node10231;
	wire [4-1:0] node10232;
	wire [4-1:0] node10235;
	wire [4-1:0] node10238;
	wire [4-1:0] node10240;
	wire [4-1:0] node10243;
	wire [4-1:0] node10244;
	wire [4-1:0] node10245;
	wire [4-1:0] node10248;
	wire [4-1:0] node10251;
	wire [4-1:0] node10252;
	wire [4-1:0] node10255;
	wire [4-1:0] node10258;
	wire [4-1:0] node10259;
	wire [4-1:0] node10261;
	wire [4-1:0] node10264;
	wire [4-1:0] node10267;
	wire [4-1:0] node10268;
	wire [4-1:0] node10269;
	wire [4-1:0] node10270;
	wire [4-1:0] node10271;
	wire [4-1:0] node10274;
	wire [4-1:0] node10277;
	wire [4-1:0] node10278;
	wire [4-1:0] node10280;
	wire [4-1:0] node10283;
	wire [4-1:0] node10285;
	wire [4-1:0] node10288;
	wire [4-1:0] node10289;
	wire [4-1:0] node10290;
	wire [4-1:0] node10293;
	wire [4-1:0] node10296;
	wire [4-1:0] node10297;
	wire [4-1:0] node10300;
	wire [4-1:0] node10303;
	wire [4-1:0] node10304;
	wire [4-1:0] node10305;
	wire [4-1:0] node10307;
	wire [4-1:0] node10310;
	wire [4-1:0] node10312;
	wire [4-1:0] node10315;
	wire [4-1:0] node10316;
	wire [4-1:0] node10317;
	wire [4-1:0] node10320;
	wire [4-1:0] node10323;
	wire [4-1:0] node10325;
	wire [4-1:0] node10328;
	wire [4-1:0] node10329;
	wire [4-1:0] node10330;
	wire [4-1:0] node10331;
	wire [4-1:0] node10332;
	wire [4-1:0] node10333;
	wire [4-1:0] node10336;
	wire [4-1:0] node10337;
	wire [4-1:0] node10339;
	wire [4-1:0] node10342;
	wire [4-1:0] node10343;
	wire [4-1:0] node10345;
	wire [4-1:0] node10349;
	wire [4-1:0] node10350;
	wire [4-1:0] node10351;
	wire [4-1:0] node10352;
	wire [4-1:0] node10353;
	wire [4-1:0] node10356;
	wire [4-1:0] node10359;
	wire [4-1:0] node10360;
	wire [4-1:0] node10363;
	wire [4-1:0] node10366;
	wire [4-1:0] node10367;
	wire [4-1:0] node10368;
	wire [4-1:0] node10372;
	wire [4-1:0] node10374;
	wire [4-1:0] node10377;
	wire [4-1:0] node10378;
	wire [4-1:0] node10379;
	wire [4-1:0] node10380;
	wire [4-1:0] node10383;
	wire [4-1:0] node10386;
	wire [4-1:0] node10387;
	wire [4-1:0] node10390;
	wire [4-1:0] node10393;
	wire [4-1:0] node10394;
	wire [4-1:0] node10395;
	wire [4-1:0] node10399;
	wire [4-1:0] node10400;
	wire [4-1:0] node10403;
	wire [4-1:0] node10406;
	wire [4-1:0] node10407;
	wire [4-1:0] node10408;
	wire [4-1:0] node10410;
	wire [4-1:0] node10412;
	wire [4-1:0] node10413;
	wire [4-1:0] node10416;
	wire [4-1:0] node10419;
	wire [4-1:0] node10421;
	wire [4-1:0] node10422;
	wire [4-1:0] node10423;
	wire [4-1:0] node10427;
	wire [4-1:0] node10430;
	wire [4-1:0] node10431;
	wire [4-1:0] node10432;
	wire [4-1:0] node10434;
	wire [4-1:0] node10436;
	wire [4-1:0] node10439;
	wire [4-1:0] node10440;
	wire [4-1:0] node10443;
	wire [4-1:0] node10446;
	wire [4-1:0] node10447;
	wire [4-1:0] node10448;
	wire [4-1:0] node10449;
	wire [4-1:0] node10452;
	wire [4-1:0] node10456;
	wire [4-1:0] node10457;
	wire [4-1:0] node10460;
	wire [4-1:0] node10462;
	wire [4-1:0] node10465;
	wire [4-1:0] node10466;
	wire [4-1:0] node10467;
	wire [4-1:0] node10468;
	wire [4-1:0] node10469;
	wire [4-1:0] node10470;
	wire [4-1:0] node10472;
	wire [4-1:0] node10475;
	wire [4-1:0] node10478;
	wire [4-1:0] node10479;
	wire [4-1:0] node10482;
	wire [4-1:0] node10483;
	wire [4-1:0] node10487;
	wire [4-1:0] node10489;
	wire [4-1:0] node10490;
	wire [4-1:0] node10493;
	wire [4-1:0] node10494;
	wire [4-1:0] node10497;
	wire [4-1:0] node10500;
	wire [4-1:0] node10501;
	wire [4-1:0] node10502;
	wire [4-1:0] node10503;
	wire [4-1:0] node10505;
	wire [4-1:0] node10509;
	wire [4-1:0] node10510;
	wire [4-1:0] node10511;
	wire [4-1:0] node10514;
	wire [4-1:0] node10517;
	wire [4-1:0] node10518;
	wire [4-1:0] node10519;
	wire [4-1:0] node10522;
	wire [4-1:0] node10525;
	wire [4-1:0] node10527;
	wire [4-1:0] node10530;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10533;
	wire [4-1:0] node10537;
	wire [4-1:0] node10539;
	wire [4-1:0] node10542;
	wire [4-1:0] node10543;
	wire [4-1:0] node10546;
	wire [4-1:0] node10548;
	wire [4-1:0] node10551;
	wire [4-1:0] node10552;
	wire [4-1:0] node10553;
	wire [4-1:0] node10554;
	wire [4-1:0] node10555;
	wire [4-1:0] node10558;
	wire [4-1:0] node10559;
	wire [4-1:0] node10562;
	wire [4-1:0] node10565;
	wire [4-1:0] node10566;
	wire [4-1:0] node10568;
	wire [4-1:0] node10572;
	wire [4-1:0] node10573;
	wire [4-1:0] node10574;
	wire [4-1:0] node10576;
	wire [4-1:0] node10579;
	wire [4-1:0] node10580;
	wire [4-1:0] node10584;
	wire [4-1:0] node10585;
	wire [4-1:0] node10588;
	wire [4-1:0] node10589;
	wire [4-1:0] node10593;
	wire [4-1:0] node10594;
	wire [4-1:0] node10595;
	wire [4-1:0] node10596;
	wire [4-1:0] node10597;
	wire [4-1:0] node10601;
	wire [4-1:0] node10604;
	wire [4-1:0] node10605;
	wire [4-1:0] node10608;
	wire [4-1:0] node10609;
	wire [4-1:0] node10613;
	wire [4-1:0] node10614;
	wire [4-1:0] node10615;
	wire [4-1:0] node10616;
	wire [4-1:0] node10619;
	wire [4-1:0] node10622;
	wire [4-1:0] node10624;
	wire [4-1:0] node10627;
	wire [4-1:0] node10628;
	wire [4-1:0] node10629;
	wire [4-1:0] node10633;
	wire [4-1:0] node10634;
	wire [4-1:0] node10637;
	wire [4-1:0] node10640;
	wire [4-1:0] node10641;
	wire [4-1:0] node10642;
	wire [4-1:0] node10643;
	wire [4-1:0] node10644;
	wire [4-1:0] node10645;
	wire [4-1:0] node10646;
	wire [4-1:0] node10649;
	wire [4-1:0] node10652;
	wire [4-1:0] node10653;
	wire [4-1:0] node10656;
	wire [4-1:0] node10659;
	wire [4-1:0] node10660;
	wire [4-1:0] node10661;
	wire [4-1:0] node10664;
	wire [4-1:0] node10667;
	wire [4-1:0] node10668;
	wire [4-1:0] node10671;
	wire [4-1:0] node10674;
	wire [4-1:0] node10675;
	wire [4-1:0] node10676;
	wire [4-1:0] node10677;
	wire [4-1:0] node10678;
	wire [4-1:0] node10681;
	wire [4-1:0] node10685;
	wire [4-1:0] node10686;
	wire [4-1:0] node10689;
	wire [4-1:0] node10692;
	wire [4-1:0] node10693;
	wire [4-1:0] node10694;
	wire [4-1:0] node10695;
	wire [4-1:0] node10699;
	wire [4-1:0] node10701;
	wire [4-1:0] node10704;
	wire [4-1:0] node10705;
	wire [4-1:0] node10708;
	wire [4-1:0] node10711;
	wire [4-1:0] node10712;
	wire [4-1:0] node10713;
	wire [4-1:0] node10714;
	wire [4-1:0] node10715;
	wire [4-1:0] node10718;
	wire [4-1:0] node10721;
	wire [4-1:0] node10722;
	wire [4-1:0] node10725;
	wire [4-1:0] node10728;
	wire [4-1:0] node10729;
	wire [4-1:0] node10730;
	wire [4-1:0] node10733;
	wire [4-1:0] node10736;
	wire [4-1:0] node10737;
	wire [4-1:0] node10739;
	wire [4-1:0] node10742;
	wire [4-1:0] node10744;
	wire [4-1:0] node10746;
	wire [4-1:0] node10749;
	wire [4-1:0] node10750;
	wire [4-1:0] node10751;
	wire [4-1:0] node10752;
	wire [4-1:0] node10755;
	wire [4-1:0] node10756;
	wire [4-1:0] node10759;
	wire [4-1:0] node10762;
	wire [4-1:0] node10763;
	wire [4-1:0] node10765;
	wire [4-1:0] node10768;
	wire [4-1:0] node10769;
	wire [4-1:0] node10773;
	wire [4-1:0] node10774;
	wire [4-1:0] node10775;
	wire [4-1:0] node10778;
	wire [4-1:0] node10781;
	wire [4-1:0] node10782;
	wire [4-1:0] node10783;
	wire [4-1:0] node10786;
	wire [4-1:0] node10789;
	wire [4-1:0] node10791;
	wire [4-1:0] node10794;
	wire [4-1:0] node10795;
	wire [4-1:0] node10796;
	wire [4-1:0] node10797;
	wire [4-1:0] node10798;
	wire [4-1:0] node10799;
	wire [4-1:0] node10802;
	wire [4-1:0] node10804;
	wire [4-1:0] node10807;
	wire [4-1:0] node10808;
	wire [4-1:0] node10810;
	wire [4-1:0] node10813;
	wire [4-1:0] node10814;
	wire [4-1:0] node10818;
	wire [4-1:0] node10819;
	wire [4-1:0] node10820;
	wire [4-1:0] node10821;
	wire [4-1:0] node10825;
	wire [4-1:0] node10826;
	wire [4-1:0] node10830;
	wire [4-1:0] node10831;
	wire [4-1:0] node10834;
	wire [4-1:0] node10836;
	wire [4-1:0] node10839;
	wire [4-1:0] node10840;
	wire [4-1:0] node10841;
	wire [4-1:0] node10842;
	wire [4-1:0] node10844;
	wire [4-1:0] node10847;
	wire [4-1:0] node10850;
	wire [4-1:0] node10851;
	wire [4-1:0] node10854;
	wire [4-1:0] node10856;
	wire [4-1:0] node10859;
	wire [4-1:0] node10860;
	wire [4-1:0] node10861;
	wire [4-1:0] node10862;
	wire [4-1:0] node10865;
	wire [4-1:0] node10868;
	wire [4-1:0] node10869;
	wire [4-1:0] node10872;
	wire [4-1:0] node10875;
	wire [4-1:0] node10876;
	wire [4-1:0] node10877;
	wire [4-1:0] node10880;
	wire [4-1:0] node10883;
	wire [4-1:0] node10886;
	wire [4-1:0] node10887;
	wire [4-1:0] node10888;
	wire [4-1:0] node10889;
	wire [4-1:0] node10890;
	wire [4-1:0] node10891;
	wire [4-1:0] node10895;
	wire [4-1:0] node10897;
	wire [4-1:0] node10900;
	wire [4-1:0] node10901;
	wire [4-1:0] node10903;
	wire [4-1:0] node10906;
	wire [4-1:0] node10909;
	wire [4-1:0] node10910;
	wire [4-1:0] node10911;
	wire [4-1:0] node10913;
	wire [4-1:0] node10916;
	wire [4-1:0] node10919;
	wire [4-1:0] node10920;
	wire [4-1:0] node10922;
	wire [4-1:0] node10925;
	wire [4-1:0] node10926;
	wire [4-1:0] node10930;
	wire [4-1:0] node10931;
	wire [4-1:0] node10932;
	wire [4-1:0] node10933;
	wire [4-1:0] node10934;
	wire [4-1:0] node10937;
	wire [4-1:0] node10940;
	wire [4-1:0] node10941;
	wire [4-1:0] node10944;
	wire [4-1:0] node10947;
	wire [4-1:0] node10948;
	wire [4-1:0] node10949;
	wire [4-1:0] node10952;
	wire [4-1:0] node10955;
	wire [4-1:0] node10956;
	wire [4-1:0] node10959;
	wire [4-1:0] node10962;
	wire [4-1:0] node10963;
	wire [4-1:0] node10964;
	wire [4-1:0] node10965;
	wire [4-1:0] node10968;
	wire [4-1:0] node10971;
	wire [4-1:0] node10972;
	wire [4-1:0] node10973;
	wire [4-1:0] node10976;
	wire [4-1:0] node10979;
	wire [4-1:0] node10980;
	wire [4-1:0] node10983;
	wire [4-1:0] node10986;
	wire [4-1:0] node10987;
	wire [4-1:0] node10988;
	wire [4-1:0] node10991;
	wire [4-1:0] node10994;
	wire [4-1:0] node10995;
	wire [4-1:0] node10998;
	wire [4-1:0] node11001;
	wire [4-1:0] node11002;
	wire [4-1:0] node11003;
	wire [4-1:0] node11004;
	wire [4-1:0] node11005;
	wire [4-1:0] node11006;
	wire [4-1:0] node11007;
	wire [4-1:0] node11008;
	wire [4-1:0] node11009;
	wire [4-1:0] node11010;
	wire [4-1:0] node11014;
	wire [4-1:0] node11018;
	wire [4-1:0] node11020;
	wire [4-1:0] node11021;
	wire [4-1:0] node11022;
	wire [4-1:0] node11025;
	wire [4-1:0] node11029;
	wire [4-1:0] node11030;
	wire [4-1:0] node11031;
	wire [4-1:0] node11032;
	wire [4-1:0] node11034;
	wire [4-1:0] node11037;
	wire [4-1:0] node11038;
	wire [4-1:0] node11039;
	wire [4-1:0] node11042;
	wire [4-1:0] node11046;
	wire [4-1:0] node11047;
	wire [4-1:0] node11049;
	wire [4-1:0] node11052;
	wire [4-1:0] node11053;
	wire [4-1:0] node11056;
	wire [4-1:0] node11059;
	wire [4-1:0] node11060;
	wire [4-1:0] node11061;
	wire [4-1:0] node11062;
	wire [4-1:0] node11065;
	wire [4-1:0] node11068;
	wire [4-1:0] node11069;
	wire [4-1:0] node11072;
	wire [4-1:0] node11075;
	wire [4-1:0] node11076;
	wire [4-1:0] node11078;
	wire [4-1:0] node11082;
	wire [4-1:0] node11083;
	wire [4-1:0] node11084;
	wire [4-1:0] node11086;
	wire [4-1:0] node11088;
	wire [4-1:0] node11089;
	wire [4-1:0] node11092;
	wire [4-1:0] node11095;
	wire [4-1:0] node11097;
	wire [4-1:0] node11098;
	wire [4-1:0] node11099;
	wire [4-1:0] node11102;
	wire [4-1:0] node11105;
	wire [4-1:0] node11106;
	wire [4-1:0] node11110;
	wire [4-1:0] node11111;
	wire [4-1:0] node11112;
	wire [4-1:0] node11114;
	wire [4-1:0] node11116;
	wire [4-1:0] node11119;
	wire [4-1:0] node11120;
	wire [4-1:0] node11121;
	wire [4-1:0] node11125;
	wire [4-1:0] node11128;
	wire [4-1:0] node11129;
	wire [4-1:0] node11130;
	wire [4-1:0] node11131;
	wire [4-1:0] node11134;
	wire [4-1:0] node11137;
	wire [4-1:0] node11138;
	wire [4-1:0] node11141;
	wire [4-1:0] node11144;
	wire [4-1:0] node11145;
	wire [4-1:0] node11147;
	wire [4-1:0] node11148;
	wire [4-1:0] node11151;
	wire [4-1:0] node11154;
	wire [4-1:0] node11156;
	wire [4-1:0] node11159;
	wire [4-1:0] node11160;
	wire [4-1:0] node11161;
	wire [4-1:0] node11162;
	wire [4-1:0] node11163;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11170;
	wire [4-1:0] node11171;
	wire [4-1:0] node11173;
	wire [4-1:0] node11176;
	wire [4-1:0] node11179;
	wire [4-1:0] node11180;
	wire [4-1:0] node11182;
	wire [4-1:0] node11183;
	wire [4-1:0] node11187;
	wire [4-1:0] node11188;
	wire [4-1:0] node11189;
	wire [4-1:0] node11192;
	wire [4-1:0] node11195;
	wire [4-1:0] node11196;
	wire [4-1:0] node11197;
	wire [4-1:0] node11200;
	wire [4-1:0] node11203;
	wire [4-1:0] node11204;
	wire [4-1:0] node11207;
	wire [4-1:0] node11210;
	wire [4-1:0] node11211;
	wire [4-1:0] node11212;
	wire [4-1:0] node11214;
	wire [4-1:0] node11215;
	wire [4-1:0] node11218;
	wire [4-1:0] node11221;
	wire [4-1:0] node11222;
	wire [4-1:0] node11223;
	wire [4-1:0] node11226;
	wire [4-1:0] node11229;
	wire [4-1:0] node11230;
	wire [4-1:0] node11234;
	wire [4-1:0] node11235;
	wire [4-1:0] node11236;
	wire [4-1:0] node11237;
	wire [4-1:0] node11241;
	wire [4-1:0] node11244;
	wire [4-1:0] node11245;
	wire [4-1:0] node11248;
	wire [4-1:0] node11249;
	wire [4-1:0] node11250;
	wire [4-1:0] node11253;
	wire [4-1:0] node11257;
	wire [4-1:0] node11258;
	wire [4-1:0] node11259;
	wire [4-1:0] node11260;
	wire [4-1:0] node11261;
	wire [4-1:0] node11265;
	wire [4-1:0] node11266;
	wire [4-1:0] node11270;
	wire [4-1:0] node11271;
	wire [4-1:0] node11272;
	wire [4-1:0] node11273;
	wire [4-1:0] node11277;
	wire [4-1:0] node11280;
	wire [4-1:0] node11281;
	wire [4-1:0] node11282;
	wire [4-1:0] node11285;
	wire [4-1:0] node11288;
	wire [4-1:0] node11289;
	wire [4-1:0] node11290;
	wire [4-1:0] node11295;
	wire [4-1:0] node11296;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11299;
	wire [4-1:0] node11302;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11310;
	wire [4-1:0] node11311;
	wire [4-1:0] node11314;
	wire [4-1:0] node11315;
	wire [4-1:0] node11319;
	wire [4-1:0] node11320;
	wire [4-1:0] node11321;
	wire [4-1:0] node11324;
	wire [4-1:0] node11327;
	wire [4-1:0] node11328;
	wire [4-1:0] node11330;
	wire [4-1:0] node11333;
	wire [4-1:0] node11334;
	wire [4-1:0] node11337;
	wire [4-1:0] node11340;
	wire [4-1:0] node11341;
	wire [4-1:0] node11342;
	wire [4-1:0] node11343;
	wire [4-1:0] node11344;
	wire [4-1:0] node11345;
	wire [4-1:0] node11346;
	wire [4-1:0] node11349;
	wire [4-1:0] node11352;
	wire [4-1:0] node11353;
	wire [4-1:0] node11354;
	wire [4-1:0] node11358;
	wire [4-1:0] node11360;
	wire [4-1:0] node11361;
	wire [4-1:0] node11364;
	wire [4-1:0] node11367;
	wire [4-1:0] node11368;
	wire [4-1:0] node11369;
	wire [4-1:0] node11371;
	wire [4-1:0] node11374;
	wire [4-1:0] node11377;
	wire [4-1:0] node11379;
	wire [4-1:0] node11381;
	wire [4-1:0] node11384;
	wire [4-1:0] node11385;
	wire [4-1:0] node11386;
	wire [4-1:0] node11387;
	wire [4-1:0] node11388;
	wire [4-1:0] node11391;
	wire [4-1:0] node11394;
	wire [4-1:0] node11395;
	wire [4-1:0] node11399;
	wire [4-1:0] node11400;
	wire [4-1:0] node11403;
	wire [4-1:0] node11404;
	wire [4-1:0] node11408;
	wire [4-1:0] node11409;
	wire [4-1:0] node11411;
	wire [4-1:0] node11414;
	wire [4-1:0] node11415;
	wire [4-1:0] node11416;
	wire [4-1:0] node11417;
	wire [4-1:0] node11420;
	wire [4-1:0] node11423;
	wire [4-1:0] node11424;
	wire [4-1:0] node11427;
	wire [4-1:0] node11431;
	wire [4-1:0] node11432;
	wire [4-1:0] node11433;
	wire [4-1:0] node11434;
	wire [4-1:0] node11435;
	wire [4-1:0] node11438;
	wire [4-1:0] node11440;
	wire [4-1:0] node11443;
	wire [4-1:0] node11444;
	wire [4-1:0] node11447;
	wire [4-1:0] node11449;
	wire [4-1:0] node11452;
	wire [4-1:0] node11453;
	wire [4-1:0] node11454;
	wire [4-1:0] node11455;
	wire [4-1:0] node11457;
	wire [4-1:0] node11460;
	wire [4-1:0] node11463;
	wire [4-1:0] node11464;
	wire [4-1:0] node11467;
	wire [4-1:0] node11470;
	wire [4-1:0] node11472;
	wire [4-1:0] node11475;
	wire [4-1:0] node11476;
	wire [4-1:0] node11477;
	wire [4-1:0] node11479;
	wire [4-1:0] node11480;
	wire [4-1:0] node11483;
	wire [4-1:0] node11486;
	wire [4-1:0] node11487;
	wire [4-1:0] node11490;
	wire [4-1:0] node11493;
	wire [4-1:0] node11494;
	wire [4-1:0] node11496;
	wire [4-1:0] node11498;
	wire [4-1:0] node11500;
	wire [4-1:0] node11503;
	wire [4-1:0] node11504;
	wire [4-1:0] node11507;
	wire [4-1:0] node11508;
	wire [4-1:0] node11512;
	wire [4-1:0] node11513;
	wire [4-1:0] node11514;
	wire [4-1:0] node11515;
	wire [4-1:0] node11516;
	wire [4-1:0] node11517;
	wire [4-1:0] node11519;
	wire [4-1:0] node11522;
	wire [4-1:0] node11523;
	wire [4-1:0] node11527;
	wire [4-1:0] node11528;
	wire [4-1:0] node11529;
	wire [4-1:0] node11532;
	wire [4-1:0] node11535;
	wire [4-1:0] node11536;
	wire [4-1:0] node11540;
	wire [4-1:0] node11541;
	wire [4-1:0] node11542;
	wire [4-1:0] node11544;
	wire [4-1:0] node11547;
	wire [4-1:0] node11550;
	wire [4-1:0] node11552;
	wire [4-1:0] node11553;
	wire [4-1:0] node11556;
	wire [4-1:0] node11559;
	wire [4-1:0] node11560;
	wire [4-1:0] node11561;
	wire [4-1:0] node11562;
	wire [4-1:0] node11563;
	wire [4-1:0] node11566;
	wire [4-1:0] node11569;
	wire [4-1:0] node11570;
	wire [4-1:0] node11574;
	wire [4-1:0] node11575;
	wire [4-1:0] node11576;
	wire [4-1:0] node11580;
	wire [4-1:0] node11581;
	wire [4-1:0] node11584;
	wire [4-1:0] node11587;
	wire [4-1:0] node11588;
	wire [4-1:0] node11589;
	wire [4-1:0] node11590;
	wire [4-1:0] node11593;
	wire [4-1:0] node11596;
	wire [4-1:0] node11597;
	wire [4-1:0] node11598;
	wire [4-1:0] node11601;
	wire [4-1:0] node11605;
	wire [4-1:0] node11606;
	wire [4-1:0] node11607;
	wire [4-1:0] node11609;
	wire [4-1:0] node11612;
	wire [4-1:0] node11613;
	wire [4-1:0] node11616;
	wire [4-1:0] node11619;
	wire [4-1:0] node11620;
	wire [4-1:0] node11621;
	wire [4-1:0] node11624;
	wire [4-1:0] node11627;
	wire [4-1:0] node11628;
	wire [4-1:0] node11632;
	wire [4-1:0] node11633;
	wire [4-1:0] node11634;
	wire [4-1:0] node11635;
	wire [4-1:0] node11636;
	wire [4-1:0] node11639;
	wire [4-1:0] node11640;
	wire [4-1:0] node11643;
	wire [4-1:0] node11646;
	wire [4-1:0] node11647;
	wire [4-1:0] node11649;
	wire [4-1:0] node11652;
	wire [4-1:0] node11654;
	wire [4-1:0] node11655;
	wire [4-1:0] node11658;
	wire [4-1:0] node11661;
	wire [4-1:0] node11662;
	wire [4-1:0] node11663;
	wire [4-1:0] node11666;
	wire [4-1:0] node11667;
	wire [4-1:0] node11670;
	wire [4-1:0] node11673;
	wire [4-1:0] node11674;
	wire [4-1:0] node11675;
	wire [4-1:0] node11678;
	wire [4-1:0] node11682;
	wire [4-1:0] node11683;
	wire [4-1:0] node11684;
	wire [4-1:0] node11685;
	wire [4-1:0] node11688;
	wire [4-1:0] node11690;
	wire [4-1:0] node11693;
	wire [4-1:0] node11694;
	wire [4-1:0] node11695;
	wire [4-1:0] node11696;
	wire [4-1:0] node11700;
	wire [4-1:0] node11702;
	wire [4-1:0] node11705;
	wire [4-1:0] node11706;
	wire [4-1:0] node11709;
	wire [4-1:0] node11712;
	wire [4-1:0] node11713;
	wire [4-1:0] node11714;
	wire [4-1:0] node11716;
	wire [4-1:0] node11719;
	wire [4-1:0] node11722;
	wire [4-1:0] node11723;
	wire [4-1:0] node11725;
	wire [4-1:0] node11728;
	wire [4-1:0] node11731;
	wire [4-1:0] node11732;
	wire [4-1:0] node11733;
	wire [4-1:0] node11734;
	wire [4-1:0] node11735;
	wire [4-1:0] node11736;
	wire [4-1:0] node11738;
	wire [4-1:0] node11739;
	wire [4-1:0] node11741;
	wire [4-1:0] node11744;
	wire [4-1:0] node11746;
	wire [4-1:0] node11749;
	wire [4-1:0] node11751;
	wire [4-1:0] node11752;
	wire [4-1:0] node11754;
	wire [4-1:0] node11757;
	wire [4-1:0] node11758;
	wire [4-1:0] node11762;
	wire [4-1:0] node11763;
	wire [4-1:0] node11764;
	wire [4-1:0] node11766;
	wire [4-1:0] node11767;
	wire [4-1:0] node11770;
	wire [4-1:0] node11773;
	wire [4-1:0] node11774;
	wire [4-1:0] node11775;
	wire [4-1:0] node11779;
	wire [4-1:0] node11780;
	wire [4-1:0] node11783;
	wire [4-1:0] node11786;
	wire [4-1:0] node11787;
	wire [4-1:0] node11788;
	wire [4-1:0] node11789;
	wire [4-1:0] node11790;
	wire [4-1:0] node11793;
	wire [4-1:0] node11797;
	wire [4-1:0] node11798;
	wire [4-1:0] node11801;
	wire [4-1:0] node11804;
	wire [4-1:0] node11805;
	wire [4-1:0] node11807;
	wire [4-1:0] node11811;
	wire [4-1:0] node11812;
	wire [4-1:0] node11813;
	wire [4-1:0] node11815;
	wire [4-1:0] node11817;
	wire [4-1:0] node11818;
	wire [4-1:0] node11821;
	wire [4-1:0] node11824;
	wire [4-1:0] node11826;
	wire [4-1:0] node11828;
	wire [4-1:0] node11829;
	wire [4-1:0] node11832;
	wire [4-1:0] node11835;
	wire [4-1:0] node11836;
	wire [4-1:0] node11837;
	wire [4-1:0] node11839;
	wire [4-1:0] node11841;
	wire [4-1:0] node11844;
	wire [4-1:0] node11845;
	wire [4-1:0] node11846;
	wire [4-1:0] node11850;
	wire [4-1:0] node11853;
	wire [4-1:0] node11854;
	wire [4-1:0] node11855;
	wire [4-1:0] node11856;
	wire [4-1:0] node11857;
	wire [4-1:0] node11860;
	wire [4-1:0] node11864;
	wire [4-1:0] node11865;
	wire [4-1:0] node11868;
	wire [4-1:0] node11871;
	wire [4-1:0] node11872;
	wire [4-1:0] node11873;
	wire [4-1:0] node11877;
	wire [4-1:0] node11879;
	wire [4-1:0] node11882;
	wire [4-1:0] node11883;
	wire [4-1:0] node11884;
	wire [4-1:0] node11885;
	wire [4-1:0] node11886;
	wire [4-1:0] node11888;
	wire [4-1:0] node11889;
	wire [4-1:0] node11893;
	wire [4-1:0] node11894;
	wire [4-1:0] node11896;
	wire [4-1:0] node11899;
	wire [4-1:0] node11901;
	wire [4-1:0] node11904;
	wire [4-1:0] node11905;
	wire [4-1:0] node11907;
	wire [4-1:0] node11909;
	wire [4-1:0] node11912;
	wire [4-1:0] node11913;
	wire [4-1:0] node11915;
	wire [4-1:0] node11918;
	wire [4-1:0] node11919;
	wire [4-1:0] node11922;
	wire [4-1:0] node11925;
	wire [4-1:0] node11926;
	wire [4-1:0] node11927;
	wire [4-1:0] node11928;
	wire [4-1:0] node11930;
	wire [4-1:0] node11933;
	wire [4-1:0] node11934;
	wire [4-1:0] node11937;
	wire [4-1:0] node11940;
	wire [4-1:0] node11941;
	wire [4-1:0] node11942;
	wire [4-1:0] node11945;
	wire [4-1:0] node11948;
	wire [4-1:0] node11949;
	wire [4-1:0] node11953;
	wire [4-1:0] node11954;
	wire [4-1:0] node11955;
	wire [4-1:0] node11956;
	wire [4-1:0] node11960;
	wire [4-1:0] node11963;
	wire [4-1:0] node11964;
	wire [4-1:0] node11967;
	wire [4-1:0] node11968;
	wire [4-1:0] node11971;
	wire [4-1:0] node11974;
	wire [4-1:0] node11975;
	wire [4-1:0] node11976;
	wire [4-1:0] node11977;
	wire [4-1:0] node11978;
	wire [4-1:0] node11982;
	wire [4-1:0] node11983;
	wire [4-1:0] node11987;
	wire [4-1:0] node11988;
	wire [4-1:0] node11989;
	wire [4-1:0] node11990;
	wire [4-1:0] node11994;
	wire [4-1:0] node11996;
	wire [4-1:0] node11999;
	wire [4-1:0] node12000;
	wire [4-1:0] node12001;
	wire [4-1:0] node12004;
	wire [4-1:0] node12007;
	wire [4-1:0] node12008;
	wire [4-1:0] node12012;
	wire [4-1:0] node12013;
	wire [4-1:0] node12014;
	wire [4-1:0] node12015;
	wire [4-1:0] node12016;
	wire [4-1:0] node12017;
	wire [4-1:0] node12020;
	wire [4-1:0] node12023;
	wire [4-1:0] node12026;
	wire [4-1:0] node12029;
	wire [4-1:0] node12030;
	wire [4-1:0] node12031;
	wire [4-1:0] node12033;
	wire [4-1:0] node12036;
	wire [4-1:0] node12039;
	wire [4-1:0] node12040;
	wire [4-1:0] node12043;
	wire [4-1:0] node12044;
	wire [4-1:0] node12048;
	wire [4-1:0] node12049;
	wire [4-1:0] node12050;
	wire [4-1:0] node12051;
	wire [4-1:0] node12053;
	wire [4-1:0] node12056;
	wire [4-1:0] node12058;
	wire [4-1:0] node12061;
	wire [4-1:0] node12062;
	wire [4-1:0] node12063;
	wire [4-1:0] node12067;
	wire [4-1:0] node12069;
	wire [4-1:0] node12072;
	wire [4-1:0] node12073;
	wire [4-1:0] node12074;
	wire [4-1:0] node12075;
	wire [4-1:0] node12079;
	wire [4-1:0] node12082;
	wire [4-1:0] node12083;
	wire [4-1:0] node12084;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12093;
	wire [4-1:0] node12094;
	wire [4-1:0] node12095;
	wire [4-1:0] node12096;
	wire [4-1:0] node12097;
	wire [4-1:0] node12098;
	wire [4-1:0] node12100;
	wire [4-1:0] node12101;
	wire [4-1:0] node12105;
	wire [4-1:0] node12106;
	wire [4-1:0] node12109;
	wire [4-1:0] node12110;
	wire [4-1:0] node12114;
	wire [4-1:0] node12115;
	wire [4-1:0] node12116;
	wire [4-1:0] node12119;
	wire [4-1:0] node12121;
	wire [4-1:0] node12124;
	wire [4-1:0] node12126;
	wire [4-1:0] node12127;
	wire [4-1:0] node12131;
	wire [4-1:0] node12132;
	wire [4-1:0] node12133;
	wire [4-1:0] node12134;
	wire [4-1:0] node12137;
	wire [4-1:0] node12140;
	wire [4-1:0] node12141;
	wire [4-1:0] node12144;
	wire [4-1:0] node12146;
	wire [4-1:0] node12149;
	wire [4-1:0] node12150;
	wire [4-1:0] node12152;
	wire [4-1:0] node12155;
	wire [4-1:0] node12156;
	wire [4-1:0] node12157;
	wire [4-1:0] node12160;
	wire [4-1:0] node12163;
	wire [4-1:0] node12164;
	wire [4-1:0] node12168;
	wire [4-1:0] node12169;
	wire [4-1:0] node12170;
	wire [4-1:0] node12171;
	wire [4-1:0] node12172;
	wire [4-1:0] node12175;
	wire [4-1:0] node12178;
	wire [4-1:0] node12179;
	wire [4-1:0] node12182;
	wire [4-1:0] node12183;
	wire [4-1:0] node12186;
	wire [4-1:0] node12189;
	wire [4-1:0] node12190;
	wire [4-1:0] node12191;
	wire [4-1:0] node12193;
	wire [4-1:0] node12196;
	wire [4-1:0] node12199;
	wire [4-1:0] node12200;
	wire [4-1:0] node12204;
	wire [4-1:0] node12205;
	wire [4-1:0] node12206;
	wire [4-1:0] node12207;
	wire [4-1:0] node12210;
	wire [4-1:0] node12212;
	wire [4-1:0] node12215;
	wire [4-1:0] node12216;
	wire [4-1:0] node12219;
	wire [4-1:0] node12222;
	wire [4-1:0] node12223;
	wire [4-1:0] node12225;
	wire [4-1:0] node12226;
	wire [4-1:0] node12230;
	wire [4-1:0] node12231;
	wire [4-1:0] node12234;
	wire [4-1:0] node12235;
	wire [4-1:0] node12239;
	wire [4-1:0] node12240;
	wire [4-1:0] node12241;
	wire [4-1:0] node12242;
	wire [4-1:0] node12243;
	wire [4-1:0] node12244;
	wire [4-1:0] node12247;
	wire [4-1:0] node12248;
	wire [4-1:0] node12252;
	wire [4-1:0] node12253;
	wire [4-1:0] node12254;
	wire [4-1:0] node12255;
	wire [4-1:0] node12258;
	wire [4-1:0] node12261;
	wire [4-1:0] node12262;
	wire [4-1:0] node12265;
	wire [4-1:0] node12268;
	wire [4-1:0] node12269;
	wire [4-1:0] node12273;
	wire [4-1:0] node12274;
	wire [4-1:0] node12275;
	wire [4-1:0] node12276;
	wire [4-1:0] node12280;
	wire [4-1:0] node12283;
	wire [4-1:0] node12285;
	wire [4-1:0] node12286;
	wire [4-1:0] node12289;
	wire [4-1:0] node12292;
	wire [4-1:0] node12293;
	wire [4-1:0] node12294;
	wire [4-1:0] node12295;
	wire [4-1:0] node12297;
	wire [4-1:0] node12300;
	wire [4-1:0] node12302;
	wire [4-1:0] node12305;
	wire [4-1:0] node12306;
	wire [4-1:0] node12309;
	wire [4-1:0] node12310;
	wire [4-1:0] node12313;
	wire [4-1:0] node12316;
	wire [4-1:0] node12317;
	wire [4-1:0] node12318;
	wire [4-1:0] node12321;
	wire [4-1:0] node12323;
	wire [4-1:0] node12326;
	wire [4-1:0] node12327;
	wire [4-1:0] node12328;
	wire [4-1:0] node12332;
	wire [4-1:0] node12333;
	wire [4-1:0] node12337;
	wire [4-1:0] node12338;
	wire [4-1:0] node12339;
	wire [4-1:0] node12340;
	wire [4-1:0] node12341;
	wire [4-1:0] node12343;
	wire [4-1:0] node12346;
	wire [4-1:0] node12347;
	wire [4-1:0] node12350;
	wire [4-1:0] node12353;
	wire [4-1:0] node12354;
	wire [4-1:0] node12355;
	wire [4-1:0] node12358;
	wire [4-1:0] node12361;
	wire [4-1:0] node12363;
	wire [4-1:0] node12366;
	wire [4-1:0] node12367;
	wire [4-1:0] node12368;
	wire [4-1:0] node12371;
	wire [4-1:0] node12373;
	wire [4-1:0] node12376;
	wire [4-1:0] node12377;
	wire [4-1:0] node12379;
	wire [4-1:0] node12382;
	wire [4-1:0] node12385;
	wire [4-1:0] node12386;
	wire [4-1:0] node12387;
	wire [4-1:0] node12388;
	wire [4-1:0] node12389;
	wire [4-1:0] node12392;
	wire [4-1:0] node12395;
	wire [4-1:0] node12396;
	wire [4-1:0] node12399;
	wire [4-1:0] node12402;
	wire [4-1:0] node12403;
	wire [4-1:0] node12404;
	wire [4-1:0] node12407;
	wire [4-1:0] node12410;
	wire [4-1:0] node12412;
	wire [4-1:0] node12415;
	wire [4-1:0] node12416;
	wire [4-1:0] node12417;
	wire [4-1:0] node12418;
	wire [4-1:0] node12421;
	wire [4-1:0] node12424;
	wire [4-1:0] node12425;
	wire [4-1:0] node12428;
	wire [4-1:0] node12431;
	wire [4-1:0] node12433;
	wire [4-1:0] node12434;
	wire [4-1:0] node12438;
	wire [4-1:0] node12439;
	wire [4-1:0] node12440;
	wire [4-1:0] node12441;
	wire [4-1:0] node12442;
	wire [4-1:0] node12443;
	wire [4-1:0] node12444;
	wire [4-1:0] node12445;
	wire [4-1:0] node12446;
	wire [4-1:0] node12447;
	wire [4-1:0] node12448;
	wire [4-1:0] node12451;
	wire [4-1:0] node12454;
	wire [4-1:0] node12455;
	wire [4-1:0] node12457;
	wire [4-1:0] node12460;
	wire [4-1:0] node12462;
	wire [4-1:0] node12465;
	wire [4-1:0] node12466;
	wire [4-1:0] node12467;
	wire [4-1:0] node12468;
	wire [4-1:0] node12471;
	wire [4-1:0] node12474;
	wire [4-1:0] node12475;
	wire [4-1:0] node12478;
	wire [4-1:0] node12481;
	wire [4-1:0] node12482;
	wire [4-1:0] node12485;
	wire [4-1:0] node12486;
	wire [4-1:0] node12490;
	wire [4-1:0] node12491;
	wire [4-1:0] node12492;
	wire [4-1:0] node12494;
	wire [4-1:0] node12495;
	wire [4-1:0] node12498;
	wire [4-1:0] node12501;
	wire [4-1:0] node12502;
	wire [4-1:0] node12505;
	wire [4-1:0] node12508;
	wire [4-1:0] node12509;
	wire [4-1:0] node12510;
	wire [4-1:0] node12511;
	wire [4-1:0] node12515;
	wire [4-1:0] node12516;
	wire [4-1:0] node12520;
	wire [4-1:0] node12522;
	wire [4-1:0] node12523;
	wire [4-1:0] node12526;
	wire [4-1:0] node12529;
	wire [4-1:0] node12530;
	wire [4-1:0] node12531;
	wire [4-1:0] node12532;
	wire [4-1:0] node12533;
	wire [4-1:0] node12536;
	wire [4-1:0] node12539;
	wire [4-1:0] node12540;
	wire [4-1:0] node12542;
	wire [4-1:0] node12546;
	wire [4-1:0] node12547;
	wire [4-1:0] node12548;
	wire [4-1:0] node12549;
	wire [4-1:0] node12552;
	wire [4-1:0] node12556;
	wire [4-1:0] node12557;
	wire [4-1:0] node12561;
	wire [4-1:0] node12562;
	wire [4-1:0] node12563;
	wire [4-1:0] node12564;
	wire [4-1:0] node12566;
	wire [4-1:0] node12569;
	wire [4-1:0] node12571;
	wire [4-1:0] node12574;
	wire [4-1:0] node12575;
	wire [4-1:0] node12576;
	wire [4-1:0] node12580;
	wire [4-1:0] node12581;
	wire [4-1:0] node12585;
	wire [4-1:0] node12586;
	wire [4-1:0] node12588;
	wire [4-1:0] node12589;
	wire [4-1:0] node12592;
	wire [4-1:0] node12595;
	wire [4-1:0] node12596;
	wire [4-1:0] node12597;
	wire [4-1:0] node12600;
	wire [4-1:0] node12603;
	wire [4-1:0] node12605;
	wire [4-1:0] node12608;
	wire [4-1:0] node12609;
	wire [4-1:0] node12610;
	wire [4-1:0] node12611;
	wire [4-1:0] node12612;
	wire [4-1:0] node12613;
	wire [4-1:0] node12615;
	wire [4-1:0] node12618;
	wire [4-1:0] node12621;
	wire [4-1:0] node12622;
	wire [4-1:0] node12625;
	wire [4-1:0] node12627;
	wire [4-1:0] node12630;
	wire [4-1:0] node12631;
	wire [4-1:0] node12633;
	wire [4-1:0] node12636;
	wire [4-1:0] node12637;
	wire [4-1:0] node12639;
	wire [4-1:0] node12642;
	wire [4-1:0] node12645;
	wire [4-1:0] node12646;
	wire [4-1:0] node12647;
	wire [4-1:0] node12648;
	wire [4-1:0] node12649;
	wire [4-1:0] node12653;
	wire [4-1:0] node12654;
	wire [4-1:0] node12658;
	wire [4-1:0] node12659;
	wire [4-1:0] node12660;
	wire [4-1:0] node12665;
	wire [4-1:0] node12666;
	wire [4-1:0] node12668;
	wire [4-1:0] node12670;
	wire [4-1:0] node12673;
	wire [4-1:0] node12675;
	wire [4-1:0] node12677;
	wire [4-1:0] node12680;
	wire [4-1:0] node12681;
	wire [4-1:0] node12682;
	wire [4-1:0] node12683;
	wire [4-1:0] node12684;
	wire [4-1:0] node12687;
	wire [4-1:0] node12690;
	wire [4-1:0] node12691;
	wire [4-1:0] node12693;
	wire [4-1:0] node12696;
	wire [4-1:0] node12698;
	wire [4-1:0] node12701;
	wire [4-1:0] node12702;
	wire [4-1:0] node12703;
	wire [4-1:0] node12707;
	wire [4-1:0] node12708;
	wire [4-1:0] node12711;
	wire [4-1:0] node12714;
	wire [4-1:0] node12715;
	wire [4-1:0] node12716;
	wire [4-1:0] node12717;
	wire [4-1:0] node12718;
	wire [4-1:0] node12721;
	wire [4-1:0] node12724;
	wire [4-1:0] node12725;
	wire [4-1:0] node12728;
	wire [4-1:0] node12731;
	wire [4-1:0] node12732;
	wire [4-1:0] node12736;
	wire [4-1:0] node12737;
	wire [4-1:0] node12738;
	wire [4-1:0] node12739;
	wire [4-1:0] node12744;
	wire [4-1:0] node12746;
	wire [4-1:0] node12747;
	wire [4-1:0] node12751;
	wire [4-1:0] node12752;
	wire [4-1:0] node12753;
	wire [4-1:0] node12754;
	wire [4-1:0] node12755;
	wire [4-1:0] node12756;
	wire [4-1:0] node12757;
	wire [4-1:0] node12760;
	wire [4-1:0] node12763;
	wire [4-1:0] node12765;
	wire [4-1:0] node12767;
	wire [4-1:0] node12770;
	wire [4-1:0] node12771;
	wire [4-1:0] node12772;
	wire [4-1:0] node12775;
	wire [4-1:0] node12776;
	wire [4-1:0] node12780;
	wire [4-1:0] node12781;
	wire [4-1:0] node12782;
	wire [4-1:0] node12786;
	wire [4-1:0] node12788;
	wire [4-1:0] node12791;
	wire [4-1:0] node12792;
	wire [4-1:0] node12793;
	wire [4-1:0] node12794;
	wire [4-1:0] node12797;
	wire [4-1:0] node12800;
	wire [4-1:0] node12801;
	wire [4-1:0] node12804;
	wire [4-1:0] node12807;
	wire [4-1:0] node12808;
	wire [4-1:0] node12810;
	wire [4-1:0] node12811;
	wire [4-1:0] node12814;
	wire [4-1:0] node12817;
	wire [4-1:0] node12818;
	wire [4-1:0] node12819;
	wire [4-1:0] node12822;
	wire [4-1:0] node12825;
	wire [4-1:0] node12826;
	wire [4-1:0] node12829;
	wire [4-1:0] node12832;
	wire [4-1:0] node12833;
	wire [4-1:0] node12834;
	wire [4-1:0] node12835;
	wire [4-1:0] node12836;
	wire [4-1:0] node12840;
	wire [4-1:0] node12841;
	wire [4-1:0] node12843;
	wire [4-1:0] node12846;
	wire [4-1:0] node12848;
	wire [4-1:0] node12851;
	wire [4-1:0] node12852;
	wire [4-1:0] node12853;
	wire [4-1:0] node12854;
	wire [4-1:0] node12857;
	wire [4-1:0] node12860;
	wire [4-1:0] node12861;
	wire [4-1:0] node12865;
	wire [4-1:0] node12866;
	wire [4-1:0] node12868;
	wire [4-1:0] node12871;
	wire [4-1:0] node12872;
	wire [4-1:0] node12876;
	wire [4-1:0] node12877;
	wire [4-1:0] node12878;
	wire [4-1:0] node12880;
	wire [4-1:0] node12881;
	wire [4-1:0] node12885;
	wire [4-1:0] node12886;
	wire [4-1:0] node12888;
	wire [4-1:0] node12891;
	wire [4-1:0] node12892;
	wire [4-1:0] node12895;
	wire [4-1:0] node12898;
	wire [4-1:0] node12899;
	wire [4-1:0] node12900;
	wire [4-1:0] node12903;
	wire [4-1:0] node12906;
	wire [4-1:0] node12907;
	wire [4-1:0] node12908;
	wire [4-1:0] node12911;
	wire [4-1:0] node12914;
	wire [4-1:0] node12915;
	wire [4-1:0] node12918;
	wire [4-1:0] node12921;
	wire [4-1:0] node12922;
	wire [4-1:0] node12923;
	wire [4-1:0] node12924;
	wire [4-1:0] node12926;
	wire [4-1:0] node12927;
	wire [4-1:0] node12929;
	wire [4-1:0] node12932;
	wire [4-1:0] node12934;
	wire [4-1:0] node12937;
	wire [4-1:0] node12938;
	wire [4-1:0] node12941;
	wire [4-1:0] node12942;
	wire [4-1:0] node12943;
	wire [4-1:0] node12946;
	wire [4-1:0] node12949;
	wire [4-1:0] node12950;
	wire [4-1:0] node12953;
	wire [4-1:0] node12956;
	wire [4-1:0] node12957;
	wire [4-1:0] node12958;
	wire [4-1:0] node12959;
	wire [4-1:0] node12961;
	wire [4-1:0] node12965;
	wire [4-1:0] node12966;
	wire [4-1:0] node12967;
	wire [4-1:0] node12970;
	wire [4-1:0] node12973;
	wire [4-1:0] node12974;
	wire [4-1:0] node12977;
	wire [4-1:0] node12980;
	wire [4-1:0] node12981;
	wire [4-1:0] node12982;
	wire [4-1:0] node12984;
	wire [4-1:0] node12987;
	wire [4-1:0] node12989;
	wire [4-1:0] node12992;
	wire [4-1:0] node12993;
	wire [4-1:0] node12995;
	wire [4-1:0] node12999;
	wire [4-1:0] node13000;
	wire [4-1:0] node13001;
	wire [4-1:0] node13002;
	wire [4-1:0] node13003;
	wire [4-1:0] node13006;
	wire [4-1:0] node13007;
	wire [4-1:0] node13011;
	wire [4-1:0] node13012;
	wire [4-1:0] node13015;
	wire [4-1:0] node13016;
	wire [4-1:0] node13020;
	wire [4-1:0] node13021;
	wire [4-1:0] node13022;
	wire [4-1:0] node13025;
	wire [4-1:0] node13028;
	wire [4-1:0] node13029;
	wire [4-1:0] node13032;
	wire [4-1:0] node13035;
	wire [4-1:0] node13036;
	wire [4-1:0] node13037;
	wire [4-1:0] node13038;
	wire [4-1:0] node13039;
	wire [4-1:0] node13042;
	wire [4-1:0] node13045;
	wire [4-1:0] node13046;
	wire [4-1:0] node13049;
	wire [4-1:0] node13052;
	wire [4-1:0] node13053;
	wire [4-1:0] node13055;
	wire [4-1:0] node13059;
	wire [4-1:0] node13060;
	wire [4-1:0] node13061;
	wire [4-1:0] node13063;
	wire [4-1:0] node13066;
	wire [4-1:0] node13067;
	wire [4-1:0] node13071;
	wire [4-1:0] node13073;
	wire [4-1:0] node13074;
	wire [4-1:0] node13077;
	wire [4-1:0] node13080;
	wire [4-1:0] node13081;
	wire [4-1:0] node13082;
	wire [4-1:0] node13083;
	wire [4-1:0] node13084;
	wire [4-1:0] node13085;
	wire [4-1:0] node13086;
	wire [4-1:0] node13087;
	wire [4-1:0] node13089;
	wire [4-1:0] node13093;
	wire [4-1:0] node13095;
	wire [4-1:0] node13098;
	wire [4-1:0] node13099;
	wire [4-1:0] node13100;
	wire [4-1:0] node13101;
	wire [4-1:0] node13104;
	wire [4-1:0] node13108;
	wire [4-1:0] node13109;
	wire [4-1:0] node13112;
	wire [4-1:0] node13115;
	wire [4-1:0] node13116;
	wire [4-1:0] node13117;
	wire [4-1:0] node13118;
	wire [4-1:0] node13119;
	wire [4-1:0] node13122;
	wire [4-1:0] node13125;
	wire [4-1:0] node13126;
	wire [4-1:0] node13130;
	wire [4-1:0] node13131;
	wire [4-1:0] node13132;
	wire [4-1:0] node13136;
	wire [4-1:0] node13137;
	wire [4-1:0] node13141;
	wire [4-1:0] node13142;
	wire [4-1:0] node13144;
	wire [4-1:0] node13145;
	wire [4-1:0] node13148;
	wire [4-1:0] node13151;
	wire [4-1:0] node13152;
	wire [4-1:0] node13153;
	wire [4-1:0] node13156;
	wire [4-1:0] node13160;
	wire [4-1:0] node13161;
	wire [4-1:0] node13162;
	wire [4-1:0] node13163;
	wire [4-1:0] node13166;
	wire [4-1:0] node13167;
	wire [4-1:0] node13169;
	wire [4-1:0] node13172;
	wire [4-1:0] node13174;
	wire [4-1:0] node13177;
	wire [4-1:0] node13178;
	wire [4-1:0] node13179;
	wire [4-1:0] node13182;
	wire [4-1:0] node13185;
	wire [4-1:0] node13186;
	wire [4-1:0] node13190;
	wire [4-1:0] node13191;
	wire [4-1:0] node13192;
	wire [4-1:0] node13194;
	wire [4-1:0] node13196;
	wire [4-1:0] node13199;
	wire [4-1:0] node13200;
	wire [4-1:0] node13203;
	wire [4-1:0] node13205;
	wire [4-1:0] node13208;
	wire [4-1:0] node13209;
	wire [4-1:0] node13210;
	wire [4-1:0] node13212;
	wire [4-1:0] node13215;
	wire [4-1:0] node13216;
	wire [4-1:0] node13220;
	wire [4-1:0] node13221;
	wire [4-1:0] node13222;
	wire [4-1:0] node13226;
	wire [4-1:0] node13227;
	wire [4-1:0] node13231;
	wire [4-1:0] node13232;
	wire [4-1:0] node13233;
	wire [4-1:0] node13234;
	wire [4-1:0] node13235;
	wire [4-1:0] node13236;
	wire [4-1:0] node13239;
	wire [4-1:0] node13242;
	wire [4-1:0] node13243;
	wire [4-1:0] node13245;
	wire [4-1:0] node13249;
	wire [4-1:0] node13250;
	wire [4-1:0] node13251;
	wire [4-1:0] node13252;
	wire [4-1:0] node13255;
	wire [4-1:0] node13259;
	wire [4-1:0] node13260;
	wire [4-1:0] node13261;
	wire [4-1:0] node13265;
	wire [4-1:0] node13266;
	wire [4-1:0] node13269;
	wire [4-1:0] node13272;
	wire [4-1:0] node13273;
	wire [4-1:0] node13274;
	wire [4-1:0] node13275;
	wire [4-1:0] node13278;
	wire [4-1:0] node13281;
	wire [4-1:0] node13282;
	wire [4-1:0] node13285;
	wire [4-1:0] node13288;
	wire [4-1:0] node13289;
	wire [4-1:0] node13290;
	wire [4-1:0] node13291;
	wire [4-1:0] node13294;
	wire [4-1:0] node13298;
	wire [4-1:0] node13299;
	wire [4-1:0] node13300;
	wire [4-1:0] node13303;
	wire [4-1:0] node13306;
	wire [4-1:0] node13307;
	wire [4-1:0] node13310;
	wire [4-1:0] node13313;
	wire [4-1:0] node13314;
	wire [4-1:0] node13315;
	wire [4-1:0] node13316;
	wire [4-1:0] node13317;
	wire [4-1:0] node13319;
	wire [4-1:0] node13322;
	wire [4-1:0] node13325;
	wire [4-1:0] node13326;
	wire [4-1:0] node13327;
	wire [4-1:0] node13331;
	wire [4-1:0] node13332;
	wire [4-1:0] node13336;
	wire [4-1:0] node13337;
	wire [4-1:0] node13338;
	wire [4-1:0] node13339;
	wire [4-1:0] node13342;
	wire [4-1:0] node13345;
	wire [4-1:0] node13348;
	wire [4-1:0] node13349;
	wire [4-1:0] node13350;
	wire [4-1:0] node13353;
	wire [4-1:0] node13356;
	wire [4-1:0] node13357;
	wire [4-1:0] node13361;
	wire [4-1:0] node13362;
	wire [4-1:0] node13363;
	wire [4-1:0] node13364;
	wire [4-1:0] node13368;
	wire [4-1:0] node13369;
	wire [4-1:0] node13372;
	wire [4-1:0] node13375;
	wire [4-1:0] node13376;
	wire [4-1:0] node13377;
	wire [4-1:0] node13378;
	wire [4-1:0] node13381;
	wire [4-1:0] node13384;
	wire [4-1:0] node13385;
	wire [4-1:0] node13388;
	wire [4-1:0] node13391;
	wire [4-1:0] node13392;
	wire [4-1:0] node13393;
	wire [4-1:0] node13396;
	wire [4-1:0] node13400;
	wire [4-1:0] node13401;
	wire [4-1:0] node13402;
	wire [4-1:0] node13403;
	wire [4-1:0] node13404;
	wire [4-1:0] node13405;
	wire [4-1:0] node13406;
	wire [4-1:0] node13409;
	wire [4-1:0] node13412;
	wire [4-1:0] node13413;
	wire [4-1:0] node13416;
	wire [4-1:0] node13419;
	wire [4-1:0] node13420;
	wire [4-1:0] node13423;
	wire [4-1:0] node13426;
	wire [4-1:0] node13427;
	wire [4-1:0] node13428;
	wire [4-1:0] node13429;
	wire [4-1:0] node13430;
	wire [4-1:0] node13433;
	wire [4-1:0] node13436;
	wire [4-1:0] node13437;
	wire [4-1:0] node13441;
	wire [4-1:0] node13442;
	wire [4-1:0] node13446;
	wire [4-1:0] node13447;
	wire [4-1:0] node13448;
	wire [4-1:0] node13451;
	wire [4-1:0] node13454;
	wire [4-1:0] node13455;
	wire [4-1:0] node13458;
	wire [4-1:0] node13461;
	wire [4-1:0] node13462;
	wire [4-1:0] node13463;
	wire [4-1:0] node13464;
	wire [4-1:0] node13465;
	wire [4-1:0] node13466;
	wire [4-1:0] node13469;
	wire [4-1:0] node13472;
	wire [4-1:0] node13473;
	wire [4-1:0] node13477;
	wire [4-1:0] node13478;
	wire [4-1:0] node13481;
	wire [4-1:0] node13484;
	wire [4-1:0] node13485;
	wire [4-1:0] node13486;
	wire [4-1:0] node13487;
	wire [4-1:0] node13490;
	wire [4-1:0] node13493;
	wire [4-1:0] node13494;
	wire [4-1:0] node13497;
	wire [4-1:0] node13500;
	wire [4-1:0] node13501;
	wire [4-1:0] node13502;
	wire [4-1:0] node13505;
	wire [4-1:0] node13509;
	wire [4-1:0] node13510;
	wire [4-1:0] node13511;
	wire [4-1:0] node13512;
	wire [4-1:0] node13514;
	wire [4-1:0] node13517;
	wire [4-1:0] node13519;
	wire [4-1:0] node13522;
	wire [4-1:0] node13523;
	wire [4-1:0] node13524;
	wire [4-1:0] node13527;
	wire [4-1:0] node13530;
	wire [4-1:0] node13531;
	wire [4-1:0] node13534;
	wire [4-1:0] node13537;
	wire [4-1:0] node13538;
	wire [4-1:0] node13539;
	wire [4-1:0] node13540;
	wire [4-1:0] node13543;
	wire [4-1:0] node13547;
	wire [4-1:0] node13549;
	wire [4-1:0] node13550;
	wire [4-1:0] node13553;
	wire [4-1:0] node13556;
	wire [4-1:0] node13557;
	wire [4-1:0] node13558;
	wire [4-1:0] node13559;
	wire [4-1:0] node13560;
	wire [4-1:0] node13561;
	wire [4-1:0] node13563;
	wire [4-1:0] node13566;
	wire [4-1:0] node13567;
	wire [4-1:0] node13570;
	wire [4-1:0] node13573;
	wire [4-1:0] node13574;
	wire [4-1:0] node13575;
	wire [4-1:0] node13578;
	wire [4-1:0] node13582;
	wire [4-1:0] node13583;
	wire [4-1:0] node13585;
	wire [4-1:0] node13588;
	wire [4-1:0] node13589;
	wire [4-1:0] node13592;
	wire [4-1:0] node13595;
	wire [4-1:0] node13596;
	wire [4-1:0] node13597;
	wire [4-1:0] node13598;
	wire [4-1:0] node13599;
	wire [4-1:0] node13603;
	wire [4-1:0] node13604;
	wire [4-1:0] node13608;
	wire [4-1:0] node13609;
	wire [4-1:0] node13610;
	wire [4-1:0] node13614;
	wire [4-1:0] node13615;
	wire [4-1:0] node13619;
	wire [4-1:0] node13620;
	wire [4-1:0] node13621;
	wire [4-1:0] node13623;
	wire [4-1:0] node13626;
	wire [4-1:0] node13627;
	wire [4-1:0] node13630;
	wire [4-1:0] node13633;
	wire [4-1:0] node13634;
	wire [4-1:0] node13635;
	wire [4-1:0] node13638;
	wire [4-1:0] node13641;
	wire [4-1:0] node13642;
	wire [4-1:0] node13646;
	wire [4-1:0] node13647;
	wire [4-1:0] node13648;
	wire [4-1:0] node13649;
	wire [4-1:0] node13650;
	wire [4-1:0] node13653;
	wire [4-1:0] node13656;
	wire [4-1:0] node13657;
	wire [4-1:0] node13658;
	wire [4-1:0] node13662;
	wire [4-1:0] node13663;
	wire [4-1:0] node13666;
	wire [4-1:0] node13669;
	wire [4-1:0] node13670;
	wire [4-1:0] node13671;
	wire [4-1:0] node13672;
	wire [4-1:0] node13675;
	wire [4-1:0] node13678;
	wire [4-1:0] node13679;
	wire [4-1:0] node13683;
	wire [4-1:0] node13684;
	wire [4-1:0] node13687;
	wire [4-1:0] node13690;
	wire [4-1:0] node13691;
	wire [4-1:0] node13692;
	wire [4-1:0] node13693;
	wire [4-1:0] node13696;
	wire [4-1:0] node13699;
	wire [4-1:0] node13700;
	wire [4-1:0] node13702;
	wire [4-1:0] node13705;
	wire [4-1:0] node13707;
	wire [4-1:0] node13710;
	wire [4-1:0] node13711;
	wire [4-1:0] node13713;
	wire [4-1:0] node13714;
	wire [4-1:0] node13717;
	wire [4-1:0] node13720;
	wire [4-1:0] node13721;
	wire [4-1:0] node13722;
	wire [4-1:0] node13727;
	wire [4-1:0] node13728;
	wire [4-1:0] node13729;
	wire [4-1:0] node13730;
	wire [4-1:0] node13731;
	wire [4-1:0] node13732;
	wire [4-1:0] node13733;
	wire [4-1:0] node13734;
	wire [4-1:0] node13736;
	wire [4-1:0] node13737;
	wire [4-1:0] node13741;
	wire [4-1:0] node13743;
	wire [4-1:0] node13746;
	wire [4-1:0] node13747;
	wire [4-1:0] node13750;
	wire [4-1:0] node13751;
	wire [4-1:0] node13755;
	wire [4-1:0] node13756;
	wire [4-1:0] node13757;
	wire [4-1:0] node13758;
	wire [4-1:0] node13761;
	wire [4-1:0] node13764;
	wire [4-1:0] node13765;
	wire [4-1:0] node13768;
	wire [4-1:0] node13771;
	wire [4-1:0] node13772;
	wire [4-1:0] node13773;
	wire [4-1:0] node13777;
	wire [4-1:0] node13778;
	wire [4-1:0] node13781;
	wire [4-1:0] node13784;
	wire [4-1:0] node13785;
	wire [4-1:0] node13786;
	wire [4-1:0] node13787;
	wire [4-1:0] node13788;
	wire [4-1:0] node13791;
	wire [4-1:0] node13792;
	wire [4-1:0] node13796;
	wire [4-1:0] node13797;
	wire [4-1:0] node13800;
	wire [4-1:0] node13802;
	wire [4-1:0] node13805;
	wire [4-1:0] node13806;
	wire [4-1:0] node13808;
	wire [4-1:0] node13810;
	wire [4-1:0] node13813;
	wire [4-1:0] node13816;
	wire [4-1:0] node13817;
	wire [4-1:0] node13818;
	wire [4-1:0] node13819;
	wire [4-1:0] node13822;
	wire [4-1:0] node13823;
	wire [4-1:0] node13826;
	wire [4-1:0] node13829;
	wire [4-1:0] node13830;
	wire [4-1:0] node13833;
	wire [4-1:0] node13836;
	wire [4-1:0] node13837;
	wire [4-1:0] node13839;
	wire [4-1:0] node13842;
	wire [4-1:0] node13843;
	wire [4-1:0] node13844;
	wire [4-1:0] node13847;
	wire [4-1:0] node13851;
	wire [4-1:0] node13852;
	wire [4-1:0] node13853;
	wire [4-1:0] node13854;
	wire [4-1:0] node13855;
	wire [4-1:0] node13856;
	wire [4-1:0] node13859;
	wire [4-1:0] node13862;
	wire [4-1:0] node13863;
	wire [4-1:0] node13866;
	wire [4-1:0] node13869;
	wire [4-1:0] node13870;
	wire [4-1:0] node13871;
	wire [4-1:0] node13874;
	wire [4-1:0] node13877;
	wire [4-1:0] node13878;
	wire [4-1:0] node13881;
	wire [4-1:0] node13884;
	wire [4-1:0] node13885;
	wire [4-1:0] node13886;
	wire [4-1:0] node13887;
	wire [4-1:0] node13890;
	wire [4-1:0] node13893;
	wire [4-1:0] node13895;
	wire [4-1:0] node13896;
	wire [4-1:0] node13900;
	wire [4-1:0] node13901;
	wire [4-1:0] node13902;
	wire [4-1:0] node13906;
	wire [4-1:0] node13907;
	wire [4-1:0] node13910;
	wire [4-1:0] node13913;
	wire [4-1:0] node13914;
	wire [4-1:0] node13915;
	wire [4-1:0] node13916;
	wire [4-1:0] node13917;
	wire [4-1:0] node13918;
	wire [4-1:0] node13922;
	wire [4-1:0] node13924;
	wire [4-1:0] node13927;
	wire [4-1:0] node13928;
	wire [4-1:0] node13929;
	wire [4-1:0] node13932;
	wire [4-1:0] node13935;
	wire [4-1:0] node13937;
	wire [4-1:0] node13940;
	wire [4-1:0] node13941;
	wire [4-1:0] node13942;
	wire [4-1:0] node13945;
	wire [4-1:0] node13948;
	wire [4-1:0] node13949;
	wire [4-1:0] node13952;
	wire [4-1:0] node13955;
	wire [4-1:0] node13956;
	wire [4-1:0] node13957;
	wire [4-1:0] node13959;
	wire [4-1:0] node13962;
	wire [4-1:0] node13963;
	wire [4-1:0] node13964;
	wire [4-1:0] node13967;
	wire [4-1:0] node13971;
	wire [4-1:0] node13972;
	wire [4-1:0] node13973;
	wire [4-1:0] node13974;
	wire [4-1:0] node13978;
	wire [4-1:0] node13979;
	wire [4-1:0] node13982;
	wire [4-1:0] node13985;
	wire [4-1:0] node13986;
	wire [4-1:0] node13989;
	wire [4-1:0] node13992;
	wire [4-1:0] node13993;
	wire [4-1:0] node13994;
	wire [4-1:0] node13995;
	wire [4-1:0] node13996;
	wire [4-1:0] node13997;
	wire [4-1:0] node13998;
	wire [4-1:0] node14001;
	wire [4-1:0] node14004;
	wire [4-1:0] node14005;
	wire [4-1:0] node14008;
	wire [4-1:0] node14011;
	wire [4-1:0] node14012;
	wire [4-1:0] node14013;
	wire [4-1:0] node14016;
	wire [4-1:0] node14019;
	wire [4-1:0] node14020;
	wire [4-1:0] node14023;
	wire [4-1:0] node14026;
	wire [4-1:0] node14027;
	wire [4-1:0] node14028;
	wire [4-1:0] node14029;
	wire [4-1:0] node14032;
	wire [4-1:0] node14035;
	wire [4-1:0] node14036;
	wire [4-1:0] node14039;
	wire [4-1:0] node14042;
	wire [4-1:0] node14043;
	wire [4-1:0] node14045;
	wire [4-1:0] node14048;
	wire [4-1:0] node14049;
	wire [4-1:0] node14052;
	wire [4-1:0] node14055;
	wire [4-1:0] node14056;
	wire [4-1:0] node14057;
	wire [4-1:0] node14058;
	wire [4-1:0] node14059;
	wire [4-1:0] node14062;
	wire [4-1:0] node14065;
	wire [4-1:0] node14066;
	wire [4-1:0] node14069;
	wire [4-1:0] node14072;
	wire [4-1:0] node14073;
	wire [4-1:0] node14074;
	wire [4-1:0] node14077;
	wire [4-1:0] node14080;
	wire [4-1:0] node14081;
	wire [4-1:0] node14085;
	wire [4-1:0] node14086;
	wire [4-1:0] node14087;
	wire [4-1:0] node14088;
	wire [4-1:0] node14091;
	wire [4-1:0] node14094;
	wire [4-1:0] node14095;
	wire [4-1:0] node14098;
	wire [4-1:0] node14101;
	wire [4-1:0] node14102;
	wire [4-1:0] node14104;
	wire [4-1:0] node14107;
	wire [4-1:0] node14108;
	wire [4-1:0] node14111;
	wire [4-1:0] node14114;
	wire [4-1:0] node14115;
	wire [4-1:0] node14116;
	wire [4-1:0] node14117;
	wire [4-1:0] node14118;
	wire [4-1:0] node14120;
	wire [4-1:0] node14122;
	wire [4-1:0] node14125;
	wire [4-1:0] node14126;
	wire [4-1:0] node14129;
	wire [4-1:0] node14132;
	wire [4-1:0] node14133;
	wire [4-1:0] node14135;
	wire [4-1:0] node14138;
	wire [4-1:0] node14139;
	wire [4-1:0] node14142;
	wire [4-1:0] node14145;
	wire [4-1:0] node14146;
	wire [4-1:0] node14147;
	wire [4-1:0] node14148;
	wire [4-1:0] node14151;
	wire [4-1:0] node14154;
	wire [4-1:0] node14156;
	wire [4-1:0] node14159;
	wire [4-1:0] node14160;
	wire [4-1:0] node14162;
	wire [4-1:0] node14163;
	wire [4-1:0] node14166;
	wire [4-1:0] node14169;
	wire [4-1:0] node14171;
	wire [4-1:0] node14174;
	wire [4-1:0] node14175;
	wire [4-1:0] node14176;
	wire [4-1:0] node14177;
	wire [4-1:0] node14178;
	wire [4-1:0] node14181;
	wire [4-1:0] node14184;
	wire [4-1:0] node14185;
	wire [4-1:0] node14188;
	wire [4-1:0] node14191;
	wire [4-1:0] node14192;
	wire [4-1:0] node14193;
	wire [4-1:0] node14194;
	wire [4-1:0] node14197;
	wire [4-1:0] node14200;
	wire [4-1:0] node14201;
	wire [4-1:0] node14205;
	wire [4-1:0] node14206;
	wire [4-1:0] node14207;
	wire [4-1:0] node14211;
	wire [4-1:0] node14212;
	wire [4-1:0] node14215;
	wire [4-1:0] node14218;
	wire [4-1:0] node14219;
	wire [4-1:0] node14220;
	wire [4-1:0] node14221;
	wire [4-1:0] node14225;
	wire [4-1:0] node14226;
	wire [4-1:0] node14229;
	wire [4-1:0] node14232;
	wire [4-1:0] node14233;
	wire [4-1:0] node14234;
	wire [4-1:0] node14237;
	wire [4-1:0] node14240;
	wire [4-1:0] node14241;
	wire [4-1:0] node14244;
	wire [4-1:0] node14247;
	wire [4-1:0] node14248;
	wire [4-1:0] node14249;
	wire [4-1:0] node14250;
	wire [4-1:0] node14251;
	wire [4-1:0] node14252;
	wire [4-1:0] node14253;
	wire [4-1:0] node14254;
	wire [4-1:0] node14257;
	wire [4-1:0] node14260;
	wire [4-1:0] node14261;
	wire [4-1:0] node14262;
	wire [4-1:0] node14266;
	wire [4-1:0] node14267;
	wire [4-1:0] node14271;
	wire [4-1:0] node14272;
	wire [4-1:0] node14273;
	wire [4-1:0] node14276;
	wire [4-1:0] node14279;
	wire [4-1:0] node14280;
	wire [4-1:0] node14283;
	wire [4-1:0] node14286;
	wire [4-1:0] node14287;
	wire [4-1:0] node14288;
	wire [4-1:0] node14289;
	wire [4-1:0] node14290;
	wire [4-1:0] node14293;
	wire [4-1:0] node14296;
	wire [4-1:0] node14297;
	wire [4-1:0] node14300;
	wire [4-1:0] node14303;
	wire [4-1:0] node14304;
	wire [4-1:0] node14307;
	wire [4-1:0] node14310;
	wire [4-1:0] node14311;
	wire [4-1:0] node14312;
	wire [4-1:0] node14315;
	wire [4-1:0] node14318;
	wire [4-1:0] node14320;
	wire [4-1:0] node14321;
	wire [4-1:0] node14324;
	wire [4-1:0] node14327;
	wire [4-1:0] node14328;
	wire [4-1:0] node14329;
	wire [4-1:0] node14330;
	wire [4-1:0] node14332;
	wire [4-1:0] node14335;
	wire [4-1:0] node14336;
	wire [4-1:0] node14339;
	wire [4-1:0] node14342;
	wire [4-1:0] node14343;
	wire [4-1:0] node14344;
	wire [4-1:0] node14346;
	wire [4-1:0] node14349;
	wire [4-1:0] node14350;
	wire [4-1:0] node14354;
	wire [4-1:0] node14355;
	wire [4-1:0] node14358;
	wire [4-1:0] node14361;
	wire [4-1:0] node14362;
	wire [4-1:0] node14364;
	wire [4-1:0] node14367;
	wire [4-1:0] node14368;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14373;
	wire [4-1:0] node14376;
	wire [4-1:0] node14378;
	wire [4-1:0] node14381;
	wire [4-1:0] node14382;
	wire [4-1:0] node14385;
	wire [4-1:0] node14388;
	wire [4-1:0] node14389;
	wire [4-1:0] node14390;
	wire [4-1:0] node14391;
	wire [4-1:0] node14392;
	wire [4-1:0] node14393;
	wire [4-1:0] node14396;
	wire [4-1:0] node14400;
	wire [4-1:0] node14401;
	wire [4-1:0] node14402;
	wire [4-1:0] node14403;
	wire [4-1:0] node14407;
	wire [4-1:0] node14411;
	wire [4-1:0] node14412;
	wire [4-1:0] node14413;
	wire [4-1:0] node14414;
	wire [4-1:0] node14415;
	wire [4-1:0] node14418;
	wire [4-1:0] node14421;
	wire [4-1:0] node14422;
	wire [4-1:0] node14425;
	wire [4-1:0] node14429;
	wire [4-1:0] node14430;
	wire [4-1:0] node14431;
	wire [4-1:0] node14434;
	wire [4-1:0] node14438;
	wire [4-1:0] node14439;
	wire [4-1:0] node14440;
	wire [4-1:0] node14441;
	wire [4-1:0] node14444;
	wire [4-1:0] node14447;
	wire [4-1:0] node14448;
	wire [4-1:0] node14451;
	wire [4-1:0] node14454;
	wire [4-1:0] node14455;
	wire [4-1:0] node14458;
	wire [4-1:0] node14461;
	wire [4-1:0] node14462;
	wire [4-1:0] node14463;
	wire [4-1:0] node14464;
	wire [4-1:0] node14465;
	wire [4-1:0] node14466;
	wire [4-1:0] node14469;
	wire [4-1:0] node14472;
	wire [4-1:0] node14473;
	wire [4-1:0] node14474;
	wire [4-1:0] node14477;
	wire [4-1:0] node14480;
	wire [4-1:0] node14481;
	wire [4-1:0] node14484;
	wire [4-1:0] node14487;
	wire [4-1:0] node14488;
	wire [4-1:0] node14489;
	wire [4-1:0] node14490;
	wire [4-1:0] node14491;
	wire [4-1:0] node14496;
	wire [4-1:0] node14497;
	wire [4-1:0] node14498;
	wire [4-1:0] node14501;
	wire [4-1:0] node14504;
	wire [4-1:0] node14506;
	wire [4-1:0] node14509;
	wire [4-1:0] node14510;
	wire [4-1:0] node14511;
	wire [4-1:0] node14512;
	wire [4-1:0] node14515;
	wire [4-1:0] node14519;
	wire [4-1:0] node14520;
	wire [4-1:0] node14521;
	wire [4-1:0] node14524;
	wire [4-1:0] node14528;
	wire [4-1:0] node14529;
	wire [4-1:0] node14530;
	wire [4-1:0] node14531;
	wire [4-1:0] node14532;
	wire [4-1:0] node14533;
	wire [4-1:0] node14537;
	wire [4-1:0] node14538;
	wire [4-1:0] node14542;
	wire [4-1:0] node14543;
	wire [4-1:0] node14544;
	wire [4-1:0] node14547;
	wire [4-1:0] node14551;
	wire [4-1:0] node14552;
	wire [4-1:0] node14553;
	wire [4-1:0] node14556;
	wire [4-1:0] node14559;
	wire [4-1:0] node14560;
	wire [4-1:0] node14564;
	wire [4-1:0] node14565;
	wire [4-1:0] node14566;
	wire [4-1:0] node14567;
	wire [4-1:0] node14570;
	wire [4-1:0] node14573;
	wire [4-1:0] node14574;
	wire [4-1:0] node14578;
	wire [4-1:0] node14579;
	wire [4-1:0] node14583;
	wire [4-1:0] node14584;
	wire [4-1:0] node14585;
	wire [4-1:0] node14586;
	wire [4-1:0] node14587;
	wire [4-1:0] node14588;
	wire [4-1:0] node14589;
	wire [4-1:0] node14593;
	wire [4-1:0] node14595;
	wire [4-1:0] node14598;
	wire [4-1:0] node14599;
	wire [4-1:0] node14600;
	wire [4-1:0] node14604;
	wire [4-1:0] node14605;
	wire [4-1:0] node14609;
	wire [4-1:0] node14610;
	wire [4-1:0] node14611;
	wire [4-1:0] node14613;
	wire [4-1:0] node14617;
	wire [4-1:0] node14618;
	wire [4-1:0] node14621;
	wire [4-1:0] node14624;
	wire [4-1:0] node14625;
	wire [4-1:0] node14626;
	wire [4-1:0] node14627;
	wire [4-1:0] node14630;
	wire [4-1:0] node14633;
	wire [4-1:0] node14634;
	wire [4-1:0] node14637;
	wire [4-1:0] node14640;
	wire [4-1:0] node14641;
	wire [4-1:0] node14644;
	wire [4-1:0] node14647;
	wire [4-1:0] node14648;
	wire [4-1:0] node14649;
	wire [4-1:0] node14650;
	wire [4-1:0] node14653;
	wire [4-1:0] node14656;
	wire [4-1:0] node14657;
	wire [4-1:0] node14658;
	wire [4-1:0] node14661;
	wire [4-1:0] node14664;
	wire [4-1:0] node14666;
	wire [4-1:0] node14669;
	wire [4-1:0] node14670;
	wire [4-1:0] node14671;
	wire [4-1:0] node14674;
	wire [4-1:0] node14677;
	wire [4-1:0] node14679;
	wire [4-1:0] node14680;
	wire [4-1:0] node14683;
	wire [4-1:0] node14686;
	wire [4-1:0] node14687;
	wire [4-1:0] node14688;
	wire [4-1:0] node14689;
	wire [4-1:0] node14690;
	wire [4-1:0] node14691;
	wire [4-1:0] node14692;
	wire [4-1:0] node14693;
	wire [4-1:0] node14694;
	wire [4-1:0] node14695;
	wire [4-1:0] node14698;
	wire [4-1:0] node14701;
	wire [4-1:0] node14702;
	wire [4-1:0] node14705;
	wire [4-1:0] node14708;
	wire [4-1:0] node14709;
	wire [4-1:0] node14710;
	wire [4-1:0] node14714;
	wire [4-1:0] node14717;
	wire [4-1:0] node14718;
	wire [4-1:0] node14719;
	wire [4-1:0] node14720;
	wire [4-1:0] node14722;
	wire [4-1:0] node14725;
	wire [4-1:0] node14728;
	wire [4-1:0] node14729;
	wire [4-1:0] node14732;
	wire [4-1:0] node14735;
	wire [4-1:0] node14736;
	wire [4-1:0] node14737;
	wire [4-1:0] node14741;
	wire [4-1:0] node14744;
	wire [4-1:0] node14745;
	wire [4-1:0] node14746;
	wire [4-1:0] node14747;
	wire [4-1:0] node14748;
	wire [4-1:0] node14751;
	wire [4-1:0] node14754;
	wire [4-1:0] node14757;
	wire [4-1:0] node14758;
	wire [4-1:0] node14759;
	wire [4-1:0] node14762;
	wire [4-1:0] node14765;
	wire [4-1:0] node14766;
	wire [4-1:0] node14769;
	wire [4-1:0] node14772;
	wire [4-1:0] node14773;
	wire [4-1:0] node14774;
	wire [4-1:0] node14776;
	wire [4-1:0] node14777;
	wire [4-1:0] node14780;
	wire [4-1:0] node14783;
	wire [4-1:0] node14784;
	wire [4-1:0] node14787;
	wire [4-1:0] node14790;
	wire [4-1:0] node14791;
	wire [4-1:0] node14792;
	wire [4-1:0] node14793;
	wire [4-1:0] node14797;
	wire [4-1:0] node14800;
	wire [4-1:0] node14801;
	wire [4-1:0] node14805;
	wire [4-1:0] node14806;
	wire [4-1:0] node14807;
	wire [4-1:0] node14808;
	wire [4-1:0] node14809;
	wire [4-1:0] node14810;
	wire [4-1:0] node14811;
	wire [4-1:0] node14815;
	wire [4-1:0] node14816;
	wire [4-1:0] node14821;
	wire [4-1:0] node14822;
	wire [4-1:0] node14823;
	wire [4-1:0] node14824;
	wire [4-1:0] node14828;
	wire [4-1:0] node14829;
	wire [4-1:0] node14833;
	wire [4-1:0] node14836;
	wire [4-1:0] node14837;
	wire [4-1:0] node14838;
	wire [4-1:0] node14841;
	wire [4-1:0] node14844;
	wire [4-1:0] node14845;
	wire [4-1:0] node14846;
	wire [4-1:0] node14849;
	wire [4-1:0] node14852;
	wire [4-1:0] node14853;
	wire [4-1:0] node14857;
	wire [4-1:0] node14858;
	wire [4-1:0] node14859;
	wire [4-1:0] node14860;
	wire [4-1:0] node14861;
	wire [4-1:0] node14864;
	wire [4-1:0] node14868;
	wire [4-1:0] node14869;
	wire [4-1:0] node14870;
	wire [4-1:0] node14872;
	wire [4-1:0] node14875;
	wire [4-1:0] node14878;
	wire [4-1:0] node14881;
	wire [4-1:0] node14882;
	wire [4-1:0] node14883;
	wire [4-1:0] node14884;
	wire [4-1:0] node14887;
	wire [4-1:0] node14890;
	wire [4-1:0] node14891;
	wire [4-1:0] node14893;
	wire [4-1:0] node14897;
	wire [4-1:0] node14898;
	wire [4-1:0] node14900;
	wire [4-1:0] node14903;
	wire [4-1:0] node14904;
	wire [4-1:0] node14907;
	wire [4-1:0] node14909;
	wire [4-1:0] node14912;
	wire [4-1:0] node14913;
	wire [4-1:0] node14914;
	wire [4-1:0] node14915;
	wire [4-1:0] node14916;
	wire [4-1:0] node14917;
	wire [4-1:0] node14918;
	wire [4-1:0] node14919;
	wire [4-1:0] node14922;
	wire [4-1:0] node14925;
	wire [4-1:0] node14926;
	wire [4-1:0] node14929;
	wire [4-1:0] node14932;
	wire [4-1:0] node14934;
	wire [4-1:0] node14935;
	wire [4-1:0] node14938;
	wire [4-1:0] node14941;
	wire [4-1:0] node14942;
	wire [4-1:0] node14945;
	wire [4-1:0] node14948;
	wire [4-1:0] node14949;
	wire [4-1:0] node14950;
	wire [4-1:0] node14951;
	wire [4-1:0] node14954;
	wire [4-1:0] node14957;
	wire [4-1:0] node14958;
	wire [4-1:0] node14961;
	wire [4-1:0] node14964;
	wire [4-1:0] node14965;
	wire [4-1:0] node14966;
	wire [4-1:0] node14967;
	wire [4-1:0] node14970;
	wire [4-1:0] node14974;
	wire [4-1:0] node14975;
	wire [4-1:0] node14976;
	wire [4-1:0] node14979;
	wire [4-1:0] node14982;
	wire [4-1:0] node14983;
	wire [4-1:0] node14986;
	wire [4-1:0] node14989;
	wire [4-1:0] node14990;
	wire [4-1:0] node14991;
	wire [4-1:0] node14992;
	wire [4-1:0] node14993;
	wire [4-1:0] node14994;
	wire [4-1:0] node14998;
	wire [4-1:0] node15000;
	wire [4-1:0] node15003;
	wire [4-1:0] node15004;
	wire [4-1:0] node15005;
	wire [4-1:0] node15008;
	wire [4-1:0] node15011;
	wire [4-1:0] node15012;
	wire [4-1:0] node15015;
	wire [4-1:0] node15018;
	wire [4-1:0] node15019;
	wire [4-1:0] node15020;
	wire [4-1:0] node15023;
	wire [4-1:0] node15026;
	wire [4-1:0] node15027;
	wire [4-1:0] node15030;
	wire [4-1:0] node15033;
	wire [4-1:0] node15034;
	wire [4-1:0] node15035;
	wire [4-1:0] node15036;
	wire [4-1:0] node15038;
	wire [4-1:0] node15041;
	wire [4-1:0] node15044;
	wire [4-1:0] node15045;
	wire [4-1:0] node15047;
	wire [4-1:0] node15050;
	wire [4-1:0] node15052;
	wire [4-1:0] node15055;
	wire [4-1:0] node15056;
	wire [4-1:0] node15057;
	wire [4-1:0] node15060;
	wire [4-1:0] node15063;
	wire [4-1:0] node15064;
	wire [4-1:0] node15065;
	wire [4-1:0] node15070;
	wire [4-1:0] node15071;
	wire [4-1:0] node15072;
	wire [4-1:0] node15073;
	wire [4-1:0] node15074;
	wire [4-1:0] node15076;
	wire [4-1:0] node15077;
	wire [4-1:0] node15080;
	wire [4-1:0] node15083;
	wire [4-1:0] node15085;
	wire [4-1:0] node15088;
	wire [4-1:0] node15089;
	wire [4-1:0] node15090;
	wire [4-1:0] node15091;
	wire [4-1:0] node15094;
	wire [4-1:0] node15098;
	wire [4-1:0] node15099;
	wire [4-1:0] node15101;
	wire [4-1:0] node15105;
	wire [4-1:0] node15106;
	wire [4-1:0] node15107;
	wire [4-1:0] node15108;
	wire [4-1:0] node15110;
	wire [4-1:0] node15114;
	wire [4-1:0] node15115;
	wire [4-1:0] node15116;
	wire [4-1:0] node15120;
	wire [4-1:0] node15121;
	wire [4-1:0] node15124;
	wire [4-1:0] node15127;
	wire [4-1:0] node15128;
	wire [4-1:0] node15129;
	wire [4-1:0] node15132;
	wire [4-1:0] node15135;
	wire [4-1:0] node15136;
	wire [4-1:0] node15140;
	wire [4-1:0] node15141;
	wire [4-1:0] node15142;
	wire [4-1:0] node15143;
	wire [4-1:0] node15144;
	wire [4-1:0] node15148;
	wire [4-1:0] node15149;
	wire [4-1:0] node15153;
	wire [4-1:0] node15154;
	wire [4-1:0] node15155;
	wire [4-1:0] node15159;
	wire [4-1:0] node15160;
	wire [4-1:0] node15164;
	wire [4-1:0] node15165;
	wire [4-1:0] node15166;
	wire [4-1:0] node15167;
	wire [4-1:0] node15168;
	wire [4-1:0] node15172;
	wire [4-1:0] node15173;
	wire [4-1:0] node15176;
	wire [4-1:0] node15179;
	wire [4-1:0] node15180;
	wire [4-1:0] node15181;
	wire [4-1:0] node15185;
	wire [4-1:0] node15187;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15192;
	wire [4-1:0] node15193;
	wire [4-1:0] node15196;
	wire [4-1:0] node15200;
	wire [4-1:0] node15201;
	wire [4-1:0] node15203;
	wire [4-1:0] node15206;
	wire [4-1:0] node15207;
	wire [4-1:0] node15211;
	wire [4-1:0] node15212;
	wire [4-1:0] node15213;
	wire [4-1:0] node15214;
	wire [4-1:0] node15215;
	wire [4-1:0] node15216;
	wire [4-1:0] node15217;
	wire [4-1:0] node15218;
	wire [4-1:0] node15222;
	wire [4-1:0] node15224;
	wire [4-1:0] node15227;
	wire [4-1:0] node15228;
	wire [4-1:0] node15229;
	wire [4-1:0] node15232;
	wire [4-1:0] node15235;
	wire [4-1:0] node15236;
	wire [4-1:0] node15240;
	wire [4-1:0] node15241;
	wire [4-1:0] node15242;
	wire [4-1:0] node15245;
	wire [4-1:0] node15246;
	wire [4-1:0] node15250;
	wire [4-1:0] node15251;
	wire [4-1:0] node15255;
	wire [4-1:0] node15256;
	wire [4-1:0] node15257;
	wire [4-1:0] node15258;
	wire [4-1:0] node15259;
	wire [4-1:0] node15263;
	wire [4-1:0] node15265;
	wire [4-1:0] node15268;
	wire [4-1:0] node15269;
	wire [4-1:0] node15271;
	wire [4-1:0] node15274;
	wire [4-1:0] node15277;
	wire [4-1:0] node15278;
	wire [4-1:0] node15279;
	wire [4-1:0] node15281;
	wire [4-1:0] node15284;
	wire [4-1:0] node15285;
	wire [4-1:0] node15289;
	wire [4-1:0] node15290;
	wire [4-1:0] node15291;
	wire [4-1:0] node15293;
	wire [4-1:0] node15297;
	wire [4-1:0] node15299;
	wire [4-1:0] node15302;
	wire [4-1:0] node15303;
	wire [4-1:0] node15304;
	wire [4-1:0] node15305;
	wire [4-1:0] node15306;
	wire [4-1:0] node15308;
	wire [4-1:0] node15310;
	wire [4-1:0] node15313;
	wire [4-1:0] node15314;
	wire [4-1:0] node15317;
	wire [4-1:0] node15320;
	wire [4-1:0] node15321;
	wire [4-1:0] node15322;
	wire [4-1:0] node15325;
	wire [4-1:0] node15328;
	wire [4-1:0] node15329;
	wire [4-1:0] node15332;
	wire [4-1:0] node15335;
	wire [4-1:0] node15336;
	wire [4-1:0] node15337;
	wire [4-1:0] node15338;
	wire [4-1:0] node15342;
	wire [4-1:0] node15344;
	wire [4-1:0] node15347;
	wire [4-1:0] node15348;
	wire [4-1:0] node15349;
	wire [4-1:0] node15350;
	wire [4-1:0] node15353;
	wire [4-1:0] node15357;
	wire [4-1:0] node15358;
	wire [4-1:0] node15361;
	wire [4-1:0] node15364;
	wire [4-1:0] node15365;
	wire [4-1:0] node15366;
	wire [4-1:0] node15367;
	wire [4-1:0] node15370;
	wire [4-1:0] node15371;
	wire [4-1:0] node15374;
	wire [4-1:0] node15377;
	wire [4-1:0] node15378;
	wire [4-1:0] node15381;
	wire [4-1:0] node15384;
	wire [4-1:0] node15385;
	wire [4-1:0] node15386;
	wire [4-1:0] node15387;
	wire [4-1:0] node15388;
	wire [4-1:0] node15392;
	wire [4-1:0] node15393;
	wire [4-1:0] node15396;
	wire [4-1:0] node15399;
	wire [4-1:0] node15401;
	wire [4-1:0] node15404;
	wire [4-1:0] node15405;
	wire [4-1:0] node15406;
	wire [4-1:0] node15409;
	wire [4-1:0] node15412;
	wire [4-1:0] node15413;
	wire [4-1:0] node15416;
	wire [4-1:0] node15419;
	wire [4-1:0] node15420;
	wire [4-1:0] node15421;
	wire [4-1:0] node15422;
	wire [4-1:0] node15423;
	wire [4-1:0] node15424;
	wire [4-1:0] node15425;
	wire [4-1:0] node15427;
	wire [4-1:0] node15431;
	wire [4-1:0] node15432;
	wire [4-1:0] node15435;
	wire [4-1:0] node15438;
	wire [4-1:0] node15439;
	wire [4-1:0] node15440;
	wire [4-1:0] node15443;
	wire [4-1:0] node15446;
	wire [4-1:0] node15447;
	wire [4-1:0] node15450;
	wire [4-1:0] node15453;
	wire [4-1:0] node15454;
	wire [4-1:0] node15455;
	wire [4-1:0] node15457;
	wire [4-1:0] node15460;
	wire [4-1:0] node15461;
	wire [4-1:0] node15464;
	wire [4-1:0] node15467;
	wire [4-1:0] node15468;
	wire [4-1:0] node15471;
	wire [4-1:0] node15472;
	wire [4-1:0] node15476;
	wire [4-1:0] node15477;
	wire [4-1:0] node15478;
	wire [4-1:0] node15479;
	wire [4-1:0] node15480;
	wire [4-1:0] node15484;
	wire [4-1:0] node15485;
	wire [4-1:0] node15488;
	wire [4-1:0] node15491;
	wire [4-1:0] node15492;
	wire [4-1:0] node15495;
	wire [4-1:0] node15498;
	wire [4-1:0] node15499;
	wire [4-1:0] node15500;
	wire [4-1:0] node15501;
	wire [4-1:0] node15504;
	wire [4-1:0] node15506;
	wire [4-1:0] node15509;
	wire [4-1:0] node15510;
	wire [4-1:0] node15511;
	wire [4-1:0] node15515;
	wire [4-1:0] node15517;
	wire [4-1:0] node15520;
	wire [4-1:0] node15521;
	wire [4-1:0] node15524;
	wire [4-1:0] node15525;
	wire [4-1:0] node15529;
	wire [4-1:0] node15530;
	wire [4-1:0] node15531;
	wire [4-1:0] node15532;
	wire [4-1:0] node15533;
	wire [4-1:0] node15534;
	wire [4-1:0] node15538;
	wire [4-1:0] node15540;
	wire [4-1:0] node15543;
	wire [4-1:0] node15545;
	wire [4-1:0] node15546;
	wire [4-1:0] node15550;
	wire [4-1:0] node15551;
	wire [4-1:0] node15552;
	wire [4-1:0] node15554;
	wire [4-1:0] node15557;
	wire [4-1:0] node15558;
	wire [4-1:0] node15562;
	wire [4-1:0] node15563;
	wire [4-1:0] node15565;
	wire [4-1:0] node15568;
	wire [4-1:0] node15569;
	wire [4-1:0] node15573;
	wire [4-1:0] node15574;
	wire [4-1:0] node15575;
	wire [4-1:0] node15576;
	wire [4-1:0] node15577;
	wire [4-1:0] node15581;
	wire [4-1:0] node15582;
	wire [4-1:0] node15586;
	wire [4-1:0] node15587;
	wire [4-1:0] node15588;
	wire [4-1:0] node15592;
	wire [4-1:0] node15594;
	wire [4-1:0] node15597;
	wire [4-1:0] node15598;
	wire [4-1:0] node15599;
	wire [4-1:0] node15601;
	wire [4-1:0] node15604;
	wire [4-1:0] node15606;
	wire [4-1:0] node15609;
	wire [4-1:0] node15610;
	wire [4-1:0] node15612;
	wire [4-1:0] node15615;
	wire [4-1:0] node15617;
	wire [4-1:0] node15620;
	wire [4-1:0] node15621;
	wire [4-1:0] node15622;
	wire [4-1:0] node15623;
	wire [4-1:0] node15624;
	wire [4-1:0] node15625;
	wire [4-1:0] node15626;
	wire [4-1:0] node15627;
	wire [4-1:0] node15630;
	wire [4-1:0] node15633;
	wire [4-1:0] node15634;
	wire [4-1:0] node15635;
	wire [4-1:0] node15636;
	wire [4-1:0] node15639;
	wire [4-1:0] node15643;
	wire [4-1:0] node15644;
	wire [4-1:0] node15648;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15653;
	wire [4-1:0] node15656;
	wire [4-1:0] node15657;
	wire [4-1:0] node15660;
	wire [4-1:0] node15663;
	wire [4-1:0] node15664;
	wire [4-1:0] node15665;
	wire [4-1:0] node15666;
	wire [4-1:0] node15667;
	wire [4-1:0] node15670;
	wire [4-1:0] node15673;
	wire [4-1:0] node15674;
	wire [4-1:0] node15675;
	wire [4-1:0] node15678;
	wire [4-1:0] node15681;
	wire [4-1:0] node15682;
	wire [4-1:0] node15685;
	wire [4-1:0] node15688;
	wire [4-1:0] node15689;
	wire [4-1:0] node15690;
	wire [4-1:0] node15691;
	wire [4-1:0] node15694;
	wire [4-1:0] node15697;
	wire [4-1:0] node15698;
	wire [4-1:0] node15702;
	wire [4-1:0] node15703;
	wire [4-1:0] node15705;
	wire [4-1:0] node15708;
	wire [4-1:0] node15709;
	wire [4-1:0] node15712;
	wire [4-1:0] node15715;
	wire [4-1:0] node15716;
	wire [4-1:0] node15717;
	wire [4-1:0] node15718;
	wire [4-1:0] node15719;
	wire [4-1:0] node15722;
	wire [4-1:0] node15725;
	wire [4-1:0] node15726;
	wire [4-1:0] node15729;
	wire [4-1:0] node15732;
	wire [4-1:0] node15733;
	wire [4-1:0] node15736;
	wire [4-1:0] node15739;
	wire [4-1:0] node15740;
	wire [4-1:0] node15741;
	wire [4-1:0] node15742;
	wire [4-1:0] node15745;
	wire [4-1:0] node15748;
	wire [4-1:0] node15749;
	wire [4-1:0] node15752;
	wire [4-1:0] node15755;
	wire [4-1:0] node15756;
	wire [4-1:0] node15759;
	wire [4-1:0] node15762;
	wire [4-1:0] node15763;
	wire [4-1:0] node15764;
	wire [4-1:0] node15765;
	wire [4-1:0] node15767;
	wire [4-1:0] node15768;
	wire [4-1:0] node15771;
	wire [4-1:0] node15774;
	wire [4-1:0] node15775;
	wire [4-1:0] node15776;
	wire [4-1:0] node15777;
	wire [4-1:0] node15781;
	wire [4-1:0] node15782;
	wire [4-1:0] node15786;
	wire [4-1:0] node15787;
	wire [4-1:0] node15790;
	wire [4-1:0] node15792;
	wire [4-1:0] node15795;
	wire [4-1:0] node15796;
	wire [4-1:0] node15797;
	wire [4-1:0] node15798;
	wire [4-1:0] node15802;
	wire [4-1:0] node15803;
	wire [4-1:0] node15807;
	wire [4-1:0] node15808;
	wire [4-1:0] node15810;
	wire [4-1:0] node15813;
	wire [4-1:0] node15816;
	wire [4-1:0] node15817;
	wire [4-1:0] node15818;
	wire [4-1:0] node15819;
	wire [4-1:0] node15822;
	wire [4-1:0] node15825;
	wire [4-1:0] node15826;
	wire [4-1:0] node15827;
	wire [4-1:0] node15828;
	wire [4-1:0] node15831;
	wire [4-1:0] node15834;
	wire [4-1:0] node15835;
	wire [4-1:0] node15838;
	wire [4-1:0] node15841;
	wire [4-1:0] node15842;
	wire [4-1:0] node15845;
	wire [4-1:0] node15848;
	wire [4-1:0] node15849;
	wire [4-1:0] node15850;
	wire [4-1:0] node15851;
	wire [4-1:0] node15855;
	wire [4-1:0] node15856;
	wire [4-1:0] node15857;
	wire [4-1:0] node15860;
	wire [4-1:0] node15863;
	wire [4-1:0] node15864;
	wire [4-1:0] node15867;
	wire [4-1:0] node15870;
	wire [4-1:0] node15871;
	wire [4-1:0] node15872;
	wire [4-1:0] node15875;
	wire [4-1:0] node15878;
	wire [4-1:0] node15879;
	wire [4-1:0] node15880;
	wire [4-1:0] node15884;
	wire [4-1:0] node15885;
	wire [4-1:0] node15888;
	wire [4-1:0] node15891;
	wire [4-1:0] node15892;
	wire [4-1:0] node15893;
	wire [4-1:0] node15894;
	wire [4-1:0] node15895;
	wire [4-1:0] node15897;
	wire [4-1:0] node15899;
	wire [4-1:0] node15902;
	wire [4-1:0] node15904;
	wire [4-1:0] node15905;
	wire [4-1:0] node15908;
	wire [4-1:0] node15911;
	wire [4-1:0] node15912;
	wire [4-1:0] node15914;
	wire [4-1:0] node15915;
	wire [4-1:0] node15918;
	wire [4-1:0] node15921;
	wire [4-1:0] node15923;
	wire [4-1:0] node15924;
	wire [4-1:0] node15928;
	wire [4-1:0] node15929;
	wire [4-1:0] node15930;
	wire [4-1:0] node15932;
	wire [4-1:0] node15933;
	wire [4-1:0] node15934;
	wire [4-1:0] node15938;
	wire [4-1:0] node15939;
	wire [4-1:0] node15942;
	wire [4-1:0] node15945;
	wire [4-1:0] node15946;
	wire [4-1:0] node15947;
	wire [4-1:0] node15950;
	wire [4-1:0] node15953;
	wire [4-1:0] node15954;
	wire [4-1:0] node15957;
	wire [4-1:0] node15960;
	wire [4-1:0] node15961;
	wire [4-1:0] node15962;
	wire [4-1:0] node15965;
	wire [4-1:0] node15968;
	wire [4-1:0] node15969;
	wire [4-1:0] node15970;
	wire [4-1:0] node15972;
	wire [4-1:0] node15976;
	wire [4-1:0] node15977;
	wire [4-1:0] node15981;
	wire [4-1:0] node15982;
	wire [4-1:0] node15983;
	wire [4-1:0] node15984;
	wire [4-1:0] node15985;
	wire [4-1:0] node15987;
	wire [4-1:0] node15988;
	wire [4-1:0] node15991;
	wire [4-1:0] node15994;
	wire [4-1:0] node15995;
	wire [4-1:0] node15996;
	wire [4-1:0] node16000;
	wire [4-1:0] node16002;
	wire [4-1:0] node16005;
	wire [4-1:0] node16006;
	wire [4-1:0] node16007;
	wire [4-1:0] node16010;
	wire [4-1:0] node16013;
	wire [4-1:0] node16014;
	wire [4-1:0] node16015;
	wire [4-1:0] node16018;
	wire [4-1:0] node16022;
	wire [4-1:0] node16023;
	wire [4-1:0] node16024;
	wire [4-1:0] node16025;
	wire [4-1:0] node16029;
	wire [4-1:0] node16030;
	wire [4-1:0] node16034;
	wire [4-1:0] node16035;
	wire [4-1:0] node16036;
	wire [4-1:0] node16039;
	wire [4-1:0] node16043;
	wire [4-1:0] node16044;
	wire [4-1:0] node16045;
	wire [4-1:0] node16046;
	wire [4-1:0] node16047;
	wire [4-1:0] node16051;
	wire [4-1:0] node16052;
	wire [4-1:0] node16054;
	wire [4-1:0] node16057;
	wire [4-1:0] node16059;
	wire [4-1:0] node16062;
	wire [4-1:0] node16063;
	wire [4-1:0] node16065;
	wire [4-1:0] node16066;
	wire [4-1:0] node16069;
	wire [4-1:0] node16073;
	wire [4-1:0] node16074;
	wire [4-1:0] node16075;
	wire [4-1:0] node16076;
	wire [4-1:0] node16078;
	wire [4-1:0] node16082;
	wire [4-1:0] node16083;
	wire [4-1:0] node16084;
	wire [4-1:0] node16089;
	wire [4-1:0] node16090;
	wire [4-1:0] node16091;
	wire [4-1:0] node16095;
	wire [4-1:0] node16096;
	wire [4-1:0] node16097;
	wire [4-1:0] node16100;
	wire [4-1:0] node16104;
	wire [4-1:0] node16105;
	wire [4-1:0] node16106;
	wire [4-1:0] node16107;
	wire [4-1:0] node16108;
	wire [4-1:0] node16109;
	wire [4-1:0] node16110;
	wire [4-1:0] node16111;
	wire [4-1:0] node16114;
	wire [4-1:0] node16117;
	wire [4-1:0] node16118;
	wire [4-1:0] node16120;
	wire [4-1:0] node16123;
	wire [4-1:0] node16124;
	wire [4-1:0] node16127;
	wire [4-1:0] node16130;
	wire [4-1:0] node16131;
	wire [4-1:0] node16133;
	wire [4-1:0] node16136;
	wire [4-1:0] node16137;
	wire [4-1:0] node16140;
	wire [4-1:0] node16143;
	wire [4-1:0] node16144;
	wire [4-1:0] node16145;
	wire [4-1:0] node16147;
	wire [4-1:0] node16149;
	wire [4-1:0] node16153;
	wire [4-1:0] node16154;
	wire [4-1:0] node16155;
	wire [4-1:0] node16159;
	wire [4-1:0] node16160;
	wire [4-1:0] node16164;
	wire [4-1:0] node16165;
	wire [4-1:0] node16166;
	wire [4-1:0] node16167;
	wire [4-1:0] node16168;
	wire [4-1:0] node16171;
	wire [4-1:0] node16174;
	wire [4-1:0] node16175;
	wire [4-1:0] node16176;
	wire [4-1:0] node16180;
	wire [4-1:0] node16182;
	wire [4-1:0] node16185;
	wire [4-1:0] node16186;
	wire [4-1:0] node16188;
	wire [4-1:0] node16191;
	wire [4-1:0] node16192;
	wire [4-1:0] node16195;
	wire [4-1:0] node16198;
	wire [4-1:0] node16199;
	wire [4-1:0] node16200;
	wire [4-1:0] node16202;
	wire [4-1:0] node16205;
	wire [4-1:0] node16208;
	wire [4-1:0] node16211;
	wire [4-1:0] node16212;
	wire [4-1:0] node16213;
	wire [4-1:0] node16214;
	wire [4-1:0] node16215;
	wire [4-1:0] node16217;
	wire [4-1:0] node16220;
	wire [4-1:0] node16221;
	wire [4-1:0] node16225;
	wire [4-1:0] node16226;
	wire [4-1:0] node16229;
	wire [4-1:0] node16230;
	wire [4-1:0] node16234;
	wire [4-1:0] node16235;
	wire [4-1:0] node16236;
	wire [4-1:0] node16237;
	wire [4-1:0] node16242;
	wire [4-1:0] node16243;
	wire [4-1:0] node16244;
	wire [4-1:0] node16248;
	wire [4-1:0] node16249;
	wire [4-1:0] node16253;
	wire [4-1:0] node16254;
	wire [4-1:0] node16255;
	wire [4-1:0] node16258;
	wire [4-1:0] node16259;
	wire [4-1:0] node16260;
	wire [4-1:0] node16264;
	wire [4-1:0] node16265;
	wire [4-1:0] node16269;
	wire [4-1:0] node16270;
	wire [4-1:0] node16271;
	wire [4-1:0] node16272;
	wire [4-1:0] node16273;
	wire [4-1:0] node16276;
	wire [4-1:0] node16279;
	wire [4-1:0] node16281;
	wire [4-1:0] node16285;
	wire [4-1:0] node16286;
	wire [4-1:0] node16287;
	wire [4-1:0] node16291;
	wire [4-1:0] node16292;
	wire [4-1:0] node16296;
	wire [4-1:0] node16297;
	wire [4-1:0] node16298;
	wire [4-1:0] node16299;
	wire [4-1:0] node16300;
	wire [4-1:0] node16301;
	wire [4-1:0] node16303;
	wire [4-1:0] node16304;
	wire [4-1:0] node16307;
	wire [4-1:0] node16310;
	wire [4-1:0] node16311;
	wire [4-1:0] node16312;
	wire [4-1:0] node16317;
	wire [4-1:0] node16318;
	wire [4-1:0] node16320;
	wire [4-1:0] node16321;
	wire [4-1:0] node16325;
	wire [4-1:0] node16326;
	wire [4-1:0] node16330;
	wire [4-1:0] node16331;
	wire [4-1:0] node16332;
	wire [4-1:0] node16334;
	wire [4-1:0] node16335;
	wire [4-1:0] node16339;
	wire [4-1:0] node16340;
	wire [4-1:0] node16343;
	wire [4-1:0] node16345;
	wire [4-1:0] node16348;
	wire [4-1:0] node16349;
	wire [4-1:0] node16350;
	wire [4-1:0] node16351;
	wire [4-1:0] node16355;
	wire [4-1:0] node16357;
	wire [4-1:0] node16360;
	wire [4-1:0] node16361;
	wire [4-1:0] node16363;
	wire [4-1:0] node16366;
	wire [4-1:0] node16369;
	wire [4-1:0] node16370;
	wire [4-1:0] node16371;
	wire [4-1:0] node16372;
	wire [4-1:0] node16375;
	wire [4-1:0] node16376;
	wire [4-1:0] node16379;
	wire [4-1:0] node16380;
	wire [4-1:0] node16384;
	wire [4-1:0] node16385;
	wire [4-1:0] node16386;
	wire [4-1:0] node16388;
	wire [4-1:0] node16392;
	wire [4-1:0] node16393;
	wire [4-1:0] node16394;
	wire [4-1:0] node16398;
	wire [4-1:0] node16400;
	wire [4-1:0] node16403;
	wire [4-1:0] node16404;
	wire [4-1:0] node16405;
	wire [4-1:0] node16406;
	wire [4-1:0] node16408;
	wire [4-1:0] node16412;
	wire [4-1:0] node16415;
	wire [4-1:0] node16416;
	wire [4-1:0] node16417;
	wire [4-1:0] node16419;
	wire [4-1:0] node16422;
	wire [4-1:0] node16423;
	wire [4-1:0] node16427;
	wire [4-1:0] node16430;
	wire [4-1:0] node16431;
	wire [4-1:0] node16432;
	wire [4-1:0] node16433;
	wire [4-1:0] node16434;
	wire [4-1:0] node16437;
	wire [4-1:0] node16440;
	wire [4-1:0] node16441;
	wire [4-1:0] node16442;
	wire [4-1:0] node16445;
	wire [4-1:0] node16448;
	wire [4-1:0] node16450;
	wire [4-1:0] node16451;
	wire [4-1:0] node16454;
	wire [4-1:0] node16457;
	wire [4-1:0] node16458;
	wire [4-1:0] node16459;
	wire [4-1:0] node16461;
	wire [4-1:0] node16462;
	wire [4-1:0] node16466;
	wire [4-1:0] node16467;
	wire [4-1:0] node16469;
	wire [4-1:0] node16472;
	wire [4-1:0] node16474;
	wire [4-1:0] node16477;
	wire [4-1:0] node16478;
	wire [4-1:0] node16479;
	wire [4-1:0] node16481;
	wire [4-1:0] node16484;
	wire [4-1:0] node16485;
	wire [4-1:0] node16489;
	wire [4-1:0] node16490;
	wire [4-1:0] node16491;
	wire [4-1:0] node16495;
	wire [4-1:0] node16496;
	wire [4-1:0] node16500;
	wire [4-1:0] node16501;
	wire [4-1:0] node16502;
	wire [4-1:0] node16503;
	wire [4-1:0] node16505;
	wire [4-1:0] node16506;
	wire [4-1:0] node16509;
	wire [4-1:0] node16513;
	wire [4-1:0] node16514;
	wire [4-1:0] node16515;
	wire [4-1:0] node16516;
	wire [4-1:0] node16519;
	wire [4-1:0] node16522;
	wire [4-1:0] node16523;
	wire [4-1:0] node16527;
	wire [4-1:0] node16529;
	wire [4-1:0] node16530;
	wire [4-1:0] node16534;
	wire [4-1:0] node16535;
	wire [4-1:0] node16536;
	wire [4-1:0] node16538;
	wire [4-1:0] node16541;
	wire [4-1:0] node16542;
	wire [4-1:0] node16546;
	wire [4-1:0] node16547;
	wire [4-1:0] node16549;
	wire [4-1:0] node16550;
	wire [4-1:0] node16554;
	wire [4-1:0] node16555;
	wire [4-1:0] node16558;
	wire [4-1:0] node16561;
	wire [4-1:0] node16562;
	wire [4-1:0] node16563;
	wire [4-1:0] node16564;
	wire [4-1:0] node16565;
	wire [4-1:0] node16566;
	wire [4-1:0] node16567;
	wire [4-1:0] node16568;
	wire [4-1:0] node16569;
	wire [4-1:0] node16570;
	wire [4-1:0] node16571;
	wire [4-1:0] node16574;
	wire [4-1:0] node16575;
	wire [4-1:0] node16577;
	wire [4-1:0] node16580;
	wire [4-1:0] node16583;
	wire [4-1:0] node16584;
	wire [4-1:0] node16585;
	wire [4-1:0] node16588;
	wire [4-1:0] node16591;
	wire [4-1:0] node16592;
	wire [4-1:0] node16595;
	wire [4-1:0] node16597;
	wire [4-1:0] node16600;
	wire [4-1:0] node16601;
	wire [4-1:0] node16602;
	wire [4-1:0] node16605;
	wire [4-1:0] node16606;
	wire [4-1:0] node16608;
	wire [4-1:0] node16611;
	wire [4-1:0] node16612;
	wire [4-1:0] node16616;
	wire [4-1:0] node16617;
	wire [4-1:0] node16618;
	wire [4-1:0] node16619;
	wire [4-1:0] node16622;
	wire [4-1:0] node16625;
	wire [4-1:0] node16626;
	wire [4-1:0] node16629;
	wire [4-1:0] node16632;
	wire [4-1:0] node16633;
	wire [4-1:0] node16634;
	wire [4-1:0] node16637;
	wire [4-1:0] node16640;
	wire [4-1:0] node16641;
	wire [4-1:0] node16644;
	wire [4-1:0] node16647;
	wire [4-1:0] node16648;
	wire [4-1:0] node16649;
	wire [4-1:0] node16650;
	wire [4-1:0] node16651;
	wire [4-1:0] node16654;
	wire [4-1:0] node16656;
	wire [4-1:0] node16659;
	wire [4-1:0] node16660;
	wire [4-1:0] node16663;
	wire [4-1:0] node16664;
	wire [4-1:0] node16667;
	wire [4-1:0] node16670;
	wire [4-1:0] node16671;
	wire [4-1:0] node16672;
	wire [4-1:0] node16675;
	wire [4-1:0] node16676;
	wire [4-1:0] node16680;
	wire [4-1:0] node16681;
	wire [4-1:0] node16682;
	wire [4-1:0] node16685;
	wire [4-1:0] node16688;
	wire [4-1:0] node16689;
	wire [4-1:0] node16692;
	wire [4-1:0] node16695;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16698;
	wire [4-1:0] node16699;
	wire [4-1:0] node16701;
	wire [4-1:0] node16704;
	wire [4-1:0] node16706;
	wire [4-1:0] node16710;
	wire [4-1:0] node16711;
	wire [4-1:0] node16714;
	wire [4-1:0] node16716;
	wire [4-1:0] node16719;
	wire [4-1:0] node16720;
	wire [4-1:0] node16721;
	wire [4-1:0] node16724;
	wire [4-1:0] node16727;
	wire [4-1:0] node16728;
	wire [4-1:0] node16729;
	wire [4-1:0] node16732;
	wire [4-1:0] node16735;
	wire [4-1:0] node16736;
	wire [4-1:0] node16739;
	wire [4-1:0] node16742;
	wire [4-1:0] node16743;
	wire [4-1:0] node16744;
	wire [4-1:0] node16745;
	wire [4-1:0] node16746;
	wire [4-1:0] node16749;
	wire [4-1:0] node16751;
	wire [4-1:0] node16754;
	wire [4-1:0] node16755;
	wire [4-1:0] node16756;
	wire [4-1:0] node16759;
	wire [4-1:0] node16761;
	wire [4-1:0] node16764;
	wire [4-1:0] node16765;
	wire [4-1:0] node16767;
	wire [4-1:0] node16770;
	wire [4-1:0] node16771;
	wire [4-1:0] node16775;
	wire [4-1:0] node16776;
	wire [4-1:0] node16777;
	wire [4-1:0] node16780;
	wire [4-1:0] node16782;
	wire [4-1:0] node16785;
	wire [4-1:0] node16786;
	wire [4-1:0] node16787;
	wire [4-1:0] node16788;
	wire [4-1:0] node16791;
	wire [4-1:0] node16794;
	wire [4-1:0] node16795;
	wire [4-1:0] node16796;
	wire [4-1:0] node16799;
	wire [4-1:0] node16802;
	wire [4-1:0] node16803;
	wire [4-1:0] node16807;
	wire [4-1:0] node16808;
	wire [4-1:0] node16810;
	wire [4-1:0] node16811;
	wire [4-1:0] node16814;
	wire [4-1:0] node16817;
	wire [4-1:0] node16818;
	wire [4-1:0] node16819;
	wire [4-1:0] node16822;
	wire [4-1:0] node16825;
	wire [4-1:0] node16826;
	wire [4-1:0] node16829;
	wire [4-1:0] node16832;
	wire [4-1:0] node16833;
	wire [4-1:0] node16834;
	wire [4-1:0] node16835;
	wire [4-1:0] node16836;
	wire [4-1:0] node16839;
	wire [4-1:0] node16842;
	wire [4-1:0] node16843;
	wire [4-1:0] node16844;
	wire [4-1:0] node16847;
	wire [4-1:0] node16850;
	wire [4-1:0] node16851;
	wire [4-1:0] node16855;
	wire [4-1:0] node16856;
	wire [4-1:0] node16857;
	wire [4-1:0] node16860;
	wire [4-1:0] node16863;
	wire [4-1:0] node16864;
	wire [4-1:0] node16865;
	wire [4-1:0] node16868;
	wire [4-1:0] node16871;
	wire [4-1:0] node16872;
	wire [4-1:0] node16875;
	wire [4-1:0] node16878;
	wire [4-1:0] node16879;
	wire [4-1:0] node16880;
	wire [4-1:0] node16881;
	wire [4-1:0] node16884;
	wire [4-1:0] node16887;
	wire [4-1:0] node16888;
	wire [4-1:0] node16891;
	wire [4-1:0] node16893;
	wire [4-1:0] node16896;
	wire [4-1:0] node16897;
	wire [4-1:0] node16898;
	wire [4-1:0] node16901;
	wire [4-1:0] node16904;
	wire [4-1:0] node16905;
	wire [4-1:0] node16906;
	wire [4-1:0] node16907;
	wire [4-1:0] node16910;
	wire [4-1:0] node16913;
	wire [4-1:0] node16915;
	wire [4-1:0] node16918;
	wire [4-1:0] node16919;
	wire [4-1:0] node16920;
	wire [4-1:0] node16923;
	wire [4-1:0] node16926;
	wire [4-1:0] node16927;
	wire [4-1:0] node16931;
	wire [4-1:0] node16932;
	wire [4-1:0] node16933;
	wire [4-1:0] node16934;
	wire [4-1:0] node16935;
	wire [4-1:0] node16936;
	wire [4-1:0] node16939;
	wire [4-1:0] node16941;
	wire [4-1:0] node16944;
	wire [4-1:0] node16945;
	wire [4-1:0] node16948;
	wire [4-1:0] node16950;
	wire [4-1:0] node16953;
	wire [4-1:0] node16954;
	wire [4-1:0] node16955;
	wire [4-1:0] node16956;
	wire [4-1:0] node16958;
	wire [4-1:0] node16961;
	wire [4-1:0] node16963;
	wire [4-1:0] node16966;
	wire [4-1:0] node16967;
	wire [4-1:0] node16970;
	wire [4-1:0] node16971;
	wire [4-1:0] node16975;
	wire [4-1:0] node16976;
	wire [4-1:0] node16977;
	wire [4-1:0] node16979;
	wire [4-1:0] node16982;
	wire [4-1:0] node16985;
	wire [4-1:0] node16986;
	wire [4-1:0] node16987;
	wire [4-1:0] node16990;
	wire [4-1:0] node16993;
	wire [4-1:0] node16995;
	wire [4-1:0] node16998;
	wire [4-1:0] node16999;
	wire [4-1:0] node17000;
	wire [4-1:0] node17001;
	wire [4-1:0] node17002;
	wire [4-1:0] node17003;
	wire [4-1:0] node17006;
	wire [4-1:0] node17009;
	wire [4-1:0] node17011;
	wire [4-1:0] node17014;
	wire [4-1:0] node17015;
	wire [4-1:0] node17017;
	wire [4-1:0] node17020;
	wire [4-1:0] node17022;
	wire [4-1:0] node17025;
	wire [4-1:0] node17026;
	wire [4-1:0] node17027;
	wire [4-1:0] node17030;
	wire [4-1:0] node17031;
	wire [4-1:0] node17034;
	wire [4-1:0] node17037;
	wire [4-1:0] node17038;
	wire [4-1:0] node17039;
	wire [4-1:0] node17042;
	wire [4-1:0] node17045;
	wire [4-1:0] node17046;
	wire [4-1:0] node17049;
	wire [4-1:0] node17052;
	wire [4-1:0] node17053;
	wire [4-1:0] node17054;
	wire [4-1:0] node17055;
	wire [4-1:0] node17058;
	wire [4-1:0] node17061;
	wire [4-1:0] node17062;
	wire [4-1:0] node17065;
	wire [4-1:0] node17067;
	wire [4-1:0] node17070;
	wire [4-1:0] node17071;
	wire [4-1:0] node17072;
	wire [4-1:0] node17075;
	wire [4-1:0] node17078;
	wire [4-1:0] node17079;
	wire [4-1:0] node17080;
	wire [4-1:0] node17083;
	wire [4-1:0] node17086;
	wire [4-1:0] node17087;
	wire [4-1:0] node17090;
	wire [4-1:0] node17093;
	wire [4-1:0] node17094;
	wire [4-1:0] node17095;
	wire [4-1:0] node17096;
	wire [4-1:0] node17097;
	wire [4-1:0] node17100;
	wire [4-1:0] node17102;
	wire [4-1:0] node17105;
	wire [4-1:0] node17106;
	wire [4-1:0] node17109;
	wire [4-1:0] node17110;
	wire [4-1:0] node17112;
	wire [4-1:0] node17115;
	wire [4-1:0] node17116;
	wire [4-1:0] node17120;
	wire [4-1:0] node17121;
	wire [4-1:0] node17122;
	wire [4-1:0] node17124;
	wire [4-1:0] node17126;
	wire [4-1:0] node17129;
	wire [4-1:0] node17131;
	wire [4-1:0] node17132;
	wire [4-1:0] node17136;
	wire [4-1:0] node17137;
	wire [4-1:0] node17138;
	wire [4-1:0] node17139;
	wire [4-1:0] node17142;
	wire [4-1:0] node17143;
	wire [4-1:0] node17146;
	wire [4-1:0] node17149;
	wire [4-1:0] node17151;
	wire [4-1:0] node17153;
	wire [4-1:0] node17156;
	wire [4-1:0] node17157;
	wire [4-1:0] node17158;
	wire [4-1:0] node17161;
	wire [4-1:0] node17164;
	wire [4-1:0] node17166;
	wire [4-1:0] node17169;
	wire [4-1:0] node17170;
	wire [4-1:0] node17171;
	wire [4-1:0] node17172;
	wire [4-1:0] node17173;
	wire [4-1:0] node17176;
	wire [4-1:0] node17179;
	wire [4-1:0] node17180;
	wire [4-1:0] node17183;
	wire [4-1:0] node17185;
	wire [4-1:0] node17188;
	wire [4-1:0] node17189;
	wire [4-1:0] node17190;
	wire [4-1:0] node17191;
	wire [4-1:0] node17194;
	wire [4-1:0] node17197;
	wire [4-1:0] node17199;
	wire [4-1:0] node17201;
	wire [4-1:0] node17204;
	wire [4-1:0] node17205;
	wire [4-1:0] node17206;
	wire [4-1:0] node17209;
	wire [4-1:0] node17210;
	wire [4-1:0] node17213;
	wire [4-1:0] node17216;
	wire [4-1:0] node17217;
	wire [4-1:0] node17220;
	wire [4-1:0] node17223;
	wire [4-1:0] node17224;
	wire [4-1:0] node17225;
	wire [4-1:0] node17226;
	wire [4-1:0] node17227;
	wire [4-1:0] node17230;
	wire [4-1:0] node17233;
	wire [4-1:0] node17234;
	wire [4-1:0] node17238;
	wire [4-1:0] node17239;
	wire [4-1:0] node17242;
	wire [4-1:0] node17245;
	wire [4-1:0] node17246;
	wire [4-1:0] node17247;
	wire [4-1:0] node17250;
	wire [4-1:0] node17252;
	wire [4-1:0] node17255;
	wire [4-1:0] node17256;
	wire [4-1:0] node17257;
	wire [4-1:0] node17259;
	wire [4-1:0] node17262;
	wire [4-1:0] node17263;
	wire [4-1:0] node17267;
	wire [4-1:0] node17268;
	wire [4-1:0] node17270;
	wire [4-1:0] node17273;
	wire [4-1:0] node17276;
	wire [4-1:0] node17277;
	wire [4-1:0] node17278;
	wire [4-1:0] node17279;
	wire [4-1:0] node17280;
	wire [4-1:0] node17281;
	wire [4-1:0] node17282;
	wire [4-1:0] node17283;
	wire [4-1:0] node17286;
	wire [4-1:0] node17289;
	wire [4-1:0] node17290;
	wire [4-1:0] node17291;
	wire [4-1:0] node17293;
	wire [4-1:0] node17296;
	wire [4-1:0] node17297;
	wire [4-1:0] node17300;
	wire [4-1:0] node17303;
	wire [4-1:0] node17304;
	wire [4-1:0] node17305;
	wire [4-1:0] node17308;
	wire [4-1:0] node17311;
	wire [4-1:0] node17312;
	wire [4-1:0] node17315;
	wire [4-1:0] node17318;
	wire [4-1:0] node17319;
	wire [4-1:0] node17320;
	wire [4-1:0] node17323;
	wire [4-1:0] node17326;
	wire [4-1:0] node17327;
	wire [4-1:0] node17328;
	wire [4-1:0] node17331;
	wire [4-1:0] node17334;
	wire [4-1:0] node17336;
	wire [4-1:0] node17339;
	wire [4-1:0] node17340;
	wire [4-1:0] node17341;
	wire [4-1:0] node17342;
	wire [4-1:0] node17345;
	wire [4-1:0] node17346;
	wire [4-1:0] node17350;
	wire [4-1:0] node17351;
	wire [4-1:0] node17353;
	wire [4-1:0] node17356;
	wire [4-1:0] node17358;
	wire [4-1:0] node17361;
	wire [4-1:0] node17362;
	wire [4-1:0] node17363;
	wire [4-1:0] node17365;
	wire [4-1:0] node17368;
	wire [4-1:0] node17371;
	wire [4-1:0] node17372;
	wire [4-1:0] node17375;
	wire [4-1:0] node17378;
	wire [4-1:0] node17379;
	wire [4-1:0] node17380;
	wire [4-1:0] node17381;
	wire [4-1:0] node17384;
	wire [4-1:0] node17385;
	wire [4-1:0] node17387;
	wire [4-1:0] node17390;
	wire [4-1:0] node17392;
	wire [4-1:0] node17395;
	wire [4-1:0] node17396;
	wire [4-1:0] node17397;
	wire [4-1:0] node17400;
	wire [4-1:0] node17402;
	wire [4-1:0] node17405;
	wire [4-1:0] node17406;
	wire [4-1:0] node17409;
	wire [4-1:0] node17412;
	wire [4-1:0] node17413;
	wire [4-1:0] node17414;
	wire [4-1:0] node17415;
	wire [4-1:0] node17418;
	wire [4-1:0] node17419;
	wire [4-1:0] node17422;
	wire [4-1:0] node17425;
	wire [4-1:0] node17426;
	wire [4-1:0] node17429;
	wire [4-1:0] node17430;
	wire [4-1:0] node17434;
	wire [4-1:0] node17435;
	wire [4-1:0] node17437;
	wire [4-1:0] node17439;
	wire [4-1:0] node17442;
	wire [4-1:0] node17445;
	wire [4-1:0] node17446;
	wire [4-1:0] node17447;
	wire [4-1:0] node17448;
	wire [4-1:0] node17449;
	wire [4-1:0] node17450;
	wire [4-1:0] node17454;
	wire [4-1:0] node17455;
	wire [4-1:0] node17458;
	wire [4-1:0] node17461;
	wire [4-1:0] node17462;
	wire [4-1:0] node17463;
	wire [4-1:0] node17464;
	wire [4-1:0] node17465;
	wire [4-1:0] node17468;
	wire [4-1:0] node17471;
	wire [4-1:0] node17472;
	wire [4-1:0] node17475;
	wire [4-1:0] node17478;
	wire [4-1:0] node17480;
	wire [4-1:0] node17482;
	wire [4-1:0] node17485;
	wire [4-1:0] node17486;
	wire [4-1:0] node17487;
	wire [4-1:0] node17490;
	wire [4-1:0] node17493;
	wire [4-1:0] node17494;
	wire [4-1:0] node17498;
	wire [4-1:0] node17499;
	wire [4-1:0] node17500;
	wire [4-1:0] node17501;
	wire [4-1:0] node17504;
	wire [4-1:0] node17507;
	wire [4-1:0] node17508;
	wire [4-1:0] node17509;
	wire [4-1:0] node17512;
	wire [4-1:0] node17515;
	wire [4-1:0] node17516;
	wire [4-1:0] node17518;
	wire [4-1:0] node17521;
	wire [4-1:0] node17522;
	wire [4-1:0] node17525;
	wire [4-1:0] node17528;
	wire [4-1:0] node17529;
	wire [4-1:0] node17530;
	wire [4-1:0] node17531;
	wire [4-1:0] node17535;
	wire [4-1:0] node17536;
	wire [4-1:0] node17540;
	wire [4-1:0] node17542;
	wire [4-1:0] node17543;
	wire [4-1:0] node17547;
	wire [4-1:0] node17548;
	wire [4-1:0] node17549;
	wire [4-1:0] node17550;
	wire [4-1:0] node17553;
	wire [4-1:0] node17554;
	wire [4-1:0] node17558;
	wire [4-1:0] node17559;
	wire [4-1:0] node17560;
	wire [4-1:0] node17561;
	wire [4-1:0] node17563;
	wire [4-1:0] node17566;
	wire [4-1:0] node17567;
	wire [4-1:0] node17570;
	wire [4-1:0] node17573;
	wire [4-1:0] node17574;
	wire [4-1:0] node17577;
	wire [4-1:0] node17580;
	wire [4-1:0] node17581;
	wire [4-1:0] node17582;
	wire [4-1:0] node17585;
	wire [4-1:0] node17588;
	wire [4-1:0] node17589;
	wire [4-1:0] node17592;
	wire [4-1:0] node17595;
	wire [4-1:0] node17596;
	wire [4-1:0] node17597;
	wire [4-1:0] node17598;
	wire [4-1:0] node17601;
	wire [4-1:0] node17602;
	wire [4-1:0] node17606;
	wire [4-1:0] node17607;
	wire [4-1:0] node17610;
	wire [4-1:0] node17613;
	wire [4-1:0] node17614;
	wire [4-1:0] node17615;
	wire [4-1:0] node17617;
	wire [4-1:0] node17620;
	wire [4-1:0] node17621;
	wire [4-1:0] node17625;
	wire [4-1:0] node17627;
	wire [4-1:0] node17630;
	wire [4-1:0] node17631;
	wire [4-1:0] node17632;
	wire [4-1:0] node17633;
	wire [4-1:0] node17634;
	wire [4-1:0] node17635;
	wire [4-1:0] node17638;
	wire [4-1:0] node17639;
	wire [4-1:0] node17641;
	wire [4-1:0] node17644;
	wire [4-1:0] node17645;
	wire [4-1:0] node17649;
	wire [4-1:0] node17650;
	wire [4-1:0] node17651;
	wire [4-1:0] node17654;
	wire [4-1:0] node17656;
	wire [4-1:0] node17659;
	wire [4-1:0] node17660;
	wire [4-1:0] node17663;
	wire [4-1:0] node17666;
	wire [4-1:0] node17667;
	wire [4-1:0] node17668;
	wire [4-1:0] node17669;
	wire [4-1:0] node17672;
	wire [4-1:0] node17675;
	wire [4-1:0] node17676;
	wire [4-1:0] node17679;
	wire [4-1:0] node17681;
	wire [4-1:0] node17684;
	wire [4-1:0] node17685;
	wire [4-1:0] node17687;
	wire [4-1:0] node17690;
	wire [4-1:0] node17692;
	wire [4-1:0] node17693;
	wire [4-1:0] node17697;
	wire [4-1:0] node17698;
	wire [4-1:0] node17699;
	wire [4-1:0] node17700;
	wire [4-1:0] node17701;
	wire [4-1:0] node17704;
	wire [4-1:0] node17707;
	wire [4-1:0] node17708;
	wire [4-1:0] node17709;
	wire [4-1:0] node17713;
	wire [4-1:0] node17714;
	wire [4-1:0] node17717;
	wire [4-1:0] node17720;
	wire [4-1:0] node17721;
	wire [4-1:0] node17722;
	wire [4-1:0] node17723;
	wire [4-1:0] node17727;
	wire [4-1:0] node17730;
	wire [4-1:0] node17731;
	wire [4-1:0] node17732;
	wire [4-1:0] node17737;
	wire [4-1:0] node17738;
	wire [4-1:0] node17739;
	wire [4-1:0] node17740;
	wire [4-1:0] node17741;
	wire [4-1:0] node17744;
	wire [4-1:0] node17747;
	wire [4-1:0] node17748;
	wire [4-1:0] node17751;
	wire [4-1:0] node17754;
	wire [4-1:0] node17755;
	wire [4-1:0] node17758;
	wire [4-1:0] node17761;
	wire [4-1:0] node17762;
	wire [4-1:0] node17763;
	wire [4-1:0] node17766;
	wire [4-1:0] node17769;
	wire [4-1:0] node17770;
	wire [4-1:0] node17772;
	wire [4-1:0] node17775;
	wire [4-1:0] node17777;
	wire [4-1:0] node17780;
	wire [4-1:0] node17781;
	wire [4-1:0] node17782;
	wire [4-1:0] node17783;
	wire [4-1:0] node17784;
	wire [4-1:0] node17785;
	wire [4-1:0] node17789;
	wire [4-1:0] node17790;
	wire [4-1:0] node17794;
	wire [4-1:0] node17795;
	wire [4-1:0] node17796;
	wire [4-1:0] node17797;
	wire [4-1:0] node17801;
	wire [4-1:0] node17804;
	wire [4-1:0] node17805;
	wire [4-1:0] node17806;
	wire [4-1:0] node17807;
	wire [4-1:0] node17812;
	wire [4-1:0] node17813;
	wire [4-1:0] node17817;
	wire [4-1:0] node17818;
	wire [4-1:0] node17819;
	wire [4-1:0] node17820;
	wire [4-1:0] node17824;
	wire [4-1:0] node17826;
	wire [4-1:0] node17829;
	wire [4-1:0] node17830;
	wire [4-1:0] node17831;
	wire [4-1:0] node17832;
	wire [4-1:0] node17836;
	wire [4-1:0] node17838;
	wire [4-1:0] node17841;
	wire [4-1:0] node17842;
	wire [4-1:0] node17843;
	wire [4-1:0] node17848;
	wire [4-1:0] node17849;
	wire [4-1:0] node17850;
	wire [4-1:0] node17851;
	wire [4-1:0] node17852;
	wire [4-1:0] node17856;
	wire [4-1:0] node17857;
	wire [4-1:0] node17858;
	wire [4-1:0] node17862;
	wire [4-1:0] node17865;
	wire [4-1:0] node17866;
	wire [4-1:0] node17868;
	wire [4-1:0] node17871;
	wire [4-1:0] node17872;
	wire [4-1:0] node17874;
	wire [4-1:0] node17877;
	wire [4-1:0] node17878;
	wire [4-1:0] node17882;
	wire [4-1:0] node17883;
	wire [4-1:0] node17884;
	wire [4-1:0] node17885;
	wire [4-1:0] node17886;
	wire [4-1:0] node17889;
	wire [4-1:0] node17892;
	wire [4-1:0] node17893;
	wire [4-1:0] node17894;
	wire [4-1:0] node17897;
	wire [4-1:0] node17900;
	wire [4-1:0] node17901;
	wire [4-1:0] node17905;
	wire [4-1:0] node17906;
	wire [4-1:0] node17907;
	wire [4-1:0] node17908;
	wire [4-1:0] node17913;
	wire [4-1:0] node17914;
	wire [4-1:0] node17915;
	wire [4-1:0] node17919;
	wire [4-1:0] node17920;
	wire [4-1:0] node17924;
	wire [4-1:0] node17925;
	wire [4-1:0] node17926;
	wire [4-1:0] node17929;
	wire [4-1:0] node17931;
	wire [4-1:0] node17934;
	wire [4-1:0] node17935;
	wire [4-1:0] node17936;
	wire [4-1:0] node17940;
	wire [4-1:0] node17942;
	wire [4-1:0] node17945;
	wire [4-1:0] node17946;
	wire [4-1:0] node17947;
	wire [4-1:0] node17948;
	wire [4-1:0] node17949;
	wire [4-1:0] node17950;
	wire [4-1:0] node17951;
	wire [4-1:0] node17952;
	wire [4-1:0] node17953;
	wire [4-1:0] node17954;
	wire [4-1:0] node17957;
	wire [4-1:0] node17960;
	wire [4-1:0] node17961;
	wire [4-1:0] node17964;
	wire [4-1:0] node17967;
	wire [4-1:0] node17968;
	wire [4-1:0] node17969;
	wire [4-1:0] node17972;
	wire [4-1:0] node17975;
	wire [4-1:0] node17976;
	wire [4-1:0] node17977;
	wire [4-1:0] node17980;
	wire [4-1:0] node17983;
	wire [4-1:0] node17984;
	wire [4-1:0] node17987;
	wire [4-1:0] node17990;
	wire [4-1:0] node17991;
	wire [4-1:0] node17992;
	wire [4-1:0] node17993;
	wire [4-1:0] node17994;
	wire [4-1:0] node17997;
	wire [4-1:0] node18000;
	wire [4-1:0] node18001;
	wire [4-1:0] node18004;
	wire [4-1:0] node18007;
	wire [4-1:0] node18008;
	wire [4-1:0] node18009;
	wire [4-1:0] node18013;
	wire [4-1:0] node18014;
	wire [4-1:0] node18018;
	wire [4-1:0] node18019;
	wire [4-1:0] node18020;
	wire [4-1:0] node18021;
	wire [4-1:0] node18024;
	wire [4-1:0] node18028;
	wire [4-1:0] node18030;
	wire [4-1:0] node18031;
	wire [4-1:0] node18034;
	wire [4-1:0] node18037;
	wire [4-1:0] node18038;
	wire [4-1:0] node18039;
	wire [4-1:0] node18040;
	wire [4-1:0] node18041;
	wire [4-1:0] node18044;
	wire [4-1:0] node18045;
	wire [4-1:0] node18048;
	wire [4-1:0] node18051;
	wire [4-1:0] node18052;
	wire [4-1:0] node18053;
	wire [4-1:0] node18057;
	wire [4-1:0] node18060;
	wire [4-1:0] node18061;
	wire [4-1:0] node18063;
	wire [4-1:0] node18064;
	wire [4-1:0] node18068;
	wire [4-1:0] node18069;
	wire [4-1:0] node18070;
	wire [4-1:0] node18073;
	wire [4-1:0] node18076;
	wire [4-1:0] node18077;
	wire [4-1:0] node18080;
	wire [4-1:0] node18083;
	wire [4-1:0] node18084;
	wire [4-1:0] node18085;
	wire [4-1:0] node18086;
	wire [4-1:0] node18089;
	wire [4-1:0] node18091;
	wire [4-1:0] node18094;
	wire [4-1:0] node18095;
	wire [4-1:0] node18098;
	wire [4-1:0] node18101;
	wire [4-1:0] node18102;
	wire [4-1:0] node18103;
	wire [4-1:0] node18105;
	wire [4-1:0] node18108;
	wire [4-1:0] node18109;
	wire [4-1:0] node18113;
	wire [4-1:0] node18115;
	wire [4-1:0] node18116;
	wire [4-1:0] node18120;
	wire [4-1:0] node18121;
	wire [4-1:0] node18122;
	wire [4-1:0] node18123;
	wire [4-1:0] node18124;
	wire [4-1:0] node18125;
	wire [4-1:0] node18128;
	wire [4-1:0] node18131;
	wire [4-1:0] node18132;
	wire [4-1:0] node18133;
	wire [4-1:0] node18137;
	wire [4-1:0] node18138;
	wire [4-1:0] node18142;
	wire [4-1:0] node18143;
	wire [4-1:0] node18144;
	wire [4-1:0] node18145;
	wire [4-1:0] node18148;
	wire [4-1:0] node18151;
	wire [4-1:0] node18152;
	wire [4-1:0] node18155;
	wire [4-1:0] node18158;
	wire [4-1:0] node18159;
	wire [4-1:0] node18162;
	wire [4-1:0] node18165;
	wire [4-1:0] node18166;
	wire [4-1:0] node18167;
	wire [4-1:0] node18169;
	wire [4-1:0] node18171;
	wire [4-1:0] node18174;
	wire [4-1:0] node18175;
	wire [4-1:0] node18178;
	wire [4-1:0] node18180;
	wire [4-1:0] node18183;
	wire [4-1:0] node18184;
	wire [4-1:0] node18186;
	wire [4-1:0] node18189;
	wire [4-1:0] node18191;
	wire [4-1:0] node18194;
	wire [4-1:0] node18195;
	wire [4-1:0] node18196;
	wire [4-1:0] node18197;
	wire [4-1:0] node18198;
	wire [4-1:0] node18201;
	wire [4-1:0] node18204;
	wire [4-1:0] node18205;
	wire [4-1:0] node18208;
	wire [4-1:0] node18209;
	wire [4-1:0] node18212;
	wire [4-1:0] node18215;
	wire [4-1:0] node18216;
	wire [4-1:0] node18217;
	wire [4-1:0] node18221;
	wire [4-1:0] node18223;
	wire [4-1:0] node18224;
	wire [4-1:0] node18228;
	wire [4-1:0] node18229;
	wire [4-1:0] node18230;
	wire [4-1:0] node18231;
	wire [4-1:0] node18232;
	wire [4-1:0] node18236;
	wire [4-1:0] node18238;
	wire [4-1:0] node18241;
	wire [4-1:0] node18242;
	wire [4-1:0] node18243;
	wire [4-1:0] node18247;
	wire [4-1:0] node18248;
	wire [4-1:0] node18251;
	wire [4-1:0] node18254;
	wire [4-1:0] node18255;
	wire [4-1:0] node18256;
	wire [4-1:0] node18259;
	wire [4-1:0] node18260;
	wire [4-1:0] node18263;
	wire [4-1:0] node18266;
	wire [4-1:0] node18267;
	wire [4-1:0] node18270;
	wire [4-1:0] node18273;
	wire [4-1:0] node18274;
	wire [4-1:0] node18275;
	wire [4-1:0] node18276;
	wire [4-1:0] node18277;
	wire [4-1:0] node18278;
	wire [4-1:0] node18281;
	wire [4-1:0] node18284;
	wire [4-1:0] node18285;
	wire [4-1:0] node18286;
	wire [4-1:0] node18290;
	wire [4-1:0] node18291;
	wire [4-1:0] node18294;
	wire [4-1:0] node18297;
	wire [4-1:0] node18298;
	wire [4-1:0] node18299;
	wire [4-1:0] node18300;
	wire [4-1:0] node18301;
	wire [4-1:0] node18304;
	wire [4-1:0] node18307;
	wire [4-1:0] node18309;
	wire [4-1:0] node18312;
	wire [4-1:0] node18314;
	wire [4-1:0] node18315;
	wire [4-1:0] node18318;
	wire [4-1:0] node18321;
	wire [4-1:0] node18322;
	wire [4-1:0] node18325;
	wire [4-1:0] node18328;
	wire [4-1:0] node18329;
	wire [4-1:0] node18330;
	wire [4-1:0] node18331;
	wire [4-1:0] node18332;
	wire [4-1:0] node18335;
	wire [4-1:0] node18338;
	wire [4-1:0] node18341;
	wire [4-1:0] node18342;
	wire [4-1:0] node18345;
	wire [4-1:0] node18346;
	wire [4-1:0] node18347;
	wire [4-1:0] node18350;
	wire [4-1:0] node18353;
	wire [4-1:0] node18355;
	wire [4-1:0] node18358;
	wire [4-1:0] node18359;
	wire [4-1:0] node18360;
	wire [4-1:0] node18361;
	wire [4-1:0] node18364;
	wire [4-1:0] node18367;
	wire [4-1:0] node18368;
	wire [4-1:0] node18369;
	wire [4-1:0] node18373;
	wire [4-1:0] node18375;
	wire [4-1:0] node18378;
	wire [4-1:0] node18379;
	wire [4-1:0] node18380;
	wire [4-1:0] node18381;
	wire [4-1:0] node18385;
	wire [4-1:0] node18386;
	wire [4-1:0] node18389;
	wire [4-1:0] node18392;
	wire [4-1:0] node18393;
	wire [4-1:0] node18394;
	wire [4-1:0] node18397;
	wire [4-1:0] node18401;
	wire [4-1:0] node18402;
	wire [4-1:0] node18403;
	wire [4-1:0] node18404;
	wire [4-1:0] node18405;
	wire [4-1:0] node18406;
	wire [4-1:0] node18410;
	wire [4-1:0] node18411;
	wire [4-1:0] node18415;
	wire [4-1:0] node18416;
	wire [4-1:0] node18419;
	wire [4-1:0] node18422;
	wire [4-1:0] node18423;
	wire [4-1:0] node18424;
	wire [4-1:0] node18425;
	wire [4-1:0] node18429;
	wire [4-1:0] node18430;
	wire [4-1:0] node18434;
	wire [4-1:0] node18435;
	wire [4-1:0] node18438;
	wire [4-1:0] node18439;
	wire [4-1:0] node18442;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18447;
	wire [4-1:0] node18448;
	wire [4-1:0] node18449;
	wire [4-1:0] node18453;
	wire [4-1:0] node18454;
	wire [4-1:0] node18458;
	wire [4-1:0] node18459;
	wire [4-1:0] node18460;
	wire [4-1:0] node18464;
	wire [4-1:0] node18465;
	wire [4-1:0] node18469;
	wire [4-1:0] node18470;
	wire [4-1:0] node18471;
	wire [4-1:0] node18472;
	wire [4-1:0] node18476;
	wire [4-1:0] node18477;
	wire [4-1:0] node18481;
	wire [4-1:0] node18482;
	wire [4-1:0] node18485;
	wire [4-1:0] node18486;
	wire [4-1:0] node18489;
	wire [4-1:0] node18492;
	wire [4-1:0] node18493;
	wire [4-1:0] node18494;
	wire [4-1:0] node18495;
	wire [4-1:0] node18496;
	wire [4-1:0] node18497;
	wire [4-1:0] node18499;
	wire [4-1:0] node18500;
	wire [4-1:0] node18502;
	wire [4-1:0] node18505;
	wire [4-1:0] node18508;
	wire [4-1:0] node18510;
	wire [4-1:0] node18511;
	wire [4-1:0] node18513;
	wire [4-1:0] node18517;
	wire [4-1:0] node18518;
	wire [4-1:0] node18520;
	wire [4-1:0] node18521;
	wire [4-1:0] node18522;
	wire [4-1:0] node18525;
	wire [4-1:0] node18528;
	wire [4-1:0] node18530;
	wire [4-1:0] node18533;
	wire [4-1:0] node18535;
	wire [4-1:0] node18536;
	wire [4-1:0] node18539;
	wire [4-1:0] node18542;
	wire [4-1:0] node18543;
	wire [4-1:0] node18544;
	wire [4-1:0] node18545;
	wire [4-1:0] node18546;
	wire [4-1:0] node18550;
	wire [4-1:0] node18551;
	wire [4-1:0] node18555;
	wire [4-1:0] node18556;
	wire [4-1:0] node18557;
	wire [4-1:0] node18561;
	wire [4-1:0] node18562;
	wire [4-1:0] node18566;
	wire [4-1:0] node18567;
	wire [4-1:0] node18568;
	wire [4-1:0] node18570;
	wire [4-1:0] node18573;
	wire [4-1:0] node18574;
	wire [4-1:0] node18578;
	wire [4-1:0] node18579;
	wire [4-1:0] node18581;
	wire [4-1:0] node18584;
	wire [4-1:0] node18586;
	wire [4-1:0] node18589;
	wire [4-1:0] node18590;
	wire [4-1:0] node18591;
	wire [4-1:0] node18592;
	wire [4-1:0] node18593;
	wire [4-1:0] node18596;
	wire [4-1:0] node18599;
	wire [4-1:0] node18600;
	wire [4-1:0] node18602;
	wire [4-1:0] node18603;
	wire [4-1:0] node18607;
	wire [4-1:0] node18608;
	wire [4-1:0] node18609;
	wire [4-1:0] node18612;
	wire [4-1:0] node18615;
	wire [4-1:0] node18616;
	wire [4-1:0] node18619;
	wire [4-1:0] node18622;
	wire [4-1:0] node18623;
	wire [4-1:0] node18624;
	wire [4-1:0] node18626;
	wire [4-1:0] node18627;
	wire [4-1:0] node18630;
	wire [4-1:0] node18633;
	wire [4-1:0] node18634;
	wire [4-1:0] node18636;
	wire [4-1:0] node18640;
	wire [4-1:0] node18641;
	wire [4-1:0] node18643;
	wire [4-1:0] node18646;
	wire [4-1:0] node18648;
	wire [4-1:0] node18651;
	wire [4-1:0] node18652;
	wire [4-1:0] node18653;
	wire [4-1:0] node18654;
	wire [4-1:0] node18657;
	wire [4-1:0] node18660;
	wire [4-1:0] node18661;
	wire [4-1:0] node18662;
	wire [4-1:0] node18663;
	wire [4-1:0] node18667;
	wire [4-1:0] node18669;
	wire [4-1:0] node18672;
	wire [4-1:0] node18674;
	wire [4-1:0] node18677;
	wire [4-1:0] node18678;
	wire [4-1:0] node18679;
	wire [4-1:0] node18682;
	wire [4-1:0] node18685;
	wire [4-1:0] node18686;
	wire [4-1:0] node18687;
	wire [4-1:0] node18688;
	wire [4-1:0] node18692;
	wire [4-1:0] node18694;
	wire [4-1:0] node18698;
	wire [4-1:0] node18699;
	wire [4-1:0] node18700;
	wire [4-1:0] node18701;
	wire [4-1:0] node18702;
	wire [4-1:0] node18703;
	wire [4-1:0] node18705;
	wire [4-1:0] node18708;
	wire [4-1:0] node18710;
	wire [4-1:0] node18713;
	wire [4-1:0] node18714;
	wire [4-1:0] node18716;
	wire [4-1:0] node18719;
	wire [4-1:0] node18721;
	wire [4-1:0] node18724;
	wire [4-1:0] node18725;
	wire [4-1:0] node18726;
	wire [4-1:0] node18728;
	wire [4-1:0] node18731;
	wire [4-1:0] node18733;
	wire [4-1:0] node18736;
	wire [4-1:0] node18737;
	wire [4-1:0] node18739;
	wire [4-1:0] node18743;
	wire [4-1:0] node18744;
	wire [4-1:0] node18745;
	wire [4-1:0] node18746;
	wire [4-1:0] node18747;
	wire [4-1:0] node18751;
	wire [4-1:0] node18752;
	wire [4-1:0] node18756;
	wire [4-1:0] node18757;
	wire [4-1:0] node18759;
	wire [4-1:0] node18762;
	wire [4-1:0] node18764;
	wire [4-1:0] node18767;
	wire [4-1:0] node18768;
	wire [4-1:0] node18769;
	wire [4-1:0] node18772;
	wire [4-1:0] node18774;
	wire [4-1:0] node18776;
	wire [4-1:0] node18779;
	wire [4-1:0] node18780;
	wire [4-1:0] node18781;
	wire [4-1:0] node18782;
	wire [4-1:0] node18786;
	wire [4-1:0] node18787;
	wire [4-1:0] node18791;
	wire [4-1:0] node18792;
	wire [4-1:0] node18793;
	wire [4-1:0] node18798;
	wire [4-1:0] node18799;
	wire [4-1:0] node18800;
	wire [4-1:0] node18801;
	wire [4-1:0] node18802;
	wire [4-1:0] node18804;
	wire [4-1:0] node18805;
	wire [4-1:0] node18809;
	wire [4-1:0] node18810;
	wire [4-1:0] node18812;
	wire [4-1:0] node18815;
	wire [4-1:0] node18816;
	wire [4-1:0] node18819;
	wire [4-1:0] node18822;
	wire [4-1:0] node18823;
	wire [4-1:0] node18825;
	wire [4-1:0] node18828;
	wire [4-1:0] node18829;
	wire [4-1:0] node18830;
	wire [4-1:0] node18835;
	wire [4-1:0] node18836;
	wire [4-1:0] node18837;
	wire [4-1:0] node18841;
	wire [4-1:0] node18842;
	wire [4-1:0] node18843;
	wire [4-1:0] node18846;
	wire [4-1:0] node18849;
	wire [4-1:0] node18850;
	wire [4-1:0] node18851;
	wire [4-1:0] node18854;
	wire [4-1:0] node18857;
	wire [4-1:0] node18858;
	wire [4-1:0] node18861;
	wire [4-1:0] node18864;
	wire [4-1:0] node18865;
	wire [4-1:0] node18866;
	wire [4-1:0] node18867;
	wire [4-1:0] node18868;
	wire [4-1:0] node18871;
	wire [4-1:0] node18874;
	wire [4-1:0] node18875;
	wire [4-1:0] node18876;
	wire [4-1:0] node18879;
	wire [4-1:0] node18882;
	wire [4-1:0] node18883;
	wire [4-1:0] node18887;
	wire [4-1:0] node18888;
	wire [4-1:0] node18890;
	wire [4-1:0] node18891;
	wire [4-1:0] node18895;
	wire [4-1:0] node18896;
	wire [4-1:0] node18899;
	wire [4-1:0] node18902;
	wire [4-1:0] node18903;
	wire [4-1:0] node18904;
	wire [4-1:0] node18905;
	wire [4-1:0] node18909;
	wire [4-1:0] node18912;
	wire [4-1:0] node18913;
	wire [4-1:0] node18914;
	wire [4-1:0] node18918;
	wire [4-1:0] node18920;
	wire [4-1:0] node18923;
	wire [4-1:0] node18924;
	wire [4-1:0] node18925;
	wire [4-1:0] node18926;
	wire [4-1:0] node18927;
	wire [4-1:0] node18928;
	wire [4-1:0] node18929;
	wire [4-1:0] node18930;
	wire [4-1:0] node18931;
	wire [4-1:0] node18934;
	wire [4-1:0] node18937;
	wire [4-1:0] node18938;
	wire [4-1:0] node18942;
	wire [4-1:0] node18944;
	wire [4-1:0] node18946;
	wire [4-1:0] node18949;
	wire [4-1:0] node18950;
	wire [4-1:0] node18951;
	wire [4-1:0] node18952;
	wire [4-1:0] node18953;
	wire [4-1:0] node18956;
	wire [4-1:0] node18959;
	wire [4-1:0] node18961;
	wire [4-1:0] node18964;
	wire [4-1:0] node18965;
	wire [4-1:0] node18967;
	wire [4-1:0] node18970;
	wire [4-1:0] node18971;
	wire [4-1:0] node18975;
	wire [4-1:0] node18976;
	wire [4-1:0] node18977;
	wire [4-1:0] node18978;
	wire [4-1:0] node18982;
	wire [4-1:0] node18984;
	wire [4-1:0] node18987;
	wire [4-1:0] node18988;
	wire [4-1:0] node18989;
	wire [4-1:0] node18992;
	wire [4-1:0] node18995;
	wire [4-1:0] node18996;
	wire [4-1:0] node18999;
	wire [4-1:0] node19002;
	wire [4-1:0] node19003;
	wire [4-1:0] node19004;
	wire [4-1:0] node19005;
	wire [4-1:0] node19006;
	wire [4-1:0] node19010;
	wire [4-1:0] node19012;
	wire [4-1:0] node19015;
	wire [4-1:0] node19017;
	wire [4-1:0] node19018;
	wire [4-1:0] node19021;
	wire [4-1:0] node19024;
	wire [4-1:0] node19025;
	wire [4-1:0] node19026;
	wire [4-1:0] node19027;
	wire [4-1:0] node19029;
	wire [4-1:0] node19032;
	wire [4-1:0] node19033;
	wire [4-1:0] node19036;
	wire [4-1:0] node19039;
	wire [4-1:0] node19040;
	wire [4-1:0] node19041;
	wire [4-1:0] node19046;
	wire [4-1:0] node19047;
	wire [4-1:0] node19048;
	wire [4-1:0] node19049;
	wire [4-1:0] node19052;
	wire [4-1:0] node19056;
	wire [4-1:0] node19057;
	wire [4-1:0] node19058;
	wire [4-1:0] node19061;
	wire [4-1:0] node19064;
	wire [4-1:0] node19065;
	wire [4-1:0] node19068;
	wire [4-1:0] node19071;
	wire [4-1:0] node19072;
	wire [4-1:0] node19073;
	wire [4-1:0] node19074;
	wire [4-1:0] node19075;
	wire [4-1:0] node19076;
	wire [4-1:0] node19079;
	wire [4-1:0] node19082;
	wire [4-1:0] node19083;
	wire [4-1:0] node19085;
	wire [4-1:0] node19089;
	wire [4-1:0] node19090;
	wire [4-1:0] node19091;
	wire [4-1:0] node19092;
	wire [4-1:0] node19096;
	wire [4-1:0] node19097;
	wire [4-1:0] node19100;
	wire [4-1:0] node19103;
	wire [4-1:0] node19106;
	wire [4-1:0] node19107;
	wire [4-1:0] node19108;
	wire [4-1:0] node19109;
	wire [4-1:0] node19112;
	wire [4-1:0] node19115;
	wire [4-1:0] node19116;
	wire [4-1:0] node19119;
	wire [4-1:0] node19122;
	wire [4-1:0] node19123;
	wire [4-1:0] node19124;
	wire [4-1:0] node19127;
	wire [4-1:0] node19130;
	wire [4-1:0] node19131;
	wire [4-1:0] node19134;
	wire [4-1:0] node19137;
	wire [4-1:0] node19138;
	wire [4-1:0] node19139;
	wire [4-1:0] node19140;
	wire [4-1:0] node19141;
	wire [4-1:0] node19144;
	wire [4-1:0] node19147;
	wire [4-1:0] node19148;
	wire [4-1:0] node19149;
	wire [4-1:0] node19153;
	wire [4-1:0] node19154;
	wire [4-1:0] node19157;
	wire [4-1:0] node19160;
	wire [4-1:0] node19161;
	wire [4-1:0] node19162;
	wire [4-1:0] node19163;
	wire [4-1:0] node19166;
	wire [4-1:0] node19170;
	wire [4-1:0] node19171;
	wire [4-1:0] node19172;
	wire [4-1:0] node19175;
	wire [4-1:0] node19178;
	wire [4-1:0] node19179;
	wire [4-1:0] node19183;
	wire [4-1:0] node19184;
	wire [4-1:0] node19185;
	wire [4-1:0] node19186;
	wire [4-1:0] node19190;
	wire [4-1:0] node19191;
	wire [4-1:0] node19194;
	wire [4-1:0] node19197;
	wire [4-1:0] node19198;
	wire [4-1:0] node19199;
	wire [4-1:0] node19200;
	wire [4-1:0] node19204;
	wire [4-1:0] node19206;
	wire [4-1:0] node19209;
	wire [4-1:0] node19210;
	wire [4-1:0] node19211;
	wire [4-1:0] node19214;
	wire [4-1:0] node19218;
	wire [4-1:0] node19219;
	wire [4-1:0] node19220;
	wire [4-1:0] node19221;
	wire [4-1:0] node19222;
	wire [4-1:0] node19223;
	wire [4-1:0] node19226;
	wire [4-1:0] node19229;
	wire [4-1:0] node19230;
	wire [4-1:0] node19231;
	wire [4-1:0] node19234;
	wire [4-1:0] node19237;
	wire [4-1:0] node19238;
	wire [4-1:0] node19242;
	wire [4-1:0] node19243;
	wire [4-1:0] node19244;
	wire [4-1:0] node19245;
	wire [4-1:0] node19246;
	wire [4-1:0] node19251;
	wire [4-1:0] node19253;
	wire [4-1:0] node19254;
	wire [4-1:0] node19257;
	wire [4-1:0] node19260;
	wire [4-1:0] node19261;
	wire [4-1:0] node19264;
	wire [4-1:0] node19267;
	wire [4-1:0] node19268;
	wire [4-1:0] node19269;
	wire [4-1:0] node19270;
	wire [4-1:0] node19271;
	wire [4-1:0] node19275;
	wire [4-1:0] node19276;
	wire [4-1:0] node19279;
	wire [4-1:0] node19282;
	wire [4-1:0] node19283;
	wire [4-1:0] node19284;
	wire [4-1:0] node19287;
	wire [4-1:0] node19290;
	wire [4-1:0] node19292;
	wire [4-1:0] node19295;
	wire [4-1:0] node19296;
	wire [4-1:0] node19297;
	wire [4-1:0] node19298;
	wire [4-1:0] node19301;
	wire [4-1:0] node19304;
	wire [4-1:0] node19306;
	wire [4-1:0] node19309;
	wire [4-1:0] node19310;
	wire [4-1:0] node19311;
	wire [4-1:0] node19314;
	wire [4-1:0] node19317;
	wire [4-1:0] node19320;
	wire [4-1:0] node19321;
	wire [4-1:0] node19322;
	wire [4-1:0] node19323;
	wire [4-1:0] node19325;
	wire [4-1:0] node19327;
	wire [4-1:0] node19330;
	wire [4-1:0] node19332;
	wire [4-1:0] node19335;
	wire [4-1:0] node19336;
	wire [4-1:0] node19337;
	wire [4-1:0] node19338;
	wire [4-1:0] node19339;
	wire [4-1:0] node19343;
	wire [4-1:0] node19344;
	wire [4-1:0] node19347;
	wire [4-1:0] node19350;
	wire [4-1:0] node19351;
	wire [4-1:0] node19352;
	wire [4-1:0] node19356;
	wire [4-1:0] node19358;
	wire [4-1:0] node19361;
	wire [4-1:0] node19362;
	wire [4-1:0] node19363;
	wire [4-1:0] node19364;
	wire [4-1:0] node19368;
	wire [4-1:0] node19369;
	wire [4-1:0] node19372;
	wire [4-1:0] node19375;
	wire [4-1:0] node19376;
	wire [4-1:0] node19379;
	wire [4-1:0] node19382;
	wire [4-1:0] node19383;
	wire [4-1:0] node19384;
	wire [4-1:0] node19385;
	wire [4-1:0] node19388;
	wire [4-1:0] node19389;
	wire [4-1:0] node19393;
	wire [4-1:0] node19394;
	wire [4-1:0] node19396;
	wire [4-1:0] node19399;
	wire [4-1:0] node19401;
	wire [4-1:0] node19404;
	wire [4-1:0] node19405;
	wire [4-1:0] node19406;
	wire [4-1:0] node19407;
	wire [4-1:0] node19408;
	wire [4-1:0] node19413;
	wire [4-1:0] node19414;
	wire [4-1:0] node19417;
	wire [4-1:0] node19420;
	wire [4-1:0] node19421;
	wire [4-1:0] node19422;
	wire [4-1:0] node19426;
	wire [4-1:0] node19427;
	wire [4-1:0] node19430;
	wire [4-1:0] node19433;
	wire [4-1:0] node19434;
	wire [4-1:0] node19435;
	wire [4-1:0] node19436;
	wire [4-1:0] node19437;
	wire [4-1:0] node19438;
	wire [4-1:0] node19439;
	wire [4-1:0] node19440;
	wire [4-1:0] node19441;
	wire [4-1:0] node19444;
	wire [4-1:0] node19447;
	wire [4-1:0] node19449;
	wire [4-1:0] node19452;
	wire [4-1:0] node19454;
	wire [4-1:0] node19457;
	wire [4-1:0] node19458;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19463;
	wire [4-1:0] node19466;
	wire [4-1:0] node19467;
	wire [4-1:0] node19470;
	wire [4-1:0] node19473;
	wire [4-1:0] node19474;
	wire [4-1:0] node19476;
	wire [4-1:0] node19479;
	wire [4-1:0] node19480;
	wire [4-1:0] node19483;
	wire [4-1:0] node19486;
	wire [4-1:0] node19487;
	wire [4-1:0] node19488;
	wire [4-1:0] node19491;
	wire [4-1:0] node19494;
	wire [4-1:0] node19495;
	wire [4-1:0] node19496;
	wire [4-1:0] node19497;
	wire [4-1:0] node19500;
	wire [4-1:0] node19503;
	wire [4-1:0] node19504;
	wire [4-1:0] node19508;
	wire [4-1:0] node19509;
	wire [4-1:0] node19512;
	wire [4-1:0] node19515;
	wire [4-1:0] node19516;
	wire [4-1:0] node19517;
	wire [4-1:0] node19518;
	wire [4-1:0] node19519;
	wire [4-1:0] node19520;
	wire [4-1:0] node19524;
	wire [4-1:0] node19525;
	wire [4-1:0] node19528;
	wire [4-1:0] node19531;
	wire [4-1:0] node19532;
	wire [4-1:0] node19535;
	wire [4-1:0] node19536;
	wire [4-1:0] node19540;
	wire [4-1:0] node19541;
	wire [4-1:0] node19542;
	wire [4-1:0] node19543;
	wire [4-1:0] node19547;
	wire [4-1:0] node19549;
	wire [4-1:0] node19552;
	wire [4-1:0] node19553;
	wire [4-1:0] node19556;
	wire [4-1:0] node19559;
	wire [4-1:0] node19560;
	wire [4-1:0] node19561;
	wire [4-1:0] node19563;
	wire [4-1:0] node19566;
	wire [4-1:0] node19569;
	wire [4-1:0] node19570;
	wire [4-1:0] node19571;
	wire [4-1:0] node19574;
	wire [4-1:0] node19577;
	wire [4-1:0] node19578;
	wire [4-1:0] node19579;
	wire [4-1:0] node19583;
	wire [4-1:0] node19585;
	wire [4-1:0] node19588;
	wire [4-1:0] node19589;
	wire [4-1:0] node19590;
	wire [4-1:0] node19591;
	wire [4-1:0] node19592;
	wire [4-1:0] node19593;
	wire [4-1:0] node19596;
	wire [4-1:0] node19599;
	wire [4-1:0] node19600;
	wire [4-1:0] node19602;
	wire [4-1:0] node19605;
	wire [4-1:0] node19606;
	wire [4-1:0] node19610;
	wire [4-1:0] node19611;
	wire [4-1:0] node19612;
	wire [4-1:0] node19613;
	wire [4-1:0] node19616;
	wire [4-1:0] node19619;
	wire [4-1:0] node19620;
	wire [4-1:0] node19624;
	wire [4-1:0] node19625;
	wire [4-1:0] node19629;
	wire [4-1:0] node19630;
	wire [4-1:0] node19631;
	wire [4-1:0] node19632;
	wire [4-1:0] node19635;
	wire [4-1:0] node19638;
	wire [4-1:0] node19639;
	wire [4-1:0] node19642;
	wire [4-1:0] node19645;
	wire [4-1:0] node19646;
	wire [4-1:0] node19648;
	wire [4-1:0] node19651;
	wire [4-1:0] node19653;
	wire [4-1:0] node19656;
	wire [4-1:0] node19657;
	wire [4-1:0] node19658;
	wire [4-1:0] node19659;
	wire [4-1:0] node19660;
	wire [4-1:0] node19663;
	wire [4-1:0] node19666;
	wire [4-1:0] node19669;
	wire [4-1:0] node19670;
	wire [4-1:0] node19671;
	wire [4-1:0] node19675;
	wire [4-1:0] node19676;
	wire [4-1:0] node19679;
	wire [4-1:0] node19682;
	wire [4-1:0] node19683;
	wire [4-1:0] node19684;
	wire [4-1:0] node19685;
	wire [4-1:0] node19686;
	wire [4-1:0] node19690;
	wire [4-1:0] node19691;
	wire [4-1:0] node19694;
	wire [4-1:0] node19697;
	wire [4-1:0] node19698;
	wire [4-1:0] node19699;
	wire [4-1:0] node19703;
	wire [4-1:0] node19704;
	wire [4-1:0] node19707;
	wire [4-1:0] node19710;
	wire [4-1:0] node19711;
	wire [4-1:0] node19712;
	wire [4-1:0] node19713;
	wire [4-1:0] node19717;
	wire [4-1:0] node19719;
	wire [4-1:0] node19722;
	wire [4-1:0] node19723;
	wire [4-1:0] node19725;
	wire [4-1:0] node19728;
	wire [4-1:0] node19729;
	wire [4-1:0] node19733;
	wire [4-1:0] node19734;
	wire [4-1:0] node19735;
	wire [4-1:0] node19736;
	wire [4-1:0] node19737;
	wire [4-1:0] node19738;
	wire [4-1:0] node19739;
	wire [4-1:0] node19742;
	wire [4-1:0] node19745;
	wire [4-1:0] node19748;
	wire [4-1:0] node19749;
	wire [4-1:0] node19750;
	wire [4-1:0] node19753;
	wire [4-1:0] node19756;
	wire [4-1:0] node19757;
	wire [4-1:0] node19760;
	wire [4-1:0] node19763;
	wire [4-1:0] node19764;
	wire [4-1:0] node19765;
	wire [4-1:0] node19767;
	wire [4-1:0] node19770;
	wire [4-1:0] node19772;
	wire [4-1:0] node19775;
	wire [4-1:0] node19777;
	wire [4-1:0] node19778;
	wire [4-1:0] node19782;
	wire [4-1:0] node19783;
	wire [4-1:0] node19784;
	wire [4-1:0] node19785;
	wire [4-1:0] node19786;
	wire [4-1:0] node19790;
	wire [4-1:0] node19791;
	wire [4-1:0] node19794;
	wire [4-1:0] node19797;
	wire [4-1:0] node19798;
	wire [4-1:0] node19799;
	wire [4-1:0] node19803;
	wire [4-1:0] node19806;
	wire [4-1:0] node19807;
	wire [4-1:0] node19808;
	wire [4-1:0] node19809;
	wire [4-1:0] node19813;
	wire [4-1:0] node19815;
	wire [4-1:0] node19818;
	wire [4-1:0] node19820;
	wire [4-1:0] node19823;
	wire [4-1:0] node19824;
	wire [4-1:0] node19825;
	wire [4-1:0] node19826;
	wire [4-1:0] node19828;
	wire [4-1:0] node19829;
	wire [4-1:0] node19830;
	wire [4-1:0] node19833;
	wire [4-1:0] node19836;
	wire [4-1:0] node19838;
	wire [4-1:0] node19841;
	wire [4-1:0] node19842;
	wire [4-1:0] node19843;
	wire [4-1:0] node19847;
	wire [4-1:0] node19850;
	wire [4-1:0] node19851;
	wire [4-1:0] node19852;
	wire [4-1:0] node19856;
	wire [4-1:0] node19857;
	wire [4-1:0] node19858;
	wire [4-1:0] node19862;
	wire [4-1:0] node19865;
	wire [4-1:0] node19866;
	wire [4-1:0] node19867;
	wire [4-1:0] node19868;
	wire [4-1:0] node19869;
	wire [4-1:0] node19872;
	wire [4-1:0] node19876;
	wire [4-1:0] node19877;
	wire [4-1:0] node19878;
	wire [4-1:0] node19879;
	wire [4-1:0] node19882;
	wire [4-1:0] node19885;
	wire [4-1:0] node19886;
	wire [4-1:0] node19891;
	wire [4-1:0] node19892;
	wire [4-1:0] node19893;
	wire [4-1:0] node19894;
	wire [4-1:0] node19897;
	wire [4-1:0] node19898;
	wire [4-1:0] node19903;
	wire [4-1:0] node19904;
	wire [4-1:0] node19905;
	wire [4-1:0] node19909;
	wire [4-1:0] node19910;
	wire [4-1:0] node19914;
	wire [4-1:0] node19915;
	wire [4-1:0] node19916;
	wire [4-1:0] node19917;
	wire [4-1:0] node19918;
	wire [4-1:0] node19919;
	wire [4-1:0] node19920;
	wire [4-1:0] node19921;
	wire [4-1:0] node19922;
	wire [4-1:0] node19923;
	wire [4-1:0] node19926;
	wire [4-1:0] node19929;
	wire [4-1:0] node19930;
	wire [4-1:0] node19931;
	wire [4-1:0] node19934;
	wire [4-1:0] node19937;
	wire [4-1:0] node19938;
	wire [4-1:0] node19941;
	wire [4-1:0] node19944;
	wire [4-1:0] node19945;
	wire [4-1:0] node19946;
	wire [4-1:0] node19949;
	wire [4-1:0] node19952;
	wire [4-1:0] node19953;
	wire [4-1:0] node19954;
	wire [4-1:0] node19957;
	wire [4-1:0] node19961;
	wire [4-1:0] node19962;
	wire [4-1:0] node19963;
	wire [4-1:0] node19964;
	wire [4-1:0] node19965;
	wire [4-1:0] node19969;
	wire [4-1:0] node19970;
	wire [4-1:0] node19971;
	wire [4-1:0] node19974;
	wire [4-1:0] node19977;
	wire [4-1:0] node19978;
	wire [4-1:0] node19982;
	wire [4-1:0] node19983;
	wire [4-1:0] node19984;
	wire [4-1:0] node19985;
	wire [4-1:0] node19988;
	wire [4-1:0] node19992;
	wire [4-1:0] node19993;
	wire [4-1:0] node19996;
	wire [4-1:0] node19999;
	wire [4-1:0] node20000;
	wire [4-1:0] node20001;
	wire [4-1:0] node20002;
	wire [4-1:0] node20005;
	wire [4-1:0] node20009;
	wire [4-1:0] node20010;
	wire [4-1:0] node20011;
	wire [4-1:0] node20014;
	wire [4-1:0] node20018;
	wire [4-1:0] node20019;
	wire [4-1:0] node20020;
	wire [4-1:0] node20021;
	wire [4-1:0] node20022;
	wire [4-1:0] node20023;
	wire [4-1:0] node20026;
	wire [4-1:0] node20029;
	wire [4-1:0] node20030;
	wire [4-1:0] node20033;
	wire [4-1:0] node20036;
	wire [4-1:0] node20037;
	wire [4-1:0] node20038;
	wire [4-1:0] node20042;
	wire [4-1:0] node20044;
	wire [4-1:0] node20045;
	wire [4-1:0] node20048;
	wire [4-1:0] node20051;
	wire [4-1:0] node20052;
	wire [4-1:0] node20053;
	wire [4-1:0] node20054;
	wire [4-1:0] node20055;
	wire [4-1:0] node20059;
	wire [4-1:0] node20061;
	wire [4-1:0] node20064;
	wire [4-1:0] node20065;
	wire [4-1:0] node20068;
	wire [4-1:0] node20071;
	wire [4-1:0] node20072;
	wire [4-1:0] node20073;
	wire [4-1:0] node20074;
	wire [4-1:0] node20077;
	wire [4-1:0] node20081;
	wire [4-1:0] node20082;
	wire [4-1:0] node20083;
	wire [4-1:0] node20087;
	wire [4-1:0] node20090;
	wire [4-1:0] node20091;
	wire [4-1:0] node20092;
	wire [4-1:0] node20093;
	wire [4-1:0] node20094;
	wire [4-1:0] node20097;
	wire [4-1:0] node20100;
	wire [4-1:0] node20101;
	wire [4-1:0] node20102;
	wire [4-1:0] node20106;
	wire [4-1:0] node20107;
	wire [4-1:0] node20111;
	wire [4-1:0] node20112;
	wire [4-1:0] node20113;
	wire [4-1:0] node20116;
	wire [4-1:0] node20119;
	wire [4-1:0] node20120;
	wire [4-1:0] node20121;
	wire [4-1:0] node20124;
	wire [4-1:0] node20127;
	wire [4-1:0] node20128;
	wire [4-1:0] node20131;
	wire [4-1:0] node20134;
	wire [4-1:0] node20135;
	wire [4-1:0] node20136;
	wire [4-1:0] node20137;
	wire [4-1:0] node20138;
	wire [4-1:0] node20142;
	wire [4-1:0] node20143;
	wire [4-1:0] node20146;
	wire [4-1:0] node20149;
	wire [4-1:0] node20151;
	wire [4-1:0] node20152;
	wire [4-1:0] node20156;
	wire [4-1:0] node20157;
	wire [4-1:0] node20159;
	wire [4-1:0] node20160;
	wire [4-1:0] node20163;
	wire [4-1:0] node20166;
	wire [4-1:0] node20167;
	wire [4-1:0] node20170;
	wire [4-1:0] node20173;
	wire [4-1:0] node20174;
	wire [4-1:0] node20175;
	wire [4-1:0] node20176;
	wire [4-1:0] node20177;
	wire [4-1:0] node20178;
	wire [4-1:0] node20181;
	wire [4-1:0] node20184;
	wire [4-1:0] node20185;
	wire [4-1:0] node20188;
	wire [4-1:0] node20191;
	wire [4-1:0] node20192;
	wire [4-1:0] node20193;
	wire [4-1:0] node20194;
	wire [4-1:0] node20197;
	wire [4-1:0] node20200;
	wire [4-1:0] node20201;
	wire [4-1:0] node20204;
	wire [4-1:0] node20207;
	wire [4-1:0] node20208;
	wire [4-1:0] node20209;
	wire [4-1:0] node20212;
	wire [4-1:0] node20215;
	wire [4-1:0] node20216;
	wire [4-1:0] node20219;
	wire [4-1:0] node20222;
	wire [4-1:0] node20223;
	wire [4-1:0] node20224;
	wire [4-1:0] node20225;
	wire [4-1:0] node20226;
	wire [4-1:0] node20229;
	wire [4-1:0] node20232;
	wire [4-1:0] node20233;
	wire [4-1:0] node20236;
	wire [4-1:0] node20239;
	wire [4-1:0] node20240;
	wire [4-1:0] node20241;
	wire [4-1:0] node20243;
	wire [4-1:0] node20246;
	wire [4-1:0] node20247;
	wire [4-1:0] node20250;
	wire [4-1:0] node20253;
	wire [4-1:0] node20254;
	wire [4-1:0] node20257;
	wire [4-1:0] node20260;
	wire [4-1:0] node20261;
	wire [4-1:0] node20262;
	wire [4-1:0] node20263;
	wire [4-1:0] node20266;
	wire [4-1:0] node20269;
	wire [4-1:0] node20270;
	wire [4-1:0] node20272;
	wire [4-1:0] node20275;
	wire [4-1:0] node20276;
	wire [4-1:0] node20279;
	wire [4-1:0] node20282;
	wire [4-1:0] node20283;
	wire [4-1:0] node20284;
	wire [4-1:0] node20288;
	wire [4-1:0] node20289;
	wire [4-1:0] node20291;
	wire [4-1:0] node20294;
	wire [4-1:0] node20296;
	wire [4-1:0] node20299;
	wire [4-1:0] node20300;
	wire [4-1:0] node20301;
	wire [4-1:0] node20302;
	wire [4-1:0] node20303;
	wire [4-1:0] node20306;
	wire [4-1:0] node20308;
	wire [4-1:0] node20311;
	wire [4-1:0] node20312;
	wire [4-1:0] node20315;
	wire [4-1:0] node20316;
	wire [4-1:0] node20319;
	wire [4-1:0] node20322;
	wire [4-1:0] node20323;
	wire [4-1:0] node20324;
	wire [4-1:0] node20325;
	wire [4-1:0] node20328;
	wire [4-1:0] node20332;
	wire [4-1:0] node20333;
	wire [4-1:0] node20334;
	wire [4-1:0] node20337;
	wire [4-1:0] node20340;
	wire [4-1:0] node20341;
	wire [4-1:0] node20344;
	wire [4-1:0] node20347;
	wire [4-1:0] node20348;
	wire [4-1:0] node20349;
	wire [4-1:0] node20350;
	wire [4-1:0] node20353;
	wire [4-1:0] node20354;
	wire [4-1:0] node20357;
	wire [4-1:0] node20360;
	wire [4-1:0] node20361;
	wire [4-1:0] node20363;
	wire [4-1:0] node20366;
	wire [4-1:0] node20367;
	wire [4-1:0] node20370;
	wire [4-1:0] node20373;
	wire [4-1:0] node20374;
	wire [4-1:0] node20375;
	wire [4-1:0] node20378;
	wire [4-1:0] node20380;
	wire [4-1:0] node20383;
	wire [4-1:0] node20384;
	wire [4-1:0] node20385;
	wire [4-1:0] node20388;
	wire [4-1:0] node20391;
	wire [4-1:0] node20392;
	wire [4-1:0] node20395;
	wire [4-1:0] node20398;
	wire [4-1:0] node20399;
	wire [4-1:0] node20400;
	wire [4-1:0] node20401;
	wire [4-1:0] node20402;
	wire [4-1:0] node20403;
	wire [4-1:0] node20404;
	wire [4-1:0] node20405;
	wire [4-1:0] node20409;
	wire [4-1:0] node20410;
	wire [4-1:0] node20413;
	wire [4-1:0] node20416;
	wire [4-1:0] node20417;
	wire [4-1:0] node20418;
	wire [4-1:0] node20419;
	wire [4-1:0] node20423;
	wire [4-1:0] node20425;
	wire [4-1:0] node20428;
	wire [4-1:0] node20429;
	wire [4-1:0] node20432;
	wire [4-1:0] node20435;
	wire [4-1:0] node20436;
	wire [4-1:0] node20437;
	wire [4-1:0] node20438;
	wire [4-1:0] node20442;
	wire [4-1:0] node20445;
	wire [4-1:0] node20446;
	wire [4-1:0] node20447;
	wire [4-1:0] node20448;
	wire [4-1:0] node20452;
	wire [4-1:0] node20453;
	wire [4-1:0] node20456;
	wire [4-1:0] node20459;
	wire [4-1:0] node20460;
	wire [4-1:0] node20463;
	wire [4-1:0] node20466;
	wire [4-1:0] node20467;
	wire [4-1:0] node20468;
	wire [4-1:0] node20469;
	wire [4-1:0] node20472;
	wire [4-1:0] node20475;
	wire [4-1:0] node20476;
	wire [4-1:0] node20479;
	wire [4-1:0] node20480;
	wire [4-1:0] node20483;
	wire [4-1:0] node20486;
	wire [4-1:0] node20487;
	wire [4-1:0] node20488;
	wire [4-1:0] node20489;
	wire [4-1:0] node20492;
	wire [4-1:0] node20495;
	wire [4-1:0] node20497;
	wire [4-1:0] node20500;
	wire [4-1:0] node20501;
	wire [4-1:0] node20502;
	wire [4-1:0] node20503;
	wire [4-1:0] node20506;
	wire [4-1:0] node20509;
	wire [4-1:0] node20510;
	wire [4-1:0] node20514;
	wire [4-1:0] node20516;
	wire [4-1:0] node20517;
	wire [4-1:0] node20520;
	wire [4-1:0] node20523;
	wire [4-1:0] node20524;
	wire [4-1:0] node20525;
	wire [4-1:0] node20526;
	wire [4-1:0] node20529;
	wire [4-1:0] node20530;
	wire [4-1:0] node20531;
	wire [4-1:0] node20532;
	wire [4-1:0] node20535;
	wire [4-1:0] node20539;
	wire [4-1:0] node20540;
	wire [4-1:0] node20541;
	wire [4-1:0] node20544;
	wire [4-1:0] node20548;
	wire [4-1:0] node20549;
	wire [4-1:0] node20550;
	wire [4-1:0] node20552;
	wire [4-1:0] node20553;
	wire [4-1:0] node20557;
	wire [4-1:0] node20560;
	wire [4-1:0] node20561;
	wire [4-1:0] node20562;
	wire [4-1:0] node20565;
	wire [4-1:0] node20568;
	wire [4-1:0] node20570;
	wire [4-1:0] node20573;
	wire [4-1:0] node20574;
	wire [4-1:0] node20575;
	wire [4-1:0] node20576;
	wire [4-1:0] node20579;
	wire [4-1:0] node20582;
	wire [4-1:0] node20583;
	wire [4-1:0] node20586;
	wire [4-1:0] node20587;
	wire [4-1:0] node20590;
	wire [4-1:0] node20593;
	wire [4-1:0] node20594;
	wire [4-1:0] node20595;
	wire [4-1:0] node20596;
	wire [4-1:0] node20599;
	wire [4-1:0] node20602;
	wire [4-1:0] node20603;
	wire [4-1:0] node20606;
	wire [4-1:0] node20609;
	wire [4-1:0] node20610;
	wire [4-1:0] node20611;
	wire [4-1:0] node20612;
	wire [4-1:0] node20615;
	wire [4-1:0] node20618;
	wire [4-1:0] node20620;
	wire [4-1:0] node20623;
	wire [4-1:0] node20624;
	wire [4-1:0] node20625;
	wire [4-1:0] node20628;
	wire [4-1:0] node20632;
	wire [4-1:0] node20633;
	wire [4-1:0] node20634;
	wire [4-1:0] node20635;
	wire [4-1:0] node20636;
	wire [4-1:0] node20637;
	wire [4-1:0] node20638;
	wire [4-1:0] node20641;
	wire [4-1:0] node20644;
	wire [4-1:0] node20645;
	wire [4-1:0] node20649;
	wire [4-1:0] node20650;
	wire [4-1:0] node20651;
	wire [4-1:0] node20655;
	wire [4-1:0] node20656;
	wire [4-1:0] node20660;
	wire [4-1:0] node20661;
	wire [4-1:0] node20662;
	wire [4-1:0] node20664;
	wire [4-1:0] node20667;
	wire [4-1:0] node20670;
	wire [4-1:0] node20671;
	wire [4-1:0] node20672;
	wire [4-1:0] node20675;
	wire [4-1:0] node20678;
	wire [4-1:0] node20679;
	wire [4-1:0] node20682;
	wire [4-1:0] node20685;
	wire [4-1:0] node20686;
	wire [4-1:0] node20687;
	wire [4-1:0] node20688;
	wire [4-1:0] node20690;
	wire [4-1:0] node20693;
	wire [4-1:0] node20694;
	wire [4-1:0] node20698;
	wire [4-1:0] node20699;
	wire [4-1:0] node20700;
	wire [4-1:0] node20703;
	wire [4-1:0] node20706;
	wire [4-1:0] node20708;
	wire [4-1:0] node20711;
	wire [4-1:0] node20712;
	wire [4-1:0] node20713;
	wire [4-1:0] node20715;
	wire [4-1:0] node20718;
	wire [4-1:0] node20720;
	wire [4-1:0] node20723;
	wire [4-1:0] node20724;
	wire [4-1:0] node20725;
	wire [4-1:0] node20728;
	wire [4-1:0] node20731;
	wire [4-1:0] node20732;
	wire [4-1:0] node20736;
	wire [4-1:0] node20737;
	wire [4-1:0] node20738;
	wire [4-1:0] node20739;
	wire [4-1:0] node20741;
	wire [4-1:0] node20743;
	wire [4-1:0] node20744;
	wire [4-1:0] node20747;
	wire [4-1:0] node20750;
	wire [4-1:0] node20751;
	wire [4-1:0] node20752;
	wire [4-1:0] node20755;
	wire [4-1:0] node20758;
	wire [4-1:0] node20759;
	wire [4-1:0] node20762;
	wire [4-1:0] node20765;
	wire [4-1:0] node20766;
	wire [4-1:0] node20767;
	wire [4-1:0] node20768;
	wire [4-1:0] node20771;
	wire [4-1:0] node20774;
	wire [4-1:0] node20775;
	wire [4-1:0] node20778;
	wire [4-1:0] node20781;
	wire [4-1:0] node20782;
	wire [4-1:0] node20783;
	wire [4-1:0] node20785;
	wire [4-1:0] node20788;
	wire [4-1:0] node20791;
	wire [4-1:0] node20792;
	wire [4-1:0] node20795;
	wire [4-1:0] node20798;
	wire [4-1:0] node20799;
	wire [4-1:0] node20800;
	wire [4-1:0] node20801;
	wire [4-1:0] node20802;
	wire [4-1:0] node20805;
	wire [4-1:0] node20808;
	wire [4-1:0] node20809;
	wire [4-1:0] node20812;
	wire [4-1:0] node20815;
	wire [4-1:0] node20816;
	wire [4-1:0] node20817;
	wire [4-1:0] node20820;
	wire [4-1:0] node20823;
	wire [4-1:0] node20824;
	wire [4-1:0] node20827;
	wire [4-1:0] node20830;
	wire [4-1:0] node20831;
	wire [4-1:0] node20832;
	wire [4-1:0] node20834;
	wire [4-1:0] node20837;
	wire [4-1:0] node20838;
	wire [4-1:0] node20842;
	wire [4-1:0] node20843;
	wire [4-1:0] node20845;
	wire [4-1:0] node20846;
	wire [4-1:0] node20849;
	wire [4-1:0] node20852;
	wire [4-1:0] node20853;
	wire [4-1:0] node20854;
	wire [4-1:0] node20857;
	wire [4-1:0] node20861;
	wire [4-1:0] node20862;
	wire [4-1:0] node20863;
	wire [4-1:0] node20864;
	wire [4-1:0] node20865;
	wire [4-1:0] node20866;
	wire [4-1:0] node20867;
	wire [4-1:0] node20868;
	wire [4-1:0] node20871;
	wire [4-1:0] node20874;
	wire [4-1:0] node20875;
	wire [4-1:0] node20879;
	wire [4-1:0] node20880;
	wire [4-1:0] node20881;
	wire [4-1:0] node20884;
	wire [4-1:0] node20887;
	wire [4-1:0] node20888;
	wire [4-1:0] node20892;
	wire [4-1:0] node20893;
	wire [4-1:0] node20894;
	wire [4-1:0] node20895;
	wire [4-1:0] node20898;
	wire [4-1:0] node20901;
	wire [4-1:0] node20902;
	wire [4-1:0] node20905;
	wire [4-1:0] node20908;
	wire [4-1:0] node20909;
	wire [4-1:0] node20910;
	wire [4-1:0] node20913;
	wire [4-1:0] node20916;
	wire [4-1:0] node20919;
	wire [4-1:0] node20920;
	wire [4-1:0] node20921;
	wire [4-1:0] node20922;
	wire [4-1:0] node20925;
	wire [4-1:0] node20927;
	wire [4-1:0] node20930;
	wire [4-1:0] node20931;
	wire [4-1:0] node20934;
	wire [4-1:0] node20935;
	wire [4-1:0] node20938;
	wire [4-1:0] node20941;
	wire [4-1:0] node20942;
	wire [4-1:0] node20943;
	wire [4-1:0] node20946;
	wire [4-1:0] node20947;
	wire [4-1:0] node20951;
	wire [4-1:0] node20953;
	wire [4-1:0] node20956;
	wire [4-1:0] node20957;
	wire [4-1:0] node20958;
	wire [4-1:0] node20959;
	wire [4-1:0] node20962;
	wire [4-1:0] node20963;
	wire [4-1:0] node20965;
	wire [4-1:0] node20968;
	wire [4-1:0] node20970;
	wire [4-1:0] node20973;
	wire [4-1:0] node20974;
	wire [4-1:0] node20975;
	wire [4-1:0] node20978;
	wire [4-1:0] node20979;
	wire [4-1:0] node20982;
	wire [4-1:0] node20985;
	wire [4-1:0] node20986;
	wire [4-1:0] node20989;
	wire [4-1:0] node20991;
	wire [4-1:0] node20994;
	wire [4-1:0] node20995;
	wire [4-1:0] node20996;
	wire [4-1:0] node20999;
	wire [4-1:0] node21000;
	wire [4-1:0] node21002;
	wire [4-1:0] node21005;
	wire [4-1:0] node21006;
	wire [4-1:0] node21009;
	wire [4-1:0] node21012;
	wire [4-1:0] node21013;
	wire [4-1:0] node21014;
	wire [4-1:0] node21017;
	wire [4-1:0] node21018;
	wire [4-1:0] node21021;
	wire [4-1:0] node21024;
	wire [4-1:0] node21025;
	wire [4-1:0] node21028;
	wire [4-1:0] node21030;
	wire [4-1:0] node21033;
	wire [4-1:0] node21034;
	wire [4-1:0] node21035;
	wire [4-1:0] node21036;
	wire [4-1:0] node21037;
	wire [4-1:0] node21038;
	wire [4-1:0] node21039;
	wire [4-1:0] node21041;
	wire [4-1:0] node21044;
	wire [4-1:0] node21045;
	wire [4-1:0] node21048;
	wire [4-1:0] node21051;
	wire [4-1:0] node21052;
	wire [4-1:0] node21054;
	wire [4-1:0] node21055;
	wire [4-1:0] node21058;
	wire [4-1:0] node21061;
	wire [4-1:0] node21062;
	wire [4-1:0] node21065;
	wire [4-1:0] node21067;
	wire [4-1:0] node21070;
	wire [4-1:0] node21071;
	wire [4-1:0] node21072;
	wire [4-1:0] node21073;
	wire [4-1:0] node21074;
	wire [4-1:0] node21078;
	wire [4-1:0] node21081;
	wire [4-1:0] node21082;
	wire [4-1:0] node21083;
	wire [4-1:0] node21086;
	wire [4-1:0] node21089;
	wire [4-1:0] node21090;
	wire [4-1:0] node21093;
	wire [4-1:0] node21096;
	wire [4-1:0] node21097;
	wire [4-1:0] node21100;
	wire [4-1:0] node21101;
	wire [4-1:0] node21105;
	wire [4-1:0] node21106;
	wire [4-1:0] node21107;
	wire [4-1:0] node21108;
	wire [4-1:0] node21109;
	wire [4-1:0] node21110;
	wire [4-1:0] node21114;
	wire [4-1:0] node21115;
	wire [4-1:0] node21119;
	wire [4-1:0] node21120;
	wire [4-1:0] node21121;
	wire [4-1:0] node21125;
	wire [4-1:0] node21126;
	wire [4-1:0] node21129;
	wire [4-1:0] node21132;
	wire [4-1:0] node21133;
	wire [4-1:0] node21134;
	wire [4-1:0] node21135;
	wire [4-1:0] node21139;
	wire [4-1:0] node21142;
	wire [4-1:0] node21143;
	wire [4-1:0] node21144;
	wire [4-1:0] node21148;
	wire [4-1:0] node21149;
	wire [4-1:0] node21153;
	wire [4-1:0] node21154;
	wire [4-1:0] node21155;
	wire [4-1:0] node21156;
	wire [4-1:0] node21157;
	wire [4-1:0] node21160;
	wire [4-1:0] node21164;
	wire [4-1:0] node21165;
	wire [4-1:0] node21166;
	wire [4-1:0] node21169;
	wire [4-1:0] node21173;
	wire [4-1:0] node21174;
	wire [4-1:0] node21175;
	wire [4-1:0] node21176;
	wire [4-1:0] node21179;
	wire [4-1:0] node21182;
	wire [4-1:0] node21185;
	wire [4-1:0] node21186;
	wire [4-1:0] node21187;
	wire [4-1:0] node21191;
	wire [4-1:0] node21192;
	wire [4-1:0] node21196;
	wire [4-1:0] node21197;
	wire [4-1:0] node21198;
	wire [4-1:0] node21199;
	wire [4-1:0] node21200;
	wire [4-1:0] node21201;
	wire [4-1:0] node21203;
	wire [4-1:0] node21208;
	wire [4-1:0] node21209;
	wire [4-1:0] node21210;
	wire [4-1:0] node21213;
	wire [4-1:0] node21216;
	wire [4-1:0] node21218;
	wire [4-1:0] node21221;
	wire [4-1:0] node21222;
	wire [4-1:0] node21223;
	wire [4-1:0] node21226;
	wire [4-1:0] node21229;
	wire [4-1:0] node21230;
	wire [4-1:0] node21233;
	wire [4-1:0] node21234;
	wire [4-1:0] node21238;
	wire [4-1:0] node21239;
	wire [4-1:0] node21240;
	wire [4-1:0] node21241;
	wire [4-1:0] node21243;
	wire [4-1:0] node21246;
	wire [4-1:0] node21249;
	wire [4-1:0] node21250;
	wire [4-1:0] node21251;
	wire [4-1:0] node21254;
	wire [4-1:0] node21257;
	wire [4-1:0] node21258;
	wire [4-1:0] node21261;
	wire [4-1:0] node21264;
	wire [4-1:0] node21265;
	wire [4-1:0] node21268;
	wire [4-1:0] node21269;
	wire [4-1:0] node21272;
	wire [4-1:0] node21275;
	wire [4-1:0] node21276;
	wire [4-1:0] node21277;
	wire [4-1:0] node21278;
	wire [4-1:0] node21279;
	wire [4-1:0] node21280;
	wire [4-1:0] node21281;
	wire [4-1:0] node21284;
	wire [4-1:0] node21287;
	wire [4-1:0] node21288;
	wire [4-1:0] node21291;
	wire [4-1:0] node21294;
	wire [4-1:0] node21295;
	wire [4-1:0] node21298;
	wire [4-1:0] node21301;
	wire [4-1:0] node21302;
	wire [4-1:0] node21303;
	wire [4-1:0] node21304;
	wire [4-1:0] node21307;
	wire [4-1:0] node21310;
	wire [4-1:0] node21311;
	wire [4-1:0] node21312;
	wire [4-1:0] node21317;
	wire [4-1:0] node21318;
	wire [4-1:0] node21319;
	wire [4-1:0] node21322;
	wire [4-1:0] node21325;
	wire [4-1:0] node21326;
	wire [4-1:0] node21329;
	wire [4-1:0] node21332;
	wire [4-1:0] node21333;
	wire [4-1:0] node21334;
	wire [4-1:0] node21335;
	wire [4-1:0] node21337;
	wire [4-1:0] node21338;
	wire [4-1:0] node21341;
	wire [4-1:0] node21344;
	wire [4-1:0] node21345;
	wire [4-1:0] node21347;
	wire [4-1:0] node21350;
	wire [4-1:0] node21351;
	wire [4-1:0] node21354;
	wire [4-1:0] node21357;
	wire [4-1:0] node21358;
	wire [4-1:0] node21359;
	wire [4-1:0] node21360;
	wire [4-1:0] node21363;
	wire [4-1:0] node21366;
	wire [4-1:0] node21367;
	wire [4-1:0] node21371;
	wire [4-1:0] node21373;
	wire [4-1:0] node21376;
	wire [4-1:0] node21377;
	wire [4-1:0] node21380;
	wire [4-1:0] node21381;
	wire [4-1:0] node21382;
	wire [4-1:0] node21385;
	wire [4-1:0] node21388;
	wire [4-1:0] node21389;
	wire [4-1:0] node21392;
	wire [4-1:0] node21395;
	wire [4-1:0] node21396;
	wire [4-1:0] node21397;
	wire [4-1:0] node21398;
	wire [4-1:0] node21399;
	wire [4-1:0] node21400;
	wire [4-1:0] node21402;
	wire [4-1:0] node21406;
	wire [4-1:0] node21407;
	wire [4-1:0] node21410;
	wire [4-1:0] node21413;
	wire [4-1:0] node21416;
	wire [4-1:0] node21417;
	wire [4-1:0] node21420;
	wire [4-1:0] node21423;
	wire [4-1:0] node21424;
	wire [4-1:0] node21425;
	wire [4-1:0] node21426;
	wire [4-1:0] node21429;
	wire [4-1:0] node21432;
	wire [4-1:0] node21433;
	wire [4-1:0] node21434;
	wire [4-1:0] node21435;
	wire [4-1:0] node21439;
	wire [4-1:0] node21441;
	wire [4-1:0] node21444;
	wire [4-1:0] node21445;
	wire [4-1:0] node21448;
	wire [4-1:0] node21451;
	wire [4-1:0] node21452;
	wire [4-1:0] node21455;
	wire [4-1:0] node21458;
	wire [4-1:0] node21459;
	wire [4-1:0] node21460;
	wire [4-1:0] node21461;
	wire [4-1:0] node21462;
	wire [4-1:0] node21463;
	wire [4-1:0] node21464;
	wire [4-1:0] node21465;
	wire [4-1:0] node21467;
	wire [4-1:0] node21470;
	wire [4-1:0] node21471;
	wire [4-1:0] node21474;
	wire [4-1:0] node21477;
	wire [4-1:0] node21478;
	wire [4-1:0] node21479;
	wire [4-1:0] node21482;
	wire [4-1:0] node21485;
	wire [4-1:0] node21486;
	wire [4-1:0] node21489;
	wire [4-1:0] node21492;
	wire [4-1:0] node21493;
	wire [4-1:0] node21494;
	wire [4-1:0] node21496;
	wire [4-1:0] node21499;
	wire [4-1:0] node21500;
	wire [4-1:0] node21503;
	wire [4-1:0] node21506;
	wire [4-1:0] node21507;
	wire [4-1:0] node21509;
	wire [4-1:0] node21512;
	wire [4-1:0] node21513;
	wire [4-1:0] node21516;
	wire [4-1:0] node21519;
	wire [4-1:0] node21520;
	wire [4-1:0] node21521;
	wire [4-1:0] node21522;
	wire [4-1:0] node21525;
	wire [4-1:0] node21526;
	wire [4-1:0] node21529;
	wire [4-1:0] node21532;
	wire [4-1:0] node21533;
	wire [4-1:0] node21534;
	wire [4-1:0] node21537;
	wire [4-1:0] node21540;
	wire [4-1:0] node21541;
	wire [4-1:0] node21544;
	wire [4-1:0] node21547;
	wire [4-1:0] node21548;
	wire [4-1:0] node21549;
	wire [4-1:0] node21551;
	wire [4-1:0] node21554;
	wire [4-1:0] node21556;
	wire [4-1:0] node21559;
	wire [4-1:0] node21560;
	wire [4-1:0] node21561;
	wire [4-1:0] node21564;
	wire [4-1:0] node21567;
	wire [4-1:0] node21568;
	wire [4-1:0] node21571;
	wire [4-1:0] node21574;
	wire [4-1:0] node21575;
	wire [4-1:0] node21576;
	wire [4-1:0] node21577;
	wire [4-1:0] node21578;
	wire [4-1:0] node21579;
	wire [4-1:0] node21582;
	wire [4-1:0] node21585;
	wire [4-1:0] node21586;
	wire [4-1:0] node21589;
	wire [4-1:0] node21592;
	wire [4-1:0] node21593;
	wire [4-1:0] node21594;
	wire [4-1:0] node21595;
	wire [4-1:0] node21599;
	wire [4-1:0] node21600;
	wire [4-1:0] node21601;
	wire [4-1:0] node21604;
	wire [4-1:0] node21607;
	wire [4-1:0] node21608;
	wire [4-1:0] node21611;
	wire [4-1:0] node21614;
	wire [4-1:0] node21617;
	wire [4-1:0] node21618;
	wire [4-1:0] node21620;
	wire [4-1:0] node21623;
	wire [4-1:0] node21625;
	wire [4-1:0] node21628;
	wire [4-1:0] node21629;
	wire [4-1:0] node21630;
	wire [4-1:0] node21631;
	wire [4-1:0] node21632;
	wire [4-1:0] node21635;
	wire [4-1:0] node21638;
	wire [4-1:0] node21639;
	wire [4-1:0] node21640;
	wire [4-1:0] node21643;
	wire [4-1:0] node21646;
	wire [4-1:0] node21647;
	wire [4-1:0] node21651;
	wire [4-1:0] node21652;
	wire [4-1:0] node21653;
	wire [4-1:0] node21654;
	wire [4-1:0] node21657;
	wire [4-1:0] node21660;
	wire [4-1:0] node21662;
	wire [4-1:0] node21665;
	wire [4-1:0] node21666;
	wire [4-1:0] node21669;
	wire [4-1:0] node21672;
	wire [4-1:0] node21673;
	wire [4-1:0] node21674;
	wire [4-1:0] node21677;
	wire [4-1:0] node21678;
	wire [4-1:0] node21679;
	wire [4-1:0] node21682;
	wire [4-1:0] node21685;
	wire [4-1:0] node21686;
	wire [4-1:0] node21689;
	wire [4-1:0] node21692;
	wire [4-1:0] node21693;
	wire [4-1:0] node21694;
	wire [4-1:0] node21695;
	wire [4-1:0] node21696;
	wire [4-1:0] node21699;
	wire [4-1:0] node21702;
	wire [4-1:0] node21703;
	wire [4-1:0] node21706;
	wire [4-1:0] node21709;
	wire [4-1:0] node21710;
	wire [4-1:0] node21711;
	wire [4-1:0] node21714;
	wire [4-1:0] node21717;
	wire [4-1:0] node21718;
	wire [4-1:0] node21722;
	wire [4-1:0] node21723;
	wire [4-1:0] node21724;
	wire [4-1:0] node21725;
	wire [4-1:0] node21729;
	wire [4-1:0] node21731;
	wire [4-1:0] node21734;
	wire [4-1:0] node21735;
	wire [4-1:0] node21737;
	wire [4-1:0] node21741;
	wire [4-1:0] node21742;
	wire [4-1:0] node21743;
	wire [4-1:0] node21744;
	wire [4-1:0] node21745;
	wire [4-1:0] node21746;
	wire [4-1:0] node21747;
	wire [4-1:0] node21748;
	wire [4-1:0] node21752;
	wire [4-1:0] node21753;
	wire [4-1:0] node21757;
	wire [4-1:0] node21758;
	wire [4-1:0] node21760;
	wire [4-1:0] node21763;
	wire [4-1:0] node21766;
	wire [4-1:0] node21767;
	wire [4-1:0] node21768;
	wire [4-1:0] node21770;
	wire [4-1:0] node21773;
	wire [4-1:0] node21774;
	wire [4-1:0] node21778;
	wire [4-1:0] node21781;
	wire [4-1:0] node21782;
	wire [4-1:0] node21783;
	wire [4-1:0] node21784;
	wire [4-1:0] node21787;
	wire [4-1:0] node21788;
	wire [4-1:0] node21791;
	wire [4-1:0] node21794;
	wire [4-1:0] node21795;
	wire [4-1:0] node21796;
	wire [4-1:0] node21799;
	wire [4-1:0] node21802;
	wire [4-1:0] node21803;
	wire [4-1:0] node21806;
	wire [4-1:0] node21809;
	wire [4-1:0] node21810;
	wire [4-1:0] node21811;
	wire [4-1:0] node21813;
	wire [4-1:0] node21816;
	wire [4-1:0] node21817;
	wire [4-1:0] node21820;
	wire [4-1:0] node21823;
	wire [4-1:0] node21824;
	wire [4-1:0] node21826;
	wire [4-1:0] node21829;
	wire [4-1:0] node21830;
	wire [4-1:0] node21833;
	wire [4-1:0] node21836;
	wire [4-1:0] node21837;
	wire [4-1:0] node21838;
	wire [4-1:0] node21839;
	wire [4-1:0] node21840;
	wire [4-1:0] node21841;
	wire [4-1:0] node21845;
	wire [4-1:0] node21846;
	wire [4-1:0] node21849;
	wire [4-1:0] node21852;
	wire [4-1:0] node21853;
	wire [4-1:0] node21854;
	wire [4-1:0] node21857;
	wire [4-1:0] node21860;
	wire [4-1:0] node21863;
	wire [4-1:0] node21864;
	wire [4-1:0] node21865;
	wire [4-1:0] node21866;
	wire [4-1:0] node21869;
	wire [4-1:0] node21872;
	wire [4-1:0] node21873;
	wire [4-1:0] node21876;
	wire [4-1:0] node21879;
	wire [4-1:0] node21880;
	wire [4-1:0] node21882;
	wire [4-1:0] node21885;
	wire [4-1:0] node21886;
	wire [4-1:0] node21889;
	wire [4-1:0] node21892;
	wire [4-1:0] node21893;
	wire [4-1:0] node21894;
	wire [4-1:0] node21895;
	wire [4-1:0] node21896;
	wire [4-1:0] node21899;
	wire [4-1:0] node21902;
	wire [4-1:0] node21904;
	wire [4-1:0] node21907;
	wire [4-1:0] node21908;
	wire [4-1:0] node21910;
	wire [4-1:0] node21913;
	wire [4-1:0] node21916;
	wire [4-1:0] node21917;
	wire [4-1:0] node21919;
	wire [4-1:0] node21920;
	wire [4-1:0] node21924;
	wire [4-1:0] node21925;
	wire [4-1:0] node21928;
	wire [4-1:0] node21931;
	wire [4-1:0] node21932;
	wire [4-1:0] node21933;
	wire [4-1:0] node21934;
	wire [4-1:0] node21935;
	wire [4-1:0] node21936;
	wire [4-1:0] node21937;
	wire [4-1:0] node21940;
	wire [4-1:0] node21943;
	wire [4-1:0] node21944;
	wire [4-1:0] node21946;
	wire [4-1:0] node21949;
	wire [4-1:0] node21950;
	wire [4-1:0] node21953;
	wire [4-1:0] node21956;
	wire [4-1:0] node21957;
	wire [4-1:0] node21958;
	wire [4-1:0] node21960;
	wire [4-1:0] node21963;
	wire [4-1:0] node21965;
	wire [4-1:0] node21968;
	wire [4-1:0] node21969;
	wire [4-1:0] node21970;
	wire [4-1:0] node21973;
	wire [4-1:0] node21976;
	wire [4-1:0] node21977;
	wire [4-1:0] node21980;
	wire [4-1:0] node21983;
	wire [4-1:0] node21984;
	wire [4-1:0] node21985;
	wire [4-1:0] node21986;
	wire [4-1:0] node21990;
	wire [4-1:0] node21991;
	wire [4-1:0] node21994;
	wire [4-1:0] node21997;
	wire [4-1:0] node21998;
	wire [4-1:0] node21999;
	wire [4-1:0] node22002;
	wire [4-1:0] node22005;
	wire [4-1:0] node22006;
	wire [4-1:0] node22009;
	wire [4-1:0] node22012;
	wire [4-1:0] node22013;
	wire [4-1:0] node22014;
	wire [4-1:0] node22015;
	wire [4-1:0] node22018;
	wire [4-1:0] node22021;
	wire [4-1:0] node22022;
	wire [4-1:0] node22023;
	wire [4-1:0] node22025;
	wire [4-1:0] node22028;
	wire [4-1:0] node22029;
	wire [4-1:0] node22032;
	wire [4-1:0] node22035;
	wire [4-1:0] node22036;
	wire [4-1:0] node22040;
	wire [4-1:0] node22041;
	wire [4-1:0] node22042;
	wire [4-1:0] node22043;
	wire [4-1:0] node22044;
	wire [4-1:0] node22047;
	wire [4-1:0] node22050;
	wire [4-1:0] node22051;
	wire [4-1:0] node22054;
	wire [4-1:0] node22057;
	wire [4-1:0] node22058;
	wire [4-1:0] node22059;
	wire [4-1:0] node22063;
	wire [4-1:0] node22064;
	wire [4-1:0] node22067;
	wire [4-1:0] node22070;
	wire [4-1:0] node22071;
	wire [4-1:0] node22072;
	wire [4-1:0] node22076;
	wire [4-1:0] node22077;
	wire [4-1:0] node22078;
	wire [4-1:0] node22081;
	wire [4-1:0] node22084;
	wire [4-1:0] node22085;
	wire [4-1:0] node22088;
	wire [4-1:0] node22091;
	wire [4-1:0] node22092;
	wire [4-1:0] node22093;
	wire [4-1:0] node22094;
	wire [4-1:0] node22095;
	wire [4-1:0] node22096;
	wire [4-1:0] node22099;
	wire [4-1:0] node22102;
	wire [4-1:0] node22105;
	wire [4-1:0] node22106;
	wire [4-1:0] node22107;
	wire [4-1:0] node22111;
	wire [4-1:0] node22112;
	wire [4-1:0] node22116;
	wire [4-1:0] node22117;
	wire [4-1:0] node22118;
	wire [4-1:0] node22120;
	wire [4-1:0] node22123;
	wire [4-1:0] node22124;
	wire [4-1:0] node22127;
	wire [4-1:0] node22130;
	wire [4-1:0] node22131;
	wire [4-1:0] node22133;
	wire [4-1:0] node22136;
	wire [4-1:0] node22137;
	wire [4-1:0] node22140;
	wire [4-1:0] node22143;
	wire [4-1:0] node22144;
	wire [4-1:0] node22145;
	wire [4-1:0] node22146;
	wire [4-1:0] node22147;
	wire [4-1:0] node22150;
	wire [4-1:0] node22153;
	wire [4-1:0] node22154;
	wire [4-1:0] node22158;
	wire [4-1:0] node22159;
	wire [4-1:0] node22160;
	wire [4-1:0] node22164;
	wire [4-1:0] node22165;
	wire [4-1:0] node22168;
	wire [4-1:0] node22171;
	wire [4-1:0] node22172;
	wire [4-1:0] node22173;
	wire [4-1:0] node22175;
	wire [4-1:0] node22178;
	wire [4-1:0] node22179;
	wire [4-1:0] node22182;
	wire [4-1:0] node22185;
	wire [4-1:0] node22186;
	wire [4-1:0] node22187;
	wire [4-1:0] node22191;
	wire [4-1:0] node22194;
	wire [4-1:0] node22195;
	wire [4-1:0] node22196;
	wire [4-1:0] node22197;
	wire [4-1:0] node22198;
	wire [4-1:0] node22199;
	wire [4-1:0] node22200;
	wire [4-1:0] node22201;
	wire [4-1:0] node22204;
	wire [4-1:0] node22207;
	wire [4-1:0] node22208;
	wire [4-1:0] node22209;
	wire [4-1:0] node22213;
	wire [4-1:0] node22216;
	wire [4-1:0] node22217;
	wire [4-1:0] node22218;
	wire [4-1:0] node22219;
	wire [4-1:0] node22222;
	wire [4-1:0] node22225;
	wire [4-1:0] node22228;
	wire [4-1:0] node22229;
	wire [4-1:0] node22230;
	wire [4-1:0] node22233;
	wire [4-1:0] node22236;
	wire [4-1:0] node22237;
	wire [4-1:0] node22240;
	wire [4-1:0] node22243;
	wire [4-1:0] node22244;
	wire [4-1:0] node22245;
	wire [4-1:0] node22246;
	wire [4-1:0] node22249;
	wire [4-1:0] node22252;
	wire [4-1:0] node22253;
	wire [4-1:0] node22254;
	wire [4-1:0] node22258;
	wire [4-1:0] node22261;
	wire [4-1:0] node22262;
	wire [4-1:0] node22263;
	wire [4-1:0] node22264;
	wire [4-1:0] node22267;
	wire [4-1:0] node22270;
	wire [4-1:0] node22273;
	wire [4-1:0] node22274;
	wire [4-1:0] node22275;
	wire [4-1:0] node22279;
	wire [4-1:0] node22282;
	wire [4-1:0] node22283;
	wire [4-1:0] node22284;
	wire [4-1:0] node22285;
	wire [4-1:0] node22286;
	wire [4-1:0] node22287;
	wire [4-1:0] node22290;
	wire [4-1:0] node22293;
	wire [4-1:0] node22294;
	wire [4-1:0] node22297;
	wire [4-1:0] node22300;
	wire [4-1:0] node22301;
	wire [4-1:0] node22302;
	wire [4-1:0] node22306;
	wire [4-1:0] node22307;
	wire [4-1:0] node22310;
	wire [4-1:0] node22313;
	wire [4-1:0] node22314;
	wire [4-1:0] node22315;
	wire [4-1:0] node22317;
	wire [4-1:0] node22320;
	wire [4-1:0] node22323;
	wire [4-1:0] node22324;
	wire [4-1:0] node22327;
	wire [4-1:0] node22330;
	wire [4-1:0] node22331;
	wire [4-1:0] node22332;
	wire [4-1:0] node22333;
	wire [4-1:0] node22334;
	wire [4-1:0] node22335;
	wire [4-1:0] node22338;
	wire [4-1:0] node22341;
	wire [4-1:0] node22342;
	wire [4-1:0] node22345;
	wire [4-1:0] node22348;
	wire [4-1:0] node22349;
	wire [4-1:0] node22350;
	wire [4-1:0] node22353;
	wire [4-1:0] node22357;
	wire [4-1:0] node22359;
	wire [4-1:0] node22360;
	wire [4-1:0] node22361;
	wire [4-1:0] node22364;
	wire [4-1:0] node22368;
	wire [4-1:0] node22369;
	wire [4-1:0] node22370;
	wire [4-1:0] node22373;
	wire [4-1:0] node22376;
	wire [4-1:0] node22377;
	wire [4-1:0] node22378;
	wire [4-1:0] node22381;
	wire [4-1:0] node22384;
	wire [4-1:0] node22385;
	wire [4-1:0] node22388;
	wire [4-1:0] node22391;
	wire [4-1:0] node22392;
	wire [4-1:0] node22393;
	wire [4-1:0] node22394;
	wire [4-1:0] node22395;
	wire [4-1:0] node22396;
	wire [4-1:0] node22397;
	wire [4-1:0] node22398;
	wire [4-1:0] node22401;
	wire [4-1:0] node22404;
	wire [4-1:0] node22405;
	wire [4-1:0] node22408;
	wire [4-1:0] node22411;
	wire [4-1:0] node22413;
	wire [4-1:0] node22414;
	wire [4-1:0] node22417;
	wire [4-1:0] node22420;
	wire [4-1:0] node22421;
	wire [4-1:0] node22422;
	wire [4-1:0] node22423;
	wire [4-1:0] node22426;
	wire [4-1:0] node22429;
	wire [4-1:0] node22430;
	wire [4-1:0] node22434;
	wire [4-1:0] node22435;
	wire [4-1:0] node22438;
	wire [4-1:0] node22439;
	wire [4-1:0] node22443;
	wire [4-1:0] node22444;
	wire [4-1:0] node22445;
	wire [4-1:0] node22447;
	wire [4-1:0] node22450;
	wire [4-1:0] node22451;
	wire [4-1:0] node22452;
	wire [4-1:0] node22455;
	wire [4-1:0] node22459;
	wire [4-1:0] node22460;
	wire [4-1:0] node22461;
	wire [4-1:0] node22465;
	wire [4-1:0] node22466;
	wire [4-1:0] node22470;
	wire [4-1:0] node22471;
	wire [4-1:0] node22472;
	wire [4-1:0] node22473;
	wire [4-1:0] node22474;
	wire [4-1:0] node22476;
	wire [4-1:0] node22479;
	wire [4-1:0] node22482;
	wire [4-1:0] node22483;
	wire [4-1:0] node22484;
	wire [4-1:0] node22489;
	wire [4-1:0] node22490;
	wire [4-1:0] node22491;
	wire [4-1:0] node22494;
	wire [4-1:0] node22496;
	wire [4-1:0] node22499;
	wire [4-1:0] node22500;
	wire [4-1:0] node22501;
	wire [4-1:0] node22505;
	wire [4-1:0] node22507;
	wire [4-1:0] node22510;
	wire [4-1:0] node22511;
	wire [4-1:0] node22512;
	wire [4-1:0] node22513;
	wire [4-1:0] node22516;
	wire [4-1:0] node22519;
	wire [4-1:0] node22520;
	wire [4-1:0] node22522;
	wire [4-1:0] node22525;
	wire [4-1:0] node22526;
	wire [4-1:0] node22530;
	wire [4-1:0] node22531;
	wire [4-1:0] node22532;
	wire [4-1:0] node22533;
	wire [4-1:0] node22536;
	wire [4-1:0] node22539;
	wire [4-1:0] node22542;
	wire [4-1:0] node22543;
	wire [4-1:0] node22544;
	wire [4-1:0] node22547;
	wire [4-1:0] node22550;
	wire [4-1:0] node22551;
	wire [4-1:0] node22554;
	wire [4-1:0] node22557;
	wire [4-1:0] node22558;
	wire [4-1:0] node22559;
	wire [4-1:0] node22560;
	wire [4-1:0] node22561;
	wire [4-1:0] node22562;
	wire [4-1:0] node22565;
	wire [4-1:0] node22568;
	wire [4-1:0] node22569;
	wire [4-1:0] node22570;
	wire [4-1:0] node22573;
	wire [4-1:0] node22577;
	wire [4-1:0] node22578;
	wire [4-1:0] node22579;
	wire [4-1:0] node22583;
	wire [4-1:0] node22586;
	wire [4-1:0] node22587;
	wire [4-1:0] node22588;
	wire [4-1:0] node22589;
	wire [4-1:0] node22592;
	wire [4-1:0] node22595;
	wire [4-1:0] node22597;
	wire [4-1:0] node22600;
	wire [4-1:0] node22601;
	wire [4-1:0] node22605;
	wire [4-1:0] node22606;
	wire [4-1:0] node22607;
	wire [4-1:0] node22608;
	wire [4-1:0] node22609;
	wire [4-1:0] node22612;
	wire [4-1:0] node22616;
	wire [4-1:0] node22617;
	wire [4-1:0] node22618;
	wire [4-1:0] node22621;
	wire [4-1:0] node22624;
	wire [4-1:0] node22627;
	wire [4-1:0] node22628;
	wire [4-1:0] node22629;
	wire [4-1:0] node22632;
	wire [4-1:0] node22633;
	wire [4-1:0] node22636;
	wire [4-1:0] node22639;
	wire [4-1:0] node22640;
	wire [4-1:0] node22642;
	wire [4-1:0] node22645;
	wire [4-1:0] node22646;
	wire [4-1:0] node22650;
	wire [4-1:0] node22651;
	wire [4-1:0] node22652;
	wire [4-1:0] node22653;
	wire [4-1:0] node22654;
	wire [4-1:0] node22655;
	wire [4-1:0] node22656;
	wire [4-1:0] node22657;
	wire [4-1:0] node22658;
	wire [4-1:0] node22661;
	wire [4-1:0] node22665;
	wire [4-1:0] node22666;
	wire [4-1:0] node22667;
	wire [4-1:0] node22670;
	wire [4-1:0] node22674;
	wire [4-1:0] node22675;
	wire [4-1:0] node22676;
	wire [4-1:0] node22679;
	wire [4-1:0] node22682;
	wire [4-1:0] node22683;
	wire [4-1:0] node22684;
	wire [4-1:0] node22687;
	wire [4-1:0] node22690;
	wire [4-1:0] node22691;
	wire [4-1:0] node22695;
	wire [4-1:0] node22696;
	wire [4-1:0] node22697;
	wire [4-1:0] node22699;
	wire [4-1:0] node22700;
	wire [4-1:0] node22704;
	wire [4-1:0] node22705;
	wire [4-1:0] node22708;
	wire [4-1:0] node22711;
	wire [4-1:0] node22712;
	wire [4-1:0] node22714;
	wire [4-1:0] node22717;
	wire [4-1:0] node22718;
	wire [4-1:0] node22721;
	wire [4-1:0] node22722;
	wire [4-1:0] node22726;
	wire [4-1:0] node22727;
	wire [4-1:0] node22728;
	wire [4-1:0] node22729;
	wire [4-1:0] node22733;
	wire [4-1:0] node22734;
	wire [4-1:0] node22737;
	wire [4-1:0] node22740;
	wire [4-1:0] node22741;
	wire [4-1:0] node22742;
	wire [4-1:0] node22743;
	wire [4-1:0] node22744;
	wire [4-1:0] node22747;
	wire [4-1:0] node22750;
	wire [4-1:0] node22751;
	wire [4-1:0] node22754;
	wire [4-1:0] node22757;
	wire [4-1:0] node22758;
	wire [4-1:0] node22759;
	wire [4-1:0] node22762;
	wire [4-1:0] node22766;
	wire [4-1:0] node22767;
	wire [4-1:0] node22768;
	wire [4-1:0] node22771;
	wire [4-1:0] node22774;
	wire [4-1:0] node22776;
	wire [4-1:0] node22779;
	wire [4-1:0] node22780;
	wire [4-1:0] node22781;
	wire [4-1:0] node22782;
	wire [4-1:0] node22783;
	wire [4-1:0] node22784;
	wire [4-1:0] node22786;
	wire [4-1:0] node22789;
	wire [4-1:0] node22790;
	wire [4-1:0] node22793;
	wire [4-1:0] node22796;
	wire [4-1:0] node22798;
	wire [4-1:0] node22799;
	wire [4-1:0] node22802;
	wire [4-1:0] node22805;
	wire [4-1:0] node22806;
	wire [4-1:0] node22807;
	wire [4-1:0] node22810;
	wire [4-1:0] node22813;
	wire [4-1:0] node22815;
	wire [4-1:0] node22818;
	wire [4-1:0] node22819;
	wire [4-1:0] node22820;
	wire [4-1:0] node22821;
	wire [4-1:0] node22824;
	wire [4-1:0] node22827;
	wire [4-1:0] node22828;
	wire [4-1:0] node22832;
	wire [4-1:0] node22833;
	wire [4-1:0] node22834;
	wire [4-1:0] node22837;
	wire [4-1:0] node22840;
	wire [4-1:0] node22841;
	wire [4-1:0] node22845;
	wire [4-1:0] node22846;
	wire [4-1:0] node22847;
	wire [4-1:0] node22848;
	wire [4-1:0] node22850;
	wire [4-1:0] node22851;
	wire [4-1:0] node22854;
	wire [4-1:0] node22857;
	wire [4-1:0] node22858;
	wire [4-1:0] node22861;
	wire [4-1:0] node22864;
	wire [4-1:0] node22865;
	wire [4-1:0] node22867;
	wire [4-1:0] node22870;
	wire [4-1:0] node22871;
	wire [4-1:0] node22874;
	wire [4-1:0] node22877;
	wire [4-1:0] node22878;
	wire [4-1:0] node22879;
	wire [4-1:0] node22880;
	wire [4-1:0] node22882;
	wire [4-1:0] node22885;
	wire [4-1:0] node22888;
	wire [4-1:0] node22889;
	wire [4-1:0] node22892;
	wire [4-1:0] node22895;
	wire [4-1:0] node22896;
	wire [4-1:0] node22898;
	wire [4-1:0] node22901;
	wire [4-1:0] node22902;
	wire [4-1:0] node22904;
	wire [4-1:0] node22907;
	wire [4-1:0] node22908;
	wire [4-1:0] node22911;
	wire [4-1:0] node22914;
	wire [4-1:0] node22915;
	wire [4-1:0] node22916;
	wire [4-1:0] node22917;
	wire [4-1:0] node22918;
	wire [4-1:0] node22919;
	wire [4-1:0] node22920;
	wire [4-1:0] node22923;
	wire [4-1:0] node22924;
	wire [4-1:0] node22928;
	wire [4-1:0] node22929;
	wire [4-1:0] node22930;
	wire [4-1:0] node22933;
	wire [4-1:0] node22936;
	wire [4-1:0] node22937;
	wire [4-1:0] node22940;
	wire [4-1:0] node22943;
	wire [4-1:0] node22944;
	wire [4-1:0] node22948;
	wire [4-1:0] node22949;
	wire [4-1:0] node22950;
	wire [4-1:0] node22953;
	wire [4-1:0] node22956;
	wire [4-1:0] node22957;
	wire [4-1:0] node22960;
	wire [4-1:0] node22963;
	wire [4-1:0] node22964;
	wire [4-1:0] node22965;
	wire [4-1:0] node22966;
	wire [4-1:0] node22969;
	wire [4-1:0] node22972;
	wire [4-1:0] node22973;
	wire [4-1:0] node22976;
	wire [4-1:0] node22979;
	wire [4-1:0] node22980;
	wire [4-1:0] node22983;
	wire [4-1:0] node22986;
	wire [4-1:0] node22987;
	wire [4-1:0] node22988;
	wire [4-1:0] node22989;
	wire [4-1:0] node22990;
	wire [4-1:0] node22991;
	wire [4-1:0] node22994;
	wire [4-1:0] node22997;
	wire [4-1:0] node22998;
	wire [4-1:0] node22999;
	wire [4-1:0] node23002;
	wire [4-1:0] node23006;
	wire [4-1:0] node23007;
	wire [4-1:0] node23008;
	wire [4-1:0] node23011;
	wire [4-1:0] node23014;
	wire [4-1:0] node23015;
	wire [4-1:0] node23018;
	wire [4-1:0] node23021;
	wire [4-1:0] node23022;
	wire [4-1:0] node23023;
	wire [4-1:0] node23024;
	wire [4-1:0] node23028;
	wire [4-1:0] node23029;
	wire [4-1:0] node23032;
	wire [4-1:0] node23035;
	wire [4-1:0] node23036;
	wire [4-1:0] node23037;
	wire [4-1:0] node23040;
	wire [4-1:0] node23043;
	wire [4-1:0] node23044;
	wire [4-1:0] node23047;
	wire [4-1:0] node23050;
	wire [4-1:0] node23051;
	wire [4-1:0] node23052;
	wire [4-1:0] node23054;
	wire [4-1:0] node23055;
	wire [4-1:0] node23058;
	wire [4-1:0] node23061;
	wire [4-1:0] node23062;
	wire [4-1:0] node23063;
	wire [4-1:0] node23064;
	wire [4-1:0] node23068;
	wire [4-1:0] node23069;
	wire [4-1:0] node23072;
	wire [4-1:0] node23075;
	wire [4-1:0] node23076;
	wire [4-1:0] node23078;
	wire [4-1:0] node23081;
	wire [4-1:0] node23082;
	wire [4-1:0] node23086;
	wire [4-1:0] node23087;
	wire [4-1:0] node23088;
	wire [4-1:0] node23091;
	wire [4-1:0] node23094;
	wire [4-1:0] node23096;
	wire [4-1:0] node23099;
	wire [4-1:0] node23100;
	wire [4-1:0] node23101;
	wire [4-1:0] node23102;
	wire [4-1:0] node23103;
	wire [4-1:0] node23104;
	wire [4-1:0] node23105;
	wire [4-1:0] node23106;
	wire [4-1:0] node23107;
	wire [4-1:0] node23109;
	wire [4-1:0] node23112;
	wire [4-1:0] node23114;
	wire [4-1:0] node23117;
	wire [4-1:0] node23118;
	wire [4-1:0] node23120;
	wire [4-1:0] node23123;
	wire [4-1:0] node23125;
	wire [4-1:0] node23128;
	wire [4-1:0] node23129;
	wire [4-1:0] node23130;
	wire [4-1:0] node23131;
	wire [4-1:0] node23132;
	wire [4-1:0] node23136;
	wire [4-1:0] node23137;
	wire [4-1:0] node23138;
	wire [4-1:0] node23139;
	wire [4-1:0] node23142;
	wire [4-1:0] node23145;
	wire [4-1:0] node23146;
	wire [4-1:0] node23149;
	wire [4-1:0] node23152;
	wire [4-1:0] node23154;
	wire [4-1:0] node23157;
	wire [4-1:0] node23158;
	wire [4-1:0] node23159;
	wire [4-1:0] node23161;
	wire [4-1:0] node23164;
	wire [4-1:0] node23167;
	wire [4-1:0] node23168;
	wire [4-1:0] node23171;
	wire [4-1:0] node23173;
	wire [4-1:0] node23176;
	wire [4-1:0] node23177;
	wire [4-1:0] node23178;
	wire [4-1:0] node23179;
	wire [4-1:0] node23182;
	wire [4-1:0] node23185;
	wire [4-1:0] node23186;
	wire [4-1:0] node23189;
	wire [4-1:0] node23192;
	wire [4-1:0] node23193;
	wire [4-1:0] node23194;
	wire [4-1:0] node23195;
	wire [4-1:0] node23198;
	wire [4-1:0] node23201;
	wire [4-1:0] node23202;
	wire [4-1:0] node23205;
	wire [4-1:0] node23208;
	wire [4-1:0] node23210;
	wire [4-1:0] node23211;
	wire [4-1:0] node23214;
	wire [4-1:0] node23217;
	wire [4-1:0] node23218;
	wire [4-1:0] node23219;
	wire [4-1:0] node23220;
	wire [4-1:0] node23221;
	wire [4-1:0] node23222;
	wire [4-1:0] node23225;
	wire [4-1:0] node23228;
	wire [4-1:0] node23229;
	wire [4-1:0] node23231;
	wire [4-1:0] node23234;
	wire [4-1:0] node23235;
	wire [4-1:0] node23238;
	wire [4-1:0] node23241;
	wire [4-1:0] node23242;
	wire [4-1:0] node23243;
	wire [4-1:0] node23246;
	wire [4-1:0] node23249;
	wire [4-1:0] node23250;
	wire [4-1:0] node23251;
	wire [4-1:0] node23255;
	wire [4-1:0] node23256;
	wire [4-1:0] node23259;
	wire [4-1:0] node23262;
	wire [4-1:0] node23263;
	wire [4-1:0] node23264;
	wire [4-1:0] node23265;
	wire [4-1:0] node23266;
	wire [4-1:0] node23269;
	wire [4-1:0] node23272;
	wire [4-1:0] node23274;
	wire [4-1:0] node23277;
	wire [4-1:0] node23278;
	wire [4-1:0] node23280;
	wire [4-1:0] node23283;
	wire [4-1:0] node23284;
	wire [4-1:0] node23286;
	wire [4-1:0] node23289;
	wire [4-1:0] node23290;
	wire [4-1:0] node23293;
	wire [4-1:0] node23296;
	wire [4-1:0] node23297;
	wire [4-1:0] node23298;
	wire [4-1:0] node23299;
	wire [4-1:0] node23302;
	wire [4-1:0] node23305;
	wire [4-1:0] node23306;
	wire [4-1:0] node23310;
	wire [4-1:0] node23311;
	wire [4-1:0] node23312;
	wire [4-1:0] node23315;
	wire [4-1:0] node23318;
	wire [4-1:0] node23320;
	wire [4-1:0] node23321;
	wire [4-1:0] node23324;
	wire [4-1:0] node23327;
	wire [4-1:0] node23328;
	wire [4-1:0] node23329;
	wire [4-1:0] node23330;
	wire [4-1:0] node23331;
	wire [4-1:0] node23332;
	wire [4-1:0] node23335;
	wire [4-1:0] node23338;
	wire [4-1:0] node23339;
	wire [4-1:0] node23342;
	wire [4-1:0] node23345;
	wire [4-1:0] node23346;
	wire [4-1:0] node23348;
	wire [4-1:0] node23351;
	wire [4-1:0] node23352;
	wire [4-1:0] node23353;
	wire [4-1:0] node23358;
	wire [4-1:0] node23359;
	wire [4-1:0] node23360;
	wire [4-1:0] node23361;
	wire [4-1:0] node23364;
	wire [4-1:0] node23367;
	wire [4-1:0] node23368;
	wire [4-1:0] node23371;
	wire [4-1:0] node23374;
	wire [4-1:0] node23375;
	wire [4-1:0] node23377;
	wire [4-1:0] node23380;
	wire [4-1:0] node23381;
	wire [4-1:0] node23385;
	wire [4-1:0] node23386;
	wire [4-1:0] node23387;
	wire [4-1:0] node23388;
	wire [4-1:0] node23392;
	wire [4-1:0] node23393;
	wire [4-1:0] node23397;
	wire [4-1:0] node23398;
	wire [4-1:0] node23399;
	wire [4-1:0] node23403;
	wire [4-1:0] node23404;
	wire [4-1:0] node23408;
	wire [4-1:0] node23409;
	wire [4-1:0] node23410;
	wire [4-1:0] node23411;
	wire [4-1:0] node23412;
	wire [4-1:0] node23413;
	wire [4-1:0] node23414;
	wire [4-1:0] node23415;
	wire [4-1:0] node23417;
	wire [4-1:0] node23420;
	wire [4-1:0] node23421;
	wire [4-1:0] node23424;
	wire [4-1:0] node23427;
	wire [4-1:0] node23428;
	wire [4-1:0] node23432;
	wire [4-1:0] node23433;
	wire [4-1:0] node23435;
	wire [4-1:0] node23438;
	wire [4-1:0] node23439;
	wire [4-1:0] node23442;
	wire [4-1:0] node23445;
	wire [4-1:0] node23446;
	wire [4-1:0] node23447;
	wire [4-1:0] node23448;
	wire [4-1:0] node23451;
	wire [4-1:0] node23454;
	wire [4-1:0] node23455;
	wire [4-1:0] node23457;
	wire [4-1:0] node23460;
	wire [4-1:0] node23461;
	wire [4-1:0] node23464;
	wire [4-1:0] node23467;
	wire [4-1:0] node23468;
	wire [4-1:0] node23469;
	wire [4-1:0] node23471;
	wire [4-1:0] node23474;
	wire [4-1:0] node23476;
	wire [4-1:0] node23479;
	wire [4-1:0] node23481;
	wire [4-1:0] node23484;
	wire [4-1:0] node23485;
	wire [4-1:0] node23486;
	wire [4-1:0] node23487;
	wire [4-1:0] node23490;
	wire [4-1:0] node23493;
	wire [4-1:0] node23494;
	wire [4-1:0] node23497;
	wire [4-1:0] node23500;
	wire [4-1:0] node23501;
	wire [4-1:0] node23502;
	wire [4-1:0] node23505;
	wire [4-1:0] node23508;
	wire [4-1:0] node23509;
	wire [4-1:0] node23512;
	wire [4-1:0] node23515;
	wire [4-1:0] node23516;
	wire [4-1:0] node23517;
	wire [4-1:0] node23518;
	wire [4-1:0] node23519;
	wire [4-1:0] node23520;
	wire [4-1:0] node23522;
	wire [4-1:0] node23525;
	wire [4-1:0] node23526;
	wire [4-1:0] node23530;
	wire [4-1:0] node23531;
	wire [4-1:0] node23532;
	wire [4-1:0] node23535;
	wire [4-1:0] node23538;
	wire [4-1:0] node23539;
	wire [4-1:0] node23542;
	wire [4-1:0] node23545;
	wire [4-1:0] node23546;
	wire [4-1:0] node23549;
	wire [4-1:0] node23552;
	wire [4-1:0] node23553;
	wire [4-1:0] node23554;
	wire [4-1:0] node23556;
	wire [4-1:0] node23557;
	wire [4-1:0] node23560;
	wire [4-1:0] node23563;
	wire [4-1:0] node23564;
	wire [4-1:0] node23567;
	wire [4-1:0] node23570;
	wire [4-1:0] node23571;
	wire [4-1:0] node23572;
	wire [4-1:0] node23574;
	wire [4-1:0] node23577;
	wire [4-1:0] node23580;
	wire [4-1:0] node23581;
	wire [4-1:0] node23582;
	wire [4-1:0] node23585;
	wire [4-1:0] node23588;
	wire [4-1:0] node23589;
	wire [4-1:0] node23592;
	wire [4-1:0] node23595;
	wire [4-1:0] node23596;
	wire [4-1:0] node23597;
	wire [4-1:0] node23598;
	wire [4-1:0] node23599;
	wire [4-1:0] node23600;
	wire [4-1:0] node23603;
	wire [4-1:0] node23606;
	wire [4-1:0] node23607;
	wire [4-1:0] node23611;
	wire [4-1:0] node23613;
	wire [4-1:0] node23614;
	wire [4-1:0] node23617;
	wire [4-1:0] node23620;
	wire [4-1:0] node23621;
	wire [4-1:0] node23622;
	wire [4-1:0] node23625;
	wire [4-1:0] node23628;
	wire [4-1:0] node23629;
	wire [4-1:0] node23632;
	wire [4-1:0] node23635;
	wire [4-1:0] node23636;
	wire [4-1:0] node23639;
	wire [4-1:0] node23642;
	wire [4-1:0] node23643;
	wire [4-1:0] node23644;
	wire [4-1:0] node23645;
	wire [4-1:0] node23646;
	wire [4-1:0] node23647;
	wire [4-1:0] node23648;
	wire [4-1:0] node23650;
	wire [4-1:0] node23653;
	wire [4-1:0] node23654;
	wire [4-1:0] node23658;
	wire [4-1:0] node23660;
	wire [4-1:0] node23663;
	wire [4-1:0] node23664;
	wire [4-1:0] node23665;
	wire [4-1:0] node23668;
	wire [4-1:0] node23671;
	wire [4-1:0] node23672;
	wire [4-1:0] node23673;
	wire [4-1:0] node23676;
	wire [4-1:0] node23680;
	wire [4-1:0] node23681;
	wire [4-1:0] node23682;
	wire [4-1:0] node23686;
	wire [4-1:0] node23687;
	wire [4-1:0] node23690;
	wire [4-1:0] node23693;
	wire [4-1:0] node23694;
	wire [4-1:0] node23695;
	wire [4-1:0] node23696;
	wire [4-1:0] node23699;
	wire [4-1:0] node23702;
	wire [4-1:0] node23703;
	wire [4-1:0] node23706;
	wire [4-1:0] node23709;
	wire [4-1:0] node23710;
	wire [4-1:0] node23713;
	wire [4-1:0] node23716;
	wire [4-1:0] node23717;
	wire [4-1:0] node23718;
	wire [4-1:0] node23719;
	wire [4-1:0] node23720;
	wire [4-1:0] node23722;
	wire [4-1:0] node23725;
	wire [4-1:0] node23727;
	wire [4-1:0] node23730;
	wire [4-1:0] node23731;
	wire [4-1:0] node23732;
	wire [4-1:0] node23734;
	wire [4-1:0] node23737;
	wire [4-1:0] node23739;
	wire [4-1:0] node23742;
	wire [4-1:0] node23744;
	wire [4-1:0] node23747;
	wire [4-1:0] node23748;
	wire [4-1:0] node23749;
	wire [4-1:0] node23751;
	wire [4-1:0] node23752;
	wire [4-1:0] node23755;
	wire [4-1:0] node23758;
	wire [4-1:0] node23759;
	wire [4-1:0] node23760;
	wire [4-1:0] node23764;
	wire [4-1:0] node23765;
	wire [4-1:0] node23769;
	wire [4-1:0] node23770;
	wire [4-1:0] node23771;
	wire [4-1:0] node23772;
	wire [4-1:0] node23776;
	wire [4-1:0] node23777;
	wire [4-1:0] node23780;
	wire [4-1:0] node23783;
	wire [4-1:0] node23784;
	wire [4-1:0] node23785;
	wire [4-1:0] node23788;
	wire [4-1:0] node23791;
	wire [4-1:0] node23792;
	wire [4-1:0] node23795;
	wire [4-1:0] node23798;
	wire [4-1:0] node23799;
	wire [4-1:0] node23800;
	wire [4-1:0] node23801;
	wire [4-1:0] node23804;
	wire [4-1:0] node23807;
	wire [4-1:0] node23808;
	wire [4-1:0] node23811;
	wire [4-1:0] node23814;
	wire [4-1:0] node23815;
	wire [4-1:0] node23816;
	wire [4-1:0] node23819;
	wire [4-1:0] node23822;
	wire [4-1:0] node23823;
	wire [4-1:0] node23826;
	wire [4-1:0] node23829;
	wire [4-1:0] node23830;
	wire [4-1:0] node23831;
	wire [4-1:0] node23832;
	wire [4-1:0] node23833;
	wire [4-1:0] node23834;
	wire [4-1:0] node23837;
	wire [4-1:0] node23838;
	wire [4-1:0] node23840;
	wire [4-1:0] node23843;
	wire [4-1:0] node23844;
	wire [4-1:0] node23848;
	wire [4-1:0] node23849;
	wire [4-1:0] node23850;
	wire [4-1:0] node23851;
	wire [4-1:0] node23854;
	wire [4-1:0] node23857;
	wire [4-1:0] node23858;
	wire [4-1:0] node23859;
	wire [4-1:0] node23863;
	wire [4-1:0] node23864;
	wire [4-1:0] node23867;
	wire [4-1:0] node23870;
	wire [4-1:0] node23871;
	wire [4-1:0] node23872;
	wire [4-1:0] node23876;
	wire [4-1:0] node23877;
	wire [4-1:0] node23881;
	wire [4-1:0] node23882;
	wire [4-1:0] node23883;
	wire [4-1:0] node23886;
	wire [4-1:0] node23887;
	wire [4-1:0] node23889;
	wire [4-1:0] node23892;
	wire [4-1:0] node23893;
	wire [4-1:0] node23897;
	wire [4-1:0] node23898;
	wire [4-1:0] node23899;
	wire [4-1:0] node23900;
	wire [4-1:0] node23902;
	wire [4-1:0] node23903;
	wire [4-1:0] node23906;
	wire [4-1:0] node23909;
	wire [4-1:0] node23910;
	wire [4-1:0] node23911;
	wire [4-1:0] node23914;
	wire [4-1:0] node23917;
	wire [4-1:0] node23919;
	wire [4-1:0] node23922;
	wire [4-1:0] node23923;
	wire [4-1:0] node23926;
	wire [4-1:0] node23929;
	wire [4-1:0] node23930;
	wire [4-1:0] node23931;
	wire [4-1:0] node23935;
	wire [4-1:0] node23936;
	wire [4-1:0] node23940;
	wire [4-1:0] node23941;
	wire [4-1:0] node23942;
	wire [4-1:0] node23943;
	wire [4-1:0] node23946;
	wire [4-1:0] node23947;
	wire [4-1:0] node23949;
	wire [4-1:0] node23952;
	wire [4-1:0] node23953;
	wire [4-1:0] node23957;
	wire [4-1:0] node23958;
	wire [4-1:0] node23959;
	wire [4-1:0] node23960;
	wire [4-1:0] node23961;
	wire [4-1:0] node23964;
	wire [4-1:0] node23967;
	wire [4-1:0] node23968;
	wire [4-1:0] node23971;
	wire [4-1:0] node23974;
	wire [4-1:0] node23975;
	wire [4-1:0] node23977;
	wire [4-1:0] node23980;
	wire [4-1:0] node23981;
	wire [4-1:0] node23982;
	wire [4-1:0] node23986;
	wire [4-1:0] node23987;
	wire [4-1:0] node23991;
	wire [4-1:0] node23992;
	wire [4-1:0] node23994;
	wire [4-1:0] node23997;
	wire [4-1:0] node23999;
	wire [4-1:0] node24002;
	wire [4-1:0] node24003;
	wire [4-1:0] node24004;
	wire [4-1:0] node24007;
	wire [4-1:0] node24008;
	wire [4-1:0] node24011;
	wire [4-1:0] node24012;
	wire [4-1:0] node24016;
	wire [4-1:0] node24017;
	wire [4-1:0] node24018;
	wire [4-1:0] node24019;
	wire [4-1:0] node24020;
	wire [4-1:0] node24023;
	wire [4-1:0] node24026;
	wire [4-1:0] node24027;
	wire [4-1:0] node24031;
	wire [4-1:0] node24032;
	wire [4-1:0] node24036;
	wire [4-1:0] node24037;
	wire [4-1:0] node24038;
	wire [4-1:0] node24041;
	wire [4-1:0] node24044;
	wire [4-1:0] node24045;
	wire [4-1:0] node24049;
	wire [4-1:0] node24050;
	wire [4-1:0] node24051;
	wire [4-1:0] node24052;
	wire [4-1:0] node24053;
	wire [4-1:0] node24056;
	wire [4-1:0] node24057;
	wire [4-1:0] node24059;
	wire [4-1:0] node24062;
	wire [4-1:0] node24063;
	wire [4-1:0] node24067;
	wire [4-1:0] node24068;
	wire [4-1:0] node24069;
	wire [4-1:0] node24070;
	wire [4-1:0] node24073;
	wire [4-1:0] node24076;
	wire [4-1:0] node24077;
	wire [4-1:0] node24078;
	wire [4-1:0] node24081;
	wire [4-1:0] node24084;
	wire [4-1:0] node24085;
	wire [4-1:0] node24086;
	wire [4-1:0] node24089;
	wire [4-1:0] node24093;
	wire [4-1:0] node24094;
	wire [4-1:0] node24096;
	wire [4-1:0] node24099;
	wire [4-1:0] node24100;
	wire [4-1:0] node24104;
	wire [4-1:0] node24105;
	wire [4-1:0] node24106;
	wire [4-1:0] node24109;
	wire [4-1:0] node24110;
	wire [4-1:0] node24112;
	wire [4-1:0] node24115;
	wire [4-1:0] node24116;
	wire [4-1:0] node24120;
	wire [4-1:0] node24121;
	wire [4-1:0] node24122;
	wire [4-1:0] node24123;
	wire [4-1:0] node24126;
	wire [4-1:0] node24129;
	wire [4-1:0] node24130;
	wire [4-1:0] node24133;
	wire [4-1:0] node24136;
	wire [4-1:0] node24137;
	wire [4-1:0] node24140;
	wire [4-1:0] node24141;
	wire [4-1:0] node24145;
	wire [4-1:0] node24146;
	wire [4-1:0] node24147;
	wire [4-1:0] node24148;
	wire [4-1:0] node24151;
	wire [4-1:0] node24152;
	wire [4-1:0] node24154;
	wire [4-1:0] node24157;
	wire [4-1:0] node24158;
	wire [4-1:0] node24162;
	wire [4-1:0] node24163;
	wire [4-1:0] node24164;
	wire [4-1:0] node24165;
	wire [4-1:0] node24168;
	wire [4-1:0] node24171;
	wire [4-1:0] node24173;
	wire [4-1:0] node24176;
	wire [4-1:0] node24177;
	wire [4-1:0] node24179;
	wire [4-1:0] node24182;
	wire [4-1:0] node24184;
	wire [4-1:0] node24187;
	wire [4-1:0] node24188;
	wire [4-1:0] node24189;
	wire [4-1:0] node24192;
	wire [4-1:0] node24193;
	wire [4-1:0] node24195;
	wire [4-1:0] node24198;
	wire [4-1:0] node24199;
	wire [4-1:0] node24203;
	wire [4-1:0] node24204;
	wire [4-1:0] node24205;
	wire [4-1:0] node24206;
	wire [4-1:0] node24207;
	wire [4-1:0] node24211;
	wire [4-1:0] node24212;
	wire [4-1:0] node24215;
	wire [4-1:0] node24218;
	wire [4-1:0] node24219;
	wire [4-1:0] node24222;
	wire [4-1:0] node24225;
	wire [4-1:0] node24226;
	wire [4-1:0] node24227;
	wire [4-1:0] node24231;
	wire [4-1:0] node24233;
	wire [4-1:0] node24236;
	wire [4-1:0] node24237;
	wire [4-1:0] node24238;
	wire [4-1:0] node24239;
	wire [4-1:0] node24240;
	wire [4-1:0] node24241;
	wire [4-1:0] node24242;
	wire [4-1:0] node24243;
	wire [4-1:0] node24247;
	wire [4-1:0] node24249;
	wire [4-1:0] node24252;
	wire [4-1:0] node24253;
	wire [4-1:0] node24255;
	wire [4-1:0] node24258;
	wire [4-1:0] node24260;
	wire [4-1:0] node24263;
	wire [4-1:0] node24264;
	wire [4-1:0] node24265;
	wire [4-1:0] node24266;
	wire [4-1:0] node24267;
	wire [4-1:0] node24269;
	wire [4-1:0] node24272;
	wire [4-1:0] node24274;
	wire [4-1:0] node24277;
	wire [4-1:0] node24278;
	wire [4-1:0] node24281;
	wire [4-1:0] node24282;
	wire [4-1:0] node24286;
	wire [4-1:0] node24287;
	wire [4-1:0] node24288;
	wire [4-1:0] node24290;
	wire [4-1:0] node24293;
	wire [4-1:0] node24294;
	wire [4-1:0] node24298;
	wire [4-1:0] node24300;
	wire [4-1:0] node24303;
	wire [4-1:0] node24304;
	wire [4-1:0] node24305;
	wire [4-1:0] node24308;
	wire [4-1:0] node24311;
	wire [4-1:0] node24312;
	wire [4-1:0] node24314;
	wire [4-1:0] node24315;
	wire [4-1:0] node24318;
	wire [4-1:0] node24321;
	wire [4-1:0] node24322;
	wire [4-1:0] node24323;
	wire [4-1:0] node24326;
	wire [4-1:0] node24329;
	wire [4-1:0] node24331;
	wire [4-1:0] node24334;
	wire [4-1:0] node24335;
	wire [4-1:0] node24336;
	wire [4-1:0] node24337;
	wire [4-1:0] node24338;
	wire [4-1:0] node24339;
	wire [4-1:0] node24342;
	wire [4-1:0] node24345;
	wire [4-1:0] node24346;
	wire [4-1:0] node24349;
	wire [4-1:0] node24352;
	wire [4-1:0] node24353;
	wire [4-1:0] node24354;
	wire [4-1:0] node24355;
	wire [4-1:0] node24359;
	wire [4-1:0] node24360;
	wire [4-1:0] node24362;
	wire [4-1:0] node24366;
	wire [4-1:0] node24368;
	wire [4-1:0] node24371;
	wire [4-1:0] node24372;
	wire [4-1:0] node24375;
	wire [4-1:0] node24378;
	wire [4-1:0] node24379;
	wire [4-1:0] node24380;
	wire [4-1:0] node24381;
	wire [4-1:0] node24384;
	wire [4-1:0] node24387;
	wire [4-1:0] node24388;
	wire [4-1:0] node24389;
	wire [4-1:0] node24392;
	wire [4-1:0] node24395;
	wire [4-1:0] node24396;
	wire [4-1:0] node24399;
	wire [4-1:0] node24400;
	wire [4-1:0] node24403;
	wire [4-1:0] node24406;
	wire [4-1:0] node24407;
	wire [4-1:0] node24408;
	wire [4-1:0] node24409;
	wire [4-1:0] node24410;
	wire [4-1:0] node24414;
	wire [4-1:0] node24416;
	wire [4-1:0] node24419;
	wire [4-1:0] node24420;
	wire [4-1:0] node24423;
	wire [4-1:0] node24426;
	wire [4-1:0] node24427;
	wire [4-1:0] node24428;
	wire [4-1:0] node24429;
	wire [4-1:0] node24432;
	wire [4-1:0] node24435;
	wire [4-1:0] node24436;
	wire [4-1:0] node24439;
	wire [4-1:0] node24442;
	wire [4-1:0] node24443;
	wire [4-1:0] node24445;
	wire [4-1:0] node24446;
	wire [4-1:0] node24449;
	wire [4-1:0] node24452;
	wire [4-1:0] node24454;
	wire [4-1:0] node24455;
	wire [4-1:0] node24458;
	wire [4-1:0] node24461;
	wire [4-1:0] node24462;
	wire [4-1:0] node24463;
	wire [4-1:0] node24464;
	wire [4-1:0] node24465;
	wire [4-1:0] node24466;
	wire [4-1:0] node24467;
	wire [4-1:0] node24471;
	wire [4-1:0] node24472;
	wire [4-1:0] node24476;
	wire [4-1:0] node24477;
	wire [4-1:0] node24479;
	wire [4-1:0] node24482;
	wire [4-1:0] node24483;
	wire [4-1:0] node24487;
	wire [4-1:0] node24488;
	wire [4-1:0] node24489;
	wire [4-1:0] node24490;
	wire [4-1:0] node24492;
	wire [4-1:0] node24495;
	wire [4-1:0] node24496;
	wire [4-1:0] node24499;
	wire [4-1:0] node24502;
	wire [4-1:0] node24503;
	wire [4-1:0] node24504;
	wire [4-1:0] node24507;
	wire [4-1:0] node24510;
	wire [4-1:0] node24511;
	wire [4-1:0] node24512;
	wire [4-1:0] node24516;
	wire [4-1:0] node24517;
	wire [4-1:0] node24520;
	wire [4-1:0] node24523;
	wire [4-1:0] node24524;
	wire [4-1:0] node24525;
	wire [4-1:0] node24527;
	wire [4-1:0] node24528;
	wire [4-1:0] node24532;
	wire [4-1:0] node24533;
	wire [4-1:0] node24534;
	wire [4-1:0] node24537;
	wire [4-1:0] node24540;
	wire [4-1:0] node24542;
	wire [4-1:0] node24545;
	wire [4-1:0] node24546;
	wire [4-1:0] node24547;
	wire [4-1:0] node24551;
	wire [4-1:0] node24552;
	wire [4-1:0] node24556;
	wire [4-1:0] node24557;
	wire [4-1:0] node24558;
	wire [4-1:0] node24559;
	wire [4-1:0] node24563;
	wire [4-1:0] node24565;
	wire [4-1:0] node24568;
	wire [4-1:0] node24569;
	wire [4-1:0] node24571;
	wire [4-1:0] node24574;
	wire [4-1:0] node24576;
	wire [4-1:0] node24579;
	wire [4-1:0] node24580;
	wire [4-1:0] node24581;
	wire [4-1:0] node24582;
	wire [4-1:0] node24583;
	wire [4-1:0] node24584;
	wire [4-1:0] node24585;
	wire [4-1:0] node24589;
	wire [4-1:0] node24590;
	wire [4-1:0] node24593;
	wire [4-1:0] node24596;
	wire [4-1:0] node24597;
	wire [4-1:0] node24599;
	wire [4-1:0] node24602;
	wire [4-1:0] node24604;
	wire [4-1:0] node24605;
	wire [4-1:0] node24608;
	wire [4-1:0] node24611;
	wire [4-1:0] node24612;
	wire [4-1:0] node24613;
	wire [4-1:0] node24616;
	wire [4-1:0] node24619;
	wire [4-1:0] node24620;
	wire [4-1:0] node24621;
	wire [4-1:0] node24622;
	wire [4-1:0] node24626;
	wire [4-1:0] node24627;
	wire [4-1:0] node24630;
	wire [4-1:0] node24633;
	wire [4-1:0] node24634;
	wire [4-1:0] node24637;
	wire [4-1:0] node24640;
	wire [4-1:0] node24641;
	wire [4-1:0] node24642;
	wire [4-1:0] node24643;
	wire [4-1:0] node24645;
	wire [4-1:0] node24646;
	wire [4-1:0] node24650;
	wire [4-1:0] node24651;
	wire [4-1:0] node24654;
	wire [4-1:0] node24657;
	wire [4-1:0] node24658;
	wire [4-1:0] node24659;
	wire [4-1:0] node24660;
	wire [4-1:0] node24664;
	wire [4-1:0] node24667;
	wire [4-1:0] node24669;
	wire [4-1:0] node24670;
	wire [4-1:0] node24674;
	wire [4-1:0] node24675;
	wire [4-1:0] node24676;
	wire [4-1:0] node24677;
	wire [4-1:0] node24681;
	wire [4-1:0] node24683;
	wire [4-1:0] node24686;
	wire [4-1:0] node24687;
	wire [4-1:0] node24689;
	wire [4-1:0] node24692;
	wire [4-1:0] node24693;
	wire [4-1:0] node24697;
	wire [4-1:0] node24698;
	wire [4-1:0] node24699;
	wire [4-1:0] node24700;
	wire [4-1:0] node24702;
	wire [4-1:0] node24703;
	wire [4-1:0] node24704;
	wire [4-1:0] node24707;
	wire [4-1:0] node24711;
	wire [4-1:0] node24712;
	wire [4-1:0] node24713;
	wire [4-1:0] node24716;
	wire [4-1:0] node24719;
	wire [4-1:0] node24720;
	wire [4-1:0] node24721;
	wire [4-1:0] node24724;
	wire [4-1:0] node24727;
	wire [4-1:0] node24729;
	wire [4-1:0] node24732;
	wire [4-1:0] node24733;
	wire [4-1:0] node24734;
	wire [4-1:0] node24735;
	wire [4-1:0] node24737;
	wire [4-1:0] node24740;
	wire [4-1:0] node24741;
	wire [4-1:0] node24744;
	wire [4-1:0] node24747;
	wire [4-1:0] node24749;
	wire [4-1:0] node24750;
	wire [4-1:0] node24753;
	wire [4-1:0] node24756;
	wire [4-1:0] node24758;
	wire [4-1:0] node24759;
	wire [4-1:0] node24760;
	wire [4-1:0] node24763;
	wire [4-1:0] node24766;
	wire [4-1:0] node24767;
	wire [4-1:0] node24770;
	wire [4-1:0] node24773;
	wire [4-1:0] node24774;
	wire [4-1:0] node24775;
	wire [4-1:0] node24776;
	wire [4-1:0] node24779;
	wire [4-1:0] node24782;
	wire [4-1:0] node24783;
	wire [4-1:0] node24785;
	wire [4-1:0] node24786;
	wire [4-1:0] node24789;
	wire [4-1:0] node24792;
	wire [4-1:0] node24793;
	wire [4-1:0] node24796;
	wire [4-1:0] node24799;
	wire [4-1:0] node24800;
	wire [4-1:0] node24801;
	wire [4-1:0] node24802;
	wire [4-1:0] node24805;
	wire [4-1:0] node24808;
	wire [4-1:0] node24809;
	wire [4-1:0] node24810;
	wire [4-1:0] node24813;
	wire [4-1:0] node24816;
	wire [4-1:0] node24817;
	wire [4-1:0] node24820;
	wire [4-1:0] node24823;
	wire [4-1:0] node24824;
	wire [4-1:0] node24825;
	wire [4-1:0] node24828;
	wire [4-1:0] node24831;
	wire [4-1:0] node24832;
	wire [4-1:0] node24835;
	wire [4-1:0] node24838;
	wire [4-1:0] node24839;
	wire [4-1:0] node24840;
	wire [4-1:0] node24841;
	wire [4-1:0] node24842;
	wire [4-1:0] node24843;
	wire [4-1:0] node24844;
	wire [4-1:0] node24845;
	wire [4-1:0] node24846;
	wire [4-1:0] node24847;
	wire [4-1:0] node24851;
	wire [4-1:0] node24853;
	wire [4-1:0] node24856;
	wire [4-1:0] node24857;
	wire [4-1:0] node24858;
	wire [4-1:0] node24862;
	wire [4-1:0] node24865;
	wire [4-1:0] node24867;
	wire [4-1:0] node24868;
	wire [4-1:0] node24870;
	wire [4-1:0] node24873;
	wire [4-1:0] node24876;
	wire [4-1:0] node24877;
	wire [4-1:0] node24878;
	wire [4-1:0] node24879;
	wire [4-1:0] node24881;
	wire [4-1:0] node24884;
	wire [4-1:0] node24886;
	wire [4-1:0] node24889;
	wire [4-1:0] node24890;
	wire [4-1:0] node24893;
	wire [4-1:0] node24896;
	wire [4-1:0] node24897;
	wire [4-1:0] node24898;
	wire [4-1:0] node24901;
	wire [4-1:0] node24904;
	wire [4-1:0] node24905;
	wire [4-1:0] node24908;
	wire [4-1:0] node24911;
	wire [4-1:0] node24912;
	wire [4-1:0] node24913;
	wire [4-1:0] node24914;
	wire [4-1:0] node24915;
	wire [4-1:0] node24916;
	wire [4-1:0] node24919;
	wire [4-1:0] node24922;
	wire [4-1:0] node24924;
	wire [4-1:0] node24927;
	wire [4-1:0] node24928;
	wire [4-1:0] node24931;
	wire [4-1:0] node24934;
	wire [4-1:0] node24935;
	wire [4-1:0] node24936;
	wire [4-1:0] node24937;
	wire [4-1:0] node24942;
	wire [4-1:0] node24943;
	wire [4-1:0] node24946;
	wire [4-1:0] node24949;
	wire [4-1:0] node24950;
	wire [4-1:0] node24951;
	wire [4-1:0] node24952;
	wire [4-1:0] node24953;
	wire [4-1:0] node24957;
	wire [4-1:0] node24958;
	wire [4-1:0] node24962;
	wire [4-1:0] node24963;
	wire [4-1:0] node24966;
	wire [4-1:0] node24969;
	wire [4-1:0] node24970;
	wire [4-1:0] node24971;
	wire [4-1:0] node24974;
	wire [4-1:0] node24978;
	wire [4-1:0] node24979;
	wire [4-1:0] node24980;
	wire [4-1:0] node24981;
	wire [4-1:0] node24983;
	wire [4-1:0] node24986;
	wire [4-1:0] node24988;
	wire [4-1:0] node24991;
	wire [4-1:0] node24992;
	wire [4-1:0] node24994;
	wire [4-1:0] node24997;
	wire [4-1:0] node24999;
	wire [4-1:0] node25002;
	wire [4-1:0] node25003;
	wire [4-1:0] node25004;
	wire [4-1:0] node25006;
	wire [4-1:0] node25009;
	wire [4-1:0] node25011;
	wire [4-1:0] node25014;
	wire [4-1:0] node25015;
	wire [4-1:0] node25017;
	wire [4-1:0] node25020;
	wire [4-1:0] node25022;
	wire [4-1:0] node25025;
	wire [4-1:0] node25026;
	wire [4-1:0] node25027;
	wire [4-1:0] node25028;
	wire [4-1:0] node25029;
	wire [4-1:0] node25030;
	wire [4-1:0] node25031;
	wire [4-1:0] node25035;
	wire [4-1:0] node25036;
	wire [4-1:0] node25039;
	wire [4-1:0] node25042;
	wire [4-1:0] node25043;
	wire [4-1:0] node25044;
	wire [4-1:0] node25045;
	wire [4-1:0] node25049;
	wire [4-1:0] node25051;
	wire [4-1:0] node25054;
	wire [4-1:0] node25055;
	wire [4-1:0] node25058;
	wire [4-1:0] node25061;
	wire [4-1:0] node25062;
	wire [4-1:0] node25063;
	wire [4-1:0] node25066;
	wire [4-1:0] node25069;
	wire [4-1:0] node25070;
	wire [4-1:0] node25071;
	wire [4-1:0] node25072;
	wire [4-1:0] node25076;
	wire [4-1:0] node25077;
	wire [4-1:0] node25080;
	wire [4-1:0] node25083;
	wire [4-1:0] node25084;
	wire [4-1:0] node25087;
	wire [4-1:0] node25090;
	wire [4-1:0] node25091;
	wire [4-1:0] node25092;
	wire [4-1:0] node25094;
	wire [4-1:0] node25097;
	wire [4-1:0] node25098;
	wire [4-1:0] node25102;
	wire [4-1:0] node25103;
	wire [4-1:0] node25105;
	wire [4-1:0] node25108;
	wire [4-1:0] node25110;
	wire [4-1:0] node25113;
	wire [4-1:0] node25114;
	wire [4-1:0] node25115;
	wire [4-1:0] node25116;
	wire [4-1:0] node25120;
	wire [4-1:0] node25121;
	wire [4-1:0] node25125;
	wire [4-1:0] node25126;
	wire [4-1:0] node25127;
	wire [4-1:0] node25131;
	wire [4-1:0] node25132;
	wire [4-1:0] node25136;
	wire [4-1:0] node25137;
	wire [4-1:0] node25138;
	wire [4-1:0] node25139;
	wire [4-1:0] node25140;
	wire [4-1:0] node25141;
	wire [4-1:0] node25142;
	wire [4-1:0] node25143;
	wire [4-1:0] node25145;
	wire [4-1:0] node25148;
	wire [4-1:0] node25149;
	wire [4-1:0] node25152;
	wire [4-1:0] node25155;
	wire [4-1:0] node25156;
	wire [4-1:0] node25159;
	wire [4-1:0] node25162;
	wire [4-1:0] node25164;
	wire [4-1:0] node25165;
	wire [4-1:0] node25166;
	wire [4-1:0] node25169;
	wire [4-1:0] node25173;
	wire [4-1:0] node25174;
	wire [4-1:0] node25175;
	wire [4-1:0] node25178;
	wire [4-1:0] node25181;
	wire [4-1:0] node25182;
	wire [4-1:0] node25183;
	wire [4-1:0] node25184;
	wire [4-1:0] node25187;
	wire [4-1:0] node25190;
	wire [4-1:0] node25191;
	wire [4-1:0] node25194;
	wire [4-1:0] node25197;
	wire [4-1:0] node25199;
	wire [4-1:0] node25200;
	wire [4-1:0] node25203;
	wire [4-1:0] node25206;
	wire [4-1:0] node25207;
	wire [4-1:0] node25208;
	wire [4-1:0] node25209;
	wire [4-1:0] node25212;
	wire [4-1:0] node25215;
	wire [4-1:0] node25216;
	wire [4-1:0] node25217;
	wire [4-1:0] node25220;
	wire [4-1:0] node25223;
	wire [4-1:0] node25224;
	wire [4-1:0] node25227;
	wire [4-1:0] node25230;
	wire [4-1:0] node25231;
	wire [4-1:0] node25232;
	wire [4-1:0] node25233;
	wire [4-1:0] node25234;
	wire [4-1:0] node25238;
	wire [4-1:0] node25239;
	wire [4-1:0] node25242;
	wire [4-1:0] node25245;
	wire [4-1:0] node25246;
	wire [4-1:0] node25250;
	wire [4-1:0] node25251;
	wire [4-1:0] node25252;
	wire [4-1:0] node25253;
	wire [4-1:0] node25258;
	wire [4-1:0] node25260;
	wire [4-1:0] node25261;
	wire [4-1:0] node25265;
	wire [4-1:0] node25266;
	wire [4-1:0] node25267;
	wire [4-1:0] node25268;
	wire [4-1:0] node25270;
	wire [4-1:0] node25273;
	wire [4-1:0] node25275;
	wire [4-1:0] node25278;
	wire [4-1:0] node25279;
	wire [4-1:0] node25280;
	wire [4-1:0] node25284;
	wire [4-1:0] node25286;
	wire [4-1:0] node25289;
	wire [4-1:0] node25290;
	wire [4-1:0] node25291;
	wire [4-1:0] node25292;
	wire [4-1:0] node25296;
	wire [4-1:0] node25297;
	wire [4-1:0] node25301;
	wire [4-1:0] node25302;
	wire [4-1:0] node25303;
	wire [4-1:0] node25307;
	wire [4-1:0] node25308;
	wire [4-1:0] node25312;
	wire [4-1:0] node25313;
	wire [4-1:0] node25314;
	wire [4-1:0] node25315;
	wire [4-1:0] node25317;
	wire [4-1:0] node25320;
	wire [4-1:0] node25323;
	wire [4-1:0] node25324;
	wire [4-1:0] node25325;
	wire [4-1:0] node25329;
	wire [4-1:0] node25332;
	wire [4-1:0] node25333;
	wire [4-1:0] node25334;
	wire [4-1:0] node25335;
	wire [4-1:0] node25340;
	wire [4-1:0] node25341;
	wire [4-1:0] node25342;
	wire [4-1:0] node25347;
	wire [4-1:0] node25348;
	wire [4-1:0] node25349;
	wire [4-1:0] node25350;
	wire [4-1:0] node25351;
	wire [4-1:0] node25352;
	wire [4-1:0] node25353;
	wire [4-1:0] node25354;
	wire [4-1:0] node25355;
	wire [4-1:0] node25356;
	wire [4-1:0] node25357;
	wire [4-1:0] node25358;
	wire [4-1:0] node25361;
	wire [4-1:0] node25365;
	wire [4-1:0] node25366;
	wire [4-1:0] node25368;
	wire [4-1:0] node25371;
	wire [4-1:0] node25372;
	wire [4-1:0] node25375;
	wire [4-1:0] node25378;
	wire [4-1:0] node25379;
	wire [4-1:0] node25382;
	wire [4-1:0] node25385;
	wire [4-1:0] node25386;
	wire [4-1:0] node25387;
	wire [4-1:0] node25391;
	wire [4-1:0] node25392;
	wire [4-1:0] node25395;
	wire [4-1:0] node25398;
	wire [4-1:0] node25399;
	wire [4-1:0] node25400;
	wire [4-1:0] node25403;
	wire [4-1:0] node25406;
	wire [4-1:0] node25407;
	wire [4-1:0] node25408;
	wire [4-1:0] node25409;
	wire [4-1:0] node25412;
	wire [4-1:0] node25415;
	wire [4-1:0] node25417;
	wire [4-1:0] node25418;
	wire [4-1:0] node25421;
	wire [4-1:0] node25424;
	wire [4-1:0] node25426;
	wire [4-1:0] node25427;
	wire [4-1:0] node25430;
	wire [4-1:0] node25433;
	wire [4-1:0] node25434;
	wire [4-1:0] node25435;
	wire [4-1:0] node25436;
	wire [4-1:0] node25437;
	wire [4-1:0] node25440;
	wire [4-1:0] node25443;
	wire [4-1:0] node25444;
	wire [4-1:0] node25447;
	wire [4-1:0] node25450;
	wire [4-1:0] node25451;
	wire [4-1:0] node25452;
	wire [4-1:0] node25455;
	wire [4-1:0] node25458;
	wire [4-1:0] node25459;
	wire [4-1:0] node25460;
	wire [4-1:0] node25463;
	wire [4-1:0] node25466;
	wire [4-1:0] node25467;
	wire [4-1:0] node25470;
	wire [4-1:0] node25473;
	wire [4-1:0] node25474;
	wire [4-1:0] node25475;
	wire [4-1:0] node25478;
	wire [4-1:0] node25481;
	wire [4-1:0] node25482;
	wire [4-1:0] node25483;
	wire [4-1:0] node25484;
	wire [4-1:0] node25485;
	wire [4-1:0] node25489;
	wire [4-1:0] node25491;
	wire [4-1:0] node25494;
	wire [4-1:0] node25495;
	wire [4-1:0] node25498;
	wire [4-1:0] node25501;
	wire [4-1:0] node25502;
	wire [4-1:0] node25505;
	wire [4-1:0] node25506;
	wire [4-1:0] node25510;
	wire [4-1:0] node25511;
	wire [4-1:0] node25512;
	wire [4-1:0] node25515;
	wire [4-1:0] node25518;
	wire [4-1:0] node25519;
	wire [4-1:0] node25520;
	wire [4-1:0] node25521;
	wire [4-1:0] node25524;
	wire [4-1:0] node25527;
	wire [4-1:0] node25528;
	wire [4-1:0] node25529;
	wire [4-1:0] node25532;
	wire [4-1:0] node25535;
	wire [4-1:0] node25536;
	wire [4-1:0] node25537;
	wire [4-1:0] node25541;
	wire [4-1:0] node25542;
	wire [4-1:0] node25545;
	wire [4-1:0] node25548;
	wire [4-1:0] node25549;
	wire [4-1:0] node25552;
	wire [4-1:0] node25555;
	wire [4-1:0] node25556;
	wire [4-1:0] node25557;
	wire [4-1:0] node25558;
	wire [4-1:0] node25559;
	wire [4-1:0] node25560;
	wire [4-1:0] node25561;
	wire [4-1:0] node25562;
	wire [4-1:0] node25563;
	wire [4-1:0] node25566;
	wire [4-1:0] node25569;
	wire [4-1:0] node25571;
	wire [4-1:0] node25574;
	wire [4-1:0] node25575;
	wire [4-1:0] node25578;
	wire [4-1:0] node25581;
	wire [4-1:0] node25582;
	wire [4-1:0] node25585;
	wire [4-1:0] node25588;
	wire [4-1:0] node25589;
	wire [4-1:0] node25590;
	wire [4-1:0] node25594;
	wire [4-1:0] node25596;
	wire [4-1:0] node25599;
	wire [4-1:0] node25600;
	wire [4-1:0] node25601;
	wire [4-1:0] node25602;
	wire [4-1:0] node25605;
	wire [4-1:0] node25608;
	wire [4-1:0] node25609;
	wire [4-1:0] node25612;
	wire [4-1:0] node25615;
	wire [4-1:0] node25616;
	wire [4-1:0] node25617;
	wire [4-1:0] node25621;
	wire [4-1:0] node25622;
	wire [4-1:0] node25626;
	wire [4-1:0] node25627;
	wire [4-1:0] node25628;
	wire [4-1:0] node25629;
	wire [4-1:0] node25630;
	wire [4-1:0] node25633;
	wire [4-1:0] node25636;
	wire [4-1:0] node25637;
	wire [4-1:0] node25638;
	wire [4-1:0] node25641;
	wire [4-1:0] node25644;
	wire [4-1:0] node25646;
	wire [4-1:0] node25649;
	wire [4-1:0] node25650;
	wire [4-1:0] node25652;
	wire [4-1:0] node25655;
	wire [4-1:0] node25657;
	wire [4-1:0] node25660;
	wire [4-1:0] node25661;
	wire [4-1:0] node25662;
	wire [4-1:0] node25663;
	wire [4-1:0] node25666;
	wire [4-1:0] node25669;
	wire [4-1:0] node25670;
	wire [4-1:0] node25673;
	wire [4-1:0] node25676;
	wire [4-1:0] node25677;
	wire [4-1:0] node25678;
	wire [4-1:0] node25682;
	wire [4-1:0] node25684;
	wire [4-1:0] node25687;
	wire [4-1:0] node25688;
	wire [4-1:0] node25689;
	wire [4-1:0] node25690;
	wire [4-1:0] node25691;
	wire [4-1:0] node25692;
	wire [4-1:0] node25694;
	wire [4-1:0] node25697;
	wire [4-1:0] node25698;
	wire [4-1:0] node25699;
	wire [4-1:0] node25702;
	wire [4-1:0] node25705;
	wire [4-1:0] node25706;
	wire [4-1:0] node25709;
	wire [4-1:0] node25712;
	wire [4-1:0] node25713;
	wire [4-1:0] node25714;
	wire [4-1:0] node25717;
	wire [4-1:0] node25720;
	wire [4-1:0] node25721;
	wire [4-1:0] node25724;
	wire [4-1:0] node25727;
	wire [4-1:0] node25728;
	wire [4-1:0] node25729;
	wire [4-1:0] node25730;
	wire [4-1:0] node25731;
	wire [4-1:0] node25735;
	wire [4-1:0] node25738;
	wire [4-1:0] node25739;
	wire [4-1:0] node25742;
	wire [4-1:0] node25745;
	wire [4-1:0] node25746;
	wire [4-1:0] node25747;
	wire [4-1:0] node25750;
	wire [4-1:0] node25751;
	wire [4-1:0] node25755;
	wire [4-1:0] node25757;
	wire [4-1:0] node25760;
	wire [4-1:0] node25761;
	wire [4-1:0] node25762;
	wire [4-1:0] node25763;
	wire [4-1:0] node25764;
	wire [4-1:0] node25768;
	wire [4-1:0] node25770;
	wire [4-1:0] node25773;
	wire [4-1:0] node25775;
	wire [4-1:0] node25776;
	wire [4-1:0] node25780;
	wire [4-1:0] node25781;
	wire [4-1:0] node25782;
	wire [4-1:0] node25783;
	wire [4-1:0] node25787;
	wire [4-1:0] node25789;
	wire [4-1:0] node25792;
	wire [4-1:0] node25793;
	wire [4-1:0] node25794;
	wire [4-1:0] node25798;
	wire [4-1:0] node25800;
	wire [4-1:0] node25803;
	wire [4-1:0] node25804;
	wire [4-1:0] node25805;
	wire [4-1:0] node25806;
	wire [4-1:0] node25807;
	wire [4-1:0] node25809;
	wire [4-1:0] node25811;
	wire [4-1:0] node25814;
	wire [4-1:0] node25815;
	wire [4-1:0] node25816;
	wire [4-1:0] node25820;
	wire [4-1:0] node25822;
	wire [4-1:0] node25825;
	wire [4-1:0] node25826;
	wire [4-1:0] node25827;
	wire [4-1:0] node25828;
	wire [4-1:0] node25832;
	wire [4-1:0] node25834;
	wire [4-1:0] node25837;
	wire [4-1:0] node25838;
	wire [4-1:0] node25842;
	wire [4-1:0] node25843;
	wire [4-1:0] node25844;
	wire [4-1:0] node25845;
	wire [4-1:0] node25846;
	wire [4-1:0] node25851;
	wire [4-1:0] node25852;
	wire [4-1:0] node25854;
	wire [4-1:0] node25857;
	wire [4-1:0] node25859;
	wire [4-1:0] node25862;
	wire [4-1:0] node25864;
	wire [4-1:0] node25865;
	wire [4-1:0] node25866;
	wire [4-1:0] node25870;
	wire [4-1:0] node25873;
	wire [4-1:0] node25874;
	wire [4-1:0] node25875;
	wire [4-1:0] node25876;
	wire [4-1:0] node25877;
	wire [4-1:0] node25878;
	wire [4-1:0] node25881;
	wire [4-1:0] node25884;
	wire [4-1:0] node25885;
	wire [4-1:0] node25889;
	wire [4-1:0] node25891;
	wire [4-1:0] node25892;
	wire [4-1:0] node25895;
	wire [4-1:0] node25898;
	wire [4-1:0] node25899;
	wire [4-1:0] node25902;
	wire [4-1:0] node25904;
	wire [4-1:0] node25906;
	wire [4-1:0] node25909;
	wire [4-1:0] node25910;
	wire [4-1:0] node25911;
	wire [4-1:0] node25912;
	wire [4-1:0] node25913;
	wire [4-1:0] node25916;
	wire [4-1:0] node25920;
	wire [4-1:0] node25922;
	wire [4-1:0] node25923;
	wire [4-1:0] node25926;
	wire [4-1:0] node25929;
	wire [4-1:0] node25930;
	wire [4-1:0] node25931;
	wire [4-1:0] node25932;
	wire [4-1:0] node25936;
	wire [4-1:0] node25939;
	wire [4-1:0] node25941;
	wire [4-1:0] node25942;
	wire [4-1:0] node25945;
	wire [4-1:0] node25948;
	wire [4-1:0] node25949;
	wire [4-1:0] node25950;
	wire [4-1:0] node25951;
	wire [4-1:0] node25952;
	wire [4-1:0] node25955;
	wire [4-1:0] node25956;
	wire [4-1:0] node25959;
	wire [4-1:0] node25962;
	wire [4-1:0] node25963;
	wire [4-1:0] node25964;
	wire [4-1:0] node25967;
	wire [4-1:0] node25970;
	wire [4-1:0] node25973;
	wire [4-1:0] node25974;
	wire [4-1:0] node25975;
	wire [4-1:0] node25977;
	wire [4-1:0] node25980;
	wire [4-1:0] node25982;
	wire [4-1:0] node25985;
	wire [4-1:0] node25986;
	wire [4-1:0] node25988;
	wire [4-1:0] node25991;
	wire [4-1:0] node25992;
	wire [4-1:0] node25996;
	wire [4-1:0] node25997;
	wire [4-1:0] node25998;
	wire [4-1:0] node25999;
	wire [4-1:0] node26000;
	wire [4-1:0] node26001;
	wire [4-1:0] node26004;
	wire [4-1:0] node26005;
	wire [4-1:0] node26008;
	wire [4-1:0] node26011;
	wire [4-1:0] node26012;
	wire [4-1:0] node26013;
	wire [4-1:0] node26016;
	wire [4-1:0] node26019;
	wire [4-1:0] node26022;
	wire [4-1:0] node26023;
	wire [4-1:0] node26024;
	wire [4-1:0] node26025;
	wire [4-1:0] node26027;
	wire [4-1:0] node26030;
	wire [4-1:0] node26032;
	wire [4-1:0] node26035;
	wire [4-1:0] node26036;
	wire [4-1:0] node26037;
	wire [4-1:0] node26041;
	wire [4-1:0] node26042;
	wire [4-1:0] node26046;
	wire [4-1:0] node26047;
	wire [4-1:0] node26048;
	wire [4-1:0] node26050;
	wire [4-1:0] node26053;
	wire [4-1:0] node26054;
	wire [4-1:0] node26058;
	wire [4-1:0] node26059;
	wire [4-1:0] node26060;
	wire [4-1:0] node26061;
	wire [4-1:0] node26066;
	wire [4-1:0] node26067;
	wire [4-1:0] node26071;
	wire [4-1:0] node26072;
	wire [4-1:0] node26073;
	wire [4-1:0] node26074;
	wire [4-1:0] node26075;
	wire [4-1:0] node26078;
	wire [4-1:0] node26079;
	wire [4-1:0] node26082;
	wire [4-1:0] node26085;
	wire [4-1:0] node26086;
	wire [4-1:0] node26089;
	wire [4-1:0] node26092;
	wire [4-1:0] node26093;
	wire [4-1:0] node26094;
	wire [4-1:0] node26095;
	wire [4-1:0] node26097;
	wire [4-1:0] node26100;
	wire [4-1:0] node26103;
	wire [4-1:0] node26104;
	wire [4-1:0] node26107;
	wire [4-1:0] node26108;
	wire [4-1:0] node26112;
	wire [4-1:0] node26113;
	wire [4-1:0] node26114;
	wire [4-1:0] node26117;
	wire [4-1:0] node26120;
	wire [4-1:0] node26121;
	wire [4-1:0] node26123;
	wire [4-1:0] node26126;
	wire [4-1:0] node26129;
	wire [4-1:0] node26130;
	wire [4-1:0] node26131;
	wire [4-1:0] node26134;
	wire [4-1:0] node26135;
	wire [4-1:0] node26138;
	wire [4-1:0] node26141;
	wire [4-1:0] node26142;
	wire [4-1:0] node26143;
	wire [4-1:0] node26146;
	wire [4-1:0] node26149;
	wire [4-1:0] node26152;
	wire [4-1:0] node26153;
	wire [4-1:0] node26154;
	wire [4-1:0] node26157;
	wire [4-1:0] node26158;
	wire [4-1:0] node26161;
	wire [4-1:0] node26164;
	wire [4-1:0] node26165;
	wire [4-1:0] node26166;
	wire [4-1:0] node26169;
	wire [4-1:0] node26172;
	wire [4-1:0] node26175;
	wire [4-1:0] node26176;
	wire [4-1:0] node26177;
	wire [4-1:0] node26178;
	wire [4-1:0] node26179;
	wire [4-1:0] node26180;
	wire [4-1:0] node26182;
	wire [4-1:0] node26185;
	wire [4-1:0] node26187;
	wire [4-1:0] node26190;
	wire [4-1:0] node26191;
	wire [4-1:0] node26193;
	wire [4-1:0] node26196;
	wire [4-1:0] node26198;
	wire [4-1:0] node26201;
	wire [4-1:0] node26202;
	wire [4-1:0] node26203;
	wire [4-1:0] node26205;
	wire [4-1:0] node26208;
	wire [4-1:0] node26210;
	wire [4-1:0] node26213;
	wire [4-1:0] node26214;
	wire [4-1:0] node26215;
	wire [4-1:0] node26219;
	wire [4-1:0] node26220;
	wire [4-1:0] node26224;
	wire [4-1:0] node26225;
	wire [4-1:0] node26226;
	wire [4-1:0] node26227;
	wire [4-1:0] node26230;
	wire [4-1:0] node26233;
	wire [4-1:0] node26234;
	wire [4-1:0] node26235;
	wire [4-1:0] node26236;
	wire [4-1:0] node26237;
	wire [4-1:0] node26240;
	wire [4-1:0] node26243;
	wire [4-1:0] node26244;
	wire [4-1:0] node26246;
	wire [4-1:0] node26249;
	wire [4-1:0] node26250;
	wire [4-1:0] node26253;
	wire [4-1:0] node26256;
	wire [4-1:0] node26257;
	wire [4-1:0] node26260;
	wire [4-1:0] node26263;
	wire [4-1:0] node26264;
	wire [4-1:0] node26265;
	wire [4-1:0] node26268;
	wire [4-1:0] node26271;
	wire [4-1:0] node26272;
	wire [4-1:0] node26273;
	wire [4-1:0] node26274;
	wire [4-1:0] node26277;
	wire [4-1:0] node26281;
	wire [4-1:0] node26282;
	wire [4-1:0] node26285;
	wire [4-1:0] node26286;
	wire [4-1:0] node26289;
	wire [4-1:0] node26292;
	wire [4-1:0] node26293;
	wire [4-1:0] node26294;
	wire [4-1:0] node26297;
	wire [4-1:0] node26300;
	wire [4-1:0] node26301;
	wire [4-1:0] node26302;
	wire [4-1:0] node26303;
	wire [4-1:0] node26304;
	wire [4-1:0] node26306;
	wire [4-1:0] node26309;
	wire [4-1:0] node26310;
	wire [4-1:0] node26313;
	wire [4-1:0] node26316;
	wire [4-1:0] node26317;
	wire [4-1:0] node26318;
	wire [4-1:0] node26321;
	wire [4-1:0] node26324;
	wire [4-1:0] node26325;
	wire [4-1:0] node26328;
	wire [4-1:0] node26331;
	wire [4-1:0] node26332;
	wire [4-1:0] node26335;
	wire [4-1:0] node26338;
	wire [4-1:0] node26339;
	wire [4-1:0] node26340;
	wire [4-1:0] node26343;
	wire [4-1:0] node26346;
	wire [4-1:0] node26347;
	wire [4-1:0] node26348;
	wire [4-1:0] node26351;
	wire [4-1:0] node26354;
	wire [4-1:0] node26355;
	wire [4-1:0] node26358;
	wire [4-1:0] node26361;
	wire [4-1:0] node26362;
	wire [4-1:0] node26363;
	wire [4-1:0] node26364;
	wire [4-1:0] node26365;
	wire [4-1:0] node26368;
	wire [4-1:0] node26371;
	wire [4-1:0] node26372;
	wire [4-1:0] node26373;
	wire [4-1:0] node26374;
	wire [4-1:0] node26375;
	wire [4-1:0] node26376;
	wire [4-1:0] node26379;
	wire [4-1:0] node26382;
	wire [4-1:0] node26383;
	wire [4-1:0] node26387;
	wire [4-1:0] node26388;
	wire [4-1:0] node26390;
	wire [4-1:0] node26394;
	wire [4-1:0] node26395;
	wire [4-1:0] node26396;
	wire [4-1:0] node26399;
	wire [4-1:0] node26402;
	wire [4-1:0] node26403;
	wire [4-1:0] node26404;
	wire [4-1:0] node26407;
	wire [4-1:0] node26410;
	wire [4-1:0] node26411;
	wire [4-1:0] node26414;
	wire [4-1:0] node26417;
	wire [4-1:0] node26418;
	wire [4-1:0] node26419;
	wire [4-1:0] node26422;
	wire [4-1:0] node26425;
	wire [4-1:0] node26426;
	wire [4-1:0] node26428;
	wire [4-1:0] node26431;
	wire [4-1:0] node26432;
	wire [4-1:0] node26434;
	wire [4-1:0] node26437;
	wire [4-1:0] node26438;
	wire [4-1:0] node26439;
	wire [4-1:0] node26442;
	wire [4-1:0] node26446;
	wire [4-1:0] node26447;
	wire [4-1:0] node26448;
	wire [4-1:0] node26449;
	wire [4-1:0] node26452;
	wire [4-1:0] node26455;
	wire [4-1:0] node26456;
	wire [4-1:0] node26457;
	wire [4-1:0] node26460;
	wire [4-1:0] node26463;
	wire [4-1:0] node26464;
	wire [4-1:0] node26465;
	wire [4-1:0] node26468;
	wire [4-1:0] node26471;
	wire [4-1:0] node26472;
	wire [4-1:0] node26475;
	wire [4-1:0] node26478;
	wire [4-1:0] node26479;
	wire [4-1:0] node26480;
	wire [4-1:0] node26483;
	wire [4-1:0] node26486;
	wire [4-1:0] node26487;
	wire [4-1:0] node26490;
	wire [4-1:0] node26493;
	wire [4-1:0] node26494;
	wire [4-1:0] node26495;
	wire [4-1:0] node26499;
	wire [4-1:0] node26500;
	wire [4-1:0] node26504;
	wire [4-1:0] node26505;
	wire [4-1:0] node26506;
	wire [4-1:0] node26507;
	wire [4-1:0] node26508;
	wire [4-1:0] node26509;
	wire [4-1:0] node26510;
	wire [4-1:0] node26511;
	wire [4-1:0] node26512;
	wire [4-1:0] node26513;
	wire [4-1:0] node26514;
	wire [4-1:0] node26515;
	wire [4-1:0] node26516;
	wire [4-1:0] node26517;
	wire [4-1:0] node26521;
	wire [4-1:0] node26522;
	wire [4-1:0] node26523;
	wire [4-1:0] node26526;
	wire [4-1:0] node26529;
	wire [4-1:0] node26530;
	wire [4-1:0] node26533;
	wire [4-1:0] node26536;
	wire [4-1:0] node26537;
	wire [4-1:0] node26538;
	wire [4-1:0] node26541;
	wire [4-1:0] node26545;
	wire [4-1:0] node26546;
	wire [4-1:0] node26547;
	wire [4-1:0] node26548;
	wire [4-1:0] node26551;
	wire [4-1:0] node26554;
	wire [4-1:0] node26555;
	wire [4-1:0] node26556;
	wire [4-1:0] node26559;
	wire [4-1:0] node26562;
	wire [4-1:0] node26563;
	wire [4-1:0] node26567;
	wire [4-1:0] node26568;
	wire [4-1:0] node26569;
	wire [4-1:0] node26572;
	wire [4-1:0] node26575;
	wire [4-1:0] node26576;
	wire [4-1:0] node26579;
	wire [4-1:0] node26582;
	wire [4-1:0] node26583;
	wire [4-1:0] node26584;
	wire [4-1:0] node26585;
	wire [4-1:0] node26586;
	wire [4-1:0] node26587;
	wire [4-1:0] node26590;
	wire [4-1:0] node26593;
	wire [4-1:0] node26594;
	wire [4-1:0] node26597;
	wire [4-1:0] node26600;
	wire [4-1:0] node26601;
	wire [4-1:0] node26604;
	wire [4-1:0] node26607;
	wire [4-1:0] node26608;
	wire [4-1:0] node26609;
	wire [4-1:0] node26613;
	wire [4-1:0] node26614;
	wire [4-1:0] node26615;
	wire [4-1:0] node26619;
	wire [4-1:0] node26620;
	wire [4-1:0] node26623;
	wire [4-1:0] node26626;
	wire [4-1:0] node26627;
	wire [4-1:0] node26628;
	wire [4-1:0] node26630;
	wire [4-1:0] node26631;
	wire [4-1:0] node26634;
	wire [4-1:0] node26637;
	wire [4-1:0] node26638;
	wire [4-1:0] node26640;
	wire [4-1:0] node26644;
	wire [4-1:0] node26645;
	wire [4-1:0] node26646;
	wire [4-1:0] node26650;
	wire [4-1:0] node26651;
	wire [4-1:0] node26654;
	wire [4-1:0] node26655;
	wire [4-1:0] node26659;
	wire [4-1:0] node26660;
	wire [4-1:0] node26661;
	wire [4-1:0] node26662;
	wire [4-1:0] node26663;
	wire [4-1:0] node26664;
	wire [4-1:0] node26667;
	wire [4-1:0] node26670;
	wire [4-1:0] node26671;
	wire [4-1:0] node26674;
	wire [4-1:0] node26676;
	wire [4-1:0] node26679;
	wire [4-1:0] node26680;
	wire [4-1:0] node26682;
	wire [4-1:0] node26684;
	wire [4-1:0] node26688;
	wire [4-1:0] node26689;
	wire [4-1:0] node26690;
	wire [4-1:0] node26691;
	wire [4-1:0] node26692;
	wire [4-1:0] node26696;
	wire [4-1:0] node26697;
	wire [4-1:0] node26700;
	wire [4-1:0] node26703;
	wire [4-1:0] node26705;
	wire [4-1:0] node26706;
	wire [4-1:0] node26709;
	wire [4-1:0] node26712;
	wire [4-1:0] node26713;
	wire [4-1:0] node26714;
	wire [4-1:0] node26715;
	wire [4-1:0] node26718;
	wire [4-1:0] node26723;
	wire [4-1:0] node26724;
	wire [4-1:0] node26725;
	wire [4-1:0] node26726;
	wire [4-1:0] node26728;
	wire [4-1:0] node26729;
	wire [4-1:0] node26733;
	wire [4-1:0] node26734;
	wire [4-1:0] node26735;
	wire [4-1:0] node26739;
	wire [4-1:0] node26741;
	wire [4-1:0] node26744;
	wire [4-1:0] node26745;
	wire [4-1:0] node26746;
	wire [4-1:0] node26750;
	wire [4-1:0] node26751;
	wire [4-1:0] node26752;
	wire [4-1:0] node26755;
	wire [4-1:0] node26759;
	wire [4-1:0] node26760;
	wire [4-1:0] node26761;
	wire [4-1:0] node26762;
	wire [4-1:0] node26763;
	wire [4-1:0] node26766;
	wire [4-1:0] node26770;
	wire [4-1:0] node26771;
	wire [4-1:0] node26775;
	wire [4-1:0] node26776;
	wire [4-1:0] node26778;
	wire [4-1:0] node26780;
	wire [4-1:0] node26783;
	wire [4-1:0] node26784;
	wire [4-1:0] node26787;
	wire [4-1:0] node26790;
	wire [4-1:0] node26791;
	wire [4-1:0] node26792;
	wire [4-1:0] node26793;
	wire [4-1:0] node26794;
	wire [4-1:0] node26795;
	wire [4-1:0] node26796;
	wire [4-1:0] node26799;
	wire [4-1:0] node26802;
	wire [4-1:0] node26803;
	wire [4-1:0] node26804;
	wire [4-1:0] node26807;
	wire [4-1:0] node26811;
	wire [4-1:0] node26812;
	wire [4-1:0] node26814;
	wire [4-1:0] node26815;
	wire [4-1:0] node26818;
	wire [4-1:0] node26821;
	wire [4-1:0] node26822;
	wire [4-1:0] node26824;
	wire [4-1:0] node26827;
	wire [4-1:0] node26828;
	wire [4-1:0] node26832;
	wire [4-1:0] node26833;
	wire [4-1:0] node26834;
	wire [4-1:0] node26835;
	wire [4-1:0] node26838;
	wire [4-1:0] node26840;
	wire [4-1:0] node26843;
	wire [4-1:0] node26844;
	wire [4-1:0] node26848;
	wire [4-1:0] node26849;
	wire [4-1:0] node26851;
	wire [4-1:0] node26854;
	wire [4-1:0] node26855;
	wire [4-1:0] node26857;
	wire [4-1:0] node26860;
	wire [4-1:0] node26861;
	wire [4-1:0] node26865;
	wire [4-1:0] node26866;
	wire [4-1:0] node26867;
	wire [4-1:0] node26868;
	wire [4-1:0] node26869;
	wire [4-1:0] node26870;
	wire [4-1:0] node26873;
	wire [4-1:0] node26876;
	wire [4-1:0] node26877;
	wire [4-1:0] node26880;
	wire [4-1:0] node26883;
	wire [4-1:0] node26885;
	wire [4-1:0] node26886;
	wire [4-1:0] node26889;
	wire [4-1:0] node26892;
	wire [4-1:0] node26893;
	wire [4-1:0] node26894;
	wire [4-1:0] node26896;
	wire [4-1:0] node26899;
	wire [4-1:0] node26900;
	wire [4-1:0] node26903;
	wire [4-1:0] node26906;
	wire [4-1:0] node26907;
	wire [4-1:0] node26909;
	wire [4-1:0] node26912;
	wire [4-1:0] node26913;
	wire [4-1:0] node26916;
	wire [4-1:0] node26919;
	wire [4-1:0] node26920;
	wire [4-1:0] node26921;
	wire [4-1:0] node26922;
	wire [4-1:0] node26923;
	wire [4-1:0] node26928;
	wire [4-1:0] node26929;
	wire [4-1:0] node26931;
	wire [4-1:0] node26934;
	wire [4-1:0] node26935;
	wire [4-1:0] node26938;
	wire [4-1:0] node26941;
	wire [4-1:0] node26942;
	wire [4-1:0] node26943;
	wire [4-1:0] node26944;
	wire [4-1:0] node26947;
	wire [4-1:0] node26950;
	wire [4-1:0] node26951;
	wire [4-1:0] node26955;
	wire [4-1:0] node26956;
	wire [4-1:0] node26959;
	wire [4-1:0] node26960;
	wire [4-1:0] node26964;
	wire [4-1:0] node26965;
	wire [4-1:0] node26966;
	wire [4-1:0] node26967;
	wire [4-1:0] node26969;
	wire [4-1:0] node26970;
	wire [4-1:0] node26972;
	wire [4-1:0] node26976;
	wire [4-1:0] node26977;
	wire [4-1:0] node26978;
	wire [4-1:0] node26982;
	wire [4-1:0] node26983;
	wire [4-1:0] node26986;
	wire [4-1:0] node26989;
	wire [4-1:0] node26990;
	wire [4-1:0] node26991;
	wire [4-1:0] node26994;
	wire [4-1:0] node26996;
	wire [4-1:0] node26998;
	wire [4-1:0] node27001;
	wire [4-1:0] node27002;
	wire [4-1:0] node27004;
	wire [4-1:0] node27007;
	wire [4-1:0] node27008;
	wire [4-1:0] node27010;
	wire [4-1:0] node27014;
	wire [4-1:0] node27015;
	wire [4-1:0] node27016;
	wire [4-1:0] node27017;
	wire [4-1:0] node27019;
	wire [4-1:0] node27021;
	wire [4-1:0] node27024;
	wire [4-1:0] node27025;
	wire [4-1:0] node27028;
	wire [4-1:0] node27031;
	wire [4-1:0] node27032;
	wire [4-1:0] node27033;
	wire [4-1:0] node27035;
	wire [4-1:0] node27038;
	wire [4-1:0] node27040;
	wire [4-1:0] node27043;
	wire [4-1:0] node27045;
	wire [4-1:0] node27047;
	wire [4-1:0] node27050;
	wire [4-1:0] node27051;
	wire [4-1:0] node27052;
	wire [4-1:0] node27054;
	wire [4-1:0] node27057;
	wire [4-1:0] node27058;
	wire [4-1:0] node27061;
	wire [4-1:0] node27063;
	wire [4-1:0] node27066;
	wire [4-1:0] node27067;
	wire [4-1:0] node27068;
	wire [4-1:0] node27069;
	wire [4-1:0] node27073;
	wire [4-1:0] node27075;
	wire [4-1:0] node27078;
	wire [4-1:0] node27079;
	wire [4-1:0] node27081;
	wire [4-1:0] node27084;
	wire [4-1:0] node27087;
	wire [4-1:0] node27088;
	wire [4-1:0] node27089;
	wire [4-1:0] node27090;
	wire [4-1:0] node27091;
	wire [4-1:0] node27092;
	wire [4-1:0] node27093;
	wire [4-1:0] node27094;
	wire [4-1:0] node27096;
	wire [4-1:0] node27099;
	wire [4-1:0] node27102;
	wire [4-1:0] node27103;
	wire [4-1:0] node27105;
	wire [4-1:0] node27108;
	wire [4-1:0] node27111;
	wire [4-1:0] node27112;
	wire [4-1:0] node27114;
	wire [4-1:0] node27118;
	wire [4-1:0] node27119;
	wire [4-1:0] node27120;
	wire [4-1:0] node27122;
	wire [4-1:0] node27125;
	wire [4-1:0] node27126;
	wire [4-1:0] node27127;
	wire [4-1:0] node27131;
	wire [4-1:0] node27134;
	wire [4-1:0] node27135;
	wire [4-1:0] node27136;
	wire [4-1:0] node27137;
	wire [4-1:0] node27141;
	wire [4-1:0] node27144;
	wire [4-1:0] node27146;
	wire [4-1:0] node27147;
	wire [4-1:0] node27151;
	wire [4-1:0] node27152;
	wire [4-1:0] node27153;
	wire [4-1:0] node27154;
	wire [4-1:0] node27155;
	wire [4-1:0] node27157;
	wire [4-1:0] node27160;
	wire [4-1:0] node27163;
	wire [4-1:0] node27164;
	wire [4-1:0] node27168;
	wire [4-1:0] node27169;
	wire [4-1:0] node27170;
	wire [4-1:0] node27171;
	wire [4-1:0] node27175;
	wire [4-1:0] node27176;
	wire [4-1:0] node27180;
	wire [4-1:0] node27181;
	wire [4-1:0] node27185;
	wire [4-1:0] node27186;
	wire [4-1:0] node27187;
	wire [4-1:0] node27188;
	wire [4-1:0] node27189;
	wire [4-1:0] node27192;
	wire [4-1:0] node27195;
	wire [4-1:0] node27196;
	wire [4-1:0] node27199;
	wire [4-1:0] node27202;
	wire [4-1:0] node27203;
	wire [4-1:0] node27204;
	wire [4-1:0] node27207;
	wire [4-1:0] node27210;
	wire [4-1:0] node27212;
	wire [4-1:0] node27215;
	wire [4-1:0] node27216;
	wire [4-1:0] node27218;
	wire [4-1:0] node27221;
	wire [4-1:0] node27222;
	wire [4-1:0] node27223;
	wire [4-1:0] node27226;
	wire [4-1:0] node27230;
	wire [4-1:0] node27231;
	wire [4-1:0] node27232;
	wire [4-1:0] node27233;
	wire [4-1:0] node27234;
	wire [4-1:0] node27235;
	wire [4-1:0] node27236;
	wire [4-1:0] node27240;
	wire [4-1:0] node27242;
	wire [4-1:0] node27245;
	wire [4-1:0] node27246;
	wire [4-1:0] node27247;
	wire [4-1:0] node27252;
	wire [4-1:0] node27253;
	wire [4-1:0] node27254;
	wire [4-1:0] node27257;
	wire [4-1:0] node27260;
	wire [4-1:0] node27261;
	wire [4-1:0] node27262;
	wire [4-1:0] node27265;
	wire [4-1:0] node27268;
	wire [4-1:0] node27269;
	wire [4-1:0] node27272;
	wire [4-1:0] node27275;
	wire [4-1:0] node27276;
	wire [4-1:0] node27277;
	wire [4-1:0] node27278;
	wire [4-1:0] node27281;
	wire [4-1:0] node27284;
	wire [4-1:0] node27285;
	wire [4-1:0] node27288;
	wire [4-1:0] node27289;
	wire [4-1:0] node27293;
	wire [4-1:0] node27294;
	wire [4-1:0] node27295;
	wire [4-1:0] node27296;
	wire [4-1:0] node27300;
	wire [4-1:0] node27303;
	wire [4-1:0] node27304;
	wire [4-1:0] node27306;
	wire [4-1:0] node27309;
	wire [4-1:0] node27312;
	wire [4-1:0] node27313;
	wire [4-1:0] node27314;
	wire [4-1:0] node27315;
	wire [4-1:0] node27317;
	wire [4-1:0] node27320;
	wire [4-1:0] node27321;
	wire [4-1:0] node27322;
	wire [4-1:0] node27325;
	wire [4-1:0] node27329;
	wire [4-1:0] node27330;
	wire [4-1:0] node27331;
	wire [4-1:0] node27333;
	wire [4-1:0] node27338;
	wire [4-1:0] node27339;
	wire [4-1:0] node27340;
	wire [4-1:0] node27341;
	wire [4-1:0] node27342;
	wire [4-1:0] node27345;
	wire [4-1:0] node27348;
	wire [4-1:0] node27349;
	wire [4-1:0] node27352;
	wire [4-1:0] node27355;
	wire [4-1:0] node27357;
	wire [4-1:0] node27360;
	wire [4-1:0] node27361;
	wire [4-1:0] node27363;
	wire [4-1:0] node27366;
	wire [4-1:0] node27368;
	wire [4-1:0] node27370;
	wire [4-1:0] node27373;
	wire [4-1:0] node27374;
	wire [4-1:0] node27375;
	wire [4-1:0] node27376;
	wire [4-1:0] node27377;
	wire [4-1:0] node27378;
	wire [4-1:0] node27379;
	wire [4-1:0] node27382;
	wire [4-1:0] node27385;
	wire [4-1:0] node27387;
	wire [4-1:0] node27389;
	wire [4-1:0] node27392;
	wire [4-1:0] node27393;
	wire [4-1:0] node27394;
	wire [4-1:0] node27398;
	wire [4-1:0] node27399;
	wire [4-1:0] node27400;
	wire [4-1:0] node27404;
	wire [4-1:0] node27405;
	wire [4-1:0] node27409;
	wire [4-1:0] node27410;
	wire [4-1:0] node27411;
	wire [4-1:0] node27412;
	wire [4-1:0] node27415;
	wire [4-1:0] node27418;
	wire [4-1:0] node27420;
	wire [4-1:0] node27423;
	wire [4-1:0] node27424;
	wire [4-1:0] node27425;
	wire [4-1:0] node27429;
	wire [4-1:0] node27430;
	wire [4-1:0] node27431;
	wire [4-1:0] node27435;
	wire [4-1:0] node27437;
	wire [4-1:0] node27440;
	wire [4-1:0] node27441;
	wire [4-1:0] node27442;
	wire [4-1:0] node27443;
	wire [4-1:0] node27444;
	wire [4-1:0] node27445;
	wire [4-1:0] node27449;
	wire [4-1:0] node27452;
	wire [4-1:0] node27454;
	wire [4-1:0] node27455;
	wire [4-1:0] node27458;
	wire [4-1:0] node27461;
	wire [4-1:0] node27462;
	wire [4-1:0] node27464;
	wire [4-1:0] node27467;
	wire [4-1:0] node27468;
	wire [4-1:0] node27470;
	wire [4-1:0] node27473;
	wire [4-1:0] node27476;
	wire [4-1:0] node27477;
	wire [4-1:0] node27478;
	wire [4-1:0] node27479;
	wire [4-1:0] node27482;
	wire [4-1:0] node27485;
	wire [4-1:0] node27486;
	wire [4-1:0] node27487;
	wire [4-1:0] node27490;
	wire [4-1:0] node27493;
	wire [4-1:0] node27494;
	wire [4-1:0] node27498;
	wire [4-1:0] node27499;
	wire [4-1:0] node27500;
	wire [4-1:0] node27503;
	wire [4-1:0] node27506;
	wire [4-1:0] node27509;
	wire [4-1:0] node27510;
	wire [4-1:0] node27511;
	wire [4-1:0] node27512;
	wire [4-1:0] node27513;
	wire [4-1:0] node27514;
	wire [4-1:0] node27515;
	wire [4-1:0] node27519;
	wire [4-1:0] node27522;
	wire [4-1:0] node27523;
	wire [4-1:0] node27524;
	wire [4-1:0] node27528;
	wire [4-1:0] node27530;
	wire [4-1:0] node27533;
	wire [4-1:0] node27534;
	wire [4-1:0] node27535;
	wire [4-1:0] node27537;
	wire [4-1:0] node27540;
	wire [4-1:0] node27541;
	wire [4-1:0] node27544;
	wire [4-1:0] node27547;
	wire [4-1:0] node27548;
	wire [4-1:0] node27550;
	wire [4-1:0] node27553;
	wire [4-1:0] node27554;
	wire [4-1:0] node27557;
	wire [4-1:0] node27560;
	wire [4-1:0] node27561;
	wire [4-1:0] node27562;
	wire [4-1:0] node27563;
	wire [4-1:0] node27564;
	wire [4-1:0] node27568;
	wire [4-1:0] node27569;
	wire [4-1:0] node27573;
	wire [4-1:0] node27574;
	wire [4-1:0] node27575;
	wire [4-1:0] node27579;
	wire [4-1:0] node27580;
	wire [4-1:0] node27584;
	wire [4-1:0] node27585;
	wire [4-1:0] node27587;
	wire [4-1:0] node27590;
	wire [4-1:0] node27591;
	wire [4-1:0] node27593;
	wire [4-1:0] node27596;
	wire [4-1:0] node27599;
	wire [4-1:0] node27600;
	wire [4-1:0] node27601;
	wire [4-1:0] node27602;
	wire [4-1:0] node27603;
	wire [4-1:0] node27605;
	wire [4-1:0] node27608;
	wire [4-1:0] node27609;
	wire [4-1:0] node27613;
	wire [4-1:0] node27614;
	wire [4-1:0] node27618;
	wire [4-1:0] node27620;
	wire [4-1:0] node27621;
	wire [4-1:0] node27624;
	wire [4-1:0] node27625;
	wire [4-1:0] node27629;
	wire [4-1:0] node27630;
	wire [4-1:0] node27631;
	wire [4-1:0] node27632;
	wire [4-1:0] node27633;
	wire [4-1:0] node27637;
	wire [4-1:0] node27639;
	wire [4-1:0] node27642;
	wire [4-1:0] node27643;
	wire [4-1:0] node27644;
	wire [4-1:0] node27648;
	wire [4-1:0] node27651;
	wire [4-1:0] node27652;
	wire [4-1:0] node27654;
	wire [4-1:0] node27657;
	wire [4-1:0] node27658;
	wire [4-1:0] node27660;
	wire [4-1:0] node27663;
	wire [4-1:0] node27664;
	wire [4-1:0] node27668;
	wire [4-1:0] node27669;
	wire [4-1:0] node27670;
	wire [4-1:0] node27671;
	wire [4-1:0] node27672;
	wire [4-1:0] node27673;
	wire [4-1:0] node27674;
	wire [4-1:0] node27675;
	wire [4-1:0] node27676;
	wire [4-1:0] node27677;
	wire [4-1:0] node27681;
	wire [4-1:0] node27685;
	wire [4-1:0] node27686;
	wire [4-1:0] node27687;
	wire [4-1:0] node27690;
	wire [4-1:0] node27693;
	wire [4-1:0] node27694;
	wire [4-1:0] node27697;
	wire [4-1:0] node27699;
	wire [4-1:0] node27702;
	wire [4-1:0] node27703;
	wire [4-1:0] node27704;
	wire [4-1:0] node27706;
	wire [4-1:0] node27707;
	wire [4-1:0] node27710;
	wire [4-1:0] node27714;
	wire [4-1:0] node27715;
	wire [4-1:0] node27717;
	wire [4-1:0] node27720;
	wire [4-1:0] node27722;
	wire [4-1:0] node27725;
	wire [4-1:0] node27726;
	wire [4-1:0] node27727;
	wire [4-1:0] node27728;
	wire [4-1:0] node27729;
	wire [4-1:0] node27733;
	wire [4-1:0] node27735;
	wire [4-1:0] node27738;
	wire [4-1:0] node27739;
	wire [4-1:0] node27741;
	wire [4-1:0] node27744;
	wire [4-1:0] node27746;
	wire [4-1:0] node27749;
	wire [4-1:0] node27750;
	wire [4-1:0] node27751;
	wire [4-1:0] node27752;
	wire [4-1:0] node27755;
	wire [4-1:0] node27757;
	wire [4-1:0] node27760;
	wire [4-1:0] node27762;
	wire [4-1:0] node27764;
	wire [4-1:0] node27767;
	wire [4-1:0] node27768;
	wire [4-1:0] node27769;
	wire [4-1:0] node27771;
	wire [4-1:0] node27774;
	wire [4-1:0] node27776;
	wire [4-1:0] node27779;
	wire [4-1:0] node27781;
	wire [4-1:0] node27783;
	wire [4-1:0] node27786;
	wire [4-1:0] node27787;
	wire [4-1:0] node27788;
	wire [4-1:0] node27789;
	wire [4-1:0] node27790;
	wire [4-1:0] node27792;
	wire [4-1:0] node27795;
	wire [4-1:0] node27796;
	wire [4-1:0] node27799;
	wire [4-1:0] node27802;
	wire [4-1:0] node27803;
	wire [4-1:0] node27804;
	wire [4-1:0] node27807;
	wire [4-1:0] node27810;
	wire [4-1:0] node27811;
	wire [4-1:0] node27815;
	wire [4-1:0] node27816;
	wire [4-1:0] node27817;
	wire [4-1:0] node27818;
	wire [4-1:0] node27822;
	wire [4-1:0] node27823;
	wire [4-1:0] node27827;
	wire [4-1:0] node27829;
	wire [4-1:0] node27830;
	wire [4-1:0] node27834;
	wire [4-1:0] node27835;
	wire [4-1:0] node27836;
	wire [4-1:0] node27837;
	wire [4-1:0] node27838;
	wire [4-1:0] node27841;
	wire [4-1:0] node27842;
	wire [4-1:0] node27846;
	wire [4-1:0] node27847;
	wire [4-1:0] node27848;
	wire [4-1:0] node27852;
	wire [4-1:0] node27855;
	wire [4-1:0] node27856;
	wire [4-1:0] node27857;
	wire [4-1:0] node27859;
	wire [4-1:0] node27862;
	wire [4-1:0] node27864;
	wire [4-1:0] node27867;
	wire [4-1:0] node27869;
	wire [4-1:0] node27870;
	wire [4-1:0] node27873;
	wire [4-1:0] node27876;
	wire [4-1:0] node27877;
	wire [4-1:0] node27878;
	wire [4-1:0] node27880;
	wire [4-1:0] node27883;
	wire [4-1:0] node27884;
	wire [4-1:0] node27886;
	wire [4-1:0] node27889;
	wire [4-1:0] node27891;
	wire [4-1:0] node27894;
	wire [4-1:0] node27895;
	wire [4-1:0] node27896;
	wire [4-1:0] node27898;
	wire [4-1:0] node27901;
	wire [4-1:0] node27903;
	wire [4-1:0] node27906;
	wire [4-1:0] node27907;
	wire [4-1:0] node27911;
	wire [4-1:0] node27912;
	wire [4-1:0] node27913;
	wire [4-1:0] node27914;
	wire [4-1:0] node27915;
	wire [4-1:0] node27916;
	wire [4-1:0] node27917;
	wire [4-1:0] node27921;
	wire [4-1:0] node27924;
	wire [4-1:0] node27925;
	wire [4-1:0] node27926;
	wire [4-1:0] node27931;
	wire [4-1:0] node27932;
	wire [4-1:0] node27933;
	wire [4-1:0] node27934;
	wire [4-1:0] node27938;
	wire [4-1:0] node27939;
	wire [4-1:0] node27943;
	wire [4-1:0] node27944;
	wire [4-1:0] node27946;
	wire [4-1:0] node27949;
	wire [4-1:0] node27950;
	wire [4-1:0] node27954;
	wire [4-1:0] node27955;
	wire [4-1:0] node27956;
	wire [4-1:0] node27957;
	wire [4-1:0] node27958;
	wire [4-1:0] node27962;
	wire [4-1:0] node27963;
	wire [4-1:0] node27967;
	wire [4-1:0] node27968;
	wire [4-1:0] node27969;
	wire [4-1:0] node27973;
	wire [4-1:0] node27974;
	wire [4-1:0] node27978;
	wire [4-1:0] node27979;
	wire [4-1:0] node27980;
	wire [4-1:0] node27981;
	wire [4-1:0] node27985;
	wire [4-1:0] node27987;
	wire [4-1:0] node27990;
	wire [4-1:0] node27991;
	wire [4-1:0] node27992;
	wire [4-1:0] node27996;
	wire [4-1:0] node27997;
	wire [4-1:0] node28001;
	wire [4-1:0] node28002;
	wire [4-1:0] node28003;
	wire [4-1:0] node28004;
	wire [4-1:0] node28005;
	wire [4-1:0] node28006;
	wire [4-1:0] node28008;
	wire [4-1:0] node28011;
	wire [4-1:0] node28012;
	wire [4-1:0] node28016;
	wire [4-1:0] node28018;
	wire [4-1:0] node28021;
	wire [4-1:0] node28022;
	wire [4-1:0] node28023;
	wire [4-1:0] node28026;
	wire [4-1:0] node28029;
	wire [4-1:0] node28031;
	wire [4-1:0] node28034;
	wire [4-1:0] node28035;
	wire [4-1:0] node28036;
	wire [4-1:0] node28038;
	wire [4-1:0] node28041;
	wire [4-1:0] node28043;
	wire [4-1:0] node28046;
	wire [4-1:0] node28047;
	wire [4-1:0] node28049;
	wire [4-1:0] node28052;
	wire [4-1:0] node28054;
	wire [4-1:0] node28057;
	wire [4-1:0] node28058;
	wire [4-1:0] node28059;
	wire [4-1:0] node28060;
	wire [4-1:0] node28061;
	wire [4-1:0] node28066;
	wire [4-1:0] node28067;
	wire [4-1:0] node28069;
	wire [4-1:0] node28072;
	wire [4-1:0] node28074;
	wire [4-1:0] node28077;
	wire [4-1:0] node28078;
	wire [4-1:0] node28079;
	wire [4-1:0] node28081;
	wire [4-1:0] node28084;
	wire [4-1:0] node28086;
	wire [4-1:0] node28089;
	wire [4-1:0] node28090;
	wire [4-1:0] node28092;
	wire [4-1:0] node28095;
	wire [4-1:0] node28097;
	wire [4-1:0] node28100;
	wire [4-1:0] node28101;
	wire [4-1:0] node28102;
	wire [4-1:0] node28103;
	wire [4-1:0] node28104;
	wire [4-1:0] node28105;
	wire [4-1:0] node28107;
	wire [4-1:0] node28109;
	wire [4-1:0] node28112;
	wire [4-1:0] node28113;
	wire [4-1:0] node28114;
	wire [4-1:0] node28118;
	wire [4-1:0] node28120;
	wire [4-1:0] node28123;
	wire [4-1:0] node28124;
	wire [4-1:0] node28125;
	wire [4-1:0] node28128;
	wire [4-1:0] node28131;
	wire [4-1:0] node28132;
	wire [4-1:0] node28133;
	wire [4-1:0] node28137;
	wire [4-1:0] node28138;
	wire [4-1:0] node28141;
	wire [4-1:0] node28144;
	wire [4-1:0] node28145;
	wire [4-1:0] node28146;
	wire [4-1:0] node28147;
	wire [4-1:0] node28149;
	wire [4-1:0] node28152;
	wire [4-1:0] node28155;
	wire [4-1:0] node28156;
	wire [4-1:0] node28158;
	wire [4-1:0] node28161;
	wire [4-1:0] node28164;
	wire [4-1:0] node28165;
	wire [4-1:0] node28166;
	wire [4-1:0] node28168;
	wire [4-1:0] node28171;
	wire [4-1:0] node28172;
	wire [4-1:0] node28175;
	wire [4-1:0] node28178;
	wire [4-1:0] node28179;
	wire [4-1:0] node28180;
	wire [4-1:0] node28181;
	wire [4-1:0] node28184;
	wire [4-1:0] node28187;
	wire [4-1:0] node28188;
	wire [4-1:0] node28191;
	wire [4-1:0] node28194;
	wire [4-1:0] node28195;
	wire [4-1:0] node28196;
	wire [4-1:0] node28199;
	wire [4-1:0] node28203;
	wire [4-1:0] node28204;
	wire [4-1:0] node28205;
	wire [4-1:0] node28206;
	wire [4-1:0] node28207;
	wire [4-1:0] node28208;
	wire [4-1:0] node28212;
	wire [4-1:0] node28214;
	wire [4-1:0] node28217;
	wire [4-1:0] node28218;
	wire [4-1:0] node28219;
	wire [4-1:0] node28223;
	wire [4-1:0] node28225;
	wire [4-1:0] node28228;
	wire [4-1:0] node28229;
	wire [4-1:0] node28230;
	wire [4-1:0] node28233;
	wire [4-1:0] node28236;
	wire [4-1:0] node28237;
	wire [4-1:0] node28239;
	wire [4-1:0] node28242;
	wire [4-1:0] node28244;
	wire [4-1:0] node28247;
	wire [4-1:0] node28248;
	wire [4-1:0] node28249;
	wire [4-1:0] node28250;
	wire [4-1:0] node28251;
	wire [4-1:0] node28255;
	wire [4-1:0] node28257;
	wire [4-1:0] node28260;
	wire [4-1:0] node28261;
	wire [4-1:0] node28262;
	wire [4-1:0] node28266;
	wire [4-1:0] node28268;
	wire [4-1:0] node28271;
	wire [4-1:0] node28272;
	wire [4-1:0] node28273;
	wire [4-1:0] node28275;
	wire [4-1:0] node28278;
	wire [4-1:0] node28279;
	wire [4-1:0] node28283;
	wire [4-1:0] node28284;
	wire [4-1:0] node28285;
	wire [4-1:0] node28289;
	wire [4-1:0] node28291;
	wire [4-1:0] node28294;
	wire [4-1:0] node28295;
	wire [4-1:0] node28296;
	wire [4-1:0] node28297;
	wire [4-1:0] node28299;
	wire [4-1:0] node28300;
	wire [4-1:0] node28301;
	wire [4-1:0] node28304;
	wire [4-1:0] node28307;
	wire [4-1:0] node28308;
	wire [4-1:0] node28309;
	wire [4-1:0] node28314;
	wire [4-1:0] node28316;
	wire [4-1:0] node28317;
	wire [4-1:0] node28320;
	wire [4-1:0] node28323;
	wire [4-1:0] node28324;
	wire [4-1:0] node28326;
	wire [4-1:0] node28327;
	wire [4-1:0] node28328;
	wire [4-1:0] node28331;
	wire [4-1:0] node28334;
	wire [4-1:0] node28335;
	wire [4-1:0] node28339;
	wire [4-1:0] node28341;
	wire [4-1:0] node28342;
	wire [4-1:0] node28343;
	wire [4-1:0] node28344;
	wire [4-1:0] node28347;
	wire [4-1:0] node28350;
	wire [4-1:0] node28351;
	wire [4-1:0] node28354;
	wire [4-1:0] node28357;
	wire [4-1:0] node28358;
	wire [4-1:0] node28361;
	wire [4-1:0] node28364;
	wire [4-1:0] node28365;
	wire [4-1:0] node28366;
	wire [4-1:0] node28368;
	wire [4-1:0] node28369;
	wire [4-1:0] node28371;
	wire [4-1:0] node28372;
	wire [4-1:0] node28376;
	wire [4-1:0] node28377;
	wire [4-1:0] node28378;
	wire [4-1:0] node28381;
	wire [4-1:0] node28384;
	wire [4-1:0] node28385;
	wire [4-1:0] node28388;
	wire [4-1:0] node28391;
	wire [4-1:0] node28393;
	wire [4-1:0] node28394;
	wire [4-1:0] node28395;
	wire [4-1:0] node28398;
	wire [4-1:0] node28401;
	wire [4-1:0] node28402;
	wire [4-1:0] node28404;
	wire [4-1:0] node28407;
	wire [4-1:0] node28409;
	wire [4-1:0] node28412;
	wire [4-1:0] node28413;
	wire [4-1:0] node28415;
	wire [4-1:0] node28416;
	wire [4-1:0] node28419;
	wire [4-1:0] node28422;
	wire [4-1:0] node28424;
	wire [4-1:0] node28425;
	wire [4-1:0] node28428;
	wire [4-1:0] node28431;
	wire [4-1:0] node28432;
	wire [4-1:0] node28433;
	wire [4-1:0] node28434;
	wire [4-1:0] node28435;
	wire [4-1:0] node28436;
	wire [4-1:0] node28437;
	wire [4-1:0] node28438;
	wire [4-1:0] node28439;
	wire [4-1:0] node28440;
	wire [4-1:0] node28443;
	wire [4-1:0] node28446;
	wire [4-1:0] node28447;
	wire [4-1:0] node28451;
	wire [4-1:0] node28452;
	wire [4-1:0] node28453;
	wire [4-1:0] node28455;
	wire [4-1:0] node28458;
	wire [4-1:0] node28459;
	wire [4-1:0] node28462;
	wire [4-1:0] node28465;
	wire [4-1:0] node28466;
	wire [4-1:0] node28467;
	wire [4-1:0] node28471;
	wire [4-1:0] node28472;
	wire [4-1:0] node28476;
	wire [4-1:0] node28477;
	wire [4-1:0] node28478;
	wire [4-1:0] node28479;
	wire [4-1:0] node28480;
	wire [4-1:0] node28483;
	wire [4-1:0] node28486;
	wire [4-1:0] node28489;
	wire [4-1:0] node28490;
	wire [4-1:0] node28493;
	wire [4-1:0] node28496;
	wire [4-1:0] node28497;
	wire [4-1:0] node28498;
	wire [4-1:0] node28499;
	wire [4-1:0] node28503;
	wire [4-1:0] node28506;
	wire [4-1:0] node28507;
	wire [4-1:0] node28510;
	wire [4-1:0] node28511;
	wire [4-1:0] node28514;
	wire [4-1:0] node28517;
	wire [4-1:0] node28518;
	wire [4-1:0] node28519;
	wire [4-1:0] node28520;
	wire [4-1:0] node28521;
	wire [4-1:0] node28522;
	wire [4-1:0] node28525;
	wire [4-1:0] node28528;
	wire [4-1:0] node28531;
	wire [4-1:0] node28532;
	wire [4-1:0] node28533;
	wire [4-1:0] node28536;
	wire [4-1:0] node28539;
	wire [4-1:0] node28542;
	wire [4-1:0] node28543;
	wire [4-1:0] node28544;
	wire [4-1:0] node28545;
	wire [4-1:0] node28548;
	wire [4-1:0] node28551;
	wire [4-1:0] node28552;
	wire [4-1:0] node28556;
	wire [4-1:0] node28557;
	wire [4-1:0] node28559;
	wire [4-1:0] node28562;
	wire [4-1:0] node28563;
	wire [4-1:0] node28567;
	wire [4-1:0] node28568;
	wire [4-1:0] node28569;
	wire [4-1:0] node28570;
	wire [4-1:0] node28572;
	wire [4-1:0] node28575;
	wire [4-1:0] node28577;
	wire [4-1:0] node28580;
	wire [4-1:0] node28581;
	wire [4-1:0] node28584;
	wire [4-1:0] node28586;
	wire [4-1:0] node28589;
	wire [4-1:0] node28590;
	wire [4-1:0] node28592;
	wire [4-1:0] node28595;
	wire [4-1:0] node28597;
	wire [4-1:0] node28599;
	wire [4-1:0] node28602;
	wire [4-1:0] node28603;
	wire [4-1:0] node28604;
	wire [4-1:0] node28605;
	wire [4-1:0] node28606;
	wire [4-1:0] node28607;
	wire [4-1:0] node28610;
	wire [4-1:0] node28613;
	wire [4-1:0] node28614;
	wire [4-1:0] node28616;
	wire [4-1:0] node28620;
	wire [4-1:0] node28621;
	wire [4-1:0] node28623;
	wire [4-1:0] node28626;
	wire [4-1:0] node28627;
	wire [4-1:0] node28630;
	wire [4-1:0] node28633;
	wire [4-1:0] node28634;
	wire [4-1:0] node28635;
	wire [4-1:0] node28636;
	wire [4-1:0] node28639;
	wire [4-1:0] node28642;
	wire [4-1:0] node28643;
	wire [4-1:0] node28646;
	wire [4-1:0] node28648;
	wire [4-1:0] node28651;
	wire [4-1:0] node28652;
	wire [4-1:0] node28653;
	wire [4-1:0] node28654;
	wire [4-1:0] node28658;
	wire [4-1:0] node28661;
	wire [4-1:0] node28663;
	wire [4-1:0] node28666;
	wire [4-1:0] node28667;
	wire [4-1:0] node28668;
	wire [4-1:0] node28669;
	wire [4-1:0] node28670;
	wire [4-1:0] node28671;
	wire [4-1:0] node28674;
	wire [4-1:0] node28678;
	wire [4-1:0] node28679;
	wire [4-1:0] node28682;
	wire [4-1:0] node28685;
	wire [4-1:0] node28686;
	wire [4-1:0] node28687;
	wire [4-1:0] node28690;
	wire [4-1:0] node28692;
	wire [4-1:0] node28695;
	wire [4-1:0] node28696;
	wire [4-1:0] node28700;
	wire [4-1:0] node28701;
	wire [4-1:0] node28702;
	wire [4-1:0] node28703;
	wire [4-1:0] node28705;
	wire [4-1:0] node28708;
	wire [4-1:0] node28709;
	wire [4-1:0] node28712;
	wire [4-1:0] node28715;
	wire [4-1:0] node28717;
	wire [4-1:0] node28720;
	wire [4-1:0] node28721;
	wire [4-1:0] node28722;
	wire [4-1:0] node28726;
	wire [4-1:0] node28729;
	wire [4-1:0] node28730;
	wire [4-1:0] node28731;
	wire [4-1:0] node28732;
	wire [4-1:0] node28733;
	wire [4-1:0] node28734;
	wire [4-1:0] node28735;
	wire [4-1:0] node28739;
	wire [4-1:0] node28740;
	wire [4-1:0] node28743;
	wire [4-1:0] node28746;
	wire [4-1:0] node28747;
	wire [4-1:0] node28748;
	wire [4-1:0] node28750;
	wire [4-1:0] node28753;
	wire [4-1:0] node28756;
	wire [4-1:0] node28757;
	wire [4-1:0] node28759;
	wire [4-1:0] node28763;
	wire [4-1:0] node28764;
	wire [4-1:0] node28765;
	wire [4-1:0] node28766;
	wire [4-1:0] node28767;
	wire [4-1:0] node28770;
	wire [4-1:0] node28774;
	wire [4-1:0] node28775;
	wire [4-1:0] node28776;
	wire [4-1:0] node28779;
	wire [4-1:0] node28782;
	wire [4-1:0] node28785;
	wire [4-1:0] node28786;
	wire [4-1:0] node28787;
	wire [4-1:0] node28789;
	wire [4-1:0] node28792;
	wire [4-1:0] node28795;
	wire [4-1:0] node28796;
	wire [4-1:0] node28799;
	wire [4-1:0] node28800;
	wire [4-1:0] node28804;
	wire [4-1:0] node28805;
	wire [4-1:0] node28806;
	wire [4-1:0] node28807;
	wire [4-1:0] node28808;
	wire [4-1:0] node28809;
	wire [4-1:0] node28813;
	wire [4-1:0] node28816;
	wire [4-1:0] node28818;
	wire [4-1:0] node28821;
	wire [4-1:0] node28822;
	wire [4-1:0] node28823;
	wire [4-1:0] node28824;
	wire [4-1:0] node28829;
	wire [4-1:0] node28832;
	wire [4-1:0] node28833;
	wire [4-1:0] node28834;
	wire [4-1:0] node28835;
	wire [4-1:0] node28836;
	wire [4-1:0] node28840;
	wire [4-1:0] node28843;
	wire [4-1:0] node28844;
	wire [4-1:0] node28846;
	wire [4-1:0] node28849;
	wire [4-1:0] node28851;
	wire [4-1:0] node28854;
	wire [4-1:0] node28855;
	wire [4-1:0] node28856;
	wire [4-1:0] node28858;
	wire [4-1:0] node28861;
	wire [4-1:0] node28864;
	wire [4-1:0] node28865;
	wire [4-1:0] node28868;
	wire [4-1:0] node28869;
	wire [4-1:0] node28872;
	wire [4-1:0] node28875;
	wire [4-1:0] node28876;
	wire [4-1:0] node28877;
	wire [4-1:0] node28878;
	wire [4-1:0] node28879;
	wire [4-1:0] node28880;
	wire [4-1:0] node28884;
	wire [4-1:0] node28885;
	wire [4-1:0] node28889;
	wire [4-1:0] node28890;
	wire [4-1:0] node28891;
	wire [4-1:0] node28894;
	wire [4-1:0] node28895;
	wire [4-1:0] node28899;
	wire [4-1:0] node28900;
	wire [4-1:0] node28902;
	wire [4-1:0] node28906;
	wire [4-1:0] node28907;
	wire [4-1:0] node28908;
	wire [4-1:0] node28909;
	wire [4-1:0] node28910;
	wire [4-1:0] node28915;
	wire [4-1:0] node28917;
	wire [4-1:0] node28920;
	wire [4-1:0] node28921;
	wire [4-1:0] node28922;
	wire [4-1:0] node28924;
	wire [4-1:0] node28927;
	wire [4-1:0] node28928;
	wire [4-1:0] node28931;
	wire [4-1:0] node28934;
	wire [4-1:0] node28935;
	wire [4-1:0] node28936;
	wire [4-1:0] node28939;
	wire [4-1:0] node28942;
	wire [4-1:0] node28943;
	wire [4-1:0] node28947;
	wire [4-1:0] node28948;
	wire [4-1:0] node28949;
	wire [4-1:0] node28950;
	wire [4-1:0] node28951;
	wire [4-1:0] node28954;
	wire [4-1:0] node28956;
	wire [4-1:0] node28959;
	wire [4-1:0] node28962;
	wire [4-1:0] node28963;
	wire [4-1:0] node28964;
	wire [4-1:0] node28967;
	wire [4-1:0] node28970;
	wire [4-1:0] node28971;
	wire [4-1:0] node28974;
	wire [4-1:0] node28975;
	wire [4-1:0] node28978;
	wire [4-1:0] node28981;
	wire [4-1:0] node28982;
	wire [4-1:0] node28983;
	wire [4-1:0] node28984;
	wire [4-1:0] node28987;
	wire [4-1:0] node28990;
	wire [4-1:0] node28991;
	wire [4-1:0] node28994;
	wire [4-1:0] node28997;
	wire [4-1:0] node28998;
	wire [4-1:0] node28999;
	wire [4-1:0] node29003;
	wire [4-1:0] node29004;
	wire [4-1:0] node29005;
	wire [4-1:0] node29009;
	wire [4-1:0] node29010;
	wire [4-1:0] node29014;
	wire [4-1:0] node29015;
	wire [4-1:0] node29016;
	wire [4-1:0] node29017;
	wire [4-1:0] node29018;
	wire [4-1:0] node29019;
	wire [4-1:0] node29020;
	wire [4-1:0] node29021;
	wire [4-1:0] node29025;
	wire [4-1:0] node29027;
	wire [4-1:0] node29030;
	wire [4-1:0] node29031;
	wire [4-1:0] node29033;
	wire [4-1:0] node29035;
	wire [4-1:0] node29038;
	wire [4-1:0] node29039;
	wire [4-1:0] node29041;
	wire [4-1:0] node29044;
	wire [4-1:0] node29046;
	wire [4-1:0] node29049;
	wire [4-1:0] node29050;
	wire [4-1:0] node29051;
	wire [4-1:0] node29052;
	wire [4-1:0] node29053;
	wire [4-1:0] node29056;
	wire [4-1:0] node29060;
	wire [4-1:0] node29061;
	wire [4-1:0] node29064;
	wire [4-1:0] node29067;
	wire [4-1:0] node29068;
	wire [4-1:0] node29069;
	wire [4-1:0] node29070;
	wire [4-1:0] node29075;
	wire [4-1:0] node29076;
	wire [4-1:0] node29078;
	wire [4-1:0] node29081;
	wire [4-1:0] node29083;
	wire [4-1:0] node29086;
	wire [4-1:0] node29087;
	wire [4-1:0] node29088;
	wire [4-1:0] node29089;
	wire [4-1:0] node29090;
	wire [4-1:0] node29091;
	wire [4-1:0] node29095;
	wire [4-1:0] node29098;
	wire [4-1:0] node29099;
	wire [4-1:0] node29102;
	wire [4-1:0] node29103;
	wire [4-1:0] node29107;
	wire [4-1:0] node29108;
	wire [4-1:0] node29109;
	wire [4-1:0] node29111;
	wire [4-1:0] node29114;
	wire [4-1:0] node29115;
	wire [4-1:0] node29118;
	wire [4-1:0] node29121;
	wire [4-1:0] node29122;
	wire [4-1:0] node29125;
	wire [4-1:0] node29126;
	wire [4-1:0] node29130;
	wire [4-1:0] node29131;
	wire [4-1:0] node29132;
	wire [4-1:0] node29134;
	wire [4-1:0] node29135;
	wire [4-1:0] node29138;
	wire [4-1:0] node29141;
	wire [4-1:0] node29142;
	wire [4-1:0] node29143;
	wire [4-1:0] node29146;
	wire [4-1:0] node29149;
	wire [4-1:0] node29150;
	wire [4-1:0] node29153;
	wire [4-1:0] node29156;
	wire [4-1:0] node29157;
	wire [4-1:0] node29158;
	wire [4-1:0] node29161;
	wire [4-1:0] node29163;
	wire [4-1:0] node29166;
	wire [4-1:0] node29167;
	wire [4-1:0] node29170;
	wire [4-1:0] node29173;
	wire [4-1:0] node29174;
	wire [4-1:0] node29175;
	wire [4-1:0] node29176;
	wire [4-1:0] node29177;
	wire [4-1:0] node29178;
	wire [4-1:0] node29180;
	wire [4-1:0] node29183;
	wire [4-1:0] node29186;
	wire [4-1:0] node29187;
	wire [4-1:0] node29190;
	wire [4-1:0] node29191;
	wire [4-1:0] node29195;
	wire [4-1:0] node29196;
	wire [4-1:0] node29197;
	wire [4-1:0] node29199;
	wire [4-1:0] node29202;
	wire [4-1:0] node29205;
	wire [4-1:0] node29206;
	wire [4-1:0] node29207;
	wire [4-1:0] node29211;
	wire [4-1:0] node29214;
	wire [4-1:0] node29215;
	wire [4-1:0] node29216;
	wire [4-1:0] node29217;
	wire [4-1:0] node29220;
	wire [4-1:0] node29222;
	wire [4-1:0] node29225;
	wire [4-1:0] node29226;
	wire [4-1:0] node29227;
	wire [4-1:0] node29231;
	wire [4-1:0] node29234;
	wire [4-1:0] node29235;
	wire [4-1:0] node29236;
	wire [4-1:0] node29239;
	wire [4-1:0] node29240;
	wire [4-1:0] node29244;
	wire [4-1:0] node29245;
	wire [4-1:0] node29246;
	wire [4-1:0] node29249;
	wire [4-1:0] node29252;
	wire [4-1:0] node29253;
	wire [4-1:0] node29257;
	wire [4-1:0] node29258;
	wire [4-1:0] node29259;
	wire [4-1:0] node29260;
	wire [4-1:0] node29261;
	wire [4-1:0] node29263;
	wire [4-1:0] node29267;
	wire [4-1:0] node29268;
	wire [4-1:0] node29271;
	wire [4-1:0] node29272;
	wire [4-1:0] node29276;
	wire [4-1:0] node29277;
	wire [4-1:0] node29279;
	wire [4-1:0] node29282;
	wire [4-1:0] node29283;
	wire [4-1:0] node29286;
	wire [4-1:0] node29288;
	wire [4-1:0] node29291;
	wire [4-1:0] node29292;
	wire [4-1:0] node29293;
	wire [4-1:0] node29295;
	wire [4-1:0] node29296;
	wire [4-1:0] node29300;
	wire [4-1:0] node29301;
	wire [4-1:0] node29305;
	wire [4-1:0] node29306;
	wire [4-1:0] node29307;
	wire [4-1:0] node29310;
	wire [4-1:0] node29313;
	wire [4-1:0] node29315;
	wire [4-1:0] node29316;
	wire [4-1:0] node29320;
	wire [4-1:0] node29321;
	wire [4-1:0] node29322;
	wire [4-1:0] node29323;
	wire [4-1:0] node29324;
	wire [4-1:0] node29325;
	wire [4-1:0] node29326;
	wire [4-1:0] node29329;
	wire [4-1:0] node29332;
	wire [4-1:0] node29333;
	wire [4-1:0] node29334;
	wire [4-1:0] node29338;
	wire [4-1:0] node29341;
	wire [4-1:0] node29342;
	wire [4-1:0] node29343;
	wire [4-1:0] node29345;
	wire [4-1:0] node29348;
	wire [4-1:0] node29349;
	wire [4-1:0] node29353;
	wire [4-1:0] node29354;
	wire [4-1:0] node29356;
	wire [4-1:0] node29359;
	wire [4-1:0] node29362;
	wire [4-1:0] node29363;
	wire [4-1:0] node29364;
	wire [4-1:0] node29365;
	wire [4-1:0] node29368;
	wire [4-1:0] node29370;
	wire [4-1:0] node29373;
	wire [4-1:0] node29374;
	wire [4-1:0] node29375;
	wire [4-1:0] node29379;
	wire [4-1:0] node29381;
	wire [4-1:0] node29384;
	wire [4-1:0] node29385;
	wire [4-1:0] node29386;
	wire [4-1:0] node29387;
	wire [4-1:0] node29391;
	wire [4-1:0] node29394;
	wire [4-1:0] node29396;
	wire [4-1:0] node29397;
	wire [4-1:0] node29401;
	wire [4-1:0] node29402;
	wire [4-1:0] node29403;
	wire [4-1:0] node29404;
	wire [4-1:0] node29405;
	wire [4-1:0] node29406;
	wire [4-1:0] node29410;
	wire [4-1:0] node29411;
	wire [4-1:0] node29415;
	wire [4-1:0] node29416;
	wire [4-1:0] node29420;
	wire [4-1:0] node29421;
	wire [4-1:0] node29422;
	wire [4-1:0] node29424;
	wire [4-1:0] node29427;
	wire [4-1:0] node29430;
	wire [4-1:0] node29431;
	wire [4-1:0] node29432;
	wire [4-1:0] node29436;
	wire [4-1:0] node29437;
	wire [4-1:0] node29441;
	wire [4-1:0] node29442;
	wire [4-1:0] node29443;
	wire [4-1:0] node29444;
	wire [4-1:0] node29445;
	wire [4-1:0] node29450;
	wire [4-1:0] node29451;
	wire [4-1:0] node29453;
	wire [4-1:0] node29457;
	wire [4-1:0] node29458;
	wire [4-1:0] node29459;
	wire [4-1:0] node29460;
	wire [4-1:0] node29464;
	wire [4-1:0] node29465;
	wire [4-1:0] node29469;
	wire [4-1:0] node29470;
	wire [4-1:0] node29472;
	wire [4-1:0] node29475;
	wire [4-1:0] node29478;
	wire [4-1:0] node29479;
	wire [4-1:0] node29480;
	wire [4-1:0] node29481;
	wire [4-1:0] node29482;
	wire [4-1:0] node29483;
	wire [4-1:0] node29486;
	wire [4-1:0] node29488;
	wire [4-1:0] node29491;
	wire [4-1:0] node29493;
	wire [4-1:0] node29496;
	wire [4-1:0] node29497;
	wire [4-1:0] node29499;
	wire [4-1:0] node29500;
	wire [4-1:0] node29504;
	wire [4-1:0] node29505;
	wire [4-1:0] node29507;
	wire [4-1:0] node29510;
	wire [4-1:0] node29512;
	wire [4-1:0] node29515;
	wire [4-1:0] node29516;
	wire [4-1:0] node29517;
	wire [4-1:0] node29518;
	wire [4-1:0] node29520;
	wire [4-1:0] node29523;
	wire [4-1:0] node29524;
	wire [4-1:0] node29528;
	wire [4-1:0] node29529;
	wire [4-1:0] node29533;
	wire [4-1:0] node29534;
	wire [4-1:0] node29537;
	wire [4-1:0] node29538;
	wire [4-1:0] node29542;
	wire [4-1:0] node29543;
	wire [4-1:0] node29544;
	wire [4-1:0] node29545;
	wire [4-1:0] node29547;
	wire [4-1:0] node29549;
	wire [4-1:0] node29552;
	wire [4-1:0] node29554;
	wire [4-1:0] node29555;
	wire [4-1:0] node29559;
	wire [4-1:0] node29560;
	wire [4-1:0] node29561;
	wire [4-1:0] node29562;
	wire [4-1:0] node29566;
	wire [4-1:0] node29568;
	wire [4-1:0] node29571;
	wire [4-1:0] node29572;
	wire [4-1:0] node29574;
	wire [4-1:0] node29577;
	wire [4-1:0] node29580;
	wire [4-1:0] node29581;
	wire [4-1:0] node29582;
	wire [4-1:0] node29583;
	wire [4-1:0] node29587;
	wire [4-1:0] node29589;
	wire [4-1:0] node29590;
	wire [4-1:0] node29593;
	wire [4-1:0] node29596;
	wire [4-1:0] node29597;
	wire [4-1:0] node29600;
	wire [4-1:0] node29601;
	wire [4-1:0] node29604;
	wire [4-1:0] node29607;
	wire [4-1:0] node29608;
	wire [4-1:0] node29609;
	wire [4-1:0] node29610;
	wire [4-1:0] node29611;
	wire [4-1:0] node29612;
	wire [4-1:0] node29613;
	wire [4-1:0] node29614;
	wire [4-1:0] node29615;
	wire [4-1:0] node29618;
	wire [4-1:0] node29621;
	wire [4-1:0] node29623;
	wire [4-1:0] node29624;
	wire [4-1:0] node29627;
	wire [4-1:0] node29630;
	wire [4-1:0] node29631;
	wire [4-1:0] node29633;
	wire [4-1:0] node29636;
	wire [4-1:0] node29637;
	wire [4-1:0] node29640;
	wire [4-1:0] node29643;
	wire [4-1:0] node29644;
	wire [4-1:0] node29645;
	wire [4-1:0] node29646;
	wire [4-1:0] node29647;
	wire [4-1:0] node29650;
	wire [4-1:0] node29653;
	wire [4-1:0] node29655;
	wire [4-1:0] node29658;
	wire [4-1:0] node29660;
	wire [4-1:0] node29662;
	wire [4-1:0] node29665;
	wire [4-1:0] node29666;
	wire [4-1:0] node29667;
	wire [4-1:0] node29670;
	wire [4-1:0] node29673;
	wire [4-1:0] node29674;
	wire [4-1:0] node29677;
	wire [4-1:0] node29680;
	wire [4-1:0] node29681;
	wire [4-1:0] node29682;
	wire [4-1:0] node29683;
	wire [4-1:0] node29684;
	wire [4-1:0] node29688;
	wire [4-1:0] node29689;
	wire [4-1:0] node29693;
	wire [4-1:0] node29695;
	wire [4-1:0] node29696;
	wire [4-1:0] node29697;
	wire [4-1:0] node29701;
	wire [4-1:0] node29704;
	wire [4-1:0] node29705;
	wire [4-1:0] node29706;
	wire [4-1:0] node29707;
	wire [4-1:0] node29710;
	wire [4-1:0] node29713;
	wire [4-1:0] node29715;
	wire [4-1:0] node29716;
	wire [4-1:0] node29720;
	wire [4-1:0] node29721;
	wire [4-1:0] node29722;
	wire [4-1:0] node29725;
	wire [4-1:0] node29728;
	wire [4-1:0] node29729;
	wire [4-1:0] node29733;
	wire [4-1:0] node29734;
	wire [4-1:0] node29735;
	wire [4-1:0] node29736;
	wire [4-1:0] node29737;
	wire [4-1:0] node29739;
	wire [4-1:0] node29742;
	wire [4-1:0] node29743;
	wire [4-1:0] node29746;
	wire [4-1:0] node29748;
	wire [4-1:0] node29751;
	wire [4-1:0] node29752;
	wire [4-1:0] node29753;
	wire [4-1:0] node29754;
	wire [4-1:0] node29758;
	wire [4-1:0] node29760;
	wire [4-1:0] node29763;
	wire [4-1:0] node29765;
	wire [4-1:0] node29766;
	wire [4-1:0] node29770;
	wire [4-1:0] node29771;
	wire [4-1:0] node29772;
	wire [4-1:0] node29773;
	wire [4-1:0] node29774;
	wire [4-1:0] node29778;
	wire [4-1:0] node29781;
	wire [4-1:0] node29782;
	wire [4-1:0] node29785;
	wire [4-1:0] node29787;
	wire [4-1:0] node29790;
	wire [4-1:0] node29791;
	wire [4-1:0] node29792;
	wire [4-1:0] node29795;
	wire [4-1:0] node29798;
	wire [4-1:0] node29800;
	wire [4-1:0] node29801;
	wire [4-1:0] node29804;
	wire [4-1:0] node29807;
	wire [4-1:0] node29808;
	wire [4-1:0] node29809;
	wire [4-1:0] node29810;
	wire [4-1:0] node29811;
	wire [4-1:0] node29813;
	wire [4-1:0] node29816;
	wire [4-1:0] node29817;
	wire [4-1:0] node29821;
	wire [4-1:0] node29822;
	wire [4-1:0] node29824;
	wire [4-1:0] node29828;
	wire [4-1:0] node29829;
	wire [4-1:0] node29830;
	wire [4-1:0] node29833;
	wire [4-1:0] node29836;
	wire [4-1:0] node29837;
	wire [4-1:0] node29838;
	wire [4-1:0] node29841;
	wire [4-1:0] node29845;
	wire [4-1:0] node29846;
	wire [4-1:0] node29847;
	wire [4-1:0] node29848;
	wire [4-1:0] node29849;
	wire [4-1:0] node29852;
	wire [4-1:0] node29855;
	wire [4-1:0] node29856;
	wire [4-1:0] node29859;
	wire [4-1:0] node29862;
	wire [4-1:0] node29864;
	wire [4-1:0] node29865;
	wire [4-1:0] node29868;
	wire [4-1:0] node29871;
	wire [4-1:0] node29872;
	wire [4-1:0] node29875;
	wire [4-1:0] node29878;
	wire [4-1:0] node29879;
	wire [4-1:0] node29880;
	wire [4-1:0] node29881;
	wire [4-1:0] node29882;
	wire [4-1:0] node29883;
	wire [4-1:0] node29885;
	wire [4-1:0] node29888;
	wire [4-1:0] node29890;
	wire [4-1:0] node29893;
	wire [4-1:0] node29894;
	wire [4-1:0] node29898;
	wire [4-1:0] node29899;
	wire [4-1:0] node29900;
	wire [4-1:0] node29901;
	wire [4-1:0] node29905;
	wire [4-1:0] node29906;
	wire [4-1:0] node29910;
	wire [4-1:0] node29911;
	wire [4-1:0] node29912;
	wire [4-1:0] node29916;
	wire [4-1:0] node29917;
	wire [4-1:0] node29921;
	wire [4-1:0] node29922;
	wire [4-1:0] node29923;
	wire [4-1:0] node29924;
	wire [4-1:0] node29925;
	wire [4-1:0] node29929;
	wire [4-1:0] node29930;
	wire [4-1:0] node29933;
	wire [4-1:0] node29936;
	wire [4-1:0] node29937;
	wire [4-1:0] node29940;
	wire [4-1:0] node29943;
	wire [4-1:0] node29944;
	wire [4-1:0] node29945;
	wire [4-1:0] node29947;
	wire [4-1:0] node29950;
	wire [4-1:0] node29953;
	wire [4-1:0] node29954;
	wire [4-1:0] node29956;
	wire [4-1:0] node29959;
	wire [4-1:0] node29961;
	wire [4-1:0] node29964;
	wire [4-1:0] node29965;
	wire [4-1:0] node29966;
	wire [4-1:0] node29967;
	wire [4-1:0] node29968;
	wire [4-1:0] node29969;
	wire [4-1:0] node29970;
	wire [4-1:0] node29973;
	wire [4-1:0] node29976;
	wire [4-1:0] node29977;
	wire [4-1:0] node29981;
	wire [4-1:0] node29982;
	wire [4-1:0] node29986;
	wire [4-1:0] node29987;
	wire [4-1:0] node29988;
	wire [4-1:0] node29989;
	wire [4-1:0] node29993;
	wire [4-1:0] node29994;
	wire [4-1:0] node29997;
	wire [4-1:0] node30000;
	wire [4-1:0] node30001;
	wire [4-1:0] node30002;
	wire [4-1:0] node30006;
	wire [4-1:0] node30007;
	wire [4-1:0] node30011;
	wire [4-1:0] node30012;
	wire [4-1:0] node30013;
	wire [4-1:0] node30014;
	wire [4-1:0] node30016;
	wire [4-1:0] node30019;
	wire [4-1:0] node30020;
	wire [4-1:0] node30024;
	wire [4-1:0] node30025;
	wire [4-1:0] node30026;
	wire [4-1:0] node30029;
	wire [4-1:0] node30032;
	wire [4-1:0] node30034;
	wire [4-1:0] node30037;
	wire [4-1:0] node30038;
	wire [4-1:0] node30040;
	wire [4-1:0] node30043;
	wire [4-1:0] node30044;
	wire [4-1:0] node30046;
	wire [4-1:0] node30049;
	wire [4-1:0] node30050;
	wire [4-1:0] node30053;
	wire [4-1:0] node30056;
	wire [4-1:0] node30057;
	wire [4-1:0] node30058;
	wire [4-1:0] node30059;
	wire [4-1:0] node30062;
	wire [4-1:0] node30065;
	wire [4-1:0] node30066;
	wire [4-1:0] node30067;
	wire [4-1:0] node30070;
	wire [4-1:0] node30073;
	wire [4-1:0] node30076;
	wire [4-1:0] node30077;
	wire [4-1:0] node30078;
	wire [4-1:0] node30080;
	wire [4-1:0] node30083;
	wire [4-1:0] node30086;
	wire [4-1:0] node30087;
	wire [4-1:0] node30088;
	wire [4-1:0] node30091;
	wire [4-1:0] node30094;
	wire [4-1:0] node30096;
	wire [4-1:0] node30099;
	wire [4-1:0] node30100;
	wire [4-1:0] node30101;
	wire [4-1:0] node30102;
	wire [4-1:0] node30103;
	wire [4-1:0] node30104;
	wire [4-1:0] node30105;
	wire [4-1:0] node30108;
	wire [4-1:0] node30110;
	wire [4-1:0] node30113;
	wire [4-1:0] node30114;
	wire [4-1:0] node30116;
	wire [4-1:0] node30118;
	wire [4-1:0] node30121;
	wire [4-1:0] node30123;
	wire [4-1:0] node30126;
	wire [4-1:0] node30127;
	wire [4-1:0] node30129;
	wire [4-1:0] node30132;
	wire [4-1:0] node30134;
	wire [4-1:0] node30135;
	wire [4-1:0] node30139;
	wire [4-1:0] node30140;
	wire [4-1:0] node30141;
	wire [4-1:0] node30142;
	wire [4-1:0] node30143;
	wire [4-1:0] node30147;
	wire [4-1:0] node30150;
	wire [4-1:0] node30151;
	wire [4-1:0] node30152;
	wire [4-1:0] node30153;
	wire [4-1:0] node30158;
	wire [4-1:0] node30160;
	wire [4-1:0] node30163;
	wire [4-1:0] node30164;
	wire [4-1:0] node30165;
	wire [4-1:0] node30166;
	wire [4-1:0] node30169;
	wire [4-1:0] node30172;
	wire [4-1:0] node30173;
	wire [4-1:0] node30174;
	wire [4-1:0] node30178;
	wire [4-1:0] node30179;
	wire [4-1:0] node30182;
	wire [4-1:0] node30185;
	wire [4-1:0] node30187;
	wire [4-1:0] node30188;
	wire [4-1:0] node30189;
	wire [4-1:0] node30192;
	wire [4-1:0] node30195;
	wire [4-1:0] node30197;
	wire [4-1:0] node30200;
	wire [4-1:0] node30201;
	wire [4-1:0] node30202;
	wire [4-1:0] node30203;
	wire [4-1:0] node30204;
	wire [4-1:0] node30206;
	wire [4-1:0] node30209;
	wire [4-1:0] node30211;
	wire [4-1:0] node30214;
	wire [4-1:0] node30215;
	wire [4-1:0] node30219;
	wire [4-1:0] node30220;
	wire [4-1:0] node30221;
	wire [4-1:0] node30222;
	wire [4-1:0] node30226;
	wire [4-1:0] node30228;
	wire [4-1:0] node30231;
	wire [4-1:0] node30232;
	wire [4-1:0] node30234;
	wire [4-1:0] node30237;
	wire [4-1:0] node30238;
	wire [4-1:0] node30242;
	wire [4-1:0] node30243;
	wire [4-1:0] node30244;
	wire [4-1:0] node30245;
	wire [4-1:0] node30248;
	wire [4-1:0] node30251;
	wire [4-1:0] node30252;
	wire [4-1:0] node30253;
	wire [4-1:0] node30256;
	wire [4-1:0] node30259;
	wire [4-1:0] node30260;
	wire [4-1:0] node30261;
	wire [4-1:0] node30264;
	wire [4-1:0] node30267;
	wire [4-1:0] node30268;
	wire [4-1:0] node30271;
	wire [4-1:0] node30274;
	wire [4-1:0] node30275;
	wire [4-1:0] node30276;
	wire [4-1:0] node30277;
	wire [4-1:0] node30281;
	wire [4-1:0] node30282;
	wire [4-1:0] node30286;
	wire [4-1:0] node30287;
	wire [4-1:0] node30288;
	wire [4-1:0] node30289;
	wire [4-1:0] node30293;
	wire [4-1:0] node30294;
	wire [4-1:0] node30297;
	wire [4-1:0] node30301;
	wire [4-1:0] node30302;
	wire [4-1:0] node30303;
	wire [4-1:0] node30304;
	wire [4-1:0] node30305;
	wire [4-1:0] node30306;
	wire [4-1:0] node30307;
	wire [4-1:0] node30310;
	wire [4-1:0] node30314;
	wire [4-1:0] node30315;
	wire [4-1:0] node30316;
	wire [4-1:0] node30317;
	wire [4-1:0] node30320;
	wire [4-1:0] node30323;
	wire [4-1:0] node30324;
	wire [4-1:0] node30327;
	wire [4-1:0] node30331;
	wire [4-1:0] node30332;
	wire [4-1:0] node30333;
	wire [4-1:0] node30334;
	wire [4-1:0] node30339;
	wire [4-1:0] node30340;
	wire [4-1:0] node30341;
	wire [4-1:0] node30344;
	wire [4-1:0] node30348;
	wire [4-1:0] node30349;
	wire [4-1:0] node30350;
	wire [4-1:0] node30351;
	wire [4-1:0] node30353;
	wire [4-1:0] node30356;
	wire [4-1:0] node30358;
	wire [4-1:0] node30360;
	wire [4-1:0] node30363;
	wire [4-1:0] node30364;
	wire [4-1:0] node30365;
	wire [4-1:0] node30366;
	wire [4-1:0] node30369;
	wire [4-1:0] node30372;
	wire [4-1:0] node30373;
	wire [4-1:0] node30377;
	wire [4-1:0] node30378;
	wire [4-1:0] node30379;
	wire [4-1:0] node30382;
	wire [4-1:0] node30386;
	wire [4-1:0] node30387;
	wire [4-1:0] node30388;
	wire [4-1:0] node30389;
	wire [4-1:0] node30391;
	wire [4-1:0] node30394;
	wire [4-1:0] node30395;
	wire [4-1:0] node30398;
	wire [4-1:0] node30401;
	wire [4-1:0] node30402;
	wire [4-1:0] node30403;
	wire [4-1:0] node30406;
	wire [4-1:0] node30409;
	wire [4-1:0] node30410;
	wire [4-1:0] node30413;
	wire [4-1:0] node30416;
	wire [4-1:0] node30417;
	wire [4-1:0] node30420;
	wire [4-1:0] node30423;
	wire [4-1:0] node30424;
	wire [4-1:0] node30425;
	wire [4-1:0] node30426;
	wire [4-1:0] node30427;
	wire [4-1:0] node30428;
	wire [4-1:0] node30431;
	wire [4-1:0] node30434;
	wire [4-1:0] node30435;
	wire [4-1:0] node30438;
	wire [4-1:0] node30441;
	wire [4-1:0] node30443;
	wire [4-1:0] node30446;
	wire [4-1:0] node30447;
	wire [4-1:0] node30448;
	wire [4-1:0] node30449;
	wire [4-1:0] node30451;
	wire [4-1:0] node30454;
	wire [4-1:0] node30456;
	wire [4-1:0] node30459;
	wire [4-1:0] node30460;
	wire [4-1:0] node30462;
	wire [4-1:0] node30465;
	wire [4-1:0] node30468;
	wire [4-1:0] node30469;
	wire [4-1:0] node30472;
	wire [4-1:0] node30475;
	wire [4-1:0] node30476;
	wire [4-1:0] node30477;
	wire [4-1:0] node30478;
	wire [4-1:0] node30479;
	wire [4-1:0] node30482;
	wire [4-1:0] node30485;
	wire [4-1:0] node30486;
	wire [4-1:0] node30490;
	wire [4-1:0] node30492;
	wire [4-1:0] node30493;
	wire [4-1:0] node30494;
	wire [4-1:0] node30497;
	wire [4-1:0] node30500;
	wire [4-1:0] node30502;
	wire [4-1:0] node30505;
	wire [4-1:0] node30506;
	wire [4-1:0] node30507;
	wire [4-1:0] node30510;
	wire [4-1:0] node30513;
	wire [4-1:0] node30514;
	wire [4-1:0] node30517;
	wire [4-1:0] node30520;
	wire [4-1:0] node30521;
	wire [4-1:0] node30522;
	wire [4-1:0] node30523;
	wire [4-1:0] node30524;
	wire [4-1:0] node30525;
	wire [4-1:0] node30526;
	wire [4-1:0] node30527;
	wire [4-1:0] node30528;
	wire [4-1:0] node30529;
	wire [4-1:0] node30531;
	wire [4-1:0] node30533;
	wire [4-1:0] node30536;
	wire [4-1:0] node30537;
	wire [4-1:0] node30538;
	wire [4-1:0] node30541;
	wire [4-1:0] node30544;
	wire [4-1:0] node30545;
	wire [4-1:0] node30548;
	wire [4-1:0] node30551;
	wire [4-1:0] node30552;
	wire [4-1:0] node30553;
	wire [4-1:0] node30555;
	wire [4-1:0] node30558;
	wire [4-1:0] node30559;
	wire [4-1:0] node30563;
	wire [4-1:0] node30564;
	wire [4-1:0] node30567;
	wire [4-1:0] node30570;
	wire [4-1:0] node30571;
	wire [4-1:0] node30572;
	wire [4-1:0] node30574;
	wire [4-1:0] node30577;
	wire [4-1:0] node30578;
	wire [4-1:0] node30579;
	wire [4-1:0] node30583;
	wire [4-1:0] node30584;
	wire [4-1:0] node30588;
	wire [4-1:0] node30589;
	wire [4-1:0] node30591;
	wire [4-1:0] node30592;
	wire [4-1:0] node30595;
	wire [4-1:0] node30598;
	wire [4-1:0] node30599;
	wire [4-1:0] node30600;
	wire [4-1:0] node30603;
	wire [4-1:0] node30606;
	wire [4-1:0] node30607;
	wire [4-1:0] node30610;
	wire [4-1:0] node30613;
	wire [4-1:0] node30614;
	wire [4-1:0] node30615;
	wire [4-1:0] node30616;
	wire [4-1:0] node30617;
	wire [4-1:0] node30618;
	wire [4-1:0] node30623;
	wire [4-1:0] node30624;
	wire [4-1:0] node30625;
	wire [4-1:0] node30629;
	wire [4-1:0] node30631;
	wire [4-1:0] node30634;
	wire [4-1:0] node30635;
	wire [4-1:0] node30636;
	wire [4-1:0] node30640;
	wire [4-1:0] node30643;
	wire [4-1:0] node30644;
	wire [4-1:0] node30645;
	wire [4-1:0] node30646;
	wire [4-1:0] node30649;
	wire [4-1:0] node30652;
	wire [4-1:0] node30653;
	wire [4-1:0] node30656;
	wire [4-1:0] node30659;
	wire [4-1:0] node30660;
	wire [4-1:0] node30661;
	wire [4-1:0] node30662;
	wire [4-1:0] node30665;
	wire [4-1:0] node30668;
	wire [4-1:0] node30669;
	wire [4-1:0] node30672;
	wire [4-1:0] node30675;
	wire [4-1:0] node30677;
	wire [4-1:0] node30678;
	wire [4-1:0] node30681;
	wire [4-1:0] node30684;
	wire [4-1:0] node30685;
	wire [4-1:0] node30686;
	wire [4-1:0] node30687;
	wire [4-1:0] node30688;
	wire [4-1:0] node30689;
	wire [4-1:0] node30691;
	wire [4-1:0] node30694;
	wire [4-1:0] node30697;
	wire [4-1:0] node30698;
	wire [4-1:0] node30699;
	wire [4-1:0] node30703;
	wire [4-1:0] node30706;
	wire [4-1:0] node30707;
	wire [4-1:0] node30708;
	wire [4-1:0] node30712;
	wire [4-1:0] node30713;
	wire [4-1:0] node30717;
	wire [4-1:0] node30718;
	wire [4-1:0] node30719;
	wire [4-1:0] node30720;
	wire [4-1:0] node30722;
	wire [4-1:0] node30725;
	wire [4-1:0] node30727;
	wire [4-1:0] node30730;
	wire [4-1:0] node30731;
	wire [4-1:0] node30732;
	wire [4-1:0] node30736;
	wire [4-1:0] node30737;
	wire [4-1:0] node30740;
	wire [4-1:0] node30743;
	wire [4-1:0] node30744;
	wire [4-1:0] node30745;
	wire [4-1:0] node30747;
	wire [4-1:0] node30750;
	wire [4-1:0] node30753;
	wire [4-1:0] node30754;
	wire [4-1:0] node30755;
	wire [4-1:0] node30758;
	wire [4-1:0] node30762;
	wire [4-1:0] node30763;
	wire [4-1:0] node30764;
	wire [4-1:0] node30765;
	wire [4-1:0] node30766;
	wire [4-1:0] node30767;
	wire [4-1:0] node30771;
	wire [4-1:0] node30772;
	wire [4-1:0] node30776;
	wire [4-1:0] node30777;
	wire [4-1:0] node30781;
	wire [4-1:0] node30782;
	wire [4-1:0] node30783;
	wire [4-1:0] node30784;
	wire [4-1:0] node30787;
	wire [4-1:0] node30790;
	wire [4-1:0] node30791;
	wire [4-1:0] node30794;
	wire [4-1:0] node30797;
	wire [4-1:0] node30798;
	wire [4-1:0] node30799;
	wire [4-1:0] node30802;
	wire [4-1:0] node30806;
	wire [4-1:0] node30807;
	wire [4-1:0] node30808;
	wire [4-1:0] node30809;
	wire [4-1:0] node30813;
	wire [4-1:0] node30814;
	wire [4-1:0] node30815;
	wire [4-1:0] node30818;
	wire [4-1:0] node30822;
	wire [4-1:0] node30823;
	wire [4-1:0] node30825;
	wire [4-1:0] node30828;
	wire [4-1:0] node30829;
	wire [4-1:0] node30830;
	wire [4-1:0] node30833;
	wire [4-1:0] node30837;
	wire [4-1:0] node30838;
	wire [4-1:0] node30839;
	wire [4-1:0] node30840;
	wire [4-1:0] node30841;
	wire [4-1:0] node30842;
	wire [4-1:0] node30843;
	wire [4-1:0] node30845;
	wire [4-1:0] node30848;
	wire [4-1:0] node30851;
	wire [4-1:0] node30852;
	wire [4-1:0] node30854;
	wire [4-1:0] node30857;
	wire [4-1:0] node30860;
	wire [4-1:0] node30861;
	wire [4-1:0] node30862;
	wire [4-1:0] node30864;
	wire [4-1:0] node30868;
	wire [4-1:0] node30869;
	wire [4-1:0] node30873;
	wire [4-1:0] node30874;
	wire [4-1:0] node30875;
	wire [4-1:0] node30876;
	wire [4-1:0] node30877;
	wire [4-1:0] node30880;
	wire [4-1:0] node30884;
	wire [4-1:0] node30885;
	wire [4-1:0] node30889;
	wire [4-1:0] node30890;
	wire [4-1:0] node30891;
	wire [4-1:0] node30892;
	wire [4-1:0] node30895;
	wire [4-1:0] node30898;
	wire [4-1:0] node30899;
	wire [4-1:0] node30903;
	wire [4-1:0] node30904;
	wire [4-1:0] node30907;
	wire [4-1:0] node30910;
	wire [4-1:0] node30911;
	wire [4-1:0] node30912;
	wire [4-1:0] node30913;
	wire [4-1:0] node30914;
	wire [4-1:0] node30915;
	wire [4-1:0] node30919;
	wire [4-1:0] node30921;
	wire [4-1:0] node30924;
	wire [4-1:0] node30925;
	wire [4-1:0] node30926;
	wire [4-1:0] node30929;
	wire [4-1:0] node30932;
	wire [4-1:0] node30933;
	wire [4-1:0] node30937;
	wire [4-1:0] node30938;
	wire [4-1:0] node30939;
	wire [4-1:0] node30940;
	wire [4-1:0] node30945;
	wire [4-1:0] node30947;
	wire [4-1:0] node30950;
	wire [4-1:0] node30951;
	wire [4-1:0] node30952;
	wire [4-1:0] node30954;
	wire [4-1:0] node30955;
	wire [4-1:0] node30958;
	wire [4-1:0] node30961;
	wire [4-1:0] node30962;
	wire [4-1:0] node30963;
	wire [4-1:0] node30966;
	wire [4-1:0] node30969;
	wire [4-1:0] node30970;
	wire [4-1:0] node30973;
	wire [4-1:0] node30976;
	wire [4-1:0] node30977;
	wire [4-1:0] node30978;
	wire [4-1:0] node30979;
	wire [4-1:0] node30983;
	wire [4-1:0] node30986;
	wire [4-1:0] node30987;
	wire [4-1:0] node30990;
	wire [4-1:0] node30992;
	wire [4-1:0] node30995;
	wire [4-1:0] node30996;
	wire [4-1:0] node30997;
	wire [4-1:0] node30998;
	wire [4-1:0] node30999;
	wire [4-1:0] node31000;
	wire [4-1:0] node31003;
	wire [4-1:0] node31006;
	wire [4-1:0] node31008;
	wire [4-1:0] node31010;
	wire [4-1:0] node31013;
	wire [4-1:0] node31014;
	wire [4-1:0] node31015;
	wire [4-1:0] node31016;
	wire [4-1:0] node31019;
	wire [4-1:0] node31022;
	wire [4-1:0] node31024;
	wire [4-1:0] node31027;
	wire [4-1:0] node31029;
	wire [4-1:0] node31032;
	wire [4-1:0] node31033;
	wire [4-1:0] node31034;
	wire [4-1:0] node31035;
	wire [4-1:0] node31036;
	wire [4-1:0] node31040;
	wire [4-1:0] node31042;
	wire [4-1:0] node31045;
	wire [4-1:0] node31046;
	wire [4-1:0] node31047;
	wire [4-1:0] node31051;
	wire [4-1:0] node31052;
	wire [4-1:0] node31056;
	wire [4-1:0] node31057;
	wire [4-1:0] node31058;
	wire [4-1:0] node31059;
	wire [4-1:0] node31063;
	wire [4-1:0] node31066;
	wire [4-1:0] node31067;
	wire [4-1:0] node31069;
	wire [4-1:0] node31073;
	wire [4-1:0] node31074;
	wire [4-1:0] node31075;
	wire [4-1:0] node31076;
	wire [4-1:0] node31077;
	wire [4-1:0] node31078;
	wire [4-1:0] node31082;
	wire [4-1:0] node31083;
	wire [4-1:0] node31087;
	wire [4-1:0] node31088;
	wire [4-1:0] node31091;
	wire [4-1:0] node31093;
	wire [4-1:0] node31096;
	wire [4-1:0] node31097;
	wire [4-1:0] node31098;
	wire [4-1:0] node31100;
	wire [4-1:0] node31103;
	wire [4-1:0] node31106;
	wire [4-1:0] node31107;
	wire [4-1:0] node31108;
	wire [4-1:0] node31112;
	wire [4-1:0] node31113;
	wire [4-1:0] node31117;
	wire [4-1:0] node31118;
	wire [4-1:0] node31119;
	wire [4-1:0] node31121;
	wire [4-1:0] node31124;
	wire [4-1:0] node31125;
	wire [4-1:0] node31128;
	wire [4-1:0] node31131;
	wire [4-1:0] node31132;
	wire [4-1:0] node31133;
	wire [4-1:0] node31136;
	wire [4-1:0] node31139;
	wire [4-1:0] node31140;
	wire [4-1:0] node31143;
	wire [4-1:0] node31146;
	wire [4-1:0] node31147;
	wire [4-1:0] node31148;
	wire [4-1:0] node31149;
	wire [4-1:0] node31150;
	wire [4-1:0] node31151;
	wire [4-1:0] node31152;
	wire [4-1:0] node31153;
	wire [4-1:0] node31154;
	wire [4-1:0] node31157;
	wire [4-1:0] node31161;
	wire [4-1:0] node31162;
	wire [4-1:0] node31164;
	wire [4-1:0] node31167;
	wire [4-1:0] node31168;
	wire [4-1:0] node31171;
	wire [4-1:0] node31174;
	wire [4-1:0] node31175;
	wire [4-1:0] node31176;
	wire [4-1:0] node31178;
	wire [4-1:0] node31181;
	wire [4-1:0] node31183;
	wire [4-1:0] node31186;
	wire [4-1:0] node31187;
	wire [4-1:0] node31190;
	wire [4-1:0] node31193;
	wire [4-1:0] node31194;
	wire [4-1:0] node31195;
	wire [4-1:0] node31196;
	wire [4-1:0] node31197;
	wire [4-1:0] node31201;
	wire [4-1:0] node31203;
	wire [4-1:0] node31206;
	wire [4-1:0] node31208;
	wire [4-1:0] node31209;
	wire [4-1:0] node31213;
	wire [4-1:0] node31214;
	wire [4-1:0] node31215;
	wire [4-1:0] node31217;
	wire [4-1:0] node31220;
	wire [4-1:0] node31221;
	wire [4-1:0] node31224;
	wire [4-1:0] node31227;
	wire [4-1:0] node31228;
	wire [4-1:0] node31230;
	wire [4-1:0] node31233;
	wire [4-1:0] node31234;
	wire [4-1:0] node31237;
	wire [4-1:0] node31240;
	wire [4-1:0] node31241;
	wire [4-1:0] node31242;
	wire [4-1:0] node31243;
	wire [4-1:0] node31245;
	wire [4-1:0] node31248;
	wire [4-1:0] node31249;
	wire [4-1:0] node31251;
	wire [4-1:0] node31254;
	wire [4-1:0] node31256;
	wire [4-1:0] node31259;
	wire [4-1:0] node31260;
	wire [4-1:0] node31261;
	wire [4-1:0] node31262;
	wire [4-1:0] node31265;
	wire [4-1:0] node31268;
	wire [4-1:0] node31269;
	wire [4-1:0] node31272;
	wire [4-1:0] node31275;
	wire [4-1:0] node31276;
	wire [4-1:0] node31279;
	wire [4-1:0] node31282;
	wire [4-1:0] node31283;
	wire [4-1:0] node31284;
	wire [4-1:0] node31285;
	wire [4-1:0] node31286;
	wire [4-1:0] node31290;
	wire [4-1:0] node31293;
	wire [4-1:0] node31294;
	wire [4-1:0] node31297;
	wire [4-1:0] node31299;
	wire [4-1:0] node31302;
	wire [4-1:0] node31303;
	wire [4-1:0] node31304;
	wire [4-1:0] node31305;
	wire [4-1:0] node31309;
	wire [4-1:0] node31311;
	wire [4-1:0] node31314;
	wire [4-1:0] node31315;
	wire [4-1:0] node31318;
	wire [4-1:0] node31319;
	wire [4-1:0] node31323;
	wire [4-1:0] node31324;
	wire [4-1:0] node31325;
	wire [4-1:0] node31326;
	wire [4-1:0] node31327;
	wire [4-1:0] node31328;
	wire [4-1:0] node31331;
	wire [4-1:0] node31332;
	wire [4-1:0] node31336;
	wire [4-1:0] node31338;
	wire [4-1:0] node31339;
	wire [4-1:0] node31342;
	wire [4-1:0] node31345;
	wire [4-1:0] node31346;
	wire [4-1:0] node31348;
	wire [4-1:0] node31349;
	wire [4-1:0] node31353;
	wire [4-1:0] node31354;
	wire [4-1:0] node31355;
	wire [4-1:0] node31358;
	wire [4-1:0] node31361;
	wire [4-1:0] node31362;
	wire [4-1:0] node31365;
	wire [4-1:0] node31368;
	wire [4-1:0] node31369;
	wire [4-1:0] node31370;
	wire [4-1:0] node31371;
	wire [4-1:0] node31373;
	wire [4-1:0] node31377;
	wire [4-1:0] node31379;
	wire [4-1:0] node31381;
	wire [4-1:0] node31384;
	wire [4-1:0] node31385;
	wire [4-1:0] node31386;
	wire [4-1:0] node31390;
	wire [4-1:0] node31391;
	wire [4-1:0] node31392;
	wire [4-1:0] node31396;
	wire [4-1:0] node31397;
	wire [4-1:0] node31401;
	wire [4-1:0] node31402;
	wire [4-1:0] node31403;
	wire [4-1:0] node31404;
	wire [4-1:0] node31405;
	wire [4-1:0] node31408;
	wire [4-1:0] node31410;
	wire [4-1:0] node31413;
	wire [4-1:0] node31414;
	wire [4-1:0] node31417;
	wire [4-1:0] node31419;
	wire [4-1:0] node31422;
	wire [4-1:0] node31423;
	wire [4-1:0] node31425;
	wire [4-1:0] node31427;
	wire [4-1:0] node31430;
	wire [4-1:0] node31431;
	wire [4-1:0] node31432;
	wire [4-1:0] node31435;
	wire [4-1:0] node31438;
	wire [4-1:0] node31439;
	wire [4-1:0] node31442;
	wire [4-1:0] node31445;
	wire [4-1:0] node31446;
	wire [4-1:0] node31447;
	wire [4-1:0] node31448;
	wire [4-1:0] node31449;
	wire [4-1:0] node31453;
	wire [4-1:0] node31454;
	wire [4-1:0] node31457;
	wire [4-1:0] node31460;
	wire [4-1:0] node31461;
	wire [4-1:0] node31463;
	wire [4-1:0] node31466;
	wire [4-1:0] node31467;
	wire [4-1:0] node31471;
	wire [4-1:0] node31472;
	wire [4-1:0] node31473;
	wire [4-1:0] node31474;
	wire [4-1:0] node31478;
	wire [4-1:0] node31481;
	wire [4-1:0] node31483;
	wire [4-1:0] node31486;
	wire [4-1:0] node31487;
	wire [4-1:0] node31488;
	wire [4-1:0] node31489;
	wire [4-1:0] node31490;
	wire [4-1:0] node31491;
	wire [4-1:0] node31492;
	wire [4-1:0] node31495;
	wire [4-1:0] node31498;
	wire [4-1:0] node31499;
	wire [4-1:0] node31500;
	wire [4-1:0] node31503;
	wire [4-1:0] node31507;
	wire [4-1:0] node31508;
	wire [4-1:0] node31511;
	wire [4-1:0] node31514;
	wire [4-1:0] node31515;
	wire [4-1:0] node31516;
	wire [4-1:0] node31517;
	wire [4-1:0] node31519;
	wire [4-1:0] node31522;
	wire [4-1:0] node31524;
	wire [4-1:0] node31527;
	wire [4-1:0] node31530;
	wire [4-1:0] node31531;
	wire [4-1:0] node31534;
	wire [4-1:0] node31535;
	wire [4-1:0] node31539;
	wire [4-1:0] node31540;
	wire [4-1:0] node31541;
	wire [4-1:0] node31543;
	wire [4-1:0] node31544;
	wire [4-1:0] node31546;
	wire [4-1:0] node31549;
	wire [4-1:0] node31550;
	wire [4-1:0] node31553;
	wire [4-1:0] node31556;
	wire [4-1:0] node31557;
	wire [4-1:0] node31558;
	wire [4-1:0] node31561;
	wire [4-1:0] node31564;
	wire [4-1:0] node31565;
	wire [4-1:0] node31566;
	wire [4-1:0] node31569;
	wire [4-1:0] node31572;
	wire [4-1:0] node31574;
	wire [4-1:0] node31577;
	wire [4-1:0] node31578;
	wire [4-1:0] node31579;
	wire [4-1:0] node31580;
	wire [4-1:0] node31585;
	wire [4-1:0] node31586;
	wire [4-1:0] node31587;
	wire [4-1:0] node31591;
	wire [4-1:0] node31593;
	wire [4-1:0] node31596;
	wire [4-1:0] node31597;
	wire [4-1:0] node31598;
	wire [4-1:0] node31599;
	wire [4-1:0] node31600;
	wire [4-1:0] node31601;
	wire [4-1:0] node31602;
	wire [4-1:0] node31606;
	wire [4-1:0] node31609;
	wire [4-1:0] node31610;
	wire [4-1:0] node31614;
	wire [4-1:0] node31615;
	wire [4-1:0] node31616;
	wire [4-1:0] node31617;
	wire [4-1:0] node31620;
	wire [4-1:0] node31624;
	wire [4-1:0] node31625;
	wire [4-1:0] node31627;
	wire [4-1:0] node31630;
	wire [4-1:0] node31632;
	wire [4-1:0] node31635;
	wire [4-1:0] node31636;
	wire [4-1:0] node31637;
	wire [4-1:0] node31639;
	wire [4-1:0] node31642;
	wire [4-1:0] node31643;
	wire [4-1:0] node31644;
	wire [4-1:0] node31648;
	wire [4-1:0] node31650;
	wire [4-1:0] node31653;
	wire [4-1:0] node31654;
	wire [4-1:0] node31656;
	wire [4-1:0] node31657;
	wire [4-1:0] node31660;
	wire [4-1:0] node31663;
	wire [4-1:0] node31664;
	wire [4-1:0] node31667;
	wire [4-1:0] node31668;
	wire [4-1:0] node31672;
	wire [4-1:0] node31673;
	wire [4-1:0] node31674;
	wire [4-1:0] node31675;
	wire [4-1:0] node31676;
	wire [4-1:0] node31679;
	wire [4-1:0] node31680;
	wire [4-1:0] node31684;
	wire [4-1:0] node31685;
	wire [4-1:0] node31688;
	wire [4-1:0] node31691;
	wire [4-1:0] node31692;
	wire [4-1:0] node31693;
	wire [4-1:0] node31695;
	wire [4-1:0] node31698;
	wire [4-1:0] node31701;
	wire [4-1:0] node31702;
	wire [4-1:0] node31704;
	wire [4-1:0] node31707;
	wire [4-1:0] node31710;
	wire [4-1:0] node31711;
	wire [4-1:0] node31712;
	wire [4-1:0] node31713;
	wire [4-1:0] node31717;
	wire [4-1:0] node31718;
	wire [4-1:0] node31722;
	wire [4-1:0] node31723;
	wire [4-1:0] node31724;
	wire [4-1:0] node31728;
	wire [4-1:0] node31731;
	wire [4-1:0] node31732;
	wire [4-1:0] node31733;
	wire [4-1:0] node31734;
	wire [4-1:0] node31735;
	wire [4-1:0] node31736;
	wire [4-1:0] node31737;
	wire [4-1:0] node31738;
	wire [4-1:0] node31740;
	wire [4-1:0] node31741;
	wire [4-1:0] node31745;
	wire [4-1:0] node31746;
	wire [4-1:0] node31747;
	wire [4-1:0] node31751;
	wire [4-1:0] node31752;
	wire [4-1:0] node31756;
	wire [4-1:0] node31757;
	wire [4-1:0] node31758;
	wire [4-1:0] node31760;
	wire [4-1:0] node31763;
	wire [4-1:0] node31764;
	wire [4-1:0] node31769;
	wire [4-1:0] node31770;
	wire [4-1:0] node31771;
	wire [4-1:0] node31774;
	wire [4-1:0] node31777;
	wire [4-1:0] node31778;
	wire [4-1:0] node31780;
	wire [4-1:0] node31781;
	wire [4-1:0] node31784;
	wire [4-1:0] node31787;
	wire [4-1:0] node31789;
	wire [4-1:0] node31790;
	wire [4-1:0] node31793;
	wire [4-1:0] node31796;
	wire [4-1:0] node31797;
	wire [4-1:0] node31798;
	wire [4-1:0] node31799;
	wire [4-1:0] node31800;
	wire [4-1:0] node31802;
	wire [4-1:0] node31805;
	wire [4-1:0] node31806;
	wire [4-1:0] node31809;
	wire [4-1:0] node31812;
	wire [4-1:0] node31813;
	wire [4-1:0] node31814;
	wire [4-1:0] node31817;
	wire [4-1:0] node31821;
	wire [4-1:0] node31822;
	wire [4-1:0] node31823;
	wire [4-1:0] node31826;
	wire [4-1:0] node31829;
	wire [4-1:0] node31830;
	wire [4-1:0] node31833;
	wire [4-1:0] node31836;
	wire [4-1:0] node31837;
	wire [4-1:0] node31838;
	wire [4-1:0] node31841;
	wire [4-1:0] node31842;
	wire [4-1:0] node31846;
	wire [4-1:0] node31847;
	wire [4-1:0] node31848;
	wire [4-1:0] node31852;
	wire [4-1:0] node31853;
	wire [4-1:0] node31857;
	wire [4-1:0] node31858;
	wire [4-1:0] node31859;
	wire [4-1:0] node31860;
	wire [4-1:0] node31861;
	wire [4-1:0] node31862;
	wire [4-1:0] node31866;
	wire [4-1:0] node31868;
	wire [4-1:0] node31871;
	wire [4-1:0] node31872;
	wire [4-1:0] node31874;
	wire [4-1:0] node31877;
	wire [4-1:0] node31880;
	wire [4-1:0] node31881;
	wire [4-1:0] node31882;
	wire [4-1:0] node31886;
	wire [4-1:0] node31887;
	wire [4-1:0] node31888;
	wire [4-1:0] node31892;
	wire [4-1:0] node31893;
	wire [4-1:0] node31897;
	wire [4-1:0] node31898;
	wire [4-1:0] node31899;
	wire [4-1:0] node31900;
	wire [4-1:0] node31901;
	wire [4-1:0] node31905;
	wire [4-1:0] node31906;
	wire [4-1:0] node31910;
	wire [4-1:0] node31911;
	wire [4-1:0] node31912;
	wire [4-1:0] node31916;
	wire [4-1:0] node31919;
	wire [4-1:0] node31920;
	wire [4-1:0] node31921;
	wire [4-1:0] node31922;
	wire [4-1:0] node31926;
	wire [4-1:0] node31927;
	wire [4-1:0] node31931;
	wire [4-1:0] node31932;
	wire [4-1:0] node31933;
	wire [4-1:0] node31937;
	wire [4-1:0] node31938;
	wire [4-1:0] node31942;
	wire [4-1:0] node31943;
	wire [4-1:0] node31944;
	wire [4-1:0] node31945;
	wire [4-1:0] node31946;
	wire [4-1:0] node31947;
	wire [4-1:0] node31950;
	wire [4-1:0] node31953;
	wire [4-1:0] node31954;
	wire [4-1:0] node31956;
	wire [4-1:0] node31959;
	wire [4-1:0] node31962;
	wire [4-1:0] node31963;
	wire [4-1:0] node31964;
	wire [4-1:0] node31965;
	wire [4-1:0] node31969;
	wire [4-1:0] node31970;
	wire [4-1:0] node31973;
	wire [4-1:0] node31976;
	wire [4-1:0] node31977;
	wire [4-1:0] node31978;
	wire [4-1:0] node31981;
	wire [4-1:0] node31984;
	wire [4-1:0] node31986;
	wire [4-1:0] node31989;
	wire [4-1:0] node31990;
	wire [4-1:0] node31991;
	wire [4-1:0] node31992;
	wire [4-1:0] node31993;
	wire [4-1:0] node31997;
	wire [4-1:0] node31998;
	wire [4-1:0] node32002;
	wire [4-1:0] node32003;
	wire [4-1:0] node32004;
	wire [4-1:0] node32008;
	wire [4-1:0] node32010;
	wire [4-1:0] node32013;
	wire [4-1:0] node32014;
	wire [4-1:0] node32016;
	wire [4-1:0] node32017;
	wire [4-1:0] node32021;
	wire [4-1:0] node32022;
	wire [4-1:0] node32023;
	wire [4-1:0] node32027;
	wire [4-1:0] node32029;
	wire [4-1:0] node32032;
	wire [4-1:0] node32033;
	wire [4-1:0] node32034;
	wire [4-1:0] node32035;
	wire [4-1:0] node32036;
	wire [4-1:0] node32037;
	wire [4-1:0] node32040;
	wire [4-1:0] node32043;
	wire [4-1:0] node32045;
	wire [4-1:0] node32048;
	wire [4-1:0] node32049;
	wire [4-1:0] node32050;
	wire [4-1:0] node32054;
	wire [4-1:0] node32055;
	wire [4-1:0] node32058;
	wire [4-1:0] node32061;
	wire [4-1:0] node32062;
	wire [4-1:0] node32063;
	wire [4-1:0] node32064;
	wire [4-1:0] node32066;
	wire [4-1:0] node32069;
	wire [4-1:0] node32070;
	wire [4-1:0] node32074;
	wire [4-1:0] node32075;
	wire [4-1:0] node32077;
	wire [4-1:0] node32081;
	wire [4-1:0] node32082;
	wire [4-1:0] node32083;
	wire [4-1:0] node32087;
	wire [4-1:0] node32089;
	wire [4-1:0] node32090;
	wire [4-1:0] node32093;
	wire [4-1:0] node32096;
	wire [4-1:0] node32097;
	wire [4-1:0] node32098;
	wire [4-1:0] node32099;
	wire [4-1:0] node32100;
	wire [4-1:0] node32102;
	wire [4-1:0] node32105;
	wire [4-1:0] node32108;
	wire [4-1:0] node32109;
	wire [4-1:0] node32112;
	wire [4-1:0] node32115;
	wire [4-1:0] node32116;
	wire [4-1:0] node32117;
	wire [4-1:0] node32119;
	wire [4-1:0] node32122;
	wire [4-1:0] node32125;
	wire [4-1:0] node32126;
	wire [4-1:0] node32128;
	wire [4-1:0] node32131;
	wire [4-1:0] node32134;
	wire [4-1:0] node32135;
	wire [4-1:0] node32136;
	wire [4-1:0] node32137;
	wire [4-1:0] node32140;
	wire [4-1:0] node32143;
	wire [4-1:0] node32144;
	wire [4-1:0] node32147;
	wire [4-1:0] node32150;
	wire [4-1:0] node32151;
	wire [4-1:0] node32152;
	wire [4-1:0] node32153;
	wire [4-1:0] node32156;
	wire [4-1:0] node32159;
	wire [4-1:0] node32160;
	wire [4-1:0] node32164;
	wire [4-1:0] node32167;
	wire [4-1:0] node32168;
	wire [4-1:0] node32169;
	wire [4-1:0] node32170;
	wire [4-1:0] node32171;
	wire [4-1:0] node32172;
	wire [4-1:0] node32173;
	wire [4-1:0] node32174;
	wire [4-1:0] node32178;
	wire [4-1:0] node32179;
	wire [4-1:0] node32183;
	wire [4-1:0] node32184;
	wire [4-1:0] node32186;
	wire [4-1:0] node32189;
	wire [4-1:0] node32191;
	wire [4-1:0] node32194;
	wire [4-1:0] node32195;
	wire [4-1:0] node32196;
	wire [4-1:0] node32199;
	wire [4-1:0] node32200;
	wire [4-1:0] node32204;
	wire [4-1:0] node32205;
	wire [4-1:0] node32207;
	wire [4-1:0] node32210;
	wire [4-1:0] node32211;
	wire [4-1:0] node32215;
	wire [4-1:0] node32216;
	wire [4-1:0] node32217;
	wire [4-1:0] node32218;
	wire [4-1:0] node32219;
	wire [4-1:0] node32222;
	wire [4-1:0] node32225;
	wire [4-1:0] node32226;
	wire [4-1:0] node32227;
	wire [4-1:0] node32230;
	wire [4-1:0] node32233;
	wire [4-1:0] node32234;
	wire [4-1:0] node32237;
	wire [4-1:0] node32240;
	wire [4-1:0] node32241;
	wire [4-1:0] node32244;
	wire [4-1:0] node32247;
	wire [4-1:0] node32248;
	wire [4-1:0] node32249;
	wire [4-1:0] node32252;
	wire [4-1:0] node32255;
	wire [4-1:0] node32256;
	wire [4-1:0] node32257;
	wire [4-1:0] node32260;
	wire [4-1:0] node32264;
	wire [4-1:0] node32265;
	wire [4-1:0] node32266;
	wire [4-1:0] node32267;
	wire [4-1:0] node32268;
	wire [4-1:0] node32269;
	wire [4-1:0] node32270;
	wire [4-1:0] node32273;
	wire [4-1:0] node32276;
	wire [4-1:0] node32277;
	wire [4-1:0] node32281;
	wire [4-1:0] node32283;
	wire [4-1:0] node32284;
	wire [4-1:0] node32288;
	wire [4-1:0] node32289;
	wire [4-1:0] node32290;
	wire [4-1:0] node32294;
	wire [4-1:0] node32295;
	wire [4-1:0] node32296;
	wire [4-1:0] node32299;
	wire [4-1:0] node32302;
	wire [4-1:0] node32304;
	wire [4-1:0] node32307;
	wire [4-1:0] node32308;
	wire [4-1:0] node32309;
	wire [4-1:0] node32313;
	wire [4-1:0] node32314;
	wire [4-1:0] node32315;
	wire [4-1:0] node32318;
	wire [4-1:0] node32321;
	wire [4-1:0] node32322;
	wire [4-1:0] node32325;
	wire [4-1:0] node32328;
	wire [4-1:0] node32329;
	wire [4-1:0] node32330;
	wire [4-1:0] node32331;
	wire [4-1:0] node32332;
	wire [4-1:0] node32334;
	wire [4-1:0] node32338;
	wire [4-1:0] node32339;
	wire [4-1:0] node32340;
	wire [4-1:0] node32343;
	wire [4-1:0] node32347;
	wire [4-1:0] node32348;
	wire [4-1:0] node32349;
	wire [4-1:0] node32353;
	wire [4-1:0] node32354;
	wire [4-1:0] node32355;
	wire [4-1:0] node32360;
	wire [4-1:0] node32361;
	wire [4-1:0] node32362;
	wire [4-1:0] node32363;
	wire [4-1:0] node32364;
	wire [4-1:0] node32369;
	wire [4-1:0] node32370;
	wire [4-1:0] node32372;
	wire [4-1:0] node32376;
	wire [4-1:0] node32377;
	wire [4-1:0] node32378;
	wire [4-1:0] node32379;
	wire [4-1:0] node32384;
	wire [4-1:0] node32385;
	wire [4-1:0] node32386;
	wire [4-1:0] node32389;
	wire [4-1:0] node32393;
	wire [4-1:0] node32394;
	wire [4-1:0] node32395;
	wire [4-1:0] node32396;
	wire [4-1:0] node32397;
	wire [4-1:0] node32398;
	wire [4-1:0] node32399;
	wire [4-1:0] node32400;
	wire [4-1:0] node32403;
	wire [4-1:0] node32406;
	wire [4-1:0] node32407;
	wire [4-1:0] node32410;
	wire [4-1:0] node32413;
	wire [4-1:0] node32414;
	wire [4-1:0] node32417;
	wire [4-1:0] node32419;
	wire [4-1:0] node32422;
	wire [4-1:0] node32423;
	wire [4-1:0] node32424;
	wire [4-1:0] node32427;
	wire [4-1:0] node32430;
	wire [4-1:0] node32431;
	wire [4-1:0] node32434;
	wire [4-1:0] node32437;
	wire [4-1:0] node32438;
	wire [4-1:0] node32439;
	wire [4-1:0] node32440;
	wire [4-1:0] node32443;
	wire [4-1:0] node32446;
	wire [4-1:0] node32448;
	wire [4-1:0] node32451;
	wire [4-1:0] node32452;
	wire [4-1:0] node32455;
	wire [4-1:0] node32458;
	wire [4-1:0] node32459;
	wire [4-1:0] node32460;
	wire [4-1:0] node32463;
	wire [4-1:0] node32466;
	wire [4-1:0] node32467;
	wire [4-1:0] node32468;
	wire [4-1:0] node32469;
	wire [4-1:0] node32472;
	wire [4-1:0] node32476;
	wire [4-1:0] node32477;
	wire [4-1:0] node32478;
	wire [4-1:0] node32481;
	wire [4-1:0] node32484;
	wire [4-1:0] node32485;
	wire [4-1:0] node32488;
	wire [4-1:0] node32491;
	wire [4-1:0] node32492;
	wire [4-1:0] node32493;
	wire [4-1:0] node32494;
	wire [4-1:0] node32496;
	wire [4-1:0] node32499;
	wire [4-1:0] node32501;
	wire [4-1:0] node32504;
	wire [4-1:0] node32505;
	wire [4-1:0] node32507;
	wire [4-1:0] node32510;
	wire [4-1:0] node32512;
	wire [4-1:0] node32515;
	wire [4-1:0] node32516;
	wire [4-1:0] node32517;
	wire [4-1:0] node32518;
	wire [4-1:0] node32522;
	wire [4-1:0] node32523;
	wire [4-1:0] node32527;
	wire [4-1:0] node32528;
	wire [4-1:0] node32529;
	wire [4-1:0] node32533;
	wire [4-1:0] node32534;
	wire [4-1:0] node32538;
	wire [4-1:0] node32539;
	wire [4-1:0] node32540;
	wire [4-1:0] node32541;
	wire [4-1:0] node32542;
	wire [4-1:0] node32543;
	wire [4-1:0] node32544;
	wire [4-1:0] node32545;
	wire [4-1:0] node32546;
	wire [4-1:0] node32547;
	wire [4-1:0] node32551;
	wire [4-1:0] node32552;
	wire [4-1:0] node32554;
	wire [4-1:0] node32558;
	wire [4-1:0] node32559;
	wire [4-1:0] node32560;
	wire [4-1:0] node32561;
	wire [4-1:0] node32565;
	wire [4-1:0] node32566;
	wire [4-1:0] node32570;
	wire [4-1:0] node32571;
	wire [4-1:0] node32574;
	wire [4-1:0] node32576;
	wire [4-1:0] node32579;
	wire [4-1:0] node32580;
	wire [4-1:0] node32581;
	wire [4-1:0] node32582;
	wire [4-1:0] node32583;
	wire [4-1:0] node32587;
	wire [4-1:0] node32590;
	wire [4-1:0] node32591;
	wire [4-1:0] node32592;
	wire [4-1:0] node32596;
	wire [4-1:0] node32597;
	wire [4-1:0] node32601;
	wire [4-1:0] node32602;
	wire [4-1:0] node32603;
	wire [4-1:0] node32607;
	wire [4-1:0] node32608;
	wire [4-1:0] node32609;
	wire [4-1:0] node32613;
	wire [4-1:0] node32615;
	wire [4-1:0] node32618;
	wire [4-1:0] node32619;
	wire [4-1:0] node32620;
	wire [4-1:0] node32621;
	wire [4-1:0] node32624;
	wire [4-1:0] node32626;
	wire [4-1:0] node32629;
	wire [4-1:0] node32630;
	wire [4-1:0] node32632;
	wire [4-1:0] node32633;
	wire [4-1:0] node32638;
	wire [4-1:0] node32639;
	wire [4-1:0] node32640;
	wire [4-1:0] node32641;
	wire [4-1:0] node32642;
	wire [4-1:0] node32645;
	wire [4-1:0] node32648;
	wire [4-1:0] node32649;
	wire [4-1:0] node32652;
	wire [4-1:0] node32655;
	wire [4-1:0] node32656;
	wire [4-1:0] node32657;
	wire [4-1:0] node32662;
	wire [4-1:0] node32663;
	wire [4-1:0] node32664;
	wire [4-1:0] node32665;
	wire [4-1:0] node32668;
	wire [4-1:0] node32673;
	wire [4-1:0] node32674;
	wire [4-1:0] node32675;
	wire [4-1:0] node32676;
	wire [4-1:0] node32677;
	wire [4-1:0] node32678;
	wire [4-1:0] node32681;
	wire [4-1:0] node32684;
	wire [4-1:0] node32686;
	wire [4-1:0] node32687;
	wire [4-1:0] node32690;
	wire [4-1:0] node32693;
	wire [4-1:0] node32694;
	wire [4-1:0] node32695;
	wire [4-1:0] node32698;
	wire [4-1:0] node32701;
	wire [4-1:0] node32702;
	wire [4-1:0] node32703;
	wire [4-1:0] node32706;
	wire [4-1:0] node32709;
	wire [4-1:0] node32711;
	wire [4-1:0] node32714;
	wire [4-1:0] node32715;
	wire [4-1:0] node32716;
	wire [4-1:0] node32717;
	wire [4-1:0] node32720;
	wire [4-1:0] node32721;
	wire [4-1:0] node32725;
	wire [4-1:0] node32726;
	wire [4-1:0] node32730;
	wire [4-1:0] node32731;
	wire [4-1:0] node32733;
	wire [4-1:0] node32734;
	wire [4-1:0] node32737;
	wire [4-1:0] node32740;
	wire [4-1:0] node32742;
	wire [4-1:0] node32745;
	wire [4-1:0] node32746;
	wire [4-1:0] node32747;
	wire [4-1:0] node32748;
	wire [4-1:0] node32749;
	wire [4-1:0] node32752;
	wire [4-1:0] node32755;
	wire [4-1:0] node32757;
	wire [4-1:0] node32758;
	wire [4-1:0] node32762;
	wire [4-1:0] node32763;
	wire [4-1:0] node32764;
	wire [4-1:0] node32765;
	wire [4-1:0] node32768;
	wire [4-1:0] node32771;
	wire [4-1:0] node32772;
	wire [4-1:0] node32775;
	wire [4-1:0] node32778;
	wire [4-1:0] node32779;
	wire [4-1:0] node32781;
	wire [4-1:0] node32785;
	wire [4-1:0] node32786;
	wire [4-1:0] node32787;
	wire [4-1:0] node32789;
	wire [4-1:0] node32791;
	wire [4-1:0] node32794;
	wire [4-1:0] node32795;
	wire [4-1:0] node32799;
	wire [4-1:0] node32800;
	wire [4-1:0] node32801;
	wire [4-1:0] node32804;
	wire [4-1:0] node32807;
	wire [4-1:0] node32809;
	wire [4-1:0] node32810;
	wire [4-1:0] node32813;
	wire [4-1:0] node32816;
	wire [4-1:0] node32817;
	wire [4-1:0] node32818;
	wire [4-1:0] node32819;
	wire [4-1:0] node32820;
	wire [4-1:0] node32821;
	wire [4-1:0] node32822;
	wire [4-1:0] node32825;
	wire [4-1:0] node32828;
	wire [4-1:0] node32829;
	wire [4-1:0] node32833;
	wire [4-1:0] node32834;
	wire [4-1:0] node32837;
	wire [4-1:0] node32840;
	wire [4-1:0] node32841;
	wire [4-1:0] node32842;
	wire [4-1:0] node32843;
	wire [4-1:0] node32844;
	wire [4-1:0] node32848;
	wire [4-1:0] node32851;
	wire [4-1:0] node32852;
	wire [4-1:0] node32853;
	wire [4-1:0] node32857;
	wire [4-1:0] node32859;
	wire [4-1:0] node32862;
	wire [4-1:0] node32863;
	wire [4-1:0] node32864;
	wire [4-1:0] node32865;
	wire [4-1:0] node32868;
	wire [4-1:0] node32871;
	wire [4-1:0] node32872;
	wire [4-1:0] node32875;
	wire [4-1:0] node32878;
	wire [4-1:0] node32879;
	wire [4-1:0] node32882;
	wire [4-1:0] node32884;
	wire [4-1:0] node32887;
	wire [4-1:0] node32888;
	wire [4-1:0] node32889;
	wire [4-1:0] node32890;
	wire [4-1:0] node32891;
	wire [4-1:0] node32895;
	wire [4-1:0] node32897;
	wire [4-1:0] node32898;
	wire [4-1:0] node32901;
	wire [4-1:0] node32904;
	wire [4-1:0] node32905;
	wire [4-1:0] node32906;
	wire [4-1:0] node32907;
	wire [4-1:0] node32912;
	wire [4-1:0] node32913;
	wire [4-1:0] node32915;
	wire [4-1:0] node32918;
	wire [4-1:0] node32919;
	wire [4-1:0] node32923;
	wire [4-1:0] node32924;
	wire [4-1:0] node32925;
	wire [4-1:0] node32926;
	wire [4-1:0] node32929;
	wire [4-1:0] node32933;
	wire [4-1:0] node32934;
	wire [4-1:0] node32935;
	wire [4-1:0] node32938;
	wire [4-1:0] node32941;
	wire [4-1:0] node32942;
	wire [4-1:0] node32944;
	wire [4-1:0] node32947;
	wire [4-1:0] node32949;
	wire [4-1:0] node32952;
	wire [4-1:0] node32953;
	wire [4-1:0] node32954;
	wire [4-1:0] node32955;
	wire [4-1:0] node32956;
	wire [4-1:0] node32958;
	wire [4-1:0] node32962;
	wire [4-1:0] node32963;
	wire [4-1:0] node32964;
	wire [4-1:0] node32967;
	wire [4-1:0] node32969;
	wire [4-1:0] node32972;
	wire [4-1:0] node32973;
	wire [4-1:0] node32974;
	wire [4-1:0] node32979;
	wire [4-1:0] node32980;
	wire [4-1:0] node32981;
	wire [4-1:0] node32982;
	wire [4-1:0] node32983;
	wire [4-1:0] node32988;
	wire [4-1:0] node32989;
	wire [4-1:0] node32993;
	wire [4-1:0] node32994;
	wire [4-1:0] node32995;
	wire [4-1:0] node32998;
	wire [4-1:0] node33001;
	wire [4-1:0] node33002;
	wire [4-1:0] node33006;
	wire [4-1:0] node33007;
	wire [4-1:0] node33008;
	wire [4-1:0] node33009;
	wire [4-1:0] node33011;
	wire [4-1:0] node33012;
	wire [4-1:0] node33015;
	wire [4-1:0] node33018;
	wire [4-1:0] node33019;
	wire [4-1:0] node33020;
	wire [4-1:0] node33024;
	wire [4-1:0] node33027;
	wire [4-1:0] node33028;
	wire [4-1:0] node33029;
	wire [4-1:0] node33031;
	wire [4-1:0] node33034;
	wire [4-1:0] node33035;
	wire [4-1:0] node33038;
	wire [4-1:0] node33041;
	wire [4-1:0] node33042;
	wire [4-1:0] node33045;
	wire [4-1:0] node33048;
	wire [4-1:0] node33049;
	wire [4-1:0] node33050;
	wire [4-1:0] node33051;
	wire [4-1:0] node33052;
	wire [4-1:0] node33055;
	wire [4-1:0] node33058;
	wire [4-1:0] node33059;
	wire [4-1:0] node33062;
	wire [4-1:0] node33065;
	wire [4-1:0] node33066;
	wire [4-1:0] node33067;
	wire [4-1:0] node33070;
	wire [4-1:0] node33073;
	wire [4-1:0] node33074;
	wire [4-1:0] node33078;
	wire [4-1:0] node33079;
	wire [4-1:0] node33080;
	wire [4-1:0] node33084;
	wire [4-1:0] node33085;
	wire [4-1:0] node33086;
	wire [4-1:0] node33090;
	wire [4-1:0] node33091;
	wire [4-1:0] node33095;
	wire [4-1:0] node33096;
	wire [4-1:0] node33097;
	wire [4-1:0] node33098;
	wire [4-1:0] node33099;
	wire [4-1:0] node33100;
	wire [4-1:0] node33101;
	wire [4-1:0] node33103;
	wire [4-1:0] node33105;
	wire [4-1:0] node33108;
	wire [4-1:0] node33109;
	wire [4-1:0] node33112;
	wire [4-1:0] node33115;
	wire [4-1:0] node33116;
	wire [4-1:0] node33117;
	wire [4-1:0] node33121;
	wire [4-1:0] node33122;
	wire [4-1:0] node33125;
	wire [4-1:0] node33128;
	wire [4-1:0] node33129;
	wire [4-1:0] node33130;
	wire [4-1:0] node33131;
	wire [4-1:0] node33132;
	wire [4-1:0] node33136;
	wire [4-1:0] node33138;
	wire [4-1:0] node33141;
	wire [4-1:0] node33142;
	wire [4-1:0] node33143;
	wire [4-1:0] node33146;
	wire [4-1:0] node33150;
	wire [4-1:0] node33151;
	wire [4-1:0] node33152;
	wire [4-1:0] node33154;
	wire [4-1:0] node33157;
	wire [4-1:0] node33159;
	wire [4-1:0] node33162;
	wire [4-1:0] node33164;
	wire [4-1:0] node33165;
	wire [4-1:0] node33169;
	wire [4-1:0] node33170;
	wire [4-1:0] node33171;
	wire [4-1:0] node33172;
	wire [4-1:0] node33173;
	wire [4-1:0] node33175;
	wire [4-1:0] node33179;
	wire [4-1:0] node33180;
	wire [4-1:0] node33183;
	wire [4-1:0] node33186;
	wire [4-1:0] node33187;
	wire [4-1:0] node33188;
	wire [4-1:0] node33191;
	wire [4-1:0] node33194;
	wire [4-1:0] node33195;
	wire [4-1:0] node33196;
	wire [4-1:0] node33200;
	wire [4-1:0] node33201;
	wire [4-1:0] node33205;
	wire [4-1:0] node33206;
	wire [4-1:0] node33207;
	wire [4-1:0] node33208;
	wire [4-1:0] node33210;
	wire [4-1:0] node33214;
	wire [4-1:0] node33215;
	wire [4-1:0] node33216;
	wire [4-1:0] node33221;
	wire [4-1:0] node33222;
	wire [4-1:0] node33224;
	wire [4-1:0] node33226;
	wire [4-1:0] node33229;
	wire [4-1:0] node33230;
	wire [4-1:0] node33232;
	wire [4-1:0] node33235;
	wire [4-1:0] node33236;
	wire [4-1:0] node33240;
	wire [4-1:0] node33241;
	wire [4-1:0] node33242;
	wire [4-1:0] node33243;
	wire [4-1:0] node33245;
	wire [4-1:0] node33246;
	wire [4-1:0] node33250;
	wire [4-1:0] node33251;
	wire [4-1:0] node33252;
	wire [4-1:0] node33254;
	wire [4-1:0] node33257;
	wire [4-1:0] node33260;
	wire [4-1:0] node33261;
	wire [4-1:0] node33263;
	wire [4-1:0] node33266;
	wire [4-1:0] node33269;
	wire [4-1:0] node33270;
	wire [4-1:0] node33271;
	wire [4-1:0] node33272;
	wire [4-1:0] node33276;
	wire [4-1:0] node33278;
	wire [4-1:0] node33279;
	wire [4-1:0] node33282;
	wire [4-1:0] node33285;
	wire [4-1:0] node33286;
	wire [4-1:0] node33289;
	wire [4-1:0] node33290;
	wire [4-1:0] node33291;
	wire [4-1:0] node33295;
	wire [4-1:0] node33297;
	wire [4-1:0] node33300;
	wire [4-1:0] node33301;
	wire [4-1:0] node33302;
	wire [4-1:0] node33305;
	wire [4-1:0] node33308;
	wire [4-1:0] node33309;
	wire [4-1:0] node33310;
	wire [4-1:0] node33313;
	wire [4-1:0] node33316;
	wire [4-1:0] node33317;
	wire [4-1:0] node33318;
	wire [4-1:0] node33321;
	wire [4-1:0] node33324;
	wire [4-1:0] node33325;
	wire [4-1:0] node33326;
	wire [4-1:0] node33329;
	wire [4-1:0] node33332;
	wire [4-1:0] node33333;
	wire [4-1:0] node33336;
	wire [4-1:0] node33339;
	wire [4-1:0] node33340;
	wire [4-1:0] node33341;
	wire [4-1:0] node33342;
	wire [4-1:0] node33343;
	wire [4-1:0] node33344;
	wire [4-1:0] node33345;
	wire [4-1:0] node33347;
	wire [4-1:0] node33350;
	wire [4-1:0] node33351;
	wire [4-1:0] node33354;
	wire [4-1:0] node33357;
	wire [4-1:0] node33359;
	wire [4-1:0] node33362;
	wire [4-1:0] node33363;
	wire [4-1:0] node33364;
	wire [4-1:0] node33365;
	wire [4-1:0] node33368;
	wire [4-1:0] node33371;
	wire [4-1:0] node33372;
	wire [4-1:0] node33375;
	wire [4-1:0] node33378;
	wire [4-1:0] node33379;
	wire [4-1:0] node33381;
	wire [4-1:0] node33384;
	wire [4-1:0] node33386;
	wire [4-1:0] node33389;
	wire [4-1:0] node33390;
	wire [4-1:0] node33391;
	wire [4-1:0] node33392;
	wire [4-1:0] node33394;
	wire [4-1:0] node33397;
	wire [4-1:0] node33398;
	wire [4-1:0] node33402;
	wire [4-1:0] node33403;
	wire [4-1:0] node33404;
	wire [4-1:0] node33407;
	wire [4-1:0] node33410;
	wire [4-1:0] node33412;
	wire [4-1:0] node33415;
	wire [4-1:0] node33416;
	wire [4-1:0] node33417;
	wire [4-1:0] node33420;
	wire [4-1:0] node33421;
	wire [4-1:0] node33425;
	wire [4-1:0] node33426;
	wire [4-1:0] node33428;
	wire [4-1:0] node33432;
	wire [4-1:0] node33433;
	wire [4-1:0] node33434;
	wire [4-1:0] node33435;
	wire [4-1:0] node33437;
	wire [4-1:0] node33438;
	wire [4-1:0] node33442;
	wire [4-1:0] node33444;
	wire [4-1:0] node33447;
	wire [4-1:0] node33448;
	wire [4-1:0] node33449;
	wire [4-1:0] node33451;
	wire [4-1:0] node33454;
	wire [4-1:0] node33456;
	wire [4-1:0] node33459;
	wire [4-1:0] node33460;
	wire [4-1:0] node33462;
	wire [4-1:0] node33465;
	wire [4-1:0] node33467;
	wire [4-1:0] node33470;
	wire [4-1:0] node33471;
	wire [4-1:0] node33472;
	wire [4-1:0] node33473;
	wire [4-1:0] node33475;
	wire [4-1:0] node33478;
	wire [4-1:0] node33479;
	wire [4-1:0] node33482;
	wire [4-1:0] node33485;
	wire [4-1:0] node33486;
	wire [4-1:0] node33489;
	wire [4-1:0] node33492;
	wire [4-1:0] node33493;
	wire [4-1:0] node33495;
	wire [4-1:0] node33496;
	wire [4-1:0] node33499;
	wire [4-1:0] node33502;
	wire [4-1:0] node33504;
	wire [4-1:0] node33507;
	wire [4-1:0] node33508;
	wire [4-1:0] node33509;
	wire [4-1:0] node33510;
	wire [4-1:0] node33511;
	wire [4-1:0] node33512;
	wire [4-1:0] node33514;
	wire [4-1:0] node33517;
	wire [4-1:0] node33518;
	wire [4-1:0] node33522;
	wire [4-1:0] node33523;
	wire [4-1:0] node33526;
	wire [4-1:0] node33529;
	wire [4-1:0] node33530;
	wire [4-1:0] node33532;
	wire [4-1:0] node33533;
	wire [4-1:0] node33537;
	wire [4-1:0] node33538;
	wire [4-1:0] node33540;
	wire [4-1:0] node33543;
	wire [4-1:0] node33546;
	wire [4-1:0] node33547;
	wire [4-1:0] node33548;
	wire [4-1:0] node33549;
	wire [4-1:0] node33551;
	wire [4-1:0] node33554;
	wire [4-1:0] node33557;
	wire [4-1:0] node33558;
	wire [4-1:0] node33562;
	wire [4-1:0] node33563;
	wire [4-1:0] node33564;
	wire [4-1:0] node33565;
	wire [4-1:0] node33568;
	wire [4-1:0] node33572;
	wire [4-1:0] node33574;
	wire [4-1:0] node33575;
	wire [4-1:0] node33578;
	wire [4-1:0] node33581;
	wire [4-1:0] node33582;
	wire [4-1:0] node33583;
	wire [4-1:0] node33584;
	wire [4-1:0] node33585;
	wire [4-1:0] node33588;
	wire [4-1:0] node33591;
	wire [4-1:0] node33593;
	wire [4-1:0] node33596;
	wire [4-1:0] node33597;
	wire [4-1:0] node33599;
	wire [4-1:0] node33600;
	wire [4-1:0] node33603;
	wire [4-1:0] node33606;
	wire [4-1:0] node33607;
	wire [4-1:0] node33608;
	wire [4-1:0] node33612;
	wire [4-1:0] node33613;
	wire [4-1:0] node33616;
	wire [4-1:0] node33619;
	wire [4-1:0] node33620;
	wire [4-1:0] node33623;
	wire [4-1:0] node33626;
	wire [4-1:0] node33627;
	wire [4-1:0] node33628;
	wire [4-1:0] node33629;
	wire [4-1:0] node33630;
	wire [4-1:0] node33631;
	wire [4-1:0] node33632;
	wire [4-1:0] node33634;
	wire [4-1:0] node33635;
	wire [4-1:0] node33638;
	wire [4-1:0] node33641;
	wire [4-1:0] node33643;
	wire [4-1:0] node33644;
	wire [4-1:0] node33647;
	wire [4-1:0] node33650;
	wire [4-1:0] node33651;
	wire [4-1:0] node33652;
	wire [4-1:0] node33653;
	wire [4-1:0] node33658;
	wire [4-1:0] node33660;
	wire [4-1:0] node33662;
	wire [4-1:0] node33663;
	wire [4-1:0] node33666;
	wire [4-1:0] node33669;
	wire [4-1:0] node33670;
	wire [4-1:0] node33671;
	wire [4-1:0] node33672;
	wire [4-1:0] node33673;
	wire [4-1:0] node33676;
	wire [4-1:0] node33679;
	wire [4-1:0] node33680;
	wire [4-1:0] node33682;
	wire [4-1:0] node33685;
	wire [4-1:0] node33687;
	wire [4-1:0] node33690;
	wire [4-1:0] node33691;
	wire [4-1:0] node33692;
	wire [4-1:0] node33693;
	wire [4-1:0] node33698;
	wire [4-1:0] node33699;
	wire [4-1:0] node33701;
	wire [4-1:0] node33704;
	wire [4-1:0] node33706;
	wire [4-1:0] node33709;
	wire [4-1:0] node33710;
	wire [4-1:0] node33711;
	wire [4-1:0] node33712;
	wire [4-1:0] node33713;
	wire [4-1:0] node33717;
	wire [4-1:0] node33720;
	wire [4-1:0] node33722;
	wire [4-1:0] node33725;
	wire [4-1:0] node33726;
	wire [4-1:0] node33729;
	wire [4-1:0] node33732;
	wire [4-1:0] node33733;
	wire [4-1:0] node33734;
	wire [4-1:0] node33735;
	wire [4-1:0] node33736;
	wire [4-1:0] node33737;
	wire [4-1:0] node33741;
	wire [4-1:0] node33742;
	wire [4-1:0] node33746;
	wire [4-1:0] node33747;
	wire [4-1:0] node33750;
	wire [4-1:0] node33752;
	wire [4-1:0] node33755;
	wire [4-1:0] node33756;
	wire [4-1:0] node33757;
	wire [4-1:0] node33760;
	wire [4-1:0] node33763;
	wire [4-1:0] node33764;
	wire [4-1:0] node33765;
	wire [4-1:0] node33766;
	wire [4-1:0] node33769;
	wire [4-1:0] node33773;
	wire [4-1:0] node33774;
	wire [4-1:0] node33775;
	wire [4-1:0] node33779;
	wire [4-1:0] node33781;
	wire [4-1:0] node33784;
	wire [4-1:0] node33785;
	wire [4-1:0] node33786;
	wire [4-1:0] node33787;
	wire [4-1:0] node33788;
	wire [4-1:0] node33791;
	wire [4-1:0] node33794;
	wire [4-1:0] node33796;
	wire [4-1:0] node33797;
	wire [4-1:0] node33800;
	wire [4-1:0] node33803;
	wire [4-1:0] node33804;
	wire [4-1:0] node33806;
	wire [4-1:0] node33807;
	wire [4-1:0] node33810;
	wire [4-1:0] node33813;
	wire [4-1:0] node33814;
	wire [4-1:0] node33815;
	wire [4-1:0] node33818;
	wire [4-1:0] node33821;
	wire [4-1:0] node33822;
	wire [4-1:0] node33825;
	wire [4-1:0] node33828;
	wire [4-1:0] node33829;
	wire [4-1:0] node33832;
	wire [4-1:0] node33835;
	wire [4-1:0] node33836;
	wire [4-1:0] node33837;
	wire [4-1:0] node33838;
	wire [4-1:0] node33839;
	wire [4-1:0] node33840;
	wire [4-1:0] node33841;
	wire [4-1:0] node33845;
	wire [4-1:0] node33846;
	wire [4-1:0] node33850;
	wire [4-1:0] node33851;
	wire [4-1:0] node33852;
	wire [4-1:0] node33856;
	wire [4-1:0] node33858;
	wire [4-1:0] node33861;
	wire [4-1:0] node33862;
	wire [4-1:0] node33863;
	wire [4-1:0] node33864;
	wire [4-1:0] node33866;
	wire [4-1:0] node33869;
	wire [4-1:0] node33871;
	wire [4-1:0] node33874;
	wire [4-1:0] node33875;
	wire [4-1:0] node33877;
	wire [4-1:0] node33881;
	wire [4-1:0] node33882;
	wire [4-1:0] node33886;
	wire [4-1:0] node33887;
	wire [4-1:0] node33888;
	wire [4-1:0] node33889;
	wire [4-1:0] node33892;
	wire [4-1:0] node33895;
	wire [4-1:0] node33896;
	wire [4-1:0] node33898;
	wire [4-1:0] node33899;
	wire [4-1:0] node33902;
	wire [4-1:0] node33905;
	wire [4-1:0] node33906;
	wire [4-1:0] node33907;
	wire [4-1:0] node33910;
	wire [4-1:0] node33913;
	wire [4-1:0] node33915;
	wire [4-1:0] node33918;
	wire [4-1:0] node33919;
	wire [4-1:0] node33920;
	wire [4-1:0] node33922;
	wire [4-1:0] node33925;
	wire [4-1:0] node33927;
	wire [4-1:0] node33930;
	wire [4-1:0] node33932;
	wire [4-1:0] node33933;
	wire [4-1:0] node33936;
	wire [4-1:0] node33939;
	wire [4-1:0] node33940;
	wire [4-1:0] node33941;
	wire [4-1:0] node33942;
	wire [4-1:0] node33943;
	wire [4-1:0] node33944;
	wire [4-1:0] node33947;
	wire [4-1:0] node33950;
	wire [4-1:0] node33951;
	wire [4-1:0] node33955;
	wire [4-1:0] node33956;
	wire [4-1:0] node33957;
	wire [4-1:0] node33960;
	wire [4-1:0] node33963;
	wire [4-1:0] node33965;
	wire [4-1:0] node33968;
	wire [4-1:0] node33969;
	wire [4-1:0] node33970;
	wire [4-1:0] node33971;
	wire [4-1:0] node33972;
	wire [4-1:0] node33977;
	wire [4-1:0] node33979;
	wire [4-1:0] node33981;
	wire [4-1:0] node33984;
	wire [4-1:0] node33985;
	wire [4-1:0] node33986;
	wire [4-1:0] node33987;
	wire [4-1:0] node33991;
	wire [4-1:0] node33993;
	wire [4-1:0] node33996;
	wire [4-1:0] node33997;
	wire [4-1:0] node33998;
	wire [4-1:0] node34002;
	wire [4-1:0] node34005;
	wire [4-1:0] node34006;
	wire [4-1:0] node34007;
	wire [4-1:0] node34008;
	wire [4-1:0] node34009;
	wire [4-1:0] node34012;
	wire [4-1:0] node34015;
	wire [4-1:0] node34016;
	wire [4-1:0] node34017;
	wire [4-1:0] node34020;
	wire [4-1:0] node34024;
	wire [4-1:0] node34025;
	wire [4-1:0] node34026;
	wire [4-1:0] node34027;
	wire [4-1:0] node34031;
	wire [4-1:0] node34032;
	wire [4-1:0] node34035;
	wire [4-1:0] node34038;
	wire [4-1:0] node34041;
	wire [4-1:0] node34042;
	wire [4-1:0] node34043;
	wire [4-1:0] node34044;
	wire [4-1:0] node34047;
	wire [4-1:0] node34050;
	wire [4-1:0] node34052;
	wire [4-1:0] node34053;
	wire [4-1:0] node34057;
	wire [4-1:0] node34058;
	wire [4-1:0] node34059;
	wire [4-1:0] node34060;
	wire [4-1:0] node34063;
	wire [4-1:0] node34066;
	wire [4-1:0] node34067;
	wire [4-1:0] node34070;
	wire [4-1:0] node34073;
	wire [4-1:0] node34074;
	wire [4-1:0] node34077;
	wire [4-1:0] node34080;
	wire [4-1:0] node34081;
	wire [4-1:0] node34082;
	wire [4-1:0] node34083;
	wire [4-1:0] node34084;
	wire [4-1:0] node34085;
	wire [4-1:0] node34086;
	wire [4-1:0] node34087;
	wire [4-1:0] node34091;
	wire [4-1:0] node34092;
	wire [4-1:0] node34096;
	wire [4-1:0] node34097;
	wire [4-1:0] node34098;
	wire [4-1:0] node34102;
	wire [4-1:0] node34103;
	wire [4-1:0] node34107;
	wire [4-1:0] node34108;
	wire [4-1:0] node34109;
	wire [4-1:0] node34111;
	wire [4-1:0] node34114;
	wire [4-1:0] node34116;
	wire [4-1:0] node34119;
	wire [4-1:0] node34120;
	wire [4-1:0] node34122;
	wire [4-1:0] node34125;
	wire [4-1:0] node34127;
	wire [4-1:0] node34130;
	wire [4-1:0] node34131;
	wire [4-1:0] node34132;
	wire [4-1:0] node34133;
	wire [4-1:0] node34134;
	wire [4-1:0] node34135;
	wire [4-1:0] node34139;
	wire [4-1:0] node34140;
	wire [4-1:0] node34144;
	wire [4-1:0] node34145;
	wire [4-1:0] node34146;
	wire [4-1:0] node34149;
	wire [4-1:0] node34153;
	wire [4-1:0] node34154;
	wire [4-1:0] node34157;
	wire [4-1:0] node34160;
	wire [4-1:0] node34161;
	wire [4-1:0] node34162;
	wire [4-1:0] node34163;
	wire [4-1:0] node34166;
	wire [4-1:0] node34167;
	wire [4-1:0] node34171;
	wire [4-1:0] node34172;
	wire [4-1:0] node34176;
	wire [4-1:0] node34178;
	wire [4-1:0] node34179;
	wire [4-1:0] node34183;
	wire [4-1:0] node34184;
	wire [4-1:0] node34185;
	wire [4-1:0] node34186;
	wire [4-1:0] node34187;
	wire [4-1:0] node34188;
	wire [4-1:0] node34189;
	wire [4-1:0] node34193;
	wire [4-1:0] node34195;
	wire [4-1:0] node34198;
	wire [4-1:0] node34200;
	wire [4-1:0] node34201;
	wire [4-1:0] node34204;
	wire [4-1:0] node34207;
	wire [4-1:0] node34208;
	wire [4-1:0] node34211;
	wire [4-1:0] node34214;
	wire [4-1:0] node34215;
	wire [4-1:0] node34216;
	wire [4-1:0] node34219;
	wire [4-1:0] node34222;
	wire [4-1:0] node34223;
	wire [4-1:0] node34225;
	wire [4-1:0] node34228;
	wire [4-1:0] node34229;
	wire [4-1:0] node34230;
	wire [4-1:0] node34234;
	wire [4-1:0] node34235;
	wire [4-1:0] node34239;
	wire [4-1:0] node34240;
	wire [4-1:0] node34241;
	wire [4-1:0] node34242;
	wire [4-1:0] node34243;
	wire [4-1:0] node34244;
	wire [4-1:0] node34247;
	wire [4-1:0] node34250;
	wire [4-1:0] node34252;
	wire [4-1:0] node34255;
	wire [4-1:0] node34256;
	wire [4-1:0] node34260;
	wire [4-1:0] node34261;
	wire [4-1:0] node34262;
	wire [4-1:0] node34263;
	wire [4-1:0] node34266;
	wire [4-1:0] node34270;
	wire [4-1:0] node34271;
	wire [4-1:0] node34274;
	wire [4-1:0] node34275;
	wire [4-1:0] node34279;
	wire [4-1:0] node34280;
	wire [4-1:0] node34281;
	wire [4-1:0] node34282;
	wire [4-1:0] node34283;
	wire [4-1:0] node34286;
	wire [4-1:0] node34290;
	wire [4-1:0] node34291;
	wire [4-1:0] node34292;
	wire [4-1:0] node34295;
	wire [4-1:0] node34298;
	wire [4-1:0] node34299;
	wire [4-1:0] node34302;
	wire [4-1:0] node34305;
	wire [4-1:0] node34306;
	wire [4-1:0] node34307;
	wire [4-1:0] node34310;
	wire [4-1:0] node34313;
	wire [4-1:0] node34315;
	wire [4-1:0] node34316;
	wire [4-1:0] node34319;
	wire [4-1:0] node34322;
	wire [4-1:0] node34323;
	wire [4-1:0] node34324;
	wire [4-1:0] node34325;
	wire [4-1:0] node34326;
	wire [4-1:0] node34327;
	wire [4-1:0] node34329;
	wire [4-1:0] node34332;
	wire [4-1:0] node34333;
	wire [4-1:0] node34336;
	wire [4-1:0] node34339;
	wire [4-1:0] node34340;
	wire [4-1:0] node34343;
	wire [4-1:0] node34346;
	wire [4-1:0] node34347;
	wire [4-1:0] node34348;
	wire [4-1:0] node34351;
	wire [4-1:0] node34354;
	wire [4-1:0] node34355;
	wire [4-1:0] node34358;
	wire [4-1:0] node34361;
	wire [4-1:0] node34362;
	wire [4-1:0] node34363;
	wire [4-1:0] node34364;
	wire [4-1:0] node34365;
	wire [4-1:0] node34366;
	wire [4-1:0] node34369;
	wire [4-1:0] node34373;
	wire [4-1:0] node34374;
	wire [4-1:0] node34375;
	wire [4-1:0] node34378;
	wire [4-1:0] node34381;
	wire [4-1:0] node34383;
	wire [4-1:0] node34386;
	wire [4-1:0] node34387;
	wire [4-1:0] node34388;
	wire [4-1:0] node34392;
	wire [4-1:0] node34393;
	wire [4-1:0] node34396;
	wire [4-1:0] node34399;
	wire [4-1:0] node34400;
	wire [4-1:0] node34403;
	wire [4-1:0] node34406;
	wire [4-1:0] node34407;
	wire [4-1:0] node34408;
	wire [4-1:0] node34409;
	wire [4-1:0] node34410;
	wire [4-1:0] node34412;
	wire [4-1:0] node34413;
	wire [4-1:0] node34416;
	wire [4-1:0] node34419;
	wire [4-1:0] node34420;
	wire [4-1:0] node34423;
	wire [4-1:0] node34426;
	wire [4-1:0] node34427;
	wire [4-1:0] node34428;
	wire [4-1:0] node34430;
	wire [4-1:0] node34433;
	wire [4-1:0] node34435;
	wire [4-1:0] node34438;
	wire [4-1:0] node34439;
	wire [4-1:0] node34440;
	wire [4-1:0] node34443;
	wire [4-1:0] node34446;
	wire [4-1:0] node34447;
	wire [4-1:0] node34450;
	wire [4-1:0] node34453;
	wire [4-1:0] node34454;
	wire [4-1:0] node34455;
	wire [4-1:0] node34456;
	wire [4-1:0] node34457;
	wire [4-1:0] node34460;
	wire [4-1:0] node34463;
	wire [4-1:0] node34464;
	wire [4-1:0] node34467;
	wire [4-1:0] node34470;
	wire [4-1:0] node34471;
	wire [4-1:0] node34473;
	wire [4-1:0] node34476;
	wire [4-1:0] node34479;
	wire [4-1:0] node34480;
	wire [4-1:0] node34481;
	wire [4-1:0] node34482;
	wire [4-1:0] node34485;
	wire [4-1:0] node34488;
	wire [4-1:0] node34490;
	wire [4-1:0] node34494;
	wire [4-1:0] node34495;
	wire [4-1:0] node34496;
	wire [4-1:0] node34499;
	wire [4-1:0] node34502;
	wire [4-1:0] node34503;
	wire [4-1:0] node34506;
	wire [4-1:0] node34509;
	wire [4-1:0] node34510;
	wire [4-1:0] node34511;
	wire [4-1:0] node34512;
	wire [4-1:0] node34513;
	wire [4-1:0] node34514;
	wire [4-1:0] node34515;
	wire [4-1:0] node34516;
	wire [4-1:0] node34517;
	wire [4-1:0] node34518;
	wire [4-1:0] node34519;
	wire [4-1:0] node34520;
	wire [4-1:0] node34523;
	wire [4-1:0] node34524;
	wire [4-1:0] node34527;
	wire [4-1:0] node34530;
	wire [4-1:0] node34531;
	wire [4-1:0] node34532;
	wire [4-1:0] node34537;
	wire [4-1:0] node34538;
	wire [4-1:0] node34539;
	wire [4-1:0] node34542;
	wire [4-1:0] node34543;
	wire [4-1:0] node34547;
	wire [4-1:0] node34548;
	wire [4-1:0] node34551;
	wire [4-1:0] node34552;
	wire [4-1:0] node34556;
	wire [4-1:0] node34557;
	wire [4-1:0] node34558;
	wire [4-1:0] node34559;
	wire [4-1:0] node34561;
	wire [4-1:0] node34564;
	wire [4-1:0] node34567;
	wire [4-1:0] node34568;
	wire [4-1:0] node34569;
	wire [4-1:0] node34574;
	wire [4-1:0] node34575;
	wire [4-1:0] node34576;
	wire [4-1:0] node34579;
	wire [4-1:0] node34580;
	wire [4-1:0] node34584;
	wire [4-1:0] node34585;
	wire [4-1:0] node34588;
	wire [4-1:0] node34589;
	wire [4-1:0] node34593;
	wire [4-1:0] node34594;
	wire [4-1:0] node34595;
	wire [4-1:0] node34596;
	wire [4-1:0] node34597;
	wire [4-1:0] node34599;
	wire [4-1:0] node34602;
	wire [4-1:0] node34605;
	wire [4-1:0] node34606;
	wire [4-1:0] node34608;
	wire [4-1:0] node34611;
	wire [4-1:0] node34614;
	wire [4-1:0] node34615;
	wire [4-1:0] node34616;
	wire [4-1:0] node34619;
	wire [4-1:0] node34622;
	wire [4-1:0] node34623;
	wire [4-1:0] node34626;
	wire [4-1:0] node34629;
	wire [4-1:0] node34630;
	wire [4-1:0] node34631;
	wire [4-1:0] node34632;
	wire [4-1:0] node34635;
	wire [4-1:0] node34637;
	wire [4-1:0] node34640;
	wire [4-1:0] node34641;
	wire [4-1:0] node34642;
	wire [4-1:0] node34645;
	wire [4-1:0] node34648;
	wire [4-1:0] node34651;
	wire [4-1:0] node34652;
	wire [4-1:0] node34653;
	wire [4-1:0] node34656;
	wire [4-1:0] node34657;
	wire [4-1:0] node34661;
	wire [4-1:0] node34662;
	wire [4-1:0] node34663;
	wire [4-1:0] node34666;
	wire [4-1:0] node34669;
	wire [4-1:0] node34672;
	wire [4-1:0] node34673;
	wire [4-1:0] node34674;
	wire [4-1:0] node34675;
	wire [4-1:0] node34676;
	wire [4-1:0] node34677;
	wire [4-1:0] node34678;
	wire [4-1:0] node34683;
	wire [4-1:0] node34684;
	wire [4-1:0] node34685;
	wire [4-1:0] node34689;
	wire [4-1:0] node34692;
	wire [4-1:0] node34693;
	wire [4-1:0] node34694;
	wire [4-1:0] node34697;
	wire [4-1:0] node34700;
	wire [4-1:0] node34701;
	wire [4-1:0] node34704;
	wire [4-1:0] node34705;
	wire [4-1:0] node34708;
	wire [4-1:0] node34711;
	wire [4-1:0] node34712;
	wire [4-1:0] node34713;
	wire [4-1:0] node34714;
	wire [4-1:0] node34715;
	wire [4-1:0] node34718;
	wire [4-1:0] node34721;
	wire [4-1:0] node34723;
	wire [4-1:0] node34726;
	wire [4-1:0] node34728;
	wire [4-1:0] node34729;
	wire [4-1:0] node34733;
	wire [4-1:0] node34734;
	wire [4-1:0] node34735;
	wire [4-1:0] node34736;
	wire [4-1:0] node34740;
	wire [4-1:0] node34743;
	wire [4-1:0] node34744;
	wire [4-1:0] node34745;
	wire [4-1:0] node34749;
	wire [4-1:0] node34751;
	wire [4-1:0] node34754;
	wire [4-1:0] node34755;
	wire [4-1:0] node34756;
	wire [4-1:0] node34757;
	wire [4-1:0] node34760;
	wire [4-1:0] node34761;
	wire [4-1:0] node34763;
	wire [4-1:0] node34767;
	wire [4-1:0] node34768;
	wire [4-1:0] node34770;
	wire [4-1:0] node34772;
	wire [4-1:0] node34775;
	wire [4-1:0] node34776;
	wire [4-1:0] node34778;
	wire [4-1:0] node34781;
	wire [4-1:0] node34783;
	wire [4-1:0] node34786;
	wire [4-1:0] node34787;
	wire [4-1:0] node34789;
	wire [4-1:0] node34790;
	wire [4-1:0] node34792;
	wire [4-1:0] node34795;
	wire [4-1:0] node34796;
	wire [4-1:0] node34799;
	wire [4-1:0] node34802;
	wire [4-1:0] node34803;
	wire [4-1:0] node34805;
	wire [4-1:0] node34806;
	wire [4-1:0] node34811;
	wire [4-1:0] node34812;
	wire [4-1:0] node34813;
	wire [4-1:0] node34814;
	wire [4-1:0] node34815;
	wire [4-1:0] node34817;
	wire [4-1:0] node34819;
	wire [4-1:0] node34820;
	wire [4-1:0] node34823;
	wire [4-1:0] node34826;
	wire [4-1:0] node34827;
	wire [4-1:0] node34829;
	wire [4-1:0] node34832;
	wire [4-1:0] node34833;
	wire [4-1:0] node34835;
	wire [4-1:0] node34838;
	wire [4-1:0] node34841;
	wire [4-1:0] node34842;
	wire [4-1:0] node34843;
	wire [4-1:0] node34845;
	wire [4-1:0] node34846;
	wire [4-1:0] node34850;
	wire [4-1:0] node34851;
	wire [4-1:0] node34852;
	wire [4-1:0] node34856;
	wire [4-1:0] node34858;
	wire [4-1:0] node34861;
	wire [4-1:0] node34862;
	wire [4-1:0] node34863;
	wire [4-1:0] node34868;
	wire [4-1:0] node34869;
	wire [4-1:0] node34870;
	wire [4-1:0] node34871;
	wire [4-1:0] node34872;
	wire [4-1:0] node34874;
	wire [4-1:0] node34878;
	wire [4-1:0] node34879;
	wire [4-1:0] node34881;
	wire [4-1:0] node34884;
	wire [4-1:0] node34887;
	wire [4-1:0] node34888;
	wire [4-1:0] node34889;
	wire [4-1:0] node34893;
	wire [4-1:0] node34894;
	wire [4-1:0] node34896;
	wire [4-1:0] node34899;
	wire [4-1:0] node34900;
	wire [4-1:0] node34904;
	wire [4-1:0] node34905;
	wire [4-1:0] node34906;
	wire [4-1:0] node34908;
	wire [4-1:0] node34911;
	wire [4-1:0] node34912;
	wire [4-1:0] node34914;
	wire [4-1:0] node34917;
	wire [4-1:0] node34919;
	wire [4-1:0] node34922;
	wire [4-1:0] node34923;
	wire [4-1:0] node34924;
	wire [4-1:0] node34925;
	wire [4-1:0] node34930;
	wire [4-1:0] node34931;
	wire [4-1:0] node34933;
	wire [4-1:0] node34936;
	wire [4-1:0] node34937;
	wire [4-1:0] node34940;
	wire [4-1:0] node34943;
	wire [4-1:0] node34944;
	wire [4-1:0] node34945;
	wire [4-1:0] node34946;
	wire [4-1:0] node34947;
	wire [4-1:0] node34948;
	wire [4-1:0] node34949;
	wire [4-1:0] node34952;
	wire [4-1:0] node34955;
	wire [4-1:0] node34958;
	wire [4-1:0] node34959;
	wire [4-1:0] node34962;
	wire [4-1:0] node34963;
	wire [4-1:0] node34966;
	wire [4-1:0] node34969;
	wire [4-1:0] node34970;
	wire [4-1:0] node34971;
	wire [4-1:0] node34975;
	wire [4-1:0] node34976;
	wire [4-1:0] node34978;
	wire [4-1:0] node34981;
	wire [4-1:0] node34984;
	wire [4-1:0] node34985;
	wire [4-1:0] node34987;
	wire [4-1:0] node34988;
	wire [4-1:0] node34989;
	wire [4-1:0] node34992;
	wire [4-1:0] node34995;
	wire [4-1:0] node34997;
	wire [4-1:0] node35000;
	wire [4-1:0] node35001;
	wire [4-1:0] node35002;
	wire [4-1:0] node35005;
	wire [4-1:0] node35007;
	wire [4-1:0] node35010;
	wire [4-1:0] node35011;
	wire [4-1:0] node35012;
	wire [4-1:0] node35015;
	wire [4-1:0] node35019;
	wire [4-1:0] node35020;
	wire [4-1:0] node35021;
	wire [4-1:0] node35022;
	wire [4-1:0] node35023;
	wire [4-1:0] node35024;
	wire [4-1:0] node35027;
	wire [4-1:0] node35030;
	wire [4-1:0] node35032;
	wire [4-1:0] node35035;
	wire [4-1:0] node35036;
	wire [4-1:0] node35039;
	wire [4-1:0] node35042;
	wire [4-1:0] node35043;
	wire [4-1:0] node35044;
	wire [4-1:0] node35045;
	wire [4-1:0] node35049;
	wire [4-1:0] node35050;
	wire [4-1:0] node35053;
	wire [4-1:0] node35056;
	wire [4-1:0] node35057;
	wire [4-1:0] node35060;
	wire [4-1:0] node35061;
	wire [4-1:0] node35065;
	wire [4-1:0] node35066;
	wire [4-1:0] node35068;
	wire [4-1:0] node35069;
	wire [4-1:0] node35073;
	wire [4-1:0] node35074;
	wire [4-1:0] node35076;
	wire [4-1:0] node35077;
	wire [4-1:0] node35080;
	wire [4-1:0] node35083;
	wire [4-1:0] node35084;
	wire [4-1:0] node35085;
	wire [4-1:0] node35090;
	wire [4-1:0] node35091;
	wire [4-1:0] node35092;
	wire [4-1:0] node35093;
	wire [4-1:0] node35094;
	wire [4-1:0] node35095;
	wire [4-1:0] node35096;
	wire [4-1:0] node35097;
	wire [4-1:0] node35099;
	wire [4-1:0] node35102;
	wire [4-1:0] node35104;
	wire [4-1:0] node35107;
	wire [4-1:0] node35108;
	wire [4-1:0] node35109;
	wire [4-1:0] node35113;
	wire [4-1:0] node35116;
	wire [4-1:0] node35117;
	wire [4-1:0] node35118;
	wire [4-1:0] node35119;
	wire [4-1:0] node35123;
	wire [4-1:0] node35124;
	wire [4-1:0] node35127;
	wire [4-1:0] node35130;
	wire [4-1:0] node35131;
	wire [4-1:0] node35132;
	wire [4-1:0] node35136;
	wire [4-1:0] node35139;
	wire [4-1:0] node35140;
	wire [4-1:0] node35141;
	wire [4-1:0] node35142;
	wire [4-1:0] node35146;
	wire [4-1:0] node35147;
	wire [4-1:0] node35149;
	wire [4-1:0] node35153;
	wire [4-1:0] node35154;
	wire [4-1:0] node35155;
	wire [4-1:0] node35156;
	wire [4-1:0] node35160;
	wire [4-1:0] node35161;
	wire [4-1:0] node35165;
	wire [4-1:0] node35166;
	wire [4-1:0] node35167;
	wire [4-1:0] node35170;
	wire [4-1:0] node35173;
	wire [4-1:0] node35174;
	wire [4-1:0] node35177;
	wire [4-1:0] node35180;
	wire [4-1:0] node35181;
	wire [4-1:0] node35182;
	wire [4-1:0] node35183;
	wire [4-1:0] node35184;
	wire [4-1:0] node35185;
	wire [4-1:0] node35189;
	wire [4-1:0] node35190;
	wire [4-1:0] node35193;
	wire [4-1:0] node35196;
	wire [4-1:0] node35197;
	wire [4-1:0] node35200;
	wire [4-1:0] node35201;
	wire [4-1:0] node35204;
	wire [4-1:0] node35207;
	wire [4-1:0] node35208;
	wire [4-1:0] node35209;
	wire [4-1:0] node35213;
	wire [4-1:0] node35214;
	wire [4-1:0] node35215;
	wire [4-1:0] node35219;
	wire [4-1:0] node35222;
	wire [4-1:0] node35223;
	wire [4-1:0] node35224;
	wire [4-1:0] node35225;
	wire [4-1:0] node35226;
	wire [4-1:0] node35230;
	wire [4-1:0] node35233;
	wire [4-1:0] node35235;
	wire [4-1:0] node35238;
	wire [4-1:0] node35239;
	wire [4-1:0] node35240;
	wire [4-1:0] node35243;
	wire [4-1:0] node35246;
	wire [4-1:0] node35247;
	wire [4-1:0] node35250;
	wire [4-1:0] node35253;
	wire [4-1:0] node35254;
	wire [4-1:0] node35255;
	wire [4-1:0] node35256;
	wire [4-1:0] node35257;
	wire [4-1:0] node35258;
	wire [4-1:0] node35259;
	wire [4-1:0] node35263;
	wire [4-1:0] node35265;
	wire [4-1:0] node35268;
	wire [4-1:0] node35269;
	wire [4-1:0] node35271;
	wire [4-1:0] node35275;
	wire [4-1:0] node35276;
	wire [4-1:0] node35277;
	wire [4-1:0] node35279;
	wire [4-1:0] node35282;
	wire [4-1:0] node35283;
	wire [4-1:0] node35286;
	wire [4-1:0] node35289;
	wire [4-1:0] node35290;
	wire [4-1:0] node35291;
	wire [4-1:0] node35294;
	wire [4-1:0] node35297;
	wire [4-1:0] node35298;
	wire [4-1:0] node35302;
	wire [4-1:0] node35303;
	wire [4-1:0] node35304;
	wire [4-1:0] node35305;
	wire [4-1:0] node35307;
	wire [4-1:0] node35311;
	wire [4-1:0] node35312;
	wire [4-1:0] node35315;
	wire [4-1:0] node35318;
	wire [4-1:0] node35319;
	wire [4-1:0] node35321;
	wire [4-1:0] node35324;
	wire [4-1:0] node35325;
	wire [4-1:0] node35327;
	wire [4-1:0] node35330;
	wire [4-1:0] node35332;
	wire [4-1:0] node35335;
	wire [4-1:0] node35336;
	wire [4-1:0] node35337;
	wire [4-1:0] node35338;
	wire [4-1:0] node35339;
	wire [4-1:0] node35341;
	wire [4-1:0] node35344;
	wire [4-1:0] node35345;
	wire [4-1:0] node35349;
	wire [4-1:0] node35350;
	wire [4-1:0] node35353;
	wire [4-1:0] node35354;
	wire [4-1:0] node35358;
	wire [4-1:0] node35359;
	wire [4-1:0] node35360;
	wire [4-1:0] node35362;
	wire [4-1:0] node35365;
	wire [4-1:0] node35366;
	wire [4-1:0] node35370;
	wire [4-1:0] node35371;
	wire [4-1:0] node35373;
	wire [4-1:0] node35376;
	wire [4-1:0] node35379;
	wire [4-1:0] node35380;
	wire [4-1:0] node35381;
	wire [4-1:0] node35382;
	wire [4-1:0] node35385;
	wire [4-1:0] node35388;
	wire [4-1:0] node35389;
	wire [4-1:0] node35392;
	wire [4-1:0] node35395;
	wire [4-1:0] node35396;
	wire [4-1:0] node35397;
	wire [4-1:0] node35398;
	wire [4-1:0] node35402;
	wire [4-1:0] node35404;
	wire [4-1:0] node35407;
	wire [4-1:0] node35408;
	wire [4-1:0] node35409;
	wire [4-1:0] node35413;
	wire [4-1:0] node35415;
	wire [4-1:0] node35418;
	wire [4-1:0] node35419;
	wire [4-1:0] node35420;
	wire [4-1:0] node35421;
	wire [4-1:0] node35422;
	wire [4-1:0] node35423;
	wire [4-1:0] node35426;
	wire [4-1:0] node35428;
	wire [4-1:0] node35429;
	wire [4-1:0] node35432;
	wire [4-1:0] node35435;
	wire [4-1:0] node35436;
	wire [4-1:0] node35437;
	wire [4-1:0] node35438;
	wire [4-1:0] node35441;
	wire [4-1:0] node35444;
	wire [4-1:0] node35447;
	wire [4-1:0] node35449;
	wire [4-1:0] node35452;
	wire [4-1:0] node35453;
	wire [4-1:0] node35454;
	wire [4-1:0] node35455;
	wire [4-1:0] node35457;
	wire [4-1:0] node35460;
	wire [4-1:0] node35461;
	wire [4-1:0] node35464;
	wire [4-1:0] node35467;
	wire [4-1:0] node35468;
	wire [4-1:0] node35469;
	wire [4-1:0] node35472;
	wire [4-1:0] node35475;
	wire [4-1:0] node35477;
	wire [4-1:0] node35480;
	wire [4-1:0] node35481;
	wire [4-1:0] node35482;
	wire [4-1:0] node35483;
	wire [4-1:0] node35486;
	wire [4-1:0] node35489;
	wire [4-1:0] node35491;
	wire [4-1:0] node35494;
	wire [4-1:0] node35496;
	wire [4-1:0] node35497;
	wire [4-1:0] node35500;
	wire [4-1:0] node35503;
	wire [4-1:0] node35504;
	wire [4-1:0] node35505;
	wire [4-1:0] node35506;
	wire [4-1:0] node35507;
	wire [4-1:0] node35508;
	wire [4-1:0] node35512;
	wire [4-1:0] node35513;
	wire [4-1:0] node35517;
	wire [4-1:0] node35518;
	wire [4-1:0] node35521;
	wire [4-1:0] node35522;
	wire [4-1:0] node35525;
	wire [4-1:0] node35528;
	wire [4-1:0] node35529;
	wire [4-1:0] node35530;
	wire [4-1:0] node35532;
	wire [4-1:0] node35535;
	wire [4-1:0] node35537;
	wire [4-1:0] node35540;
	wire [4-1:0] node35541;
	wire [4-1:0] node35543;
	wire [4-1:0] node35546;
	wire [4-1:0] node35549;
	wire [4-1:0] node35550;
	wire [4-1:0] node35551;
	wire [4-1:0] node35553;
	wire [4-1:0] node35556;
	wire [4-1:0] node35557;
	wire [4-1:0] node35558;
	wire [4-1:0] node35562;
	wire [4-1:0] node35565;
	wire [4-1:0] node35566;
	wire [4-1:0] node35567;
	wire [4-1:0] node35570;
	wire [4-1:0] node35573;
	wire [4-1:0] node35574;
	wire [4-1:0] node35578;
	wire [4-1:0] node35579;
	wire [4-1:0] node35580;
	wire [4-1:0] node35581;
	wire [4-1:0] node35582;
	wire [4-1:0] node35584;
	wire [4-1:0] node35585;
	wire [4-1:0] node35589;
	wire [4-1:0] node35590;
	wire [4-1:0] node35591;
	wire [4-1:0] node35595;
	wire [4-1:0] node35598;
	wire [4-1:0] node35599;
	wire [4-1:0] node35600;
	wire [4-1:0] node35604;
	wire [4-1:0] node35605;
	wire [4-1:0] node35608;
	wire [4-1:0] node35610;
	wire [4-1:0] node35613;
	wire [4-1:0] node35614;
	wire [4-1:0] node35615;
	wire [4-1:0] node35616;
	wire [4-1:0] node35619;
	wire [4-1:0] node35621;
	wire [4-1:0] node35624;
	wire [4-1:0] node35627;
	wire [4-1:0] node35628;
	wire [4-1:0] node35629;
	wire [4-1:0] node35630;
	wire [4-1:0] node35634;
	wire [4-1:0] node35637;
	wire [4-1:0] node35638;
	wire [4-1:0] node35641;
	wire [4-1:0] node35642;
	wire [4-1:0] node35646;
	wire [4-1:0] node35647;
	wire [4-1:0] node35648;
	wire [4-1:0] node35649;
	wire [4-1:0] node35651;
	wire [4-1:0] node35652;
	wire [4-1:0] node35655;
	wire [4-1:0] node35658;
	wire [4-1:0] node35659;
	wire [4-1:0] node35662;
	wire [4-1:0] node35663;
	wire [4-1:0] node35666;
	wire [4-1:0] node35669;
	wire [4-1:0] node35670;
	wire [4-1:0] node35671;
	wire [4-1:0] node35674;
	wire [4-1:0] node35676;
	wire [4-1:0] node35679;
	wire [4-1:0] node35682;
	wire [4-1:0] node35683;
	wire [4-1:0] node35684;
	wire [4-1:0] node35686;
	wire [4-1:0] node35687;
	wire [4-1:0] node35690;
	wire [4-1:0] node35693;
	wire [4-1:0] node35694;
	wire [4-1:0] node35697;
	wire [4-1:0] node35698;
	wire [4-1:0] node35702;
	wire [4-1:0] node35703;
	wire [4-1:0] node35704;
	wire [4-1:0] node35705;
	wire [4-1:0] node35708;
	wire [4-1:0] node35711;
	wire [4-1:0] node35713;
	wire [4-1:0] node35716;
	wire [4-1:0] node35717;
	wire [4-1:0] node35719;
	wire [4-1:0] node35723;
	wire [4-1:0] node35724;
	wire [4-1:0] node35725;
	wire [4-1:0] node35726;
	wire [4-1:0] node35727;
	wire [4-1:0] node35728;
	wire [4-1:0] node35729;
	wire [4-1:0] node35730;
	wire [4-1:0] node35731;
	wire [4-1:0] node35732;
	wire [4-1:0] node35735;
	wire [4-1:0] node35739;
	wire [4-1:0] node35740;
	wire [4-1:0] node35742;
	wire [4-1:0] node35745;
	wire [4-1:0] node35747;
	wire [4-1:0] node35750;
	wire [4-1:0] node35751;
	wire [4-1:0] node35752;
	wire [4-1:0] node35755;
	wire [4-1:0] node35756;
	wire [4-1:0] node35759;
	wire [4-1:0] node35762;
	wire [4-1:0] node35763;
	wire [4-1:0] node35764;
	wire [4-1:0] node35767;
	wire [4-1:0] node35770;
	wire [4-1:0] node35771;
	wire [4-1:0] node35775;
	wire [4-1:0] node35776;
	wire [4-1:0] node35777;
	wire [4-1:0] node35778;
	wire [4-1:0] node35779;
	wire [4-1:0] node35782;
	wire [4-1:0] node35786;
	wire [4-1:0] node35787;
	wire [4-1:0] node35788;
	wire [4-1:0] node35793;
	wire [4-1:0] node35794;
	wire [4-1:0] node35795;
	wire [4-1:0] node35798;
	wire [4-1:0] node35799;
	wire [4-1:0] node35802;
	wire [4-1:0] node35805;
	wire [4-1:0] node35806;
	wire [4-1:0] node35807;
	wire [4-1:0] node35811;
	wire [4-1:0] node35813;
	wire [4-1:0] node35816;
	wire [4-1:0] node35817;
	wire [4-1:0] node35818;
	wire [4-1:0] node35819;
	wire [4-1:0] node35820;
	wire [4-1:0] node35823;
	wire [4-1:0] node35824;
	wire [4-1:0] node35828;
	wire [4-1:0] node35829;
	wire [4-1:0] node35832;
	wire [4-1:0] node35835;
	wire [4-1:0] node35836;
	wire [4-1:0] node35837;
	wire [4-1:0] node35838;
	wire [4-1:0] node35841;
	wire [4-1:0] node35844;
	wire [4-1:0] node35845;
	wire [4-1:0] node35848;
	wire [4-1:0] node35851;
	wire [4-1:0] node35852;
	wire [4-1:0] node35853;
	wire [4-1:0] node35856;
	wire [4-1:0] node35860;
	wire [4-1:0] node35861;
	wire [4-1:0] node35862;
	wire [4-1:0] node35863;
	wire [4-1:0] node35865;
	wire [4-1:0] node35868;
	wire [4-1:0] node35870;
	wire [4-1:0] node35873;
	wire [4-1:0] node35875;
	wire [4-1:0] node35878;
	wire [4-1:0] node35879;
	wire [4-1:0] node35880;
	wire [4-1:0] node35883;
	wire [4-1:0] node35886;
	wire [4-1:0] node35887;
	wire [4-1:0] node35888;
	wire [4-1:0] node35891;
	wire [4-1:0] node35894;
	wire [4-1:0] node35895;
	wire [4-1:0] node35898;
	wire [4-1:0] node35901;
	wire [4-1:0] node35902;
	wire [4-1:0] node35903;
	wire [4-1:0] node35904;
	wire [4-1:0] node35905;
	wire [4-1:0] node35906;
	wire [4-1:0] node35908;
	wire [4-1:0] node35911;
	wire [4-1:0] node35913;
	wire [4-1:0] node35916;
	wire [4-1:0] node35917;
	wire [4-1:0] node35919;
	wire [4-1:0] node35922;
	wire [4-1:0] node35925;
	wire [4-1:0] node35927;
	wire [4-1:0] node35928;
	wire [4-1:0] node35931;
	wire [4-1:0] node35934;
	wire [4-1:0] node35935;
	wire [4-1:0] node35937;
	wire [4-1:0] node35939;
	wire [4-1:0] node35940;
	wire [4-1:0] node35943;
	wire [4-1:0] node35946;
	wire [4-1:0] node35947;
	wire [4-1:0] node35948;
	wire [4-1:0] node35949;
	wire [4-1:0] node35954;
	wire [4-1:0] node35955;
	wire [4-1:0] node35958;
	wire [4-1:0] node35959;
	wire [4-1:0] node35962;
	wire [4-1:0] node35965;
	wire [4-1:0] node35966;
	wire [4-1:0] node35967;
	wire [4-1:0] node35968;
	wire [4-1:0] node35969;
	wire [4-1:0] node35972;
	wire [4-1:0] node35974;
	wire [4-1:0] node35977;
	wire [4-1:0] node35978;
	wire [4-1:0] node35981;
	wire [4-1:0] node35982;
	wire [4-1:0] node35986;
	wire [4-1:0] node35987;
	wire [4-1:0] node35988;
	wire [4-1:0] node35992;
	wire [4-1:0] node35993;
	wire [4-1:0] node35997;
	wire [4-1:0] node35998;
	wire [4-1:0] node35999;
	wire [4-1:0] node36000;
	wire [4-1:0] node36003;
	wire [4-1:0] node36006;
	wire [4-1:0] node36009;
	wire [4-1:0] node36010;
	wire [4-1:0] node36011;
	wire [4-1:0] node36013;
	wire [4-1:0] node36017;
	wire [4-1:0] node36019;
	wire [4-1:0] node36020;
	wire [4-1:0] node36024;
	wire [4-1:0] node36025;
	wire [4-1:0] node36026;
	wire [4-1:0] node36027;
	wire [4-1:0] node36028;
	wire [4-1:0] node36029;
	wire [4-1:0] node36030;
	wire [4-1:0] node36034;
	wire [4-1:0] node36036;
	wire [4-1:0] node36039;
	wire [4-1:0] node36040;
	wire [4-1:0] node36041;
	wire [4-1:0] node36045;
	wire [4-1:0] node36046;
	wire [4-1:0] node36048;
	wire [4-1:0] node36051;
	wire [4-1:0] node36053;
	wire [4-1:0] node36056;
	wire [4-1:0] node36057;
	wire [4-1:0] node36058;
	wire [4-1:0] node36059;
	wire [4-1:0] node36060;
	wire [4-1:0] node36063;
	wire [4-1:0] node36067;
	wire [4-1:0] node36069;
	wire [4-1:0] node36070;
	wire [4-1:0] node36073;
	wire [4-1:0] node36076;
	wire [4-1:0] node36077;
	wire [4-1:0] node36078;
	wire [4-1:0] node36082;
	wire [4-1:0] node36083;
	wire [4-1:0] node36087;
	wire [4-1:0] node36088;
	wire [4-1:0] node36089;
	wire [4-1:0] node36090;
	wire [4-1:0] node36091;
	wire [4-1:0] node36095;
	wire [4-1:0] node36096;
	wire [4-1:0] node36100;
	wire [4-1:0] node36101;
	wire [4-1:0] node36103;
	wire [4-1:0] node36106;
	wire [4-1:0] node36107;
	wire [4-1:0] node36109;
	wire [4-1:0] node36112;
	wire [4-1:0] node36114;
	wire [4-1:0] node36117;
	wire [4-1:0] node36118;
	wire [4-1:0] node36119;
	wire [4-1:0] node36120;
	wire [4-1:0] node36123;
	wire [4-1:0] node36125;
	wire [4-1:0] node36128;
	wire [4-1:0] node36129;
	wire [4-1:0] node36132;
	wire [4-1:0] node36135;
	wire [4-1:0] node36136;
	wire [4-1:0] node36137;
	wire [4-1:0] node36140;
	wire [4-1:0] node36141;
	wire [4-1:0] node36145;
	wire [4-1:0] node36147;
	wire [4-1:0] node36150;
	wire [4-1:0] node36151;
	wire [4-1:0] node36152;
	wire [4-1:0] node36153;
	wire [4-1:0] node36154;
	wire [4-1:0] node36156;
	wire [4-1:0] node36157;
	wire [4-1:0] node36162;
	wire [4-1:0] node36163;
	wire [4-1:0] node36164;
	wire [4-1:0] node36165;
	wire [4-1:0] node36169;
	wire [4-1:0] node36170;
	wire [4-1:0] node36174;
	wire [4-1:0] node36175;
	wire [4-1:0] node36178;
	wire [4-1:0] node36180;
	wire [4-1:0] node36183;
	wire [4-1:0] node36184;
	wire [4-1:0] node36185;
	wire [4-1:0] node36186;
	wire [4-1:0] node36187;
	wire [4-1:0] node36192;
	wire [4-1:0] node36193;
	wire [4-1:0] node36196;
	wire [4-1:0] node36197;
	wire [4-1:0] node36201;
	wire [4-1:0] node36202;
	wire [4-1:0] node36203;
	wire [4-1:0] node36205;
	wire [4-1:0] node36209;
	wire [4-1:0] node36210;
	wire [4-1:0] node36212;
	wire [4-1:0] node36215;
	wire [4-1:0] node36216;
	wire [4-1:0] node36220;
	wire [4-1:0] node36221;
	wire [4-1:0] node36222;
	wire [4-1:0] node36223;
	wire [4-1:0] node36224;
	wire [4-1:0] node36225;
	wire [4-1:0] node36230;
	wire [4-1:0] node36231;
	wire [4-1:0] node36233;
	wire [4-1:0] node36236;
	wire [4-1:0] node36237;
	wire [4-1:0] node36241;
	wire [4-1:0] node36242;
	wire [4-1:0] node36243;
	wire [4-1:0] node36244;
	wire [4-1:0] node36248;
	wire [4-1:0] node36249;
	wire [4-1:0] node36254;
	wire [4-1:0] node36255;
	wire [4-1:0] node36256;
	wire [4-1:0] node36257;
	wire [4-1:0] node36258;
	wire [4-1:0] node36262;
	wire [4-1:0] node36265;
	wire [4-1:0] node36267;
	wire [4-1:0] node36270;
	wire [4-1:0] node36271;
	wire [4-1:0] node36272;
	wire [4-1:0] node36274;
	wire [4-1:0] node36278;
	wire [4-1:0] node36279;
	wire [4-1:0] node36283;
	wire [4-1:0] node36284;
	wire [4-1:0] node36285;
	wire [4-1:0] node36286;
	wire [4-1:0] node36287;
	wire [4-1:0] node36288;
	wire [4-1:0] node36289;
	wire [4-1:0] node36290;
	wire [4-1:0] node36292;
	wire [4-1:0] node36295;
	wire [4-1:0] node36296;
	wire [4-1:0] node36299;
	wire [4-1:0] node36302;
	wire [4-1:0] node36303;
	wire [4-1:0] node36305;
	wire [4-1:0] node36308;
	wire [4-1:0] node36309;
	wire [4-1:0] node36313;
	wire [4-1:0] node36314;
	wire [4-1:0] node36315;
	wire [4-1:0] node36317;
	wire [4-1:0] node36321;
	wire [4-1:0] node36322;
	wire [4-1:0] node36323;
	wire [4-1:0] node36326;
	wire [4-1:0] node36330;
	wire [4-1:0] node36331;
	wire [4-1:0] node36332;
	wire [4-1:0] node36333;
	wire [4-1:0] node36334;
	wire [4-1:0] node36338;
	wire [4-1:0] node36341;
	wire [4-1:0] node36342;
	wire [4-1:0] node36343;
	wire [4-1:0] node36347;
	wire [4-1:0] node36348;
	wire [4-1:0] node36351;
	wire [4-1:0] node36354;
	wire [4-1:0] node36355;
	wire [4-1:0] node36357;
	wire [4-1:0] node36358;
	wire [4-1:0] node36361;
	wire [4-1:0] node36364;
	wire [4-1:0] node36365;
	wire [4-1:0] node36367;
	wire [4-1:0] node36370;
	wire [4-1:0] node36371;
	wire [4-1:0] node36374;
	wire [4-1:0] node36377;
	wire [4-1:0] node36378;
	wire [4-1:0] node36379;
	wire [4-1:0] node36380;
	wire [4-1:0] node36381;
	wire [4-1:0] node36383;
	wire [4-1:0] node36386;
	wire [4-1:0] node36387;
	wire [4-1:0] node36391;
	wire [4-1:0] node36392;
	wire [4-1:0] node36393;
	wire [4-1:0] node36396;
	wire [4-1:0] node36399;
	wire [4-1:0] node36400;
	wire [4-1:0] node36403;
	wire [4-1:0] node36406;
	wire [4-1:0] node36407;
	wire [4-1:0] node36408;
	wire [4-1:0] node36411;
	wire [4-1:0] node36412;
	wire [4-1:0] node36415;
	wire [4-1:0] node36418;
	wire [4-1:0] node36419;
	wire [4-1:0] node36420;
	wire [4-1:0] node36423;
	wire [4-1:0] node36426;
	wire [4-1:0] node36427;
	wire [4-1:0] node36431;
	wire [4-1:0] node36432;
	wire [4-1:0] node36433;
	wire [4-1:0] node36435;
	wire [4-1:0] node36437;
	wire [4-1:0] node36440;
	wire [4-1:0] node36441;
	wire [4-1:0] node36442;
	wire [4-1:0] node36445;
	wire [4-1:0] node36448;
	wire [4-1:0] node36449;
	wire [4-1:0] node36452;
	wire [4-1:0] node36455;
	wire [4-1:0] node36456;
	wire [4-1:0] node36457;
	wire [4-1:0] node36458;
	wire [4-1:0] node36462;
	wire [4-1:0] node36464;
	wire [4-1:0] node36467;
	wire [4-1:0] node36468;
	wire [4-1:0] node36469;
	wire [4-1:0] node36472;
	wire [4-1:0] node36476;
	wire [4-1:0] node36477;
	wire [4-1:0] node36478;
	wire [4-1:0] node36479;
	wire [4-1:0] node36480;
	wire [4-1:0] node36481;
	wire [4-1:0] node36482;
	wire [4-1:0] node36485;
	wire [4-1:0] node36488;
	wire [4-1:0] node36491;
	wire [4-1:0] node36492;
	wire [4-1:0] node36495;
	wire [4-1:0] node36498;
	wire [4-1:0] node36499;
	wire [4-1:0] node36500;
	wire [4-1:0] node36502;
	wire [4-1:0] node36505;
	wire [4-1:0] node36506;
	wire [4-1:0] node36510;
	wire [4-1:0] node36511;
	wire [4-1:0] node36514;
	wire [4-1:0] node36515;
	wire [4-1:0] node36519;
	wire [4-1:0] node36520;
	wire [4-1:0] node36521;
	wire [4-1:0] node36522;
	wire [4-1:0] node36523;
	wire [4-1:0] node36526;
	wire [4-1:0] node36529;
	wire [4-1:0] node36530;
	wire [4-1:0] node36534;
	wire [4-1:0] node36535;
	wire [4-1:0] node36538;
	wire [4-1:0] node36540;
	wire [4-1:0] node36543;
	wire [4-1:0] node36544;
	wire [4-1:0] node36545;
	wire [4-1:0] node36547;
	wire [4-1:0] node36551;
	wire [4-1:0] node36554;
	wire [4-1:0] node36555;
	wire [4-1:0] node36556;
	wire [4-1:0] node36557;
	wire [4-1:0] node36558;
	wire [4-1:0] node36559;
	wire [4-1:0] node36562;
	wire [4-1:0] node36566;
	wire [4-1:0] node36567;
	wire [4-1:0] node36570;
	wire [4-1:0] node36573;
	wire [4-1:0] node36574;
	wire [4-1:0] node36575;
	wire [4-1:0] node36577;
	wire [4-1:0] node36580;
	wire [4-1:0] node36582;
	wire [4-1:0] node36585;
	wire [4-1:0] node36587;
	wire [4-1:0] node36588;
	wire [4-1:0] node36592;
	wire [4-1:0] node36593;
	wire [4-1:0] node36594;
	wire [4-1:0] node36595;
	wire [4-1:0] node36596;
	wire [4-1:0] node36599;
	wire [4-1:0] node36602;
	wire [4-1:0] node36603;
	wire [4-1:0] node36607;
	wire [4-1:0] node36608;
	wire [4-1:0] node36610;
	wire [4-1:0] node36613;
	wire [4-1:0] node36616;
	wire [4-1:0] node36617;
	wire [4-1:0] node36618;
	wire [4-1:0] node36621;
	wire [4-1:0] node36622;
	wire [4-1:0] node36626;
	wire [4-1:0] node36629;
	wire [4-1:0] node36630;
	wire [4-1:0] node36631;
	wire [4-1:0] node36632;
	wire [4-1:0] node36633;
	wire [4-1:0] node36634;
	wire [4-1:0] node36635;
	wire [4-1:0] node36636;
	wire [4-1:0] node36639;
	wire [4-1:0] node36643;
	wire [4-1:0] node36644;
	wire [4-1:0] node36645;
	wire [4-1:0] node36648;
	wire [4-1:0] node36652;
	wire [4-1:0] node36653;
	wire [4-1:0] node36654;
	wire [4-1:0] node36656;
	wire [4-1:0] node36659;
	wire [4-1:0] node36660;
	wire [4-1:0] node36663;
	wire [4-1:0] node36666;
	wire [4-1:0] node36667;
	wire [4-1:0] node36669;
	wire [4-1:0] node36672;
	wire [4-1:0] node36673;
	wire [4-1:0] node36677;
	wire [4-1:0] node36678;
	wire [4-1:0] node36679;
	wire [4-1:0] node36680;
	wire [4-1:0] node36683;
	wire [4-1:0] node36686;
	wire [4-1:0] node36687;
	wire [4-1:0] node36688;
	wire [4-1:0] node36691;
	wire [4-1:0] node36695;
	wire [4-1:0] node36696;
	wire [4-1:0] node36698;
	wire [4-1:0] node36701;
	wire [4-1:0] node36702;
	wire [4-1:0] node36704;
	wire [4-1:0] node36707;
	wire [4-1:0] node36708;
	wire [4-1:0] node36712;
	wire [4-1:0] node36713;
	wire [4-1:0] node36714;
	wire [4-1:0] node36715;
	wire [4-1:0] node36716;
	wire [4-1:0] node36719;
	wire [4-1:0] node36722;
	wire [4-1:0] node36723;
	wire [4-1:0] node36724;
	wire [4-1:0] node36728;
	wire [4-1:0] node36729;
	wire [4-1:0] node36733;
	wire [4-1:0] node36734;
	wire [4-1:0] node36735;
	wire [4-1:0] node36736;
	wire [4-1:0] node36739;
	wire [4-1:0] node36742;
	wire [4-1:0] node36745;
	wire [4-1:0] node36746;
	wire [4-1:0] node36747;
	wire [4-1:0] node36751;
	wire [4-1:0] node36754;
	wire [4-1:0] node36755;
	wire [4-1:0] node36756;
	wire [4-1:0] node36757;
	wire [4-1:0] node36760;
	wire [4-1:0] node36763;
	wire [4-1:0] node36764;
	wire [4-1:0] node36767;
	wire [4-1:0] node36770;
	wire [4-1:0] node36771;
	wire [4-1:0] node36772;
	wire [4-1:0] node36775;
	wire [4-1:0] node36778;
	wire [4-1:0] node36780;
	wire [4-1:0] node36781;
	wire [4-1:0] node36784;
	wire [4-1:0] node36787;
	wire [4-1:0] node36788;
	wire [4-1:0] node36789;
	wire [4-1:0] node36790;
	wire [4-1:0] node36791;
	wire [4-1:0] node36792;
	wire [4-1:0] node36794;
	wire [4-1:0] node36797;
	wire [4-1:0] node36799;
	wire [4-1:0] node36802;
	wire [4-1:0] node36803;
	wire [4-1:0] node36804;
	wire [4-1:0] node36807;
	wire [4-1:0] node36811;
	wire [4-1:0] node36812;
	wire [4-1:0] node36813;
	wire [4-1:0] node36815;
	wire [4-1:0] node36818;
	wire [4-1:0] node36819;
	wire [4-1:0] node36823;
	wire [4-1:0] node36824;
	wire [4-1:0] node36826;
	wire [4-1:0] node36830;
	wire [4-1:0] node36831;
	wire [4-1:0] node36832;
	wire [4-1:0] node36833;
	wire [4-1:0] node36834;
	wire [4-1:0] node36837;
	wire [4-1:0] node36841;
	wire [4-1:0] node36842;
	wire [4-1:0] node36845;
	wire [4-1:0] node36846;
	wire [4-1:0] node36850;
	wire [4-1:0] node36852;
	wire [4-1:0] node36853;
	wire [4-1:0] node36856;
	wire [4-1:0] node36859;
	wire [4-1:0] node36860;
	wire [4-1:0] node36861;
	wire [4-1:0] node36862;
	wire [4-1:0] node36863;
	wire [4-1:0] node36866;
	wire [4-1:0] node36868;
	wire [4-1:0] node36871;
	wire [4-1:0] node36872;
	wire [4-1:0] node36873;
	wire [4-1:0] node36876;
	wire [4-1:0] node36880;
	wire [4-1:0] node36881;
	wire [4-1:0] node36882;
	wire [4-1:0] node36883;
	wire [4-1:0] node36886;
	wire [4-1:0] node36890;
	wire [4-1:0] node36891;
	wire [4-1:0] node36894;
	wire [4-1:0] node36897;
	wire [4-1:0] node36898;
	wire [4-1:0] node36899;
	wire [4-1:0] node36900;
	wire [4-1:0] node36903;
	wire [4-1:0] node36905;
	wire [4-1:0] node36908;
	wire [4-1:0] node36910;
	wire [4-1:0] node36913;
	wire [4-1:0] node36914;
	wire [4-1:0] node36915;
	wire [4-1:0] node36916;
	wire [4-1:0] node36920;
	wire [4-1:0] node36922;
	wire [4-1:0] node36925;
	wire [4-1:0] node36926;
	wire [4-1:0] node36929;
	wire [4-1:0] node36932;
	wire [4-1:0] node36933;
	wire [4-1:0] node36934;
	wire [4-1:0] node36935;
	wire [4-1:0] node36936;
	wire [4-1:0] node36937;
	wire [4-1:0] node36938;
	wire [4-1:0] node36939;
	wire [4-1:0] node36942;
	wire [4-1:0] node36943;
	wire [4-1:0] node36946;
	wire [4-1:0] node36949;
	wire [4-1:0] node36950;
	wire [4-1:0] node36951;
	wire [4-1:0] node36954;
	wire [4-1:0] node36957;
	wire [4-1:0] node36958;
	wire [4-1:0] node36961;
	wire [4-1:0] node36964;
	wire [4-1:0] node36965;
	wire [4-1:0] node36966;
	wire [4-1:0] node36967;
	wire [4-1:0] node36970;
	wire [4-1:0] node36973;
	wire [4-1:0] node36974;
	wire [4-1:0] node36977;
	wire [4-1:0] node36980;
	wire [4-1:0] node36981;
	wire [4-1:0] node36983;
	wire [4-1:0] node36986;
	wire [4-1:0] node36987;
	wire [4-1:0] node36991;
	wire [4-1:0] node36992;
	wire [4-1:0] node36993;
	wire [4-1:0] node36994;
	wire [4-1:0] node36997;
	wire [4-1:0] node37000;
	wire [4-1:0] node37001;
	wire [4-1:0] node37002;
	wire [4-1:0] node37005;
	wire [4-1:0] node37008;
	wire [4-1:0] node37010;
	wire [4-1:0] node37013;
	wire [4-1:0] node37014;
	wire [4-1:0] node37016;
	wire [4-1:0] node37017;
	wire [4-1:0] node37021;
	wire [4-1:0] node37022;
	wire [4-1:0] node37026;
	wire [4-1:0] node37027;
	wire [4-1:0] node37028;
	wire [4-1:0] node37029;
	wire [4-1:0] node37030;
	wire [4-1:0] node37032;
	wire [4-1:0] node37035;
	wire [4-1:0] node37037;
	wire [4-1:0] node37040;
	wire [4-1:0] node37041;
	wire [4-1:0] node37042;
	wire [4-1:0] node37043;
	wire [4-1:0] node37046;
	wire [4-1:0] node37049;
	wire [4-1:0] node37050;
	wire [4-1:0] node37053;
	wire [4-1:0] node37056;
	wire [4-1:0] node37057;
	wire [4-1:0] node37058;
	wire [4-1:0] node37061;
	wire [4-1:0] node37064;
	wire [4-1:0] node37066;
	wire [4-1:0] node37069;
	wire [4-1:0] node37070;
	wire [4-1:0] node37071;
	wire [4-1:0] node37073;
	wire [4-1:0] node37076;
	wire [4-1:0] node37077;
	wire [4-1:0] node37081;
	wire [4-1:0] node37084;
	wire [4-1:0] node37085;
	wire [4-1:0] node37086;
	wire [4-1:0] node37087;
	wire [4-1:0] node37089;
	wire [4-1:0] node37092;
	wire [4-1:0] node37094;
	wire [4-1:0] node37097;
	wire [4-1:0] node37098;
	wire [4-1:0] node37099;
	wire [4-1:0] node37100;
	wire [4-1:0] node37101;
	wire [4-1:0] node37105;
	wire [4-1:0] node37106;
	wire [4-1:0] node37109;
	wire [4-1:0] node37112;
	wire [4-1:0] node37114;
	wire [4-1:0] node37117;
	wire [4-1:0] node37118;
	wire [4-1:0] node37119;
	wire [4-1:0] node37122;
	wire [4-1:0] node37125;
	wire [4-1:0] node37127;
	wire [4-1:0] node37130;
	wire [4-1:0] node37131;
	wire [4-1:0] node37132;
	wire [4-1:0] node37134;
	wire [4-1:0] node37137;
	wire [4-1:0] node37138;
	wire [4-1:0] node37142;
	wire [4-1:0] node37145;
	wire [4-1:0] node37146;
	wire [4-1:0] node37147;
	wire [4-1:0] node37148;
	wire [4-1:0] node37149;
	wire [4-1:0] node37150;
	wire [4-1:0] node37153;
	wire [4-1:0] node37154;
	wire [4-1:0] node37158;
	wire [4-1:0] node37159;
	wire [4-1:0] node37160;
	wire [4-1:0] node37163;
	wire [4-1:0] node37166;
	wire [4-1:0] node37167;
	wire [4-1:0] node37170;
	wire [4-1:0] node37173;
	wire [4-1:0] node37174;
	wire [4-1:0] node37175;
	wire [4-1:0] node37177;
	wire [4-1:0] node37180;
	wire [4-1:0] node37181;
	wire [4-1:0] node37185;
	wire [4-1:0] node37186;
	wire [4-1:0] node37187;
	wire [4-1:0] node37190;
	wire [4-1:0] node37193;
	wire [4-1:0] node37194;
	wire [4-1:0] node37198;
	wire [4-1:0] node37199;
	wire [4-1:0] node37200;
	wire [4-1:0] node37201;
	wire [4-1:0] node37202;
	wire [4-1:0] node37206;
	wire [4-1:0] node37208;
	wire [4-1:0] node37211;
	wire [4-1:0] node37212;
	wire [4-1:0] node37214;
	wire [4-1:0] node37215;
	wire [4-1:0] node37218;
	wire [4-1:0] node37219;
	wire [4-1:0] node37223;
	wire [4-1:0] node37224;
	wire [4-1:0] node37225;
	wire [4-1:0] node37226;
	wire [4-1:0] node37230;
	wire [4-1:0] node37231;
	wire [4-1:0] node37234;
	wire [4-1:0] node37237;
	wire [4-1:0] node37238;
	wire [4-1:0] node37239;
	wire [4-1:0] node37242;
	wire [4-1:0] node37246;
	wire [4-1:0] node37247;
	wire [4-1:0] node37248;
	wire [4-1:0] node37250;
	wire [4-1:0] node37253;
	wire [4-1:0] node37254;
	wire [4-1:0] node37258;
	wire [4-1:0] node37261;
	wire [4-1:0] node37262;
	wire [4-1:0] node37263;
	wire [4-1:0] node37264;
	wire [4-1:0] node37266;
	wire [4-1:0] node37269;
	wire [4-1:0] node37270;
	wire [4-1:0] node37272;
	wire [4-1:0] node37276;
	wire [4-1:0] node37277;
	wire [4-1:0] node37278;
	wire [4-1:0] node37279;
	wire [4-1:0] node37283;
	wire [4-1:0] node37284;
	wire [4-1:0] node37285;
	wire [4-1:0] node37289;
	wire [4-1:0] node37290;
	wire [4-1:0] node37293;
	wire [4-1:0] node37296;
	wire [4-1:0] node37297;
	wire [4-1:0] node37301;
	wire [4-1:0] node37302;
	wire [4-1:0] node37303;
	wire [4-1:0] node37304;
	wire [4-1:0] node37305;
	wire [4-1:0] node37309;
	wire [4-1:0] node37310;
	wire [4-1:0] node37314;
	wire [4-1:0] node37315;
	wire [4-1:0] node37317;
	wire [4-1:0] node37318;
	wire [4-1:0] node37320;
	wire [4-1:0] node37323;
	wire [4-1:0] node37325;
	wire [4-1:0] node37328;
	wire [4-1:0] node37329;
	wire [4-1:0] node37332;
	wire [4-1:0] node37335;
	wire [4-1:0] node37336;
	wire [4-1:0] node37337;
	wire [4-1:0] node37339;
	wire [4-1:0] node37342;
	wire [4-1:0] node37343;
	wire [4-1:0] node37347;
	wire [4-1:0] node37350;
	wire [4-1:0] node37351;
	wire [4-1:0] node37352;
	wire [4-1:0] node37353;
	wire [4-1:0] node37354;
	wire [4-1:0] node37355;
	wire [4-1:0] node37356;
	wire [4-1:0] node37359;
	wire [4-1:0] node37360;
	wire [4-1:0] node37363;
	wire [4-1:0] node37366;
	wire [4-1:0] node37367;
	wire [4-1:0] node37368;
	wire [4-1:0] node37371;
	wire [4-1:0] node37374;
	wire [4-1:0] node37375;
	wire [4-1:0] node37378;
	wire [4-1:0] node37381;
	wire [4-1:0] node37382;
	wire [4-1:0] node37383;
	wire [4-1:0] node37384;
	wire [4-1:0] node37387;
	wire [4-1:0] node37390;
	wire [4-1:0] node37391;
	wire [4-1:0] node37394;
	wire [4-1:0] node37397;
	wire [4-1:0] node37398;
	wire [4-1:0] node37400;
	wire [4-1:0] node37403;
	wire [4-1:0] node37404;
	wire [4-1:0] node37407;
	wire [4-1:0] node37410;
	wire [4-1:0] node37411;
	wire [4-1:0] node37412;
	wire [4-1:0] node37413;
	wire [4-1:0] node37415;
	wire [4-1:0] node37418;
	wire [4-1:0] node37419;
	wire [4-1:0] node37423;
	wire [4-1:0] node37424;
	wire [4-1:0] node37425;
	wire [4-1:0] node37427;
	wire [4-1:0] node37430;
	wire [4-1:0] node37431;
	wire [4-1:0] node37434;
	wire [4-1:0] node37437;
	wire [4-1:0] node37438;
	wire [4-1:0] node37439;
	wire [4-1:0] node37443;
	wire [4-1:0] node37444;
	wire [4-1:0] node37447;
	wire [4-1:0] node37450;
	wire [4-1:0] node37451;
	wire [4-1:0] node37452;
	wire [4-1:0] node37454;
	wire [4-1:0] node37457;
	wire [4-1:0] node37458;
	wire [4-1:0] node37462;
	wire [4-1:0] node37465;
	wire [4-1:0] node37466;
	wire [4-1:0] node37467;
	wire [4-1:0] node37468;
	wire [4-1:0] node37469;
	wire [4-1:0] node37471;
	wire [4-1:0] node37474;
	wire [4-1:0] node37477;
	wire [4-1:0] node37478;
	wire [4-1:0] node37481;
	wire [4-1:0] node37482;
	wire [4-1:0] node37485;
	wire [4-1:0] node37488;
	wire [4-1:0] node37489;
	wire [4-1:0] node37490;
	wire [4-1:0] node37491;
	wire [4-1:0] node37495;
	wire [4-1:0] node37496;
	wire [4-1:0] node37499;
	wire [4-1:0] node37502;
	wire [4-1:0] node37503;
	wire [4-1:0] node37504;
	wire [4-1:0] node37505;
	wire [4-1:0] node37508;
	wire [4-1:0] node37511;
	wire [4-1:0] node37512;
	wire [4-1:0] node37514;
	wire [4-1:0] node37518;
	wire [4-1:0] node37519;
	wire [4-1:0] node37522;
	wire [4-1:0] node37525;
	wire [4-1:0] node37526;
	wire [4-1:0] node37527;
	wire [4-1:0] node37528;
	wire [4-1:0] node37531;
	wire [4-1:0] node37534;
	wire [4-1:0] node37535;
	wire [4-1:0] node37537;
	wire [4-1:0] node37541;
	wire [4-1:0] node37544;
	wire [4-1:0] node37545;
	wire [4-1:0] node37546;
	wire [4-1:0] node37547;
	wire [4-1:0] node37548;
	wire [4-1:0] node37549;
	wire [4-1:0] node37552;
	wire [4-1:0] node37553;
	wire [4-1:0] node37556;
	wire [4-1:0] node37559;
	wire [4-1:0] node37560;
	wire [4-1:0] node37561;
	wire [4-1:0] node37562;
	wire [4-1:0] node37565;
	wire [4-1:0] node37568;
	wire [4-1:0] node37569;
	wire [4-1:0] node37573;
	wire [4-1:0] node37574;
	wire [4-1:0] node37575;
	wire [4-1:0] node37578;
	wire [4-1:0] node37581;
	wire [4-1:0] node37582;
	wire [4-1:0] node37585;
	wire [4-1:0] node37588;
	wire [4-1:0] node37589;
	wire [4-1:0] node37590;
	wire [4-1:0] node37592;
	wire [4-1:0] node37595;
	wire [4-1:0] node37596;
	wire [4-1:0] node37599;
	wire [4-1:0] node37602;
	wire [4-1:0] node37603;
	wire [4-1:0] node37604;
	wire [4-1:0] node37608;
	wire [4-1:0] node37609;
	wire [4-1:0] node37613;
	wire [4-1:0] node37614;
	wire [4-1:0] node37615;
	wire [4-1:0] node37616;
	wire [4-1:0] node37617;
	wire [4-1:0] node37621;
	wire [4-1:0] node37623;
	wire [4-1:0] node37626;
	wire [4-1:0] node37627;
	wire [4-1:0] node37628;
	wire [4-1:0] node37629;
	wire [4-1:0] node37632;
	wire [4-1:0] node37635;
	wire [4-1:0] node37636;
	wire [4-1:0] node37639;
	wire [4-1:0] node37642;
	wire [4-1:0] node37643;
	wire [4-1:0] node37645;
	wire [4-1:0] node37648;
	wire [4-1:0] node37649;
	wire [4-1:0] node37650;
	wire [4-1:0] node37653;
	wire [4-1:0] node37657;
	wire [4-1:0] node37658;
	wire [4-1:0] node37659;
	wire [4-1:0] node37661;
	wire [4-1:0] node37664;
	wire [4-1:0] node37665;
	wire [4-1:0] node37669;
	wire [4-1:0] node37672;
	wire [4-1:0] node37673;
	wire [4-1:0] node37674;
	wire [4-1:0] node37675;
	wire [4-1:0] node37676;
	wire [4-1:0] node37679;
	wire [4-1:0] node37680;
	wire [4-1:0] node37684;
	wire [4-1:0] node37685;
	wire [4-1:0] node37688;
	wire [4-1:0] node37689;
	wire [4-1:0] node37691;
	wire [4-1:0] node37694;
	wire [4-1:0] node37695;
	wire [4-1:0] node37699;
	wire [4-1:0] node37700;
	wire [4-1:0] node37701;
	wire [4-1:0] node37702;
	wire [4-1:0] node37704;
	wire [4-1:0] node37707;
	wire [4-1:0] node37708;
	wire [4-1:0] node37711;
	wire [4-1:0] node37714;
	wire [4-1:0] node37716;
	wire [4-1:0] node37719;
	wire [4-1:0] node37720;
	wire [4-1:0] node37721;
	wire [4-1:0] node37725;
	wire [4-1:0] node37726;
	wire [4-1:0] node37729;
	wire [4-1:0] node37732;
	wire [4-1:0] node37733;
	wire [4-1:0] node37734;
	wire [4-1:0] node37735;
	wire [4-1:0] node37738;
	wire [4-1:0] node37741;
	wire [4-1:0] node37742;
	wire [4-1:0] node37744;
	wire [4-1:0] node37748;
	wire [4-1:0] node37751;
	wire [4-1:0] node37752;
	wire [4-1:0] node37753;
	wire [4-1:0] node37754;
	wire [4-1:0] node37755;
	wire [4-1:0] node37756;
	wire [4-1:0] node37757;
	wire [4-1:0] node37758;
	wire [4-1:0] node37759;
	wire [4-1:0] node37760;
	wire [4-1:0] node37761;
	wire [4-1:0] node37763;
	wire [4-1:0] node37766;
	wire [4-1:0] node37769;
	wire [4-1:0] node37770;
	wire [4-1:0] node37771;
	wire [4-1:0] node37775;
	wire [4-1:0] node37777;
	wire [4-1:0] node37780;
	wire [4-1:0] node37781;
	wire [4-1:0] node37782;
	wire [4-1:0] node37783;
	wire [4-1:0] node37786;
	wire [4-1:0] node37789;
	wire [4-1:0] node37792;
	wire [4-1:0] node37793;
	wire [4-1:0] node37794;
	wire [4-1:0] node37798;
	wire [4-1:0] node37799;
	wire [4-1:0] node37803;
	wire [4-1:0] node37804;
	wire [4-1:0] node37805;
	wire [4-1:0] node37807;
	wire [4-1:0] node37809;
	wire [4-1:0] node37812;
	wire [4-1:0] node37813;
	wire [4-1:0] node37816;
	wire [4-1:0] node37817;
	wire [4-1:0] node37821;
	wire [4-1:0] node37822;
	wire [4-1:0] node37823;
	wire [4-1:0] node37827;
	wire [4-1:0] node37828;
	wire [4-1:0] node37831;
	wire [4-1:0] node37832;
	wire [4-1:0] node37836;
	wire [4-1:0] node37837;
	wire [4-1:0] node37838;
	wire [4-1:0] node37839;
	wire [4-1:0] node37840;
	wire [4-1:0] node37843;
	wire [4-1:0] node37846;
	wire [4-1:0] node37847;
	wire [4-1:0] node37850;
	wire [4-1:0] node37853;
	wire [4-1:0] node37854;
	wire [4-1:0] node37855;
	wire [4-1:0] node37857;
	wire [4-1:0] node37860;
	wire [4-1:0] node37863;
	wire [4-1:0] node37864;
	wire [4-1:0] node37867;
	wire [4-1:0] node37868;
	wire [4-1:0] node37872;
	wire [4-1:0] node37873;
	wire [4-1:0] node37874;
	wire [4-1:0] node37875;
	wire [4-1:0] node37878;
	wire [4-1:0] node37881;
	wire [4-1:0] node37882;
	wire [4-1:0] node37885;
	wire [4-1:0] node37886;
	wire [4-1:0] node37890;
	wire [4-1:0] node37891;
	wire [4-1:0] node37892;
	wire [4-1:0] node37894;
	wire [4-1:0] node37897;
	wire [4-1:0] node37898;
	wire [4-1:0] node37902;
	wire [4-1:0] node37903;
	wire [4-1:0] node37905;
	wire [4-1:0] node37909;
	wire [4-1:0] node37910;
	wire [4-1:0] node37911;
	wire [4-1:0] node37912;
	wire [4-1:0] node37914;
	wire [4-1:0] node37916;
	wire [4-1:0] node37919;
	wire [4-1:0] node37920;
	wire [4-1:0] node37922;
	wire [4-1:0] node37925;
	wire [4-1:0] node37926;
	wire [4-1:0] node37929;
	wire [4-1:0] node37930;
	wire [4-1:0] node37934;
	wire [4-1:0] node37935;
	wire [4-1:0] node37936;
	wire [4-1:0] node37937;
	wire [4-1:0] node37938;
	wire [4-1:0] node37942;
	wire [4-1:0] node37945;
	wire [4-1:0] node37948;
	wire [4-1:0] node37949;
	wire [4-1:0] node37950;
	wire [4-1:0] node37951;
	wire [4-1:0] node37955;
	wire [4-1:0] node37958;
	wire [4-1:0] node37960;
	wire [4-1:0] node37963;
	wire [4-1:0] node37964;
	wire [4-1:0] node37965;
	wire [4-1:0] node37966;
	wire [4-1:0] node37968;
	wire [4-1:0] node37969;
	wire [4-1:0] node37973;
	wire [4-1:0] node37975;
	wire [4-1:0] node37978;
	wire [4-1:0] node37979;
	wire [4-1:0] node37980;
	wire [4-1:0] node37981;
	wire [4-1:0] node37985;
	wire [4-1:0] node37987;
	wire [4-1:0] node37990;
	wire [4-1:0] node37992;
	wire [4-1:0] node37995;
	wire [4-1:0] node37996;
	wire [4-1:0] node37997;
	wire [4-1:0] node37999;
	wire [4-1:0] node38001;
	wire [4-1:0] node38004;
	wire [4-1:0] node38007;
	wire [4-1:0] node38008;
	wire [4-1:0] node38009;
	wire [4-1:0] node38010;
	wire [4-1:0] node38014;
	wire [4-1:0] node38016;
	wire [4-1:0] node38019;
	wire [4-1:0] node38020;
	wire [4-1:0] node38024;
	wire [4-1:0] node38025;
	wire [4-1:0] node38026;
	wire [4-1:0] node38027;
	wire [4-1:0] node38028;
	wire [4-1:0] node38029;
	wire [4-1:0] node38031;
	wire [4-1:0] node38034;
	wire [4-1:0] node38035;
	wire [4-1:0] node38036;
	wire [4-1:0] node38040;
	wire [4-1:0] node38041;
	wire [4-1:0] node38045;
	wire [4-1:0] node38046;
	wire [4-1:0] node38047;
	wire [4-1:0] node38050;
	wire [4-1:0] node38053;
	wire [4-1:0] node38055;
	wire [4-1:0] node38056;
	wire [4-1:0] node38060;
	wire [4-1:0] node38061;
	wire [4-1:0] node38062;
	wire [4-1:0] node38063;
	wire [4-1:0] node38065;
	wire [4-1:0] node38068;
	wire [4-1:0] node38071;
	wire [4-1:0] node38073;
	wire [4-1:0] node38075;
	wire [4-1:0] node38078;
	wire [4-1:0] node38079;
	wire [4-1:0] node38081;
	wire [4-1:0] node38084;
	wire [4-1:0] node38086;
	wire [4-1:0] node38089;
	wire [4-1:0] node38090;
	wire [4-1:0] node38091;
	wire [4-1:0] node38092;
	wire [4-1:0] node38094;
	wire [4-1:0] node38097;
	wire [4-1:0] node38098;
	wire [4-1:0] node38099;
	wire [4-1:0] node38103;
	wire [4-1:0] node38104;
	wire [4-1:0] node38108;
	wire [4-1:0] node38109;
	wire [4-1:0] node38110;
	wire [4-1:0] node38112;
	wire [4-1:0] node38115;
	wire [4-1:0] node38117;
	wire [4-1:0] node38120;
	wire [4-1:0] node38122;
	wire [4-1:0] node38125;
	wire [4-1:0] node38126;
	wire [4-1:0] node38127;
	wire [4-1:0] node38128;
	wire [4-1:0] node38132;
	wire [4-1:0] node38133;
	wire [4-1:0] node38137;
	wire [4-1:0] node38138;
	wire [4-1:0] node38139;
	wire [4-1:0] node38143;
	wire [4-1:0] node38144;
	wire [4-1:0] node38148;
	wire [4-1:0] node38149;
	wire [4-1:0] node38150;
	wire [4-1:0] node38151;
	wire [4-1:0] node38152;
	wire [4-1:0] node38153;
	wire [4-1:0] node38154;
	wire [4-1:0] node38157;
	wire [4-1:0] node38161;
	wire [4-1:0] node38162;
	wire [4-1:0] node38163;
	wire [4-1:0] node38167;
	wire [4-1:0] node38168;
	wire [4-1:0] node38172;
	wire [4-1:0] node38173;
	wire [4-1:0] node38174;
	wire [4-1:0] node38177;
	wire [4-1:0] node38178;
	wire [4-1:0] node38182;
	wire [4-1:0] node38183;
	wire [4-1:0] node38187;
	wire [4-1:0] node38188;
	wire [4-1:0] node38189;
	wire [4-1:0] node38190;
	wire [4-1:0] node38194;
	wire [4-1:0] node38195;
	wire [4-1:0] node38199;
	wire [4-1:0] node38200;
	wire [4-1:0] node38201;
	wire [4-1:0] node38205;
	wire [4-1:0] node38208;
	wire [4-1:0] node38209;
	wire [4-1:0] node38210;
	wire [4-1:0] node38211;
	wire [4-1:0] node38213;
	wire [4-1:0] node38216;
	wire [4-1:0] node38217;
	wire [4-1:0] node38220;
	wire [4-1:0] node38222;
	wire [4-1:0] node38225;
	wire [4-1:0] node38226;
	wire [4-1:0] node38227;
	wire [4-1:0] node38230;
	wire [4-1:0] node38233;
	wire [4-1:0] node38234;
	wire [4-1:0] node38236;
	wire [4-1:0] node38240;
	wire [4-1:0] node38241;
	wire [4-1:0] node38242;
	wire [4-1:0] node38243;
	wire [4-1:0] node38247;
	wire [4-1:0] node38250;
	wire [4-1:0] node38251;
	wire [4-1:0] node38252;
	wire [4-1:0] node38256;
	wire [4-1:0] node38257;
	wire [4-1:0] node38261;
	wire [4-1:0] node38262;
	wire [4-1:0] node38263;
	wire [4-1:0] node38264;
	wire [4-1:0] node38265;
	wire [4-1:0] node38266;
	wire [4-1:0] node38267;
	wire [4-1:0] node38268;
	wire [4-1:0] node38271;
	wire [4-1:0] node38274;
	wire [4-1:0] node38276;
	wire [4-1:0] node38277;
	wire [4-1:0] node38281;
	wire [4-1:0] node38282;
	wire [4-1:0] node38283;
	wire [4-1:0] node38285;
	wire [4-1:0] node38288;
	wire [4-1:0] node38289;
	wire [4-1:0] node38293;
	wire [4-1:0] node38294;
	wire [4-1:0] node38297;
	wire [4-1:0] node38300;
	wire [4-1:0] node38301;
	wire [4-1:0] node38302;
	wire [4-1:0] node38303;
	wire [4-1:0] node38306;
	wire [4-1:0] node38309;
	wire [4-1:0] node38310;
	wire [4-1:0] node38313;
	wire [4-1:0] node38315;
	wire [4-1:0] node38318;
	wire [4-1:0] node38319;
	wire [4-1:0] node38320;
	wire [4-1:0] node38323;
	wire [4-1:0] node38325;
	wire [4-1:0] node38328;
	wire [4-1:0] node38329;
	wire [4-1:0] node38332;
	wire [4-1:0] node38335;
	wire [4-1:0] node38336;
	wire [4-1:0] node38337;
	wire [4-1:0] node38338;
	wire [4-1:0] node38339;
	wire [4-1:0] node38340;
	wire [4-1:0] node38343;
	wire [4-1:0] node38346;
	wire [4-1:0] node38348;
	wire [4-1:0] node38351;
	wire [4-1:0] node38352;
	wire [4-1:0] node38353;
	wire [4-1:0] node38357;
	wire [4-1:0] node38359;
	wire [4-1:0] node38362;
	wire [4-1:0] node38363;
	wire [4-1:0] node38364;
	wire [4-1:0] node38365;
	wire [4-1:0] node38370;
	wire [4-1:0] node38372;
	wire [4-1:0] node38375;
	wire [4-1:0] node38376;
	wire [4-1:0] node38377;
	wire [4-1:0] node38378;
	wire [4-1:0] node38380;
	wire [4-1:0] node38383;
	wire [4-1:0] node38385;
	wire [4-1:0] node38388;
	wire [4-1:0] node38389;
	wire [4-1:0] node38390;
	wire [4-1:0] node38393;
	wire [4-1:0] node38396;
	wire [4-1:0] node38397;
	wire [4-1:0] node38400;
	wire [4-1:0] node38403;
	wire [4-1:0] node38404;
	wire [4-1:0] node38406;
	wire [4-1:0] node38407;
	wire [4-1:0] node38411;
	wire [4-1:0] node38412;
	wire [4-1:0] node38415;
	wire [4-1:0] node38418;
	wire [4-1:0] node38419;
	wire [4-1:0] node38420;
	wire [4-1:0] node38421;
	wire [4-1:0] node38422;
	wire [4-1:0] node38423;
	wire [4-1:0] node38424;
	wire [4-1:0] node38427;
	wire [4-1:0] node38430;
	wire [4-1:0] node38431;
	wire [4-1:0] node38434;
	wire [4-1:0] node38437;
	wire [4-1:0] node38438;
	wire [4-1:0] node38439;
	wire [4-1:0] node38442;
	wire [4-1:0] node38446;
	wire [4-1:0] node38447;
	wire [4-1:0] node38448;
	wire [4-1:0] node38451;
	wire [4-1:0] node38454;
	wire [4-1:0] node38455;
	wire [4-1:0] node38457;
	wire [4-1:0] node38460;
	wire [4-1:0] node38462;
	wire [4-1:0] node38465;
	wire [4-1:0] node38466;
	wire [4-1:0] node38467;
	wire [4-1:0] node38468;
	wire [4-1:0] node38471;
	wire [4-1:0] node38474;
	wire [4-1:0] node38476;
	wire [4-1:0] node38479;
	wire [4-1:0] node38480;
	wire [4-1:0] node38481;
	wire [4-1:0] node38484;
	wire [4-1:0] node38487;
	wire [4-1:0] node38488;
	wire [4-1:0] node38491;
	wire [4-1:0] node38493;
	wire [4-1:0] node38496;
	wire [4-1:0] node38497;
	wire [4-1:0] node38498;
	wire [4-1:0] node38499;
	wire [4-1:0] node38500;
	wire [4-1:0] node38503;
	wire [4-1:0] node38506;
	wire [4-1:0] node38507;
	wire [4-1:0] node38509;
	wire [4-1:0] node38512;
	wire [4-1:0] node38513;
	wire [4-1:0] node38517;
	wire [4-1:0] node38518;
	wire [4-1:0] node38519;
	wire [4-1:0] node38522;
	wire [4-1:0] node38525;
	wire [4-1:0] node38528;
	wire [4-1:0] node38529;
	wire [4-1:0] node38530;
	wire [4-1:0] node38531;
	wire [4-1:0] node38534;
	wire [4-1:0] node38537;
	wire [4-1:0] node38538;
	wire [4-1:0] node38542;
	wire [4-1:0] node38543;
	wire [4-1:0] node38544;
	wire [4-1:0] node38546;
	wire [4-1:0] node38549;
	wire [4-1:0] node38552;
	wire [4-1:0] node38553;
	wire [4-1:0] node38554;
	wire [4-1:0] node38557;
	wire [4-1:0] node38560;
	wire [4-1:0] node38561;
	wire [4-1:0] node38565;
	wire [4-1:0] node38566;
	wire [4-1:0] node38567;
	wire [4-1:0] node38568;
	wire [4-1:0] node38569;
	wire [4-1:0] node38570;
	wire [4-1:0] node38571;
	wire [4-1:0] node38574;
	wire [4-1:0] node38575;
	wire [4-1:0] node38579;
	wire [4-1:0] node38582;
	wire [4-1:0] node38583;
	wire [4-1:0] node38584;
	wire [4-1:0] node38585;
	wire [4-1:0] node38589;
	wire [4-1:0] node38590;
	wire [4-1:0] node38593;
	wire [4-1:0] node38596;
	wire [4-1:0] node38597;
	wire [4-1:0] node38598;
	wire [4-1:0] node38602;
	wire [4-1:0] node38605;
	wire [4-1:0] node38606;
	wire [4-1:0] node38607;
	wire [4-1:0] node38608;
	wire [4-1:0] node38609;
	wire [4-1:0] node38613;
	wire [4-1:0] node38616;
	wire [4-1:0] node38617;
	wire [4-1:0] node38618;
	wire [4-1:0] node38621;
	wire [4-1:0] node38624;
	wire [4-1:0] node38627;
	wire [4-1:0] node38628;
	wire [4-1:0] node38630;
	wire [4-1:0] node38631;
	wire [4-1:0] node38634;
	wire [4-1:0] node38637;
	wire [4-1:0] node38639;
	wire [4-1:0] node38642;
	wire [4-1:0] node38643;
	wire [4-1:0] node38644;
	wire [4-1:0] node38645;
	wire [4-1:0] node38646;
	wire [4-1:0] node38647;
	wire [4-1:0] node38651;
	wire [4-1:0] node38652;
	wire [4-1:0] node38656;
	wire [4-1:0] node38658;
	wire [4-1:0] node38659;
	wire [4-1:0] node38663;
	wire [4-1:0] node38664;
	wire [4-1:0] node38665;
	wire [4-1:0] node38667;
	wire [4-1:0] node38671;
	wire [4-1:0] node38672;
	wire [4-1:0] node38674;
	wire [4-1:0] node38677;
	wire [4-1:0] node38678;
	wire [4-1:0] node38681;
	wire [4-1:0] node38684;
	wire [4-1:0] node38685;
	wire [4-1:0] node38686;
	wire [4-1:0] node38687;
	wire [4-1:0] node38688;
	wire [4-1:0] node38692;
	wire [4-1:0] node38695;
	wire [4-1:0] node38697;
	wire [4-1:0] node38700;
	wire [4-1:0] node38701;
	wire [4-1:0] node38702;
	wire [4-1:0] node38705;
	wire [4-1:0] node38707;
	wire [4-1:0] node38710;
	wire [4-1:0] node38711;
	wire [4-1:0] node38713;
	wire [4-1:0] node38716;
	wire [4-1:0] node38719;
	wire [4-1:0] node38720;
	wire [4-1:0] node38721;
	wire [4-1:0] node38722;
	wire [4-1:0] node38723;
	wire [4-1:0] node38725;
	wire [4-1:0] node38726;
	wire [4-1:0] node38730;
	wire [4-1:0] node38731;
	wire [4-1:0] node38732;
	wire [4-1:0] node38735;
	wire [4-1:0] node38738;
	wire [4-1:0] node38739;
	wire [4-1:0] node38743;
	wire [4-1:0] node38744;
	wire [4-1:0] node38745;
	wire [4-1:0] node38748;
	wire [4-1:0] node38751;
	wire [4-1:0] node38752;
	wire [4-1:0] node38755;
	wire [4-1:0] node38758;
	wire [4-1:0] node38759;
	wire [4-1:0] node38760;
	wire [4-1:0] node38761;
	wire [4-1:0] node38762;
	wire [4-1:0] node38765;
	wire [4-1:0] node38768;
	wire [4-1:0] node38770;
	wire [4-1:0] node38773;
	wire [4-1:0] node38775;
	wire [4-1:0] node38778;
	wire [4-1:0] node38779;
	wire [4-1:0] node38780;
	wire [4-1:0] node38783;
	wire [4-1:0] node38786;
	wire [4-1:0] node38787;
	wire [4-1:0] node38790;
	wire [4-1:0] node38793;
	wire [4-1:0] node38794;
	wire [4-1:0] node38795;
	wire [4-1:0] node38796;
	wire [4-1:0] node38797;
	wire [4-1:0] node38800;
	wire [4-1:0] node38801;
	wire [4-1:0] node38804;
	wire [4-1:0] node38807;
	wire [4-1:0] node38808;
	wire [4-1:0] node38812;
	wire [4-1:0] node38813;
	wire [4-1:0] node38814;
	wire [4-1:0] node38815;
	wire [4-1:0] node38818;
	wire [4-1:0] node38821;
	wire [4-1:0] node38822;
	wire [4-1:0] node38825;
	wire [4-1:0] node38828;
	wire [4-1:0] node38830;
	wire [4-1:0] node38833;
	wire [4-1:0] node38834;
	wire [4-1:0] node38835;
	wire [4-1:0] node38836;
	wire [4-1:0] node38837;
	wire [4-1:0] node38840;
	wire [4-1:0] node38843;
	wire [4-1:0] node38845;
	wire [4-1:0] node38848;
	wire [4-1:0] node38849;
	wire [4-1:0] node38852;
	wire [4-1:0] node38855;
	wire [4-1:0] node38856;
	wire [4-1:0] node38857;
	wire [4-1:0] node38858;
	wire [4-1:0] node38861;
	wire [4-1:0] node38864;
	wire [4-1:0] node38866;
	wire [4-1:0] node38869;
	wire [4-1:0] node38870;
	wire [4-1:0] node38873;
	wire [4-1:0] node38876;
	wire [4-1:0] node38877;
	wire [4-1:0] node38878;
	wire [4-1:0] node38879;
	wire [4-1:0] node38880;
	wire [4-1:0] node38881;
	wire [4-1:0] node38882;
	wire [4-1:0] node38883;
	wire [4-1:0] node38885;
	wire [4-1:0] node38887;
	wire [4-1:0] node38890;
	wire [4-1:0] node38891;
	wire [4-1:0] node38892;
	wire [4-1:0] node38895;
	wire [4-1:0] node38899;
	wire [4-1:0] node38900;
	wire [4-1:0] node38901;
	wire [4-1:0] node38903;
	wire [4-1:0] node38906;
	wire [4-1:0] node38908;
	wire [4-1:0] node38911;
	wire [4-1:0] node38913;
	wire [4-1:0] node38916;
	wire [4-1:0] node38917;
	wire [4-1:0] node38918;
	wire [4-1:0] node38920;
	wire [4-1:0] node38922;
	wire [4-1:0] node38925;
	wire [4-1:0] node38926;
	wire [4-1:0] node38929;
	wire [4-1:0] node38932;
	wire [4-1:0] node38933;
	wire [4-1:0] node38934;
	wire [4-1:0] node38937;
	wire [4-1:0] node38939;
	wire [4-1:0] node38942;
	wire [4-1:0] node38944;
	wire [4-1:0] node38945;
	wire [4-1:0] node38948;
	wire [4-1:0] node38951;
	wire [4-1:0] node38952;
	wire [4-1:0] node38953;
	wire [4-1:0] node38954;
	wire [4-1:0] node38955;
	wire [4-1:0] node38957;
	wire [4-1:0] node38960;
	wire [4-1:0] node38961;
	wire [4-1:0] node38965;
	wire [4-1:0] node38966;
	wire [4-1:0] node38968;
	wire [4-1:0] node38971;
	wire [4-1:0] node38972;
	wire [4-1:0] node38976;
	wire [4-1:0] node38977;
	wire [4-1:0] node38979;
	wire [4-1:0] node38980;
	wire [4-1:0] node38983;
	wire [4-1:0] node38986;
	wire [4-1:0] node38987;
	wire [4-1:0] node38991;
	wire [4-1:0] node38992;
	wire [4-1:0] node38993;
	wire [4-1:0] node38994;
	wire [4-1:0] node38995;
	wire [4-1:0] node39000;
	wire [4-1:0] node39001;
	wire [4-1:0] node39004;
	wire [4-1:0] node39007;
	wire [4-1:0] node39008;
	wire [4-1:0] node39009;
	wire [4-1:0] node39010;
	wire [4-1:0] node39014;
	wire [4-1:0] node39015;
	wire [4-1:0] node39019;
	wire [4-1:0] node39020;
	wire [4-1:0] node39021;
	wire [4-1:0] node39026;
	wire [4-1:0] node39027;
	wire [4-1:0] node39028;
	wire [4-1:0] node39029;
	wire [4-1:0] node39030;
	wire [4-1:0] node39031;
	wire [4-1:0] node39035;
	wire [4-1:0] node39036;
	wire [4-1:0] node39037;
	wire [4-1:0] node39040;
	wire [4-1:0] node39044;
	wire [4-1:0] node39045;
	wire [4-1:0] node39048;
	wire [4-1:0] node39049;
	wire [4-1:0] node39050;
	wire [4-1:0] node39054;
	wire [4-1:0] node39055;
	wire [4-1:0] node39059;
	wire [4-1:0] node39060;
	wire [4-1:0] node39061;
	wire [4-1:0] node39062;
	wire [4-1:0] node39063;
	wire [4-1:0] node39066;
	wire [4-1:0] node39069;
	wire [4-1:0] node39070;
	wire [4-1:0] node39073;
	wire [4-1:0] node39076;
	wire [4-1:0] node39078;
	wire [4-1:0] node39081;
	wire [4-1:0] node39082;
	wire [4-1:0] node39084;
	wire [4-1:0] node39086;
	wire [4-1:0] node39089;
	wire [4-1:0] node39090;
	wire [4-1:0] node39093;
	wire [4-1:0] node39096;
	wire [4-1:0] node39097;
	wire [4-1:0] node39098;
	wire [4-1:0] node39099;
	wire [4-1:0] node39100;
	wire [4-1:0] node39101;
	wire [4-1:0] node39104;
	wire [4-1:0] node39108;
	wire [4-1:0] node39110;
	wire [4-1:0] node39113;
	wire [4-1:0] node39114;
	wire [4-1:0] node39115;
	wire [4-1:0] node39117;
	wire [4-1:0] node39121;
	wire [4-1:0] node39122;
	wire [4-1:0] node39124;
	wire [4-1:0] node39127;
	wire [4-1:0] node39129;
	wire [4-1:0] node39132;
	wire [4-1:0] node39133;
	wire [4-1:0] node39134;
	wire [4-1:0] node39135;
	wire [4-1:0] node39139;
	wire [4-1:0] node39140;
	wire [4-1:0] node39142;
	wire [4-1:0] node39146;
	wire [4-1:0] node39147;
	wire [4-1:0] node39148;
	wire [4-1:0] node39151;
	wire [4-1:0] node39152;
	wire [4-1:0] node39156;
	wire [4-1:0] node39157;
	wire [4-1:0] node39158;
	wire [4-1:0] node39162;
	wire [4-1:0] node39163;
	wire [4-1:0] node39167;
	wire [4-1:0] node39168;
	wire [4-1:0] node39169;
	wire [4-1:0] node39170;
	wire [4-1:0] node39171;
	wire [4-1:0] node39172;
	wire [4-1:0] node39173;
	wire [4-1:0] node39174;
	wire [4-1:0] node39177;
	wire [4-1:0] node39181;
	wire [4-1:0] node39182;
	wire [4-1:0] node39184;
	wire [4-1:0] node39187;
	wire [4-1:0] node39188;
	wire [4-1:0] node39192;
	wire [4-1:0] node39193;
	wire [4-1:0] node39196;
	wire [4-1:0] node39197;
	wire [4-1:0] node39200;
	wire [4-1:0] node39203;
	wire [4-1:0] node39204;
	wire [4-1:0] node39205;
	wire [4-1:0] node39206;
	wire [4-1:0] node39209;
	wire [4-1:0] node39212;
	wire [4-1:0] node39213;
	wire [4-1:0] node39215;
	wire [4-1:0] node39219;
	wire [4-1:0] node39220;
	wire [4-1:0] node39221;
	wire [4-1:0] node39225;
	wire [4-1:0] node39228;
	wire [4-1:0] node39229;
	wire [4-1:0] node39230;
	wire [4-1:0] node39231;
	wire [4-1:0] node39232;
	wire [4-1:0] node39236;
	wire [4-1:0] node39237;
	wire [4-1:0] node39240;
	wire [4-1:0] node39242;
	wire [4-1:0] node39245;
	wire [4-1:0] node39246;
	wire [4-1:0] node39247;
	wire [4-1:0] node39248;
	wire [4-1:0] node39252;
	wire [4-1:0] node39255;
	wire [4-1:0] node39256;
	wire [4-1:0] node39259;
	wire [4-1:0] node39262;
	wire [4-1:0] node39263;
	wire [4-1:0] node39264;
	wire [4-1:0] node39265;
	wire [4-1:0] node39268;
	wire [4-1:0] node39271;
	wire [4-1:0] node39272;
	wire [4-1:0] node39274;
	wire [4-1:0] node39278;
	wire [4-1:0] node39279;
	wire [4-1:0] node39281;
	wire [4-1:0] node39284;
	wire [4-1:0] node39285;
	wire [4-1:0] node39287;
	wire [4-1:0] node39291;
	wire [4-1:0] node39292;
	wire [4-1:0] node39293;
	wire [4-1:0] node39294;
	wire [4-1:0] node39295;
	wire [4-1:0] node39296;
	wire [4-1:0] node39297;
	wire [4-1:0] node39302;
	wire [4-1:0] node39303;
	wire [4-1:0] node39304;
	wire [4-1:0] node39309;
	wire [4-1:0] node39310;
	wire [4-1:0] node39311;
	wire [4-1:0] node39312;
	wire [4-1:0] node39316;
	wire [4-1:0] node39319;
	wire [4-1:0] node39320;
	wire [4-1:0] node39324;
	wire [4-1:0] node39325;
	wire [4-1:0] node39326;
	wire [4-1:0] node39328;
	wire [4-1:0] node39332;
	wire [4-1:0] node39333;
	wire [4-1:0] node39334;
	wire [4-1:0] node39338;
	wire [4-1:0] node39341;
	wire [4-1:0] node39342;
	wire [4-1:0] node39343;
	wire [4-1:0] node39344;
	wire [4-1:0] node39345;
	wire [4-1:0] node39346;
	wire [4-1:0] node39351;
	wire [4-1:0] node39353;
	wire [4-1:0] node39355;
	wire [4-1:0] node39358;
	wire [4-1:0] node39359;
	wire [4-1:0] node39360;
	wire [4-1:0] node39362;
	wire [4-1:0] node39366;
	wire [4-1:0] node39367;
	wire [4-1:0] node39371;
	wire [4-1:0] node39372;
	wire [4-1:0] node39373;
	wire [4-1:0] node39374;
	wire [4-1:0] node39375;
	wire [4-1:0] node39378;
	wire [4-1:0] node39382;
	wire [4-1:0] node39385;
	wire [4-1:0] node39386;
	wire [4-1:0] node39387;
	wire [4-1:0] node39391;
	wire [4-1:0] node39392;
	wire [4-1:0] node39394;
	wire [4-1:0] node39398;
	wire [4-1:0] node39399;
	wire [4-1:0] node39400;
	wire [4-1:0] node39401;
	wire [4-1:0] node39402;
	wire [4-1:0] node39403;
	wire [4-1:0] node39404;
	wire [4-1:0] node39405;
	wire [4-1:0] node39406;
	wire [4-1:0] node39409;
	wire [4-1:0] node39412;
	wire [4-1:0] node39415;
	wire [4-1:0] node39417;
	wire [4-1:0] node39418;
	wire [4-1:0] node39422;
	wire [4-1:0] node39423;
	wire [4-1:0] node39424;
	wire [4-1:0] node39425;
	wire [4-1:0] node39430;
	wire [4-1:0] node39431;
	wire [4-1:0] node39432;
	wire [4-1:0] node39435;
	wire [4-1:0] node39439;
	wire [4-1:0] node39440;
	wire [4-1:0] node39441;
	wire [4-1:0] node39442;
	wire [4-1:0] node39445;
	wire [4-1:0] node39448;
	wire [4-1:0] node39449;
	wire [4-1:0] node39450;
	wire [4-1:0] node39454;
	wire [4-1:0] node39457;
	wire [4-1:0] node39458;
	wire [4-1:0] node39459;
	wire [4-1:0] node39461;
	wire [4-1:0] node39464;
	wire [4-1:0] node39465;
	wire [4-1:0] node39469;
	wire [4-1:0] node39470;
	wire [4-1:0] node39472;
	wire [4-1:0] node39476;
	wire [4-1:0] node39477;
	wire [4-1:0] node39478;
	wire [4-1:0] node39479;
	wire [4-1:0] node39480;
	wire [4-1:0] node39482;
	wire [4-1:0] node39485;
	wire [4-1:0] node39486;
	wire [4-1:0] node39489;
	wire [4-1:0] node39492;
	wire [4-1:0] node39493;
	wire [4-1:0] node39494;
	wire [4-1:0] node39497;
	wire [4-1:0] node39501;
	wire [4-1:0] node39502;
	wire [4-1:0] node39503;
	wire [4-1:0] node39506;
	wire [4-1:0] node39509;
	wire [4-1:0] node39512;
	wire [4-1:0] node39513;
	wire [4-1:0] node39514;
	wire [4-1:0] node39515;
	wire [4-1:0] node39517;
	wire [4-1:0] node39521;
	wire [4-1:0] node39523;
	wire [4-1:0] node39526;
	wire [4-1:0] node39527;
	wire [4-1:0] node39528;
	wire [4-1:0] node39529;
	wire [4-1:0] node39533;
	wire [4-1:0] node39534;
	wire [4-1:0] node39538;
	wire [4-1:0] node39539;
	wire [4-1:0] node39540;
	wire [4-1:0] node39545;
	wire [4-1:0] node39546;
	wire [4-1:0] node39547;
	wire [4-1:0] node39548;
	wire [4-1:0] node39549;
	wire [4-1:0] node39550;
	wire [4-1:0] node39551;
	wire [4-1:0] node39554;
	wire [4-1:0] node39558;
	wire [4-1:0] node39559;
	wire [4-1:0] node39561;
	wire [4-1:0] node39564;
	wire [4-1:0] node39567;
	wire [4-1:0] node39568;
	wire [4-1:0] node39570;
	wire [4-1:0] node39571;
	wire [4-1:0] node39575;
	wire [4-1:0] node39577;
	wire [4-1:0] node39578;
	wire [4-1:0] node39582;
	wire [4-1:0] node39583;
	wire [4-1:0] node39584;
	wire [4-1:0] node39587;
	wire [4-1:0] node39588;
	wire [4-1:0] node39590;
	wire [4-1:0] node39594;
	wire [4-1:0] node39595;
	wire [4-1:0] node39596;
	wire [4-1:0] node39599;
	wire [4-1:0] node39600;
	wire [4-1:0] node39604;
	wire [4-1:0] node39605;
	wire [4-1:0] node39606;
	wire [4-1:0] node39611;
	wire [4-1:0] node39612;
	wire [4-1:0] node39613;
	wire [4-1:0] node39614;
	wire [4-1:0] node39615;
	wire [4-1:0] node39616;
	wire [4-1:0] node39620;
	wire [4-1:0] node39621;
	wire [4-1:0] node39625;
	wire [4-1:0] node39626;
	wire [4-1:0] node39627;
	wire [4-1:0] node39630;
	wire [4-1:0] node39634;
	wire [4-1:0] node39635;
	wire [4-1:0] node39636;
	wire [4-1:0] node39637;
	wire [4-1:0] node39641;
	wire [4-1:0] node39643;
	wire [4-1:0] node39646;
	wire [4-1:0] node39649;
	wire [4-1:0] node39650;
	wire [4-1:0] node39651;
	wire [4-1:0] node39652;
	wire [4-1:0] node39655;
	wire [4-1:0] node39659;
	wire [4-1:0] node39660;
	wire [4-1:0] node39661;
	wire [4-1:0] node39662;
	wire [4-1:0] node39668;
	wire [4-1:0] node39669;
	wire [4-1:0] node39670;
	wire [4-1:0] node39671;
	wire [4-1:0] node39672;
	wire [4-1:0] node39673;
	wire [4-1:0] node39674;
	wire [4-1:0] node39675;
	wire [4-1:0] node39678;
	wire [4-1:0] node39681;
	wire [4-1:0] node39684;
	wire [4-1:0] node39685;
	wire [4-1:0] node39686;
	wire [4-1:0] node39690;
	wire [4-1:0] node39693;
	wire [4-1:0] node39694;
	wire [4-1:0] node39695;
	wire [4-1:0] node39696;
	wire [4-1:0] node39700;
	wire [4-1:0] node39701;
	wire [4-1:0] node39705;
	wire [4-1:0] node39706;
	wire [4-1:0] node39709;
	wire [4-1:0] node39710;
	wire [4-1:0] node39714;
	wire [4-1:0] node39715;
	wire [4-1:0] node39716;
	wire [4-1:0] node39717;
	wire [4-1:0] node39718;
	wire [4-1:0] node39722;
	wire [4-1:0] node39723;
	wire [4-1:0] node39726;
	wire [4-1:0] node39729;
	wire [4-1:0] node39730;
	wire [4-1:0] node39732;
	wire [4-1:0] node39735;
	wire [4-1:0] node39736;
	wire [4-1:0] node39739;
	wire [4-1:0] node39742;
	wire [4-1:0] node39743;
	wire [4-1:0] node39744;
	wire [4-1:0] node39747;
	wire [4-1:0] node39750;
	wire [4-1:0] node39753;
	wire [4-1:0] node39754;
	wire [4-1:0] node39755;
	wire [4-1:0] node39756;
	wire [4-1:0] node39757;
	wire [4-1:0] node39758;
	wire [4-1:0] node39761;
	wire [4-1:0] node39764;
	wire [4-1:0] node39765;
	wire [4-1:0] node39769;
	wire [4-1:0] node39770;
	wire [4-1:0] node39771;
	wire [4-1:0] node39774;
	wire [4-1:0] node39778;
	wire [4-1:0] node39779;
	wire [4-1:0] node39780;
	wire [4-1:0] node39783;
	wire [4-1:0] node39786;
	wire [4-1:0] node39789;
	wire [4-1:0] node39790;
	wire [4-1:0] node39791;
	wire [4-1:0] node39792;
	wire [4-1:0] node39793;
	wire [4-1:0] node39798;
	wire [4-1:0] node39799;
	wire [4-1:0] node39800;
	wire [4-1:0] node39804;
	wire [4-1:0] node39807;
	wire [4-1:0] node39808;
	wire [4-1:0] node39809;
	wire [4-1:0] node39810;
	wire [4-1:0] node39814;
	wire [4-1:0] node39815;
	wire [4-1:0] node39819;
	wire [4-1:0] node39820;
	wire [4-1:0] node39824;
	wire [4-1:0] node39825;
	wire [4-1:0] node39826;
	wire [4-1:0] node39827;
	wire [4-1:0] node39828;
	wire [4-1:0] node39829;
	wire [4-1:0] node39830;
	wire [4-1:0] node39834;
	wire [4-1:0] node39837;
	wire [4-1:0] node39838;
	wire [4-1:0] node39839;
	wire [4-1:0] node39843;
	wire [4-1:0] node39844;
	wire [4-1:0] node39848;
	wire [4-1:0] node39850;
	wire [4-1:0] node39852;
	wire [4-1:0] node39853;
	wire [4-1:0] node39856;
	wire [4-1:0] node39859;
	wire [4-1:0] node39860;
	wire [4-1:0] node39861;
	wire [4-1:0] node39862;
	wire [4-1:0] node39863;
	wire [4-1:0] node39867;
	wire [4-1:0] node39869;
	wire [4-1:0] node39872;
	wire [4-1:0] node39873;
	wire [4-1:0] node39874;
	wire [4-1:0] node39877;
	wire [4-1:0] node39880;
	wire [4-1:0] node39883;
	wire [4-1:0] node39884;
	wire [4-1:0] node39885;
	wire [4-1:0] node39888;
	wire [4-1:0] node39891;
	wire [4-1:0] node39894;
	wire [4-1:0] node39895;
	wire [4-1:0] node39896;
	wire [4-1:0] node39897;
	wire [4-1:0] node39898;
	wire [4-1:0] node39899;
	wire [4-1:0] node39903;
	wire [4-1:0] node39904;
	wire [4-1:0] node39908;
	wire [4-1:0] node39910;
	wire [4-1:0] node39913;
	wire [4-1:0] node39914;
	wire [4-1:0] node39915;
	wire [4-1:0] node39916;
	wire [4-1:0] node39919;
	wire [4-1:0] node39922;
	wire [4-1:0] node39925;
	wire [4-1:0] node39926;
	wire [4-1:0] node39927;
	wire [4-1:0] node39931;
	wire [4-1:0] node39932;
	wire [4-1:0] node39936;
	wire [4-1:0] node39937;
	wire [4-1:0] node39938;
	wire [4-1:0] node39940;
	wire [4-1:0] node39941;
	wire [4-1:0] node39945;
	wire [4-1:0] node39946;
	wire [4-1:0] node39947;
	wire [4-1:0] node39951;
	wire [4-1:0] node39952;
	wire [4-1:0] node39956;
	wire [4-1:0] node39957;
	wire [4-1:0] node39959;
	wire [4-1:0] node39960;
	wire [4-1:0] node39963;
	wire [4-1:0] node39966;
	wire [4-1:0] node39967;
	wire [4-1:0] node39970;
	wire [4-1:0] node39973;
	wire [4-1:0] node39974;
	wire [4-1:0] node39975;
	wire [4-1:0] node39976;
	wire [4-1:0] node39977;
	wire [4-1:0] node39978;
	wire [4-1:0] node39979;
	wire [4-1:0] node39980;
	wire [4-1:0] node39981;
	wire [4-1:0] node39982;
	wire [4-1:0] node39985;
	wire [4-1:0] node39988;
	wire [4-1:0] node39989;
	wire [4-1:0] node39990;
	wire [4-1:0] node39993;
	wire [4-1:0] node39996;
	wire [4-1:0] node39997;
	wire [4-1:0] node40000;
	wire [4-1:0] node40003;
	wire [4-1:0] node40004;
	wire [4-1:0] node40007;
	wire [4-1:0] node40010;
	wire [4-1:0] node40011;
	wire [4-1:0] node40012;
	wire [4-1:0] node40015;
	wire [4-1:0] node40018;
	wire [4-1:0] node40019;
	wire [4-1:0] node40022;
	wire [4-1:0] node40025;
	wire [4-1:0] node40026;
	wire [4-1:0] node40027;
	wire [4-1:0] node40029;
	wire [4-1:0] node40032;
	wire [4-1:0] node40034;
	wire [4-1:0] node40037;
	wire [4-1:0] node40038;
	wire [4-1:0] node40040;
	wire [4-1:0] node40043;
	wire [4-1:0] node40045;
	wire [4-1:0] node40048;
	wire [4-1:0] node40049;
	wire [4-1:0] node40050;
	wire [4-1:0] node40051;
	wire [4-1:0] node40052;
	wire [4-1:0] node40055;
	wire [4-1:0] node40058;
	wire [4-1:0] node40059;
	wire [4-1:0] node40060;
	wire [4-1:0] node40064;
	wire [4-1:0] node40065;
	wire [4-1:0] node40068;
	wire [4-1:0] node40071;
	wire [4-1:0] node40072;
	wire [4-1:0] node40075;
	wire [4-1:0] node40078;
	wire [4-1:0] node40079;
	wire [4-1:0] node40080;
	wire [4-1:0] node40081;
	wire [4-1:0] node40082;
	wire [4-1:0] node40083;
	wire [4-1:0] node40087;
	wire [4-1:0] node40089;
	wire [4-1:0] node40092;
	wire [4-1:0] node40093;
	wire [4-1:0] node40096;
	wire [4-1:0] node40099;
	wire [4-1:0] node40100;
	wire [4-1:0] node40101;
	wire [4-1:0] node40104;
	wire [4-1:0] node40107;
	wire [4-1:0] node40108;
	wire [4-1:0] node40111;
	wire [4-1:0] node40114;
	wire [4-1:0] node40115;
	wire [4-1:0] node40116;
	wire [4-1:0] node40117;
	wire [4-1:0] node40118;
	wire [4-1:0] node40121;
	wire [4-1:0] node40124;
	wire [4-1:0] node40125;
	wire [4-1:0] node40128;
	wire [4-1:0] node40131;
	wire [4-1:0] node40132;
	wire [4-1:0] node40133;
	wire [4-1:0] node40136;
	wire [4-1:0] node40140;
	wire [4-1:0] node40142;
	wire [4-1:0] node40143;
	wire [4-1:0] node40145;
	wire [4-1:0] node40148;
	wire [4-1:0] node40150;
	wire [4-1:0] node40153;
	wire [4-1:0] node40154;
	wire [4-1:0] node40155;
	wire [4-1:0] node40156;
	wire [4-1:0] node40157;
	wire [4-1:0] node40158;
	wire [4-1:0] node40162;
	wire [4-1:0] node40163;
	wire [4-1:0] node40167;
	wire [4-1:0] node40168;
	wire [4-1:0] node40169;
	wire [4-1:0] node40173;
	wire [4-1:0] node40174;
	wire [4-1:0] node40178;
	wire [4-1:0] node40179;
	wire [4-1:0] node40180;
	wire [4-1:0] node40181;
	wire [4-1:0] node40183;
	wire [4-1:0] node40184;
	wire [4-1:0] node40188;
	wire [4-1:0] node40189;
	wire [4-1:0] node40190;
	wire [4-1:0] node40194;
	wire [4-1:0] node40197;
	wire [4-1:0] node40198;
	wire [4-1:0] node40199;
	wire [4-1:0] node40200;
	wire [4-1:0] node40204;
	wire [4-1:0] node40205;
	wire [4-1:0] node40208;
	wire [4-1:0] node40211;
	wire [4-1:0] node40213;
	wire [4-1:0] node40214;
	wire [4-1:0] node40217;
	wire [4-1:0] node40220;
	wire [4-1:0] node40221;
	wire [4-1:0] node40222;
	wire [4-1:0] node40225;
	wire [4-1:0] node40226;
	wire [4-1:0] node40230;
	wire [4-1:0] node40231;
	wire [4-1:0] node40232;
	wire [4-1:0] node40236;
	wire [4-1:0] node40237;
	wire [4-1:0] node40241;
	wire [4-1:0] node40242;
	wire [4-1:0] node40243;
	wire [4-1:0] node40244;
	wire [4-1:0] node40245;
	wire [4-1:0] node40247;
	wire [4-1:0] node40249;
	wire [4-1:0] node40252;
	wire [4-1:0] node40253;
	wire [4-1:0] node40254;
	wire [4-1:0] node40257;
	wire [4-1:0] node40261;
	wire [4-1:0] node40262;
	wire [4-1:0] node40263;
	wire [4-1:0] node40267;
	wire [4-1:0] node40268;
	wire [4-1:0] node40271;
	wire [4-1:0] node40274;
	wire [4-1:0] node40275;
	wire [4-1:0] node40276;
	wire [4-1:0] node40277;
	wire [4-1:0] node40278;
	wire [4-1:0] node40282;
	wire [4-1:0] node40283;
	wire [4-1:0] node40287;
	wire [4-1:0] node40288;
	wire [4-1:0] node40289;
	wire [4-1:0] node40293;
	wire [4-1:0] node40294;
	wire [4-1:0] node40298;
	wire [4-1:0] node40299;
	wire [4-1:0] node40300;
	wire [4-1:0] node40301;
	wire [4-1:0] node40304;
	wire [4-1:0] node40308;
	wire [4-1:0] node40309;
	wire [4-1:0] node40312;
	wire [4-1:0] node40315;
	wire [4-1:0] node40316;
	wire [4-1:0] node40317;
	wire [4-1:0] node40318;
	wire [4-1:0] node40319;
	wire [4-1:0] node40320;
	wire [4-1:0] node40324;
	wire [4-1:0] node40325;
	wire [4-1:0] node40329;
	wire [4-1:0] node40331;
	wire [4-1:0] node40332;
	wire [4-1:0] node40336;
	wire [4-1:0] node40337;
	wire [4-1:0] node40338;
	wire [4-1:0] node40340;
	wire [4-1:0] node40343;
	wire [4-1:0] node40344;
	wire [4-1:0] node40347;
	wire [4-1:0] node40351;
	wire [4-1:0] node40352;
	wire [4-1:0] node40353;
	wire [4-1:0] node40354;
	wire [4-1:0] node40355;
	wire [4-1:0] node40359;
	wire [4-1:0] node40360;
	wire [4-1:0] node40364;
	wire [4-1:0] node40365;
	wire [4-1:0] node40366;
	wire [4-1:0] node40370;
	wire [4-1:0] node40373;
	wire [4-1:0] node40374;
	wire [4-1:0] node40376;
	wire [4-1:0] node40377;
	wire [4-1:0] node40380;
	wire [4-1:0] node40383;
	wire [4-1:0] node40384;
	wire [4-1:0] node40387;
	wire [4-1:0] node40390;
	wire [4-1:0] node40391;
	wire [4-1:0] node40392;
	wire [4-1:0] node40393;
	wire [4-1:0] node40394;
	wire [4-1:0] node40395;
	wire [4-1:0] node40397;
	wire [4-1:0] node40398;
	wire [4-1:0] node40402;
	wire [4-1:0] node40404;
	wire [4-1:0] node40405;
	wire [4-1:0] node40409;
	wire [4-1:0] node40410;
	wire [4-1:0] node40411;
	wire [4-1:0] node40412;
	wire [4-1:0] node40416;
	wire [4-1:0] node40418;
	wire [4-1:0] node40421;
	wire [4-1:0] node40422;
	wire [4-1:0] node40424;
	wire [4-1:0] node40425;
	wire [4-1:0] node40428;
	wire [4-1:0] node40431;
	wire [4-1:0] node40433;
	wire [4-1:0] node40434;
	wire [4-1:0] node40438;
	wire [4-1:0] node40439;
	wire [4-1:0] node40440;
	wire [4-1:0] node40441;
	wire [4-1:0] node40442;
	wire [4-1:0] node40443;
	wire [4-1:0] node40447;
	wire [4-1:0] node40448;
	wire [4-1:0] node40452;
	wire [4-1:0] node40453;
	wire [4-1:0] node40454;
	wire [4-1:0] node40457;
	wire [4-1:0] node40461;
	wire [4-1:0] node40462;
	wire [4-1:0] node40463;
	wire [4-1:0] node40464;
	wire [4-1:0] node40468;
	wire [4-1:0] node40472;
	wire [4-1:0] node40473;
	wire [4-1:0] node40474;
	wire [4-1:0] node40476;
	wire [4-1:0] node40477;
	wire [4-1:0] node40480;
	wire [4-1:0] node40483;
	wire [4-1:0] node40484;
	wire [4-1:0] node40487;
	wire [4-1:0] node40490;
	wire [4-1:0] node40491;
	wire [4-1:0] node40493;
	wire [4-1:0] node40494;
	wire [4-1:0] node40497;
	wire [4-1:0] node40500;
	wire [4-1:0] node40501;
	wire [4-1:0] node40502;
	wire [4-1:0] node40506;
	wire [4-1:0] node40507;
	wire [4-1:0] node40510;
	wire [4-1:0] node40513;
	wire [4-1:0] node40514;
	wire [4-1:0] node40515;
	wire [4-1:0] node40516;
	wire [4-1:0] node40517;
	wire [4-1:0] node40518;
	wire [4-1:0] node40522;
	wire [4-1:0] node40523;
	wire [4-1:0] node40525;
	wire [4-1:0] node40528;
	wire [4-1:0] node40530;
	wire [4-1:0] node40534;
	wire [4-1:0] node40535;
	wire [4-1:0] node40539;
	wire [4-1:0] node40540;
	wire [4-1:0] node40541;
	wire [4-1:0] node40542;
	wire [4-1:0] node40545;
	wire [4-1:0] node40549;
	wire [4-1:0] node40550;
	wire [4-1:0] node40554;
	wire [4-1:0] node40555;
	wire [4-1:0] node40556;
	wire [4-1:0] node40557;
	wire [4-1:0] node40559;
	wire [4-1:0] node40562;
	wire [4-1:0] node40565;
	wire [4-1:0] node40566;
	wire [4-1:0] node40567;
	wire [4-1:0] node40571;
	wire [4-1:0] node40574;
	wire [4-1:0] node40575;
	wire [4-1:0] node40576;
	wire [4-1:0] node40577;
	wire [4-1:0] node40582;
	wire [4-1:0] node40583;
	wire [4-1:0] node40584;
	wire [4-1:0] node40589;
	wire [4-1:0] node40590;
	wire [4-1:0] node40591;
	wire [4-1:0] node40592;
	wire [4-1:0] node40593;
	wire [4-1:0] node40594;
	wire [4-1:0] node40595;
	wire [4-1:0] node40596;
	wire [4-1:0] node40597;
	wire [4-1:0] node40600;
	wire [4-1:0] node40603;
	wire [4-1:0] node40604;
	wire [4-1:0] node40607;
	wire [4-1:0] node40610;
	wire [4-1:0] node40611;
	wire [4-1:0] node40612;
	wire [4-1:0] node40615;
	wire [4-1:0] node40619;
	wire [4-1:0] node40620;
	wire [4-1:0] node40621;
	wire [4-1:0] node40622;
	wire [4-1:0] node40625;
	wire [4-1:0] node40628;
	wire [4-1:0] node40629;
	wire [4-1:0] node40632;
	wire [4-1:0] node40635;
	wire [4-1:0] node40636;
	wire [4-1:0] node40637;
	wire [4-1:0] node40640;
	wire [4-1:0] node40643;
	wire [4-1:0] node40645;
	wire [4-1:0] node40646;
	wire [4-1:0] node40650;
	wire [4-1:0] node40651;
	wire [4-1:0] node40652;
	wire [4-1:0] node40653;
	wire [4-1:0] node40657;
	wire [4-1:0] node40658;
	wire [4-1:0] node40659;
	wire [4-1:0] node40662;
	wire [4-1:0] node40665;
	wire [4-1:0] node40666;
	wire [4-1:0] node40667;
	wire [4-1:0] node40671;
	wire [4-1:0] node40672;
	wire [4-1:0] node40675;
	wire [4-1:0] node40678;
	wire [4-1:0] node40679;
	wire [4-1:0] node40680;
	wire [4-1:0] node40683;
	wire [4-1:0] node40686;
	wire [4-1:0] node40687;
	wire [4-1:0] node40690;
	wire [4-1:0] node40693;
	wire [4-1:0] node40694;
	wire [4-1:0] node40695;
	wire [4-1:0] node40696;
	wire [4-1:0] node40697;
	wire [4-1:0] node40698;
	wire [4-1:0] node40701;
	wire [4-1:0] node40704;
	wire [4-1:0] node40705;
	wire [4-1:0] node40708;
	wire [4-1:0] node40711;
	wire [4-1:0] node40712;
	wire [4-1:0] node40713;
	wire [4-1:0] node40717;
	wire [4-1:0] node40718;
	wire [4-1:0] node40721;
	wire [4-1:0] node40722;
	wire [4-1:0] node40726;
	wire [4-1:0] node40727;
	wire [4-1:0] node40728;
	wire [4-1:0] node40732;
	wire [4-1:0] node40733;
	wire [4-1:0] node40734;
	wire [4-1:0] node40738;
	wire [4-1:0] node40739;
	wire [4-1:0] node40743;
	wire [4-1:0] node40744;
	wire [4-1:0] node40745;
	wire [4-1:0] node40746;
	wire [4-1:0] node40749;
	wire [4-1:0] node40750;
	wire [4-1:0] node40751;
	wire [4-1:0] node40755;
	wire [4-1:0] node40756;
	wire [4-1:0] node40760;
	wire [4-1:0] node40762;
	wire [4-1:0] node40763;
	wire [4-1:0] node40766;
	wire [4-1:0] node40769;
	wire [4-1:0] node40770;
	wire [4-1:0] node40771;
	wire [4-1:0] node40772;
	wire [4-1:0] node40776;
	wire [4-1:0] node40777;
	wire [4-1:0] node40781;
	wire [4-1:0] node40782;
	wire [4-1:0] node40783;
	wire [4-1:0] node40787;
	wire [4-1:0] node40788;
	wire [4-1:0] node40792;
	wire [4-1:0] node40793;
	wire [4-1:0] node40794;
	wire [4-1:0] node40795;
	wire [4-1:0] node40796;
	wire [4-1:0] node40798;
	wire [4-1:0] node40801;
	wire [4-1:0] node40803;
	wire [4-1:0] node40806;
	wire [4-1:0] node40807;
	wire [4-1:0] node40809;
	wire [4-1:0] node40812;
	wire [4-1:0] node40814;
	wire [4-1:0] node40817;
	wire [4-1:0] node40818;
	wire [4-1:0] node40819;
	wire [4-1:0] node40820;
	wire [4-1:0] node40824;
	wire [4-1:0] node40825;
	wire [4-1:0] node40829;
	wire [4-1:0] node40830;
	wire [4-1:0] node40831;
	wire [4-1:0] node40835;
	wire [4-1:0] node40836;
	wire [4-1:0] node40840;
	wire [4-1:0] node40841;
	wire [4-1:0] node40842;
	wire [4-1:0] node40843;
	wire [4-1:0] node40844;
	wire [4-1:0] node40845;
	wire [4-1:0] node40848;
	wire [4-1:0] node40851;
	wire [4-1:0] node40852;
	wire [4-1:0] node40855;
	wire [4-1:0] node40858;
	wire [4-1:0] node40859;
	wire [4-1:0] node40860;
	wire [4-1:0] node40863;
	wire [4-1:0] node40866;
	wire [4-1:0] node40867;
	wire [4-1:0] node40868;
	wire [4-1:0] node40871;
	wire [4-1:0] node40874;
	wire [4-1:0] node40875;
	wire [4-1:0] node40878;
	wire [4-1:0] node40881;
	wire [4-1:0] node40882;
	wire [4-1:0] node40885;
	wire [4-1:0] node40888;
	wire [4-1:0] node40889;
	wire [4-1:0] node40890;
	wire [4-1:0] node40891;
	wire [4-1:0] node40895;
	wire [4-1:0] node40896;
	wire [4-1:0] node40900;
	wire [4-1:0] node40901;
	wire [4-1:0] node40902;
	wire [4-1:0] node40906;
	wire [4-1:0] node40907;
	wire [4-1:0] node40911;
	wire [4-1:0] node40912;
	wire [4-1:0] node40913;
	wire [4-1:0] node40914;
	wire [4-1:0] node40915;
	wire [4-1:0] node40919;
	wire [4-1:0] node40920;
	wire [4-1:0] node40925;
	wire [4-1:0] node40926;
	wire [4-1:0] node40927;
	wire [4-1:0] node40928;
	wire [4-1:0] node40932;
	wire [4-1:0] node40933;
	wire [4-1:0] node40938;
	wire [4-1:0] node40939;
	wire [4-1:0] node40940;
	wire [4-1:0] node40941;
	wire [4-1:0] node40942;
	wire [4-1:0] node40943;
	wire [4-1:0] node40944;
	wire [4-1:0] node40945;
	wire [4-1:0] node40946;
	wire [4-1:0] node40947;
	wire [4-1:0] node40948;
	wire [4-1:0] node40949;
	wire [4-1:0] node40950;
	wire [4-1:0] node40954;
	wire [4-1:0] node40955;
	wire [4-1:0] node40958;
	wire [4-1:0] node40961;
	wire [4-1:0] node40962;
	wire [4-1:0] node40963;
	wire [4-1:0] node40964;
	wire [4-1:0] node40967;
	wire [4-1:0] node40970;
	wire [4-1:0] node40971;
	wire [4-1:0] node40974;
	wire [4-1:0] node40977;
	wire [4-1:0] node40979;
	wire [4-1:0] node40980;
	wire [4-1:0] node40983;
	wire [4-1:0] node40986;
	wire [4-1:0] node40987;
	wire [4-1:0] node40988;
	wire [4-1:0] node40991;
	wire [4-1:0] node40994;
	wire [4-1:0] node40995;
	wire [4-1:0] node40996;
	wire [4-1:0] node40997;
	wire [4-1:0] node41000;
	wire [4-1:0] node41004;
	wire [4-1:0] node41005;
	wire [4-1:0] node41006;
	wire [4-1:0] node41010;
	wire [4-1:0] node41011;
	wire [4-1:0] node41014;
	wire [4-1:0] node41017;
	wire [4-1:0] node41018;
	wire [4-1:0] node41019;
	wire [4-1:0] node41021;
	wire [4-1:0] node41024;
	wire [4-1:0] node41026;
	wire [4-1:0] node41029;
	wire [4-1:0] node41030;
	wire [4-1:0] node41032;
	wire [4-1:0] node41035;
	wire [4-1:0] node41037;
	wire [4-1:0] node41040;
	wire [4-1:0] node41041;
	wire [4-1:0] node41042;
	wire [4-1:0] node41043;
	wire [4-1:0] node41044;
	wire [4-1:0] node41045;
	wire [4-1:0] node41046;
	wire [4-1:0] node41049;
	wire [4-1:0] node41052;
	wire [4-1:0] node41054;
	wire [4-1:0] node41057;
	wire [4-1:0] node41058;
	wire [4-1:0] node41061;
	wire [4-1:0] node41064;
	wire [4-1:0] node41065;
	wire [4-1:0] node41066;
	wire [4-1:0] node41070;
	wire [4-1:0] node41071;
	wire [4-1:0] node41074;
	wire [4-1:0] node41077;
	wire [4-1:0] node41078;
	wire [4-1:0] node41079;
	wire [4-1:0] node41082;
	wire [4-1:0] node41085;
	wire [4-1:0] node41087;
	wire [4-1:0] node41088;
	wire [4-1:0] node41091;
	wire [4-1:0] node41094;
	wire [4-1:0] node41095;
	wire [4-1:0] node41096;
	wire [4-1:0] node41097;
	wire [4-1:0] node41100;
	wire [4-1:0] node41101;
	wire [4-1:0] node41102;
	wire [4-1:0] node41106;
	wire [4-1:0] node41107;
	wire [4-1:0] node41111;
	wire [4-1:0] node41112;
	wire [4-1:0] node41113;
	wire [4-1:0] node41114;
	wire [4-1:0] node41117;
	wire [4-1:0] node41120;
	wire [4-1:0] node41121;
	wire [4-1:0] node41124;
	wire [4-1:0] node41127;
	wire [4-1:0] node41128;
	wire [4-1:0] node41131;
	wire [4-1:0] node41134;
	wire [4-1:0] node41135;
	wire [4-1:0] node41136;
	wire [4-1:0] node41137;
	wire [4-1:0] node41140;
	wire [4-1:0] node41143;
	wire [4-1:0] node41144;
	wire [4-1:0] node41147;
	wire [4-1:0] node41150;
	wire [4-1:0] node41151;
	wire [4-1:0] node41154;
	wire [4-1:0] node41157;
	wire [4-1:0] node41158;
	wire [4-1:0] node41159;
	wire [4-1:0] node41160;
	wire [4-1:0] node41161;
	wire [4-1:0] node41162;
	wire [4-1:0] node41165;
	wire [4-1:0] node41168;
	wire [4-1:0] node41169;
	wire [4-1:0] node41172;
	wire [4-1:0] node41175;
	wire [4-1:0] node41176;
	wire [4-1:0] node41177;
	wire [4-1:0] node41178;
	wire [4-1:0] node41181;
	wire [4-1:0] node41184;
	wire [4-1:0] node41185;
	wire [4-1:0] node41188;
	wire [4-1:0] node41191;
	wire [4-1:0] node41192;
	wire [4-1:0] node41195;
	wire [4-1:0] node41198;
	wire [4-1:0] node41199;
	wire [4-1:0] node41200;
	wire [4-1:0] node41201;
	wire [4-1:0] node41204;
	wire [4-1:0] node41206;
	wire [4-1:0] node41209;
	wire [4-1:0] node41210;
	wire [4-1:0] node41212;
	wire [4-1:0] node41215;
	wire [4-1:0] node41217;
	wire [4-1:0] node41220;
	wire [4-1:0] node41221;
	wire [4-1:0] node41222;
	wire [4-1:0] node41225;
	wire [4-1:0] node41228;
	wire [4-1:0] node41229;
	wire [4-1:0] node41230;
	wire [4-1:0] node41232;
	wire [4-1:0] node41235;
	wire [4-1:0] node41238;
	wire [4-1:0] node41239;
	wire [4-1:0] node41240;
	wire [4-1:0] node41243;
	wire [4-1:0] node41246;
	wire [4-1:0] node41248;
	wire [4-1:0] node41251;
	wire [4-1:0] node41252;
	wire [4-1:0] node41253;
	wire [4-1:0] node41254;
	wire [4-1:0] node41257;
	wire [4-1:0] node41260;
	wire [4-1:0] node41261;
	wire [4-1:0] node41262;
	wire [4-1:0] node41264;
	wire [4-1:0] node41265;
	wire [4-1:0] node41270;
	wire [4-1:0] node41271;
	wire [4-1:0] node41273;
	wire [4-1:0] node41274;
	wire [4-1:0] node41277;
	wire [4-1:0] node41280;
	wire [4-1:0] node41281;
	wire [4-1:0] node41282;
	wire [4-1:0] node41285;
	wire [4-1:0] node41288;
	wire [4-1:0] node41290;
	wire [4-1:0] node41293;
	wire [4-1:0] node41294;
	wire [4-1:0] node41295;
	wire [4-1:0] node41297;
	wire [4-1:0] node41300;
	wire [4-1:0] node41302;
	wire [4-1:0] node41305;
	wire [4-1:0] node41306;
	wire [4-1:0] node41308;
	wire [4-1:0] node41311;
	wire [4-1:0] node41313;
	wire [4-1:0] node41316;
	wire [4-1:0] node41317;
	wire [4-1:0] node41318;
	wire [4-1:0] node41319;
	wire [4-1:0] node41320;
	wire [4-1:0] node41321;
	wire [4-1:0] node41322;
	wire [4-1:0] node41323;
	wire [4-1:0] node41324;
	wire [4-1:0] node41328;
	wire [4-1:0] node41330;
	wire [4-1:0] node41333;
	wire [4-1:0] node41334;
	wire [4-1:0] node41337;
	wire [4-1:0] node41340;
	wire [4-1:0] node41341;
	wire [4-1:0] node41342;
	wire [4-1:0] node41345;
	wire [4-1:0] node41348;
	wire [4-1:0] node41349;
	wire [4-1:0] node41352;
	wire [4-1:0] node41355;
	wire [4-1:0] node41356;
	wire [4-1:0] node41357;
	wire [4-1:0] node41358;
	wire [4-1:0] node41361;
	wire [4-1:0] node41364;
	wire [4-1:0] node41366;
	wire [4-1:0] node41369;
	wire [4-1:0] node41370;
	wire [4-1:0] node41371;
	wire [4-1:0] node41374;
	wire [4-1:0] node41377;
	wire [4-1:0] node41378;
	wire [4-1:0] node41382;
	wire [4-1:0] node41383;
	wire [4-1:0] node41384;
	wire [4-1:0] node41385;
	wire [4-1:0] node41386;
	wire [4-1:0] node41388;
	wire [4-1:0] node41391;
	wire [4-1:0] node41393;
	wire [4-1:0] node41396;
	wire [4-1:0] node41397;
	wire [4-1:0] node41399;
	wire [4-1:0] node41402;
	wire [4-1:0] node41403;
	wire [4-1:0] node41407;
	wire [4-1:0] node41408;
	wire [4-1:0] node41409;
	wire [4-1:0] node41410;
	wire [4-1:0] node41413;
	wire [4-1:0] node41416;
	wire [4-1:0] node41417;
	wire [4-1:0] node41420;
	wire [4-1:0] node41423;
	wire [4-1:0] node41425;
	wire [4-1:0] node41428;
	wire [4-1:0] node41429;
	wire [4-1:0] node41430;
	wire [4-1:0] node41431;
	wire [4-1:0] node41432;
	wire [4-1:0] node41435;
	wire [4-1:0] node41438;
	wire [4-1:0] node41439;
	wire [4-1:0] node41443;
	wire [4-1:0] node41444;
	wire [4-1:0] node41446;
	wire [4-1:0] node41450;
	wire [4-1:0] node41451;
	wire [4-1:0] node41452;
	wire [4-1:0] node41454;
	wire [4-1:0] node41457;
	wire [4-1:0] node41458;
	wire [4-1:0] node41461;
	wire [4-1:0] node41464;
	wire [4-1:0] node41465;
	wire [4-1:0] node41468;
	wire [4-1:0] node41471;
	wire [4-1:0] node41472;
	wire [4-1:0] node41473;
	wire [4-1:0] node41474;
	wire [4-1:0] node41477;
	wire [4-1:0] node41480;
	wire [4-1:0] node41481;
	wire [4-1:0] node41482;
	wire [4-1:0] node41485;
	wire [4-1:0] node41488;
	wire [4-1:0] node41489;
	wire [4-1:0] node41490;
	wire [4-1:0] node41491;
	wire [4-1:0] node41494;
	wire [4-1:0] node41498;
	wire [4-1:0] node41499;
	wire [4-1:0] node41500;
	wire [4-1:0] node41503;
	wire [4-1:0] node41506;
	wire [4-1:0] node41507;
	wire [4-1:0] node41511;
	wire [4-1:0] node41512;
	wire [4-1:0] node41513;
	wire [4-1:0] node41514;
	wire [4-1:0] node41517;
	wire [4-1:0] node41520;
	wire [4-1:0] node41521;
	wire [4-1:0] node41523;
	wire [4-1:0] node41524;
	wire [4-1:0] node41528;
	wire [4-1:0] node41529;
	wire [4-1:0] node41532;
	wire [4-1:0] node41535;
	wire [4-1:0] node41536;
	wire [4-1:0] node41537;
	wire [4-1:0] node41538;
	wire [4-1:0] node41541;
	wire [4-1:0] node41544;
	wire [4-1:0] node41545;
	wire [4-1:0] node41548;
	wire [4-1:0] node41551;
	wire [4-1:0] node41552;
	wire [4-1:0] node41555;
	wire [4-1:0] node41558;
	wire [4-1:0] node41559;
	wire [4-1:0] node41560;
	wire [4-1:0] node41561;
	wire [4-1:0] node41562;
	wire [4-1:0] node41563;
	wire [4-1:0] node41566;
	wire [4-1:0] node41569;
	wire [4-1:0] node41570;
	wire [4-1:0] node41571;
	wire [4-1:0] node41572;
	wire [4-1:0] node41575;
	wire [4-1:0] node41578;
	wire [4-1:0] node41579;
	wire [4-1:0] node41582;
	wire [4-1:0] node41585;
	wire [4-1:0] node41586;
	wire [4-1:0] node41589;
	wire [4-1:0] node41592;
	wire [4-1:0] node41593;
	wire [4-1:0] node41594;
	wire [4-1:0] node41596;
	wire [4-1:0] node41600;
	wire [4-1:0] node41601;
	wire [4-1:0] node41604;
	wire [4-1:0] node41607;
	wire [4-1:0] node41608;
	wire [4-1:0] node41609;
	wire [4-1:0] node41612;
	wire [4-1:0] node41615;
	wire [4-1:0] node41616;
	wire [4-1:0] node41617;
	wire [4-1:0] node41618;
	wire [4-1:0] node41621;
	wire [4-1:0] node41624;
	wire [4-1:0] node41625;
	wire [4-1:0] node41626;
	wire [4-1:0] node41629;
	wire [4-1:0] node41632;
	wire [4-1:0] node41633;
	wire [4-1:0] node41637;
	wire [4-1:0] node41638;
	wire [4-1:0] node41639;
	wire [4-1:0] node41642;
	wire [4-1:0] node41645;
	wire [4-1:0] node41646;
	wire [4-1:0] node41649;
	wire [4-1:0] node41652;
	wire [4-1:0] node41653;
	wire [4-1:0] node41654;
	wire [4-1:0] node41655;
	wire [4-1:0] node41656;
	wire [4-1:0] node41660;
	wire [4-1:0] node41661;
	wire [4-1:0] node41665;
	wire [4-1:0] node41666;
	wire [4-1:0] node41667;
	wire [4-1:0] node41671;
	wire [4-1:0] node41672;
	wire [4-1:0] node41676;
	wire [4-1:0] node41677;
	wire [4-1:0] node41678;
	wire [4-1:0] node41679;
	wire [4-1:0] node41681;
	wire [4-1:0] node41684;
	wire [4-1:0] node41685;
	wire [4-1:0] node41686;
	wire [4-1:0] node41689;
	wire [4-1:0] node41692;
	wire [4-1:0] node41694;
	wire [4-1:0] node41697;
	wire [4-1:0] node41698;
	wire [4-1:0] node41699;
	wire [4-1:0] node41701;
	wire [4-1:0] node41704;
	wire [4-1:0] node41705;
	wire [4-1:0] node41708;
	wire [4-1:0] node41711;
	wire [4-1:0] node41712;
	wire [4-1:0] node41714;
	wire [4-1:0] node41717;
	wire [4-1:0] node41718;
	wire [4-1:0] node41721;
	wire [4-1:0] node41724;
	wire [4-1:0] node41725;
	wire [4-1:0] node41726;
	wire [4-1:0] node41729;
	wire [4-1:0] node41732;
	wire [4-1:0] node41733;
	wire [4-1:0] node41734;
	wire [4-1:0] node41736;
	wire [4-1:0] node41740;
	wire [4-1:0] node41741;
	wire [4-1:0] node41742;
	wire [4-1:0] node41746;
	wire [4-1:0] node41747;
	wire [4-1:0] node41751;
	wire [4-1:0] node41752;
	wire [4-1:0] node41753;
	wire [4-1:0] node41754;
	wire [4-1:0] node41755;
	wire [4-1:0] node41756;
	wire [4-1:0] node41757;
	wire [4-1:0] node41761;
	wire [4-1:0] node41762;
	wire [4-1:0] node41766;
	wire [4-1:0] node41767;
	wire [4-1:0] node41768;
	wire [4-1:0] node41770;
	wire [4-1:0] node41773;
	wire [4-1:0] node41775;
	wire [4-1:0] node41778;
	wire [4-1:0] node41779;
	wire [4-1:0] node41781;
	wire [4-1:0] node41784;
	wire [4-1:0] node41786;
	wire [4-1:0] node41789;
	wire [4-1:0] node41790;
	wire [4-1:0] node41791;
	wire [4-1:0] node41794;
	wire [4-1:0] node41795;
	wire [4-1:0] node41796;
	wire [4-1:0] node41799;
	wire [4-1:0] node41802;
	wire [4-1:0] node41805;
	wire [4-1:0] node41806;
	wire [4-1:0] node41807;
	wire [4-1:0] node41810;
	wire [4-1:0] node41811;
	wire [4-1:0] node41814;
	wire [4-1:0] node41817;
	wire [4-1:0] node41818;
	wire [4-1:0] node41821;
	wire [4-1:0] node41822;
	wire [4-1:0] node41825;
	wire [4-1:0] node41828;
	wire [4-1:0] node41829;
	wire [4-1:0] node41830;
	wire [4-1:0] node41831;
	wire [4-1:0] node41832;
	wire [4-1:0] node41835;
	wire [4-1:0] node41836;
	wire [4-1:0] node41839;
	wire [4-1:0] node41842;
	wire [4-1:0] node41843;
	wire [4-1:0] node41846;
	wire [4-1:0] node41847;
	wire [4-1:0] node41851;
	wire [4-1:0] node41852;
	wire [4-1:0] node41855;
	wire [4-1:0] node41856;
	wire [4-1:0] node41857;
	wire [4-1:0] node41858;
	wire [4-1:0] node41862;
	wire [4-1:0] node41863;
	wire [4-1:0] node41864;
	wire [4-1:0] node41867;
	wire [4-1:0] node41870;
	wire [4-1:0] node41871;
	wire [4-1:0] node41875;
	wire [4-1:0] node41878;
	wire [4-1:0] node41879;
	wire [4-1:0] node41880;
	wire [4-1:0] node41882;
	wire [4-1:0] node41883;
	wire [4-1:0] node41884;
	wire [4-1:0] node41886;
	wire [4-1:0] node41890;
	wire [4-1:0] node41892;
	wire [4-1:0] node41894;
	wire [4-1:0] node41897;
	wire [4-1:0] node41899;
	wire [4-1:0] node41902;
	wire [4-1:0] node41903;
	wire [4-1:0] node41904;
	wire [4-1:0] node41907;
	wire [4-1:0] node41908;
	wire [4-1:0] node41911;
	wire [4-1:0] node41914;
	wire [4-1:0] node41915;
	wire [4-1:0] node41918;
	wire [4-1:0] node41919;
	wire [4-1:0] node41922;
	wire [4-1:0] node41925;
	wire [4-1:0] node41926;
	wire [4-1:0] node41927;
	wire [4-1:0] node41928;
	wire [4-1:0] node41929;
	wire [4-1:0] node41930;
	wire [4-1:0] node41931;
	wire [4-1:0] node41932;
	wire [4-1:0] node41937;
	wire [4-1:0] node41938;
	wire [4-1:0] node41939;
	wire [4-1:0] node41940;
	wire [4-1:0] node41945;
	wire [4-1:0] node41946;
	wire [4-1:0] node41948;
	wire [4-1:0] node41952;
	wire [4-1:0] node41953;
	wire [4-1:0] node41954;
	wire [4-1:0] node41955;
	wire [4-1:0] node41957;
	wire [4-1:0] node41960;
	wire [4-1:0] node41963;
	wire [4-1:0] node41964;
	wire [4-1:0] node41965;
	wire [4-1:0] node41968;
	wire [4-1:0] node41972;
	wire [4-1:0] node41973;
	wire [4-1:0] node41975;
	wire [4-1:0] node41978;
	wire [4-1:0] node41980;
	wire [4-1:0] node41982;
	wire [4-1:0] node41985;
	wire [4-1:0] node41986;
	wire [4-1:0] node41987;
	wire [4-1:0] node41988;
	wire [4-1:0] node41990;
	wire [4-1:0] node41994;
	wire [4-1:0] node41995;
	wire [4-1:0] node41996;
	wire [4-1:0] node42000;
	wire [4-1:0] node42001;
	wire [4-1:0] node42005;
	wire [4-1:0] node42006;
	wire [4-1:0] node42007;
	wire [4-1:0] node42008;
	wire [4-1:0] node42009;
	wire [4-1:0] node42012;
	wire [4-1:0] node42016;
	wire [4-1:0] node42017;
	wire [4-1:0] node42018;
	wire [4-1:0] node42021;
	wire [4-1:0] node42024;
	wire [4-1:0] node42025;
	wire [4-1:0] node42028;
	wire [4-1:0] node42031;
	wire [4-1:0] node42032;
	wire [4-1:0] node42035;
	wire [4-1:0] node42038;
	wire [4-1:0] node42039;
	wire [4-1:0] node42040;
	wire [4-1:0] node42041;
	wire [4-1:0] node42042;
	wire [4-1:0] node42043;
	wire [4-1:0] node42045;
	wire [4-1:0] node42049;
	wire [4-1:0] node42052;
	wire [4-1:0] node42053;
	wire [4-1:0] node42054;
	wire [4-1:0] node42055;
	wire [4-1:0] node42060;
	wire [4-1:0] node42061;
	wire [4-1:0] node42064;
	wire [4-1:0] node42067;
	wire [4-1:0] node42068;
	wire [4-1:0] node42069;
	wire [4-1:0] node42070;
	wire [4-1:0] node42071;
	wire [4-1:0] node42075;
	wire [4-1:0] node42076;
	wire [4-1:0] node42080;
	wire [4-1:0] node42082;
	wire [4-1:0] node42085;
	wire [4-1:0] node42086;
	wire [4-1:0] node42088;
	wire [4-1:0] node42091;
	wire [4-1:0] node42093;
	wire [4-1:0] node42096;
	wire [4-1:0] node42097;
	wire [4-1:0] node42098;
	wire [4-1:0] node42099;
	wire [4-1:0] node42101;
	wire [4-1:0] node42104;
	wire [4-1:0] node42106;
	wire [4-1:0] node42107;
	wire [4-1:0] node42110;
	wire [4-1:0] node42113;
	wire [4-1:0] node42114;
	wire [4-1:0] node42115;
	wire [4-1:0] node42116;
	wire [4-1:0] node42119;
	wire [4-1:0] node42122;
	wire [4-1:0] node42123;
	wire [4-1:0] node42127;
	wire [4-1:0] node42128;
	wire [4-1:0] node42129;
	wire [4-1:0] node42132;
	wire [4-1:0] node42135;
	wire [4-1:0] node42136;
	wire [4-1:0] node42139;
	wire [4-1:0] node42142;
	wire [4-1:0] node42143;
	wire [4-1:0] node42144;
	wire [4-1:0] node42146;
	wire [4-1:0] node42147;
	wire [4-1:0] node42151;
	wire [4-1:0] node42152;
	wire [4-1:0] node42153;
	wire [4-1:0] node42158;
	wire [4-1:0] node42159;
	wire [4-1:0] node42160;
	wire [4-1:0] node42162;
	wire [4-1:0] node42166;
	wire [4-1:0] node42167;
	wire [4-1:0] node42170;
	wire [4-1:0] node42173;
	wire [4-1:0] node42174;
	wire [4-1:0] node42175;
	wire [4-1:0] node42176;
	wire [4-1:0] node42177;
	wire [4-1:0] node42178;
	wire [4-1:0] node42181;
	wire [4-1:0] node42184;
	wire [4-1:0] node42185;
	wire [4-1:0] node42188;
	wire [4-1:0] node42191;
	wire [4-1:0] node42192;
	wire [4-1:0] node42193;
	wire [4-1:0] node42196;
	wire [4-1:0] node42199;
	wire [4-1:0] node42200;
	wire [4-1:0] node42201;
	wire [4-1:0] node42204;
	wire [4-1:0] node42208;
	wire [4-1:0] node42209;
	wire [4-1:0] node42210;
	wire [4-1:0] node42211;
	wire [4-1:0] node42214;
	wire [4-1:0] node42217;
	wire [4-1:0] node42218;
	wire [4-1:0] node42221;
	wire [4-1:0] node42224;
	wire [4-1:0] node42225;
	wire [4-1:0] node42227;
	wire [4-1:0] node42228;
	wire [4-1:0] node42231;
	wire [4-1:0] node42234;
	wire [4-1:0] node42235;
	wire [4-1:0] node42238;
	wire [4-1:0] node42241;
	wire [4-1:0] node42242;
	wire [4-1:0] node42243;
	wire [4-1:0] node42244;
	wire [4-1:0] node42245;
	wire [4-1:0] node42249;
	wire [4-1:0] node42252;
	wire [4-1:0] node42253;
	wire [4-1:0] node42254;
	wire [4-1:0] node42258;
	wire [4-1:0] node42261;
	wire [4-1:0] node42262;
	wire [4-1:0] node42263;
	wire [4-1:0] node42264;
	wire [4-1:0] node42268;
	wire [4-1:0] node42271;
	wire [4-1:0] node42272;
	wire [4-1:0] node42273;
	wire [4-1:0] node42277;
	wire [4-1:0] node42280;
	wire [4-1:0] node42281;
	wire [4-1:0] node42282;
	wire [4-1:0] node42283;
	wire [4-1:0] node42284;
	wire [4-1:0] node42285;
	wire [4-1:0] node42286;
	wire [4-1:0] node42287;
	wire [4-1:0] node42288;
	wire [4-1:0] node42290;
	wire [4-1:0] node42291;
	wire [4-1:0] node42294;
	wire [4-1:0] node42298;
	wire [4-1:0] node42299;
	wire [4-1:0] node42301;
	wire [4-1:0] node42304;
	wire [4-1:0] node42305;
	wire [4-1:0] node42307;
	wire [4-1:0] node42311;
	wire [4-1:0] node42312;
	wire [4-1:0] node42313;
	wire [4-1:0] node42314;
	wire [4-1:0] node42317;
	wire [4-1:0] node42320;
	wire [4-1:0] node42321;
	wire [4-1:0] node42322;
	wire [4-1:0] node42325;
	wire [4-1:0] node42328;
	wire [4-1:0] node42330;
	wire [4-1:0] node42333;
	wire [4-1:0] node42334;
	wire [4-1:0] node42335;
	wire [4-1:0] node42337;
	wire [4-1:0] node42340;
	wire [4-1:0] node42341;
	wire [4-1:0] node42344;
	wire [4-1:0] node42347;
	wire [4-1:0] node42348;
	wire [4-1:0] node42349;
	wire [4-1:0] node42352;
	wire [4-1:0] node42355;
	wire [4-1:0] node42356;
	wire [4-1:0] node42359;
	wire [4-1:0] node42362;
	wire [4-1:0] node42363;
	wire [4-1:0] node42364;
	wire [4-1:0] node42365;
	wire [4-1:0] node42366;
	wire [4-1:0] node42369;
	wire [4-1:0] node42372;
	wire [4-1:0] node42374;
	wire [4-1:0] node42375;
	wire [4-1:0] node42378;
	wire [4-1:0] node42381;
	wire [4-1:0] node42382;
	wire [4-1:0] node42383;
	wire [4-1:0] node42384;
	wire [4-1:0] node42387;
	wire [4-1:0] node42390;
	wire [4-1:0] node42391;
	wire [4-1:0] node42394;
	wire [4-1:0] node42397;
	wire [4-1:0] node42398;
	wire [4-1:0] node42399;
	wire [4-1:0] node42402;
	wire [4-1:0] node42405;
	wire [4-1:0] node42406;
	wire [4-1:0] node42409;
	wire [4-1:0] node42412;
	wire [4-1:0] node42413;
	wire [4-1:0] node42414;
	wire [4-1:0] node42416;
	wire [4-1:0] node42417;
	wire [4-1:0] node42421;
	wire [4-1:0] node42423;
	wire [4-1:0] node42424;
	wire [4-1:0] node42427;
	wire [4-1:0] node42430;
	wire [4-1:0] node42431;
	wire [4-1:0] node42433;
	wire [4-1:0] node42435;
	wire [4-1:0] node42438;
	wire [4-1:0] node42440;
	wire [4-1:0] node42442;
	wire [4-1:0] node42445;
	wire [4-1:0] node42446;
	wire [4-1:0] node42447;
	wire [4-1:0] node42448;
	wire [4-1:0] node42450;
	wire [4-1:0] node42451;
	wire [4-1:0] node42455;
	wire [4-1:0] node42456;
	wire [4-1:0] node42457;
	wire [4-1:0] node42458;
	wire [4-1:0] node42461;
	wire [4-1:0] node42464;
	wire [4-1:0] node42465;
	wire [4-1:0] node42469;
	wire [4-1:0] node42471;
	wire [4-1:0] node42474;
	wire [4-1:0] node42475;
	wire [4-1:0] node42477;
	wire [4-1:0] node42479;
	wire [4-1:0] node42481;
	wire [4-1:0] node42484;
	wire [4-1:0] node42485;
	wire [4-1:0] node42486;
	wire [4-1:0] node42489;
	wire [4-1:0] node42492;
	wire [4-1:0] node42494;
	wire [4-1:0] node42497;
	wire [4-1:0] node42498;
	wire [4-1:0] node42499;
	wire [4-1:0] node42501;
	wire [4-1:0] node42503;
	wire [4-1:0] node42505;
	wire [4-1:0] node42508;
	wire [4-1:0] node42509;
	wire [4-1:0] node42510;
	wire [4-1:0] node42513;
	wire [4-1:0] node42516;
	wire [4-1:0] node42519;
	wire [4-1:0] node42520;
	wire [4-1:0] node42521;
	wire [4-1:0] node42523;
	wire [4-1:0] node42527;
	wire [4-1:0] node42528;
	wire [4-1:0] node42529;
	wire [4-1:0] node42532;
	wire [4-1:0] node42535;
	wire [4-1:0] node42537;
	wire [4-1:0] node42540;
	wire [4-1:0] node42541;
	wire [4-1:0] node42542;
	wire [4-1:0] node42543;
	wire [4-1:0] node42545;
	wire [4-1:0] node42546;
	wire [4-1:0] node42548;
	wire [4-1:0] node42549;
	wire [4-1:0] node42552;
	wire [4-1:0] node42555;
	wire [4-1:0] node42556;
	wire [4-1:0] node42559;
	wire [4-1:0] node42562;
	wire [4-1:0] node42564;
	wire [4-1:0] node42565;
	wire [4-1:0] node42568;
	wire [4-1:0] node42571;
	wire [4-1:0] node42572;
	wire [4-1:0] node42574;
	wire [4-1:0] node42575;
	wire [4-1:0] node42576;
	wire [4-1:0] node42579;
	wire [4-1:0] node42582;
	wire [4-1:0] node42583;
	wire [4-1:0] node42586;
	wire [4-1:0] node42589;
	wire [4-1:0] node42591;
	wire [4-1:0] node42592;
	wire [4-1:0] node42593;
	wire [4-1:0] node42595;
	wire [4-1:0] node42598;
	wire [4-1:0] node42599;
	wire [4-1:0] node42603;
	wire [4-1:0] node42604;
	wire [4-1:0] node42605;
	wire [4-1:0] node42609;
	wire [4-1:0] node42612;
	wire [4-1:0] node42613;
	wire [4-1:0] node42614;
	wire [4-1:0] node42615;
	wire [4-1:0] node42616;
	wire [4-1:0] node42617;
	wire [4-1:0] node42620;
	wire [4-1:0] node42623;
	wire [4-1:0] node42624;
	wire [4-1:0] node42627;
	wire [4-1:0] node42630;
	wire [4-1:0] node42631;
	wire [4-1:0] node42632;
	wire [4-1:0] node42635;
	wire [4-1:0] node42638;
	wire [4-1:0] node42639;
	wire [4-1:0] node42643;
	wire [4-1:0] node42644;
	wire [4-1:0] node42645;
	wire [4-1:0] node42647;
	wire [4-1:0] node42648;
	wire [4-1:0] node42651;
	wire [4-1:0] node42654;
	wire [4-1:0] node42655;
	wire [4-1:0] node42658;
	wire [4-1:0] node42661;
	wire [4-1:0] node42662;
	wire [4-1:0] node42664;
	wire [4-1:0] node42667;
	wire [4-1:0] node42668;
	wire [4-1:0] node42672;
	wire [4-1:0] node42673;
	wire [4-1:0] node42674;
	wire [4-1:0] node42675;
	wire [4-1:0] node42676;
	wire [4-1:0] node42677;
	wire [4-1:0] node42681;
	wire [4-1:0] node42682;
	wire [4-1:0] node42686;
	wire [4-1:0] node42687;
	wire [4-1:0] node42690;
	wire [4-1:0] node42691;
	wire [4-1:0] node42695;
	wire [4-1:0] node42696;
	wire [4-1:0] node42697;
	wire [4-1:0] node42700;
	wire [4-1:0] node42703;
	wire [4-1:0] node42704;
	wire [4-1:0] node42705;
	wire [4-1:0] node42709;
	wire [4-1:0] node42712;
	wire [4-1:0] node42713;
	wire [4-1:0] node42714;
	wire [4-1:0] node42716;
	wire [4-1:0] node42719;
	wire [4-1:0] node42720;
	wire [4-1:0] node42721;
	wire [4-1:0] node42724;
	wire [4-1:0] node42727;
	wire [4-1:0] node42729;
	wire [4-1:0] node42732;
	wire [4-1:0] node42733;
	wire [4-1:0] node42734;
	wire [4-1:0] node42737;
	wire [4-1:0] node42740;
	wire [4-1:0] node42741;
	wire [4-1:0] node42744;
	wire [4-1:0] node42746;
	wire [4-1:0] node42749;
	wire [4-1:0] node42750;
	wire [4-1:0] node42751;
	wire [4-1:0] node42752;
	wire [4-1:0] node42753;
	wire [4-1:0] node42754;
	wire [4-1:0] node42756;
	wire [4-1:0] node42759;
	wire [4-1:0] node42761;
	wire [4-1:0] node42764;
	wire [4-1:0] node42765;
	wire [4-1:0] node42767;
	wire [4-1:0] node42770;
	wire [4-1:0] node42772;
	wire [4-1:0] node42775;
	wire [4-1:0] node42776;
	wire [4-1:0] node42779;
	wire [4-1:0] node42782;
	wire [4-1:0] node42783;
	wire [4-1:0] node42784;
	wire [4-1:0] node42785;
	wire [4-1:0] node42786;
	wire [4-1:0] node42789;
	wire [4-1:0] node42792;
	wire [4-1:0] node42793;
	wire [4-1:0] node42797;
	wire [4-1:0] node42798;
	wire [4-1:0] node42799;
	wire [4-1:0] node42800;
	wire [4-1:0] node42803;
	wire [4-1:0] node42806;
	wire [4-1:0] node42807;
	wire [4-1:0] node42808;
	wire [4-1:0] node42812;
	wire [4-1:0] node42813;
	wire [4-1:0] node42816;
	wire [4-1:0] node42819;
	wire [4-1:0] node42820;
	wire [4-1:0] node42824;
	wire [4-1:0] node42825;
	wire [4-1:0] node42826;
	wire [4-1:0] node42827;
	wire [4-1:0] node42828;
	wire [4-1:0] node42829;
	wire [4-1:0] node42833;
	wire [4-1:0] node42834;
	wire [4-1:0] node42838;
	wire [4-1:0] node42839;
	wire [4-1:0] node42842;
	wire [4-1:0] node42845;
	wire [4-1:0] node42846;
	wire [4-1:0] node42850;
	wire [4-1:0] node42851;
	wire [4-1:0] node42852;
	wire [4-1:0] node42855;
	wire [4-1:0] node42858;
	wire [4-1:0] node42859;
	wire [4-1:0] node42863;
	wire [4-1:0] node42864;
	wire [4-1:0] node42865;
	wire [4-1:0] node42866;
	wire [4-1:0] node42867;
	wire [4-1:0] node42868;
	wire [4-1:0] node42869;
	wire [4-1:0] node42873;
	wire [4-1:0] node42874;
	wire [4-1:0] node42878;
	wire [4-1:0] node42879;
	wire [4-1:0] node42880;
	wire [4-1:0] node42883;
	wire [4-1:0] node42886;
	wire [4-1:0] node42887;
	wire [4-1:0] node42888;
	wire [4-1:0] node42891;
	wire [4-1:0] node42894;
	wire [4-1:0] node42895;
	wire [4-1:0] node42898;
	wire [4-1:0] node42901;
	wire [4-1:0] node42902;
	wire [4-1:0] node42904;
	wire [4-1:0] node42905;
	wire [4-1:0] node42908;
	wire [4-1:0] node42911;
	wire [4-1:0] node42912;
	wire [4-1:0] node42915;
	wire [4-1:0] node42918;
	wire [4-1:0] node42919;
	wire [4-1:0] node42920;
	wire [4-1:0] node42921;
	wire [4-1:0] node42922;
	wire [4-1:0] node42925;
	wire [4-1:0] node42928;
	wire [4-1:0] node42929;
	wire [4-1:0] node42932;
	wire [4-1:0] node42935;
	wire [4-1:0] node42936;
	wire [4-1:0] node42937;
	wire [4-1:0] node42938;
	wire [4-1:0] node42942;
	wire [4-1:0] node42943;
	wire [4-1:0] node42946;
	wire [4-1:0] node42949;
	wire [4-1:0] node42950;
	wire [4-1:0] node42951;
	wire [4-1:0] node42955;
	wire [4-1:0] node42956;
	wire [4-1:0] node42959;
	wire [4-1:0] node42962;
	wire [4-1:0] node42963;
	wire [4-1:0] node42964;
	wire [4-1:0] node42965;
	wire [4-1:0] node42969;
	wire [4-1:0] node42970;
	wire [4-1:0] node42974;
	wire [4-1:0] node42975;
	wire [4-1:0] node42977;
	wire [4-1:0] node42978;
	wire [4-1:0] node42981;
	wire [4-1:0] node42984;
	wire [4-1:0] node42985;
	wire [4-1:0] node42988;
	wire [4-1:0] node42991;
	wire [4-1:0] node42992;
	wire [4-1:0] node42993;
	wire [4-1:0] node42995;
	wire [4-1:0] node42996;
	wire [4-1:0] node43000;
	wire [4-1:0] node43002;
	wire [4-1:0] node43003;
	wire [4-1:0] node43007;
	wire [4-1:0] node43008;
	wire [4-1:0] node43009;
	wire [4-1:0] node43010;
	wire [4-1:0] node43015;
	wire [4-1:0] node43016;
	wire [4-1:0] node43018;
	wire [4-1:0] node43022;
	wire [4-1:0] node43023;
	wire [4-1:0] node43024;
	wire [4-1:0] node43025;
	wire [4-1:0] node43026;
	wire [4-1:0] node43027;
	wire [4-1:0] node43029;
	wire [4-1:0] node43031;
	wire [4-1:0] node43034;
	wire [4-1:0] node43035;
	wire [4-1:0] node43037;
	wire [4-1:0] node43040;
	wire [4-1:0] node43041;
	wire [4-1:0] node43042;
	wire [4-1:0] node43044;
	wire [4-1:0] node43048;
	wire [4-1:0] node43049;
	wire [4-1:0] node43052;
	wire [4-1:0] node43055;
	wire [4-1:0] node43056;
	wire [4-1:0] node43058;
	wire [4-1:0] node43059;
	wire [4-1:0] node43063;
	wire [4-1:0] node43064;
	wire [4-1:0] node43065;
	wire [4-1:0] node43069;
	wire [4-1:0] node43070;
	wire [4-1:0] node43071;
	wire [4-1:0] node43072;
	wire [4-1:0] node43075;
	wire [4-1:0] node43078;
	wire [4-1:0] node43079;
	wire [4-1:0] node43083;
	wire [4-1:0] node43085;
	wire [4-1:0] node43088;
	wire [4-1:0] node43089;
	wire [4-1:0] node43090;
	wire [4-1:0] node43092;
	wire [4-1:0] node43094;
	wire [4-1:0] node43097;
	wire [4-1:0] node43098;
	wire [4-1:0] node43099;
	wire [4-1:0] node43100;
	wire [4-1:0] node43103;
	wire [4-1:0] node43106;
	wire [4-1:0] node43107;
	wire [4-1:0] node43110;
	wire [4-1:0] node43113;
	wire [4-1:0] node43115;
	wire [4-1:0] node43118;
	wire [4-1:0] node43119;
	wire [4-1:0] node43121;
	wire [4-1:0] node43123;
	wire [4-1:0] node43126;
	wire [4-1:0] node43127;
	wire [4-1:0] node43129;
	wire [4-1:0] node43132;
	wire [4-1:0] node43133;
	wire [4-1:0] node43134;
	wire [4-1:0] node43135;
	wire [4-1:0] node43138;
	wire [4-1:0] node43141;
	wire [4-1:0] node43142;
	wire [4-1:0] node43146;
	wire [4-1:0] node43148;
	wire [4-1:0] node43151;
	wire [4-1:0] node43152;
	wire [4-1:0] node43153;
	wire [4-1:0] node43154;
	wire [4-1:0] node43155;
	wire [4-1:0] node43157;
	wire [4-1:0] node43158;
	wire [4-1:0] node43161;
	wire [4-1:0] node43163;
	wire [4-1:0] node43166;
	wire [4-1:0] node43168;
	wire [4-1:0] node43170;
	wire [4-1:0] node43173;
	wire [4-1:0] node43174;
	wire [4-1:0] node43176;
	wire [4-1:0] node43177;
	wire [4-1:0] node43180;
	wire [4-1:0] node43183;
	wire [4-1:0] node43185;
	wire [4-1:0] node43186;
	wire [4-1:0] node43190;
	wire [4-1:0] node43191;
	wire [4-1:0] node43192;
	wire [4-1:0] node43193;
	wire [4-1:0] node43194;
	wire [4-1:0] node43195;
	wire [4-1:0] node43198;
	wire [4-1:0] node43201;
	wire [4-1:0] node43202;
	wire [4-1:0] node43206;
	wire [4-1:0] node43207;
	wire [4-1:0] node43210;
	wire [4-1:0] node43213;
	wire [4-1:0] node43214;
	wire [4-1:0] node43215;
	wire [4-1:0] node43217;
	wire [4-1:0] node43220;
	wire [4-1:0] node43223;
	wire [4-1:0] node43224;
	wire [4-1:0] node43227;
	wire [4-1:0] node43230;
	wire [4-1:0] node43231;
	wire [4-1:0] node43233;
	wire [4-1:0] node43234;
	wire [4-1:0] node43237;
	wire [4-1:0] node43240;
	wire [4-1:0] node43241;
	wire [4-1:0] node43242;
	wire [4-1:0] node43245;
	wire [4-1:0] node43248;
	wire [4-1:0] node43249;
	wire [4-1:0] node43251;
	wire [4-1:0] node43254;
	wire [4-1:0] node43257;
	wire [4-1:0] node43258;
	wire [4-1:0] node43259;
	wire [4-1:0] node43260;
	wire [4-1:0] node43261;
	wire [4-1:0] node43262;
	wire [4-1:0] node43266;
	wire [4-1:0] node43267;
	wire [4-1:0] node43269;
	wire [4-1:0] node43272;
	wire [4-1:0] node43273;
	wire [4-1:0] node43276;
	wire [4-1:0] node43279;
	wire [4-1:0] node43280;
	wire [4-1:0] node43281;
	wire [4-1:0] node43284;
	wire [4-1:0] node43287;
	wire [4-1:0] node43288;
	wire [4-1:0] node43290;
	wire [4-1:0] node43293;
	wire [4-1:0] node43294;
	wire [4-1:0] node43298;
	wire [4-1:0] node43299;
	wire [4-1:0] node43300;
	wire [4-1:0] node43301;
	wire [4-1:0] node43304;
	wire [4-1:0] node43307;
	wire [4-1:0] node43308;
	wire [4-1:0] node43311;
	wire [4-1:0] node43314;
	wire [4-1:0] node43315;
	wire [4-1:0] node43316;
	wire [4-1:0] node43319;
	wire [4-1:0] node43322;
	wire [4-1:0] node43323;
	wire [4-1:0] node43326;
	wire [4-1:0] node43329;
	wire [4-1:0] node43330;
	wire [4-1:0] node43331;
	wire [4-1:0] node43333;
	wire [4-1:0] node43334;
	wire [4-1:0] node43336;
	wire [4-1:0] node43339;
	wire [4-1:0] node43341;
	wire [4-1:0] node43344;
	wire [4-1:0] node43345;
	wire [4-1:0] node43346;
	wire [4-1:0] node43349;
	wire [4-1:0] node43352;
	wire [4-1:0] node43353;
	wire [4-1:0] node43356;
	wire [4-1:0] node43359;
	wire [4-1:0] node43360;
	wire [4-1:0] node43363;
	wire [4-1:0] node43366;
	wire [4-1:0] node43367;
	wire [4-1:0] node43368;
	wire [4-1:0] node43369;
	wire [4-1:0] node43370;
	wire [4-1:0] node43373;
	wire [4-1:0] node43376;
	wire [4-1:0] node43377;
	wire [4-1:0] node43378;
	wire [4-1:0] node43379;
	wire [4-1:0] node43381;
	wire [4-1:0] node43382;
	wire [4-1:0] node43387;
	wire [4-1:0] node43388;
	wire [4-1:0] node43390;
	wire [4-1:0] node43393;
	wire [4-1:0] node43394;
	wire [4-1:0] node43397;
	wire [4-1:0] node43400;
	wire [4-1:0] node43401;
	wire [4-1:0] node43402;
	wire [4-1:0] node43403;
	wire [4-1:0] node43404;
	wire [4-1:0] node43407;
	wire [4-1:0] node43410;
	wire [4-1:0] node43411;
	wire [4-1:0] node43414;
	wire [4-1:0] node43417;
	wire [4-1:0] node43419;
	wire [4-1:0] node43420;
	wire [4-1:0] node43424;
	wire [4-1:0] node43425;
	wire [4-1:0] node43426;
	wire [4-1:0] node43429;
	wire [4-1:0] node43432;
	wire [4-1:0] node43433;
	wire [4-1:0] node43435;
	wire [4-1:0] node43438;
	wire [4-1:0] node43439;
	wire [4-1:0] node43442;
	wire [4-1:0] node43445;
	wire [4-1:0] node43446;
	wire [4-1:0] node43447;
	wire [4-1:0] node43448;
	wire [4-1:0] node43449;
	wire [4-1:0] node43450;
	wire [4-1:0] node43451;
	wire [4-1:0] node43454;
	wire [4-1:0] node43457;
	wire [4-1:0] node43459;
	wire [4-1:0] node43463;
	wire [4-1:0] node43464;
	wire [4-1:0] node43465;
	wire [4-1:0] node43466;
	wire [4-1:0] node43469;
	wire [4-1:0] node43473;
	wire [4-1:0] node43474;
	wire [4-1:0] node43475;
	wire [4-1:0] node43478;
	wire [4-1:0] node43481;
	wire [4-1:0] node43483;
	wire [4-1:0] node43486;
	wire [4-1:0] node43487;
	wire [4-1:0] node43488;
	wire [4-1:0] node43489;
	wire [4-1:0] node43494;
	wire [4-1:0] node43495;
	wire [4-1:0] node43496;
	wire [4-1:0] node43500;
	wire [4-1:0] node43501;
	wire [4-1:0] node43505;
	wire [4-1:0] node43506;
	wire [4-1:0] node43507;
	wire [4-1:0] node43508;
	wire [4-1:0] node43509;
	wire [4-1:0] node43510;
	wire [4-1:0] node43513;
	wire [4-1:0] node43517;
	wire [4-1:0] node43519;
	wire [4-1:0] node43521;
	wire [4-1:0] node43524;
	wire [4-1:0] node43525;
	wire [4-1:0] node43526;
	wire [4-1:0] node43527;
	wire [4-1:0] node43530;
	wire [4-1:0] node43534;
	wire [4-1:0] node43535;
	wire [4-1:0] node43536;
	wire [4-1:0] node43539;
	wire [4-1:0] node43543;
	wire [4-1:0] node43544;
	wire [4-1:0] node43545;
	wire [4-1:0] node43546;
	wire [4-1:0] node43550;
	wire [4-1:0] node43551;
	wire [4-1:0] node43555;
	wire [4-1:0] node43556;
	wire [4-1:0] node43557;
	wire [4-1:0] node43561;
	wire [4-1:0] node43562;
	wire [4-1:0] node43566;
	wire [4-1:0] node43567;
	wire [4-1:0] node43568;
	wire [4-1:0] node43569;
	wire [4-1:0] node43570;
	wire [4-1:0] node43571;
	wire [4-1:0] node43572;
	wire [4-1:0] node43577;
	wire [4-1:0] node43578;
	wire [4-1:0] node43579;
	wire [4-1:0] node43582;
	wire [4-1:0] node43585;
	wire [4-1:0] node43586;
	wire [4-1:0] node43589;
	wire [4-1:0] node43592;
	wire [4-1:0] node43594;
	wire [4-1:0] node43595;
	wire [4-1:0] node43599;
	wire [4-1:0] node43600;
	wire [4-1:0] node43601;
	wire [4-1:0] node43602;
	wire [4-1:0] node43605;
	wire [4-1:0] node43608;
	wire [4-1:0] node43610;
	wire [4-1:0] node43613;
	wire [4-1:0] node43615;
	wire [4-1:0] node43616;
	wire [4-1:0] node43620;
	wire [4-1:0] node43621;
	wire [4-1:0] node43622;
	wire [4-1:0] node43623;
	wire [4-1:0] node43624;
	wire [4-1:0] node43628;
	wire [4-1:0] node43629;
	wire [4-1:0] node43630;
	wire [4-1:0] node43631;
	wire [4-1:0] node43634;
	wire [4-1:0] node43637;
	wire [4-1:0] node43638;
	wire [4-1:0] node43641;
	wire [4-1:0] node43644;
	wire [4-1:0] node43645;
	wire [4-1:0] node43648;
	wire [4-1:0] node43651;
	wire [4-1:0] node43652;
	wire [4-1:0] node43653;
	wire [4-1:0] node43658;
	wire [4-1:0] node43659;
	wire [4-1:0] node43660;
	wire [4-1:0] node43661;
	wire [4-1:0] node43662;
	wire [4-1:0] node43665;
	wire [4-1:0] node43668;
	wire [4-1:0] node43670;
	wire [4-1:0] node43671;
	wire [4-1:0] node43674;
	wire [4-1:0] node43677;
	wire [4-1:0] node43679;
	wire [4-1:0] node43682;
	wire [4-1:0] node43683;
	wire [4-1:0] node43684;
	wire [4-1:0] node43689;
	wire [4-1:0] node43690;
	wire [4-1:0] node43691;
	wire [4-1:0] node43692;
	wire [4-1:0] node43693;
	wire [4-1:0] node43694;
	wire [4-1:0] node43695;
	wire [4-1:0] node43696;
	wire [4-1:0] node43699;
	wire [4-1:0] node43702;
	wire [4-1:0] node43703;
	wire [4-1:0] node43704;
	wire [4-1:0] node43707;
	wire [4-1:0] node43710;
	wire [4-1:0] node43711;
	wire [4-1:0] node43714;
	wire [4-1:0] node43717;
	wire [4-1:0] node43718;
	wire [4-1:0] node43719;
	wire [4-1:0] node43721;
	wire [4-1:0] node43724;
	wire [4-1:0] node43726;
	wire [4-1:0] node43729;
	wire [4-1:0] node43730;
	wire [4-1:0] node43732;
	wire [4-1:0] node43735;
	wire [4-1:0] node43737;
	wire [4-1:0] node43740;
	wire [4-1:0] node43741;
	wire [4-1:0] node43742;
	wire [4-1:0] node43743;
	wire [4-1:0] node43744;
	wire [4-1:0] node43745;
	wire [4-1:0] node43746;
	wire [4-1:0] node43748;
	wire [4-1:0] node43751;
	wire [4-1:0] node43754;
	wire [4-1:0] node43755;
	wire [4-1:0] node43758;
	wire [4-1:0] node43761;
	wire [4-1:0] node43762;
	wire [4-1:0] node43764;
	wire [4-1:0] node43767;
	wire [4-1:0] node43768;
	wire [4-1:0] node43769;
	wire [4-1:0] node43773;
	wire [4-1:0] node43774;
	wire [4-1:0] node43777;
	wire [4-1:0] node43780;
	wire [4-1:0] node43781;
	wire [4-1:0] node43782;
	wire [4-1:0] node43785;
	wire [4-1:0] node43788;
	wire [4-1:0] node43789;
	wire [4-1:0] node43792;
	wire [4-1:0] node43795;
	wire [4-1:0] node43796;
	wire [4-1:0] node43797;
	wire [4-1:0] node43800;
	wire [4-1:0] node43803;
	wire [4-1:0] node43804;
	wire [4-1:0] node43805;
	wire [4-1:0] node43806;
	wire [4-1:0] node43807;
	wire [4-1:0] node43810;
	wire [4-1:0] node43813;
	wire [4-1:0] node43814;
	wire [4-1:0] node43817;
	wire [4-1:0] node43820;
	wire [4-1:0] node43822;
	wire [4-1:0] node43823;
	wire [4-1:0] node43826;
	wire [4-1:0] node43829;
	wire [4-1:0] node43830;
	wire [4-1:0] node43831;
	wire [4-1:0] node43834;
	wire [4-1:0] node43838;
	wire [4-1:0] node43839;
	wire [4-1:0] node43840;
	wire [4-1:0] node43841;
	wire [4-1:0] node43845;
	wire [4-1:0] node43846;
	wire [4-1:0] node43850;
	wire [4-1:0] node43851;
	wire [4-1:0] node43852;
	wire [4-1:0] node43856;
	wire [4-1:0] node43857;
	wire [4-1:0] node43861;
	wire [4-1:0] node43862;
	wire [4-1:0] node43863;
	wire [4-1:0] node43864;
	wire [4-1:0] node43865;
	wire [4-1:0] node43866;
	wire [4-1:0] node43867;
	wire [4-1:0] node43868;
	wire [4-1:0] node43871;
	wire [4-1:0] node43874;
	wire [4-1:0] node43875;
	wire [4-1:0] node43878;
	wire [4-1:0] node43881;
	wire [4-1:0] node43882;
	wire [4-1:0] node43885;
	wire [4-1:0] node43888;
	wire [4-1:0] node43889;
	wire [4-1:0] node43890;
	wire [4-1:0] node43891;
	wire [4-1:0] node43892;
	wire [4-1:0] node43895;
	wire [4-1:0] node43899;
	wire [4-1:0] node43900;
	wire [4-1:0] node43902;
	wire [4-1:0] node43905;
	wire [4-1:0] node43906;
	wire [4-1:0] node43909;
	wire [4-1:0] node43912;
	wire [4-1:0] node43913;
	wire [4-1:0] node43914;
	wire [4-1:0] node43918;
	wire [4-1:0] node43919;
	wire [4-1:0] node43922;
	wire [4-1:0] node43925;
	wire [4-1:0] node43926;
	wire [4-1:0] node43927;
	wire [4-1:0] node43928;
	wire [4-1:0] node43929;
	wire [4-1:0] node43932;
	wire [4-1:0] node43935;
	wire [4-1:0] node43936;
	wire [4-1:0] node43939;
	wire [4-1:0] node43942;
	wire [4-1:0] node43943;
	wire [4-1:0] node43944;
	wire [4-1:0] node43948;
	wire [4-1:0] node43949;
	wire [4-1:0] node43950;
	wire [4-1:0] node43954;
	wire [4-1:0] node43956;
	wire [4-1:0] node43959;
	wire [4-1:0] node43960;
	wire [4-1:0] node43963;
	wire [4-1:0] node43966;
	wire [4-1:0] node43967;
	wire [4-1:0] node43968;
	wire [4-1:0] node43969;
	wire [4-1:0] node43970;
	wire [4-1:0] node43973;
	wire [4-1:0] node43976;
	wire [4-1:0] node43977;
	wire [4-1:0] node43980;
	wire [4-1:0] node43983;
	wire [4-1:0] node43984;
	wire [4-1:0] node43985;
	wire [4-1:0] node43986;
	wire [4-1:0] node43987;
	wire [4-1:0] node43991;
	wire [4-1:0] node43994;
	wire [4-1:0] node43995;
	wire [4-1:0] node43996;
	wire [4-1:0] node43999;
	wire [4-1:0] node44002;
	wire [4-1:0] node44003;
	wire [4-1:0] node44006;
	wire [4-1:0] node44009;
	wire [4-1:0] node44010;
	wire [4-1:0] node44011;
	wire [4-1:0] node44014;
	wire [4-1:0] node44017;
	wire [4-1:0] node44018;
	wire [4-1:0] node44021;
	wire [4-1:0] node44024;
	wire [4-1:0] node44025;
	wire [4-1:0] node44026;
	wire [4-1:0] node44027;
	wire [4-1:0] node44028;
	wire [4-1:0] node44032;
	wire [4-1:0] node44033;
	wire [4-1:0] node44034;
	wire [4-1:0] node44037;
	wire [4-1:0] node44040;
	wire [4-1:0] node44041;
	wire [4-1:0] node44044;
	wire [4-1:0] node44047;
	wire [4-1:0] node44048;
	wire [4-1:0] node44049;
	wire [4-1:0] node44052;
	wire [4-1:0] node44055;
	wire [4-1:0] node44056;
	wire [4-1:0] node44060;
	wire [4-1:0] node44061;
	wire [4-1:0] node44062;
	wire [4-1:0] node44063;
	wire [4-1:0] node44064;
	wire [4-1:0] node44067;
	wire [4-1:0] node44070;
	wire [4-1:0] node44071;
	wire [4-1:0] node44074;
	wire [4-1:0] node44078;
	wire [4-1:0] node44079;
	wire [4-1:0] node44081;
	wire [4-1:0] node44082;
	wire [4-1:0] node44085;
	wire [4-1:0] node44088;
	wire [4-1:0] node44089;
	wire [4-1:0] node44090;
	wire [4-1:0] node44093;
	wire [4-1:0] node44096;
	wire [4-1:0] node44097;
	wire [4-1:0] node44100;
	wire [4-1:0] node44103;
	wire [4-1:0] node44104;
	wire [4-1:0] node44105;
	wire [4-1:0] node44106;
	wire [4-1:0] node44107;
	wire [4-1:0] node44110;
	wire [4-1:0] node44113;
	wire [4-1:0] node44114;
	wire [4-1:0] node44115;
	wire [4-1:0] node44116;
	wire [4-1:0] node44119;
	wire [4-1:0] node44122;
	wire [4-1:0] node44123;
	wire [4-1:0] node44126;
	wire [4-1:0] node44129;
	wire [4-1:0] node44130;
	wire [4-1:0] node44132;
	wire [4-1:0] node44135;
	wire [4-1:0] node44136;
	wire [4-1:0] node44138;
	wire [4-1:0] node44141;
	wire [4-1:0] node44142;
	wire [4-1:0] node44145;
	wire [4-1:0] node44148;
	wire [4-1:0] node44149;
	wire [4-1:0] node44150;
	wire [4-1:0] node44151;
	wire [4-1:0] node44154;
	wire [4-1:0] node44157;
	wire [4-1:0] node44158;
	wire [4-1:0] node44159;
	wire [4-1:0] node44162;
	wire [4-1:0] node44165;
	wire [4-1:0] node44167;
	wire [4-1:0] node44168;
	wire [4-1:0] node44171;
	wire [4-1:0] node44174;
	wire [4-1:0] node44175;
	wire [4-1:0] node44176;
	wire [4-1:0] node44179;
	wire [4-1:0] node44182;
	wire [4-1:0] node44183;
	wire [4-1:0] node44186;
	wire [4-1:0] node44189;
	wire [4-1:0] node44190;
	wire [4-1:0] node44191;
	wire [4-1:0] node44192;
	wire [4-1:0] node44193;
	wire [4-1:0] node44196;
	wire [4-1:0] node44199;
	wire [4-1:0] node44200;
	wire [4-1:0] node44201;
	wire [4-1:0] node44204;
	wire [4-1:0] node44207;
	wire [4-1:0] node44208;
	wire [4-1:0] node44211;
	wire [4-1:0] node44213;
	wire [4-1:0] node44216;
	wire [4-1:0] node44217;
	wire [4-1:0] node44219;
	wire [4-1:0] node44222;
	wire [4-1:0] node44223;
	wire [4-1:0] node44226;
	wire [4-1:0] node44229;
	wire [4-1:0] node44230;
	wire [4-1:0] node44231;
	wire [4-1:0] node44232;
	wire [4-1:0] node44235;
	wire [4-1:0] node44238;
	wire [4-1:0] node44239;
	wire [4-1:0] node44240;
	wire [4-1:0] node44243;
	wire [4-1:0] node44246;
	wire [4-1:0] node44248;
	wire [4-1:0] node44251;
	wire [4-1:0] node44252;
	wire [4-1:0] node44253;
	wire [4-1:0] node44256;
	wire [4-1:0] node44259;
	wire [4-1:0] node44260;
	wire [4-1:0] node44261;
	wire [4-1:0] node44263;
	wire [4-1:0] node44266;
	wire [4-1:0] node44267;
	wire [4-1:0] node44270;
	wire [4-1:0] node44273;
	wire [4-1:0] node44274;
	wire [4-1:0] node44277;
	wire [4-1:0] node44280;
	wire [4-1:0] node44281;
	wire [4-1:0] node44282;
	wire [4-1:0] node44283;
	wire [4-1:0] node44284;
	wire [4-1:0] node44285;
	wire [4-1:0] node44286;
	wire [4-1:0] node44289;
	wire [4-1:0] node44292;
	wire [4-1:0] node44295;
	wire [4-1:0] node44296;
	wire [4-1:0] node44297;
	wire [4-1:0] node44301;
	wire [4-1:0] node44302;
	wire [4-1:0] node44306;
	wire [4-1:0] node44307;
	wire [4-1:0] node44308;
	wire [4-1:0] node44309;
	wire [4-1:0] node44312;
	wire [4-1:0] node44315;
	wire [4-1:0] node44316;
	wire [4-1:0] node44319;
	wire [4-1:0] node44322;
	wire [4-1:0] node44323;
	wire [4-1:0] node44324;
	wire [4-1:0] node44328;
	wire [4-1:0] node44329;
	wire [4-1:0] node44333;
	wire [4-1:0] node44334;
	wire [4-1:0] node44335;
	wire [4-1:0] node44336;
	wire [4-1:0] node44337;
	wire [4-1:0] node44341;
	wire [4-1:0] node44342;
	wire [4-1:0] node44346;
	wire [4-1:0] node44347;
	wire [4-1:0] node44348;
	wire [4-1:0] node44351;
	wire [4-1:0] node44354;
	wire [4-1:0] node44357;
	wire [4-1:0] node44358;
	wire [4-1:0] node44359;
	wire [4-1:0] node44360;
	wire [4-1:0] node44361;
	wire [4-1:0] node44364;
	wire [4-1:0] node44367;
	wire [4-1:0] node44368;
	wire [4-1:0] node44369;
	wire [4-1:0] node44370;
	wire [4-1:0] node44373;
	wire [4-1:0] node44376;
	wire [4-1:0] node44377;
	wire [4-1:0] node44380;
	wire [4-1:0] node44383;
	wire [4-1:0] node44384;
	wire [4-1:0] node44385;
	wire [4-1:0] node44388;
	wire [4-1:0] node44391;
	wire [4-1:0] node44392;
	wire [4-1:0] node44395;
	wire [4-1:0] node44398;
	wire [4-1:0] node44401;
	wire [4-1:0] node44402;
	wire [4-1:0] node44406;
	wire [4-1:0] node44407;
	wire [4-1:0] node44408;
	wire [4-1:0] node44409;
	wire [4-1:0] node44410;
	wire [4-1:0] node44411;
	wire [4-1:0] node44414;
	wire [4-1:0] node44417;
	wire [4-1:0] node44420;
	wire [4-1:0] node44421;
	wire [4-1:0] node44422;
	wire [4-1:0] node44426;
	wire [4-1:0] node44427;
	wire [4-1:0] node44431;
	wire [4-1:0] node44432;
	wire [4-1:0] node44433;
	wire [4-1:0] node44436;
	wire [4-1:0] node44437;
	wire [4-1:0] node44438;
	wire [4-1:0] node44441;
	wire [4-1:0] node44444;
	wire [4-1:0] node44445;
	wire [4-1:0] node44446;
	wire [4-1:0] node44448;
	wire [4-1:0] node44451;
	wire [4-1:0] node44452;
	wire [4-1:0] node44455;
	wire [4-1:0] node44458;
	wire [4-1:0] node44460;
	wire [4-1:0] node44463;
	wire [4-1:0] node44464;
	wire [4-1:0] node44468;
	wire [4-1:0] node44469;
	wire [4-1:0] node44470;
	wire [4-1:0] node44471;
	wire [4-1:0] node44472;
	wire [4-1:0] node44476;
	wire [4-1:0] node44477;
	wire [4-1:0] node44481;
	wire [4-1:0] node44482;
	wire [4-1:0] node44483;
	wire [4-1:0] node44486;
	wire [4-1:0] node44489;
	wire [4-1:0] node44492;
	wire [4-1:0] node44493;
	wire [4-1:0] node44494;
	wire [4-1:0] node44495;
	wire [4-1:0] node44496;
	wire [4-1:0] node44499;
	wire [4-1:0] node44502;
	wire [4-1:0] node44503;
	wire [4-1:0] node44504;
	wire [4-1:0] node44508;
	wire [4-1:0] node44509;
	wire [4-1:0] node44512;
	wire [4-1:0] node44515;
	wire [4-1:0] node44518;
	wire [4-1:0] node44519;
	wire [4-1:0] node44523;
	wire [4-1:0] node44524;
	wire [4-1:0] node44525;
	wire [4-1:0] node44526;
	wire [4-1:0] node44527;
	wire [4-1:0] node44528;
	wire [4-1:0] node44530;
	wire [4-1:0] node44533;
	wire [4-1:0] node44535;
	wire [4-1:0] node44538;
	wire [4-1:0] node44539;
	wire [4-1:0] node44541;
	wire [4-1:0] node44544;
	wire [4-1:0] node44546;
	wire [4-1:0] node44549;
	wire [4-1:0] node44550;
	wire [4-1:0] node44551;
	wire [4-1:0] node44552;
	wire [4-1:0] node44553;
	wire [4-1:0] node44554;
	wire [4-1:0] node44557;
	wire [4-1:0] node44560;
	wire [4-1:0] node44561;
	wire [4-1:0] node44562;
	wire [4-1:0] node44565;
	wire [4-1:0] node44569;
	wire [4-1:0] node44570;
	wire [4-1:0] node44573;
	wire [4-1:0] node44576;
	wire [4-1:0] node44577;
	wire [4-1:0] node44578;
	wire [4-1:0] node44579;
	wire [4-1:0] node44580;
	wire [4-1:0] node44583;
	wire [4-1:0] node44586;
	wire [4-1:0] node44587;
	wire [4-1:0] node44590;
	wire [4-1:0] node44593;
	wire [4-1:0] node44594;
	wire [4-1:0] node44596;
	wire [4-1:0] node44599;
	wire [4-1:0] node44600;
	wire [4-1:0] node44603;
	wire [4-1:0] node44606;
	wire [4-1:0] node44607;
	wire [4-1:0] node44608;
	wire [4-1:0] node44609;
	wire [4-1:0] node44610;
	wire [4-1:0] node44614;
	wire [4-1:0] node44615;
	wire [4-1:0] node44618;
	wire [4-1:0] node44621;
	wire [4-1:0] node44622;
	wire [4-1:0] node44625;
	wire [4-1:0] node44628;
	wire [4-1:0] node44629;
	wire [4-1:0] node44631;
	wire [4-1:0] node44632;
	wire [4-1:0] node44635;
	wire [4-1:0] node44638;
	wire [4-1:0] node44639;
	wire [4-1:0] node44642;
	wire [4-1:0] node44645;
	wire [4-1:0] node44646;
	wire [4-1:0] node44647;
	wire [4-1:0] node44648;
	wire [4-1:0] node44649;
	wire [4-1:0] node44653;
	wire [4-1:0] node44654;
	wire [4-1:0] node44657;
	wire [4-1:0] node44660;
	wire [4-1:0] node44661;
	wire [4-1:0] node44662;
	wire [4-1:0] node44663;
	wire [4-1:0] node44666;
	wire [4-1:0] node44669;
	wire [4-1:0] node44670;
	wire [4-1:0] node44674;
	wire [4-1:0] node44675;
	wire [4-1:0] node44678;
	wire [4-1:0] node44681;
	wire [4-1:0] node44682;
	wire [4-1:0] node44683;
	wire [4-1:0] node44684;
	wire [4-1:0] node44687;
	wire [4-1:0] node44690;
	wire [4-1:0] node44691;
	wire [4-1:0] node44694;
	wire [4-1:0] node44695;
	wire [4-1:0] node44698;
	wire [4-1:0] node44701;
	wire [4-1:0] node44702;
	wire [4-1:0] node44705;
	wire [4-1:0] node44708;
	wire [4-1:0] node44709;
	wire [4-1:0] node44710;
	wire [4-1:0] node44711;
	wire [4-1:0] node44712;
	wire [4-1:0] node44713;
	wire [4-1:0] node44714;
	wire [4-1:0] node44717;
	wire [4-1:0] node44721;
	wire [4-1:0] node44722;
	wire [4-1:0] node44723;
	wire [4-1:0] node44725;
	wire [4-1:0] node44728;
	wire [4-1:0] node44729;
	wire [4-1:0] node44730;
	wire [4-1:0] node44733;
	wire [4-1:0] node44738;
	wire [4-1:0] node44739;
	wire [4-1:0] node44740;
	wire [4-1:0] node44744;
	wire [4-1:0] node44745;
	wire [4-1:0] node44749;
	wire [4-1:0] node44750;
	wire [4-1:0] node44751;
	wire [4-1:0] node44752;
	wire [4-1:0] node44754;
	wire [4-1:0] node44757;
	wire [4-1:0] node44758;
	wire [4-1:0] node44762;
	wire [4-1:0] node44763;
	wire [4-1:0] node44765;
	wire [4-1:0] node44768;
	wire [4-1:0] node44769;
	wire [4-1:0] node44773;
	wire [4-1:0] node44774;
	wire [4-1:0] node44777;
	wire [4-1:0] node44780;
	wire [4-1:0] node44781;
	wire [4-1:0] node44782;
	wire [4-1:0] node44783;
	wire [4-1:0] node44785;
	wire [4-1:0] node44788;
	wire [4-1:0] node44791;
	wire [4-1:0] node44792;
	wire [4-1:0] node44794;
	wire [4-1:0] node44797;
	wire [4-1:0] node44798;
	wire [4-1:0] node44799;
	wire [4-1:0] node44801;
	wire [4-1:0] node44804;
	wire [4-1:0] node44805;
	wire [4-1:0] node44808;
	wire [4-1:0] node44811;
	wire [4-1:0] node44812;
	wire [4-1:0] node44813;
	wire [4-1:0] node44816;
	wire [4-1:0] node44819;
	wire [4-1:0] node44820;
	wire [4-1:0] node44824;
	wire [4-1:0] node44825;
	wire [4-1:0] node44826;
	wire [4-1:0] node44827;
	wire [4-1:0] node44832;
	wire [4-1:0] node44833;
	wire [4-1:0] node44834;
	wire [4-1:0] node44839;
	wire [4-1:0] node44840;
	wire [4-1:0] node44841;
	wire [4-1:0] node44842;
	wire [4-1:0] node44843;
	wire [4-1:0] node44844;
	wire [4-1:0] node44845;
	wire [4-1:0] node44846;
	wire [4-1:0] node44847;
	wire [4-1:0] node44848;
	wire [4-1:0] node44851;
	wire [4-1:0] node44854;
	wire [4-1:0] node44856;
	wire [4-1:0] node44859;
	wire [4-1:0] node44861;
	wire [4-1:0] node44864;
	wire [4-1:0] node44865;
	wire [4-1:0] node44866;
	wire [4-1:0] node44869;
	wire [4-1:0] node44872;
	wire [4-1:0] node44873;
	wire [4-1:0] node44874;
	wire [4-1:0] node44877;
	wire [4-1:0] node44880;
	wire [4-1:0] node44881;
	wire [4-1:0] node44885;
	wire [4-1:0] node44886;
	wire [4-1:0] node44887;
	wire [4-1:0] node44890;
	wire [4-1:0] node44893;
	wire [4-1:0] node44894;
	wire [4-1:0] node44895;
	wire [4-1:0] node44899;
	wire [4-1:0] node44900;
	wire [4-1:0] node44902;
	wire [4-1:0] node44905;
	wire [4-1:0] node44907;
	wire [4-1:0] node44910;
	wire [4-1:0] node44911;
	wire [4-1:0] node44912;
	wire [4-1:0] node44913;
	wire [4-1:0] node44916;
	wire [4-1:0] node44919;
	wire [4-1:0] node44920;
	wire [4-1:0] node44922;
	wire [4-1:0] node44925;
	wire [4-1:0] node44926;
	wire [4-1:0] node44927;
	wire [4-1:0] node44930;
	wire [4-1:0] node44933;
	wire [4-1:0] node44934;
	wire [4-1:0] node44938;
	wire [4-1:0] node44939;
	wire [4-1:0] node44940;
	wire [4-1:0] node44943;
	wire [4-1:0] node44946;
	wire [4-1:0] node44947;
	wire [4-1:0] node44950;
	wire [4-1:0] node44953;
	wire [4-1:0] node44954;
	wire [4-1:0] node44955;
	wire [4-1:0] node44958;
	wire [4-1:0] node44961;
	wire [4-1:0] node44962;
	wire [4-1:0] node44963;
	wire [4-1:0] node44964;
	wire [4-1:0] node44965;
	wire [4-1:0] node44966;
	wire [4-1:0] node44969;
	wire [4-1:0] node44972;
	wire [4-1:0] node44973;
	wire [4-1:0] node44976;
	wire [4-1:0] node44979;
	wire [4-1:0] node44980;
	wire [4-1:0] node44983;
	wire [4-1:0] node44986;
	wire [4-1:0] node44987;
	wire [4-1:0] node44990;
	wire [4-1:0] node44993;
	wire [4-1:0] node44994;
	wire [4-1:0] node44997;
	wire [4-1:0] node45000;
	wire [4-1:0] node45001;
	wire [4-1:0] node45004;
	wire [4-1:0] node45007;
	wire [4-1:0] node45008;
	wire [4-1:0] node45009;
	wire [4-1:0] node45010;
	wire [4-1:0] node45011;
	wire [4-1:0] node45015;
	wire [4-1:0] node45016;
	wire [4-1:0] node45021;
	wire [4-1:0] node45022;
	wire [4-1:0] node45023;
	wire [4-1:0] node45024;
	wire [4-1:0] node45028;
	wire [4-1:0] node45029;
	wire [4-1:0] node45034;
	wire [4-1:0] node45035;
	wire [4-1:0] node45036;
	wire [4-1:0] node45037;
	wire [4-1:0] node45038;
	wire [4-1:0] node45039;
	wire [4-1:0] node45040;
	wire [4-1:0] node45041;
	wire [4-1:0] node45042;
	wire [4-1:0] node45043;
	wire [4-1:0] node45044;
	wire [4-1:0] node45045;
	wire [4-1:0] node45048;
	wire [4-1:0] node45051;
	wire [4-1:0] node45052;
	wire [4-1:0] node45055;
	wire [4-1:0] node45058;
	wire [4-1:0] node45059;
	wire [4-1:0] node45060;
	wire [4-1:0] node45064;
	wire [4-1:0] node45066;
	wire [4-1:0] node45067;
	wire [4-1:0] node45070;
	wire [4-1:0] node45073;
	wire [4-1:0] node45074;
	wire [4-1:0] node45075;
	wire [4-1:0] node45077;
	wire [4-1:0] node45080;
	wire [4-1:0] node45081;
	wire [4-1:0] node45083;
	wire [4-1:0] node45086;
	wire [4-1:0] node45087;
	wire [4-1:0] node45091;
	wire [4-1:0] node45092;
	wire [4-1:0] node45093;
	wire [4-1:0] node45097;
	wire [4-1:0] node45098;
	wire [4-1:0] node45101;
	wire [4-1:0] node45104;
	wire [4-1:0] node45105;
	wire [4-1:0] node45106;
	wire [4-1:0] node45107;
	wire [4-1:0] node45110;
	wire [4-1:0] node45113;
	wire [4-1:0] node45114;
	wire [4-1:0] node45117;
	wire [4-1:0] node45120;
	wire [4-1:0] node45121;
	wire [4-1:0] node45122;
	wire [4-1:0] node45125;
	wire [4-1:0] node45128;
	wire [4-1:0] node45129;
	wire [4-1:0] node45132;
	wire [4-1:0] node45135;
	wire [4-1:0] node45136;
	wire [4-1:0] node45137;
	wire [4-1:0] node45138;
	wire [4-1:0] node45139;
	wire [4-1:0] node45140;
	wire [4-1:0] node45144;
	wire [4-1:0] node45145;
	wire [4-1:0] node45148;
	wire [4-1:0] node45151;
	wire [4-1:0] node45152;
	wire [4-1:0] node45153;
	wire [4-1:0] node45155;
	wire [4-1:0] node45158;
	wire [4-1:0] node45160;
	wire [4-1:0] node45163;
	wire [4-1:0] node45164;
	wire [4-1:0] node45167;
	wire [4-1:0] node45170;
	wire [4-1:0] node45171;
	wire [4-1:0] node45172;
	wire [4-1:0] node45173;
	wire [4-1:0] node45175;
	wire [4-1:0] node45178;
	wire [4-1:0] node45179;
	wire [4-1:0] node45182;
	wire [4-1:0] node45185;
	wire [4-1:0] node45188;
	wire [4-1:0] node45189;
	wire [4-1:0] node45190;
	wire [4-1:0] node45192;
	wire [4-1:0] node45195;
	wire [4-1:0] node45196;
	wire [4-1:0] node45199;
	wire [4-1:0] node45202;
	wire [4-1:0] node45203;
	wire [4-1:0] node45205;
	wire [4-1:0] node45208;
	wire [4-1:0] node45209;
	wire [4-1:0] node45213;
	wire [4-1:0] node45214;
	wire [4-1:0] node45215;
	wire [4-1:0] node45216;
	wire [4-1:0] node45217;
	wire [4-1:0] node45218;
	wire [4-1:0] node45223;
	wire [4-1:0] node45224;
	wire [4-1:0] node45225;
	wire [4-1:0] node45228;
	wire [4-1:0] node45231;
	wire [4-1:0] node45232;
	wire [4-1:0] node45236;
	wire [4-1:0] node45237;
	wire [4-1:0] node45238;
	wire [4-1:0] node45241;
	wire [4-1:0] node45244;
	wire [4-1:0] node45245;
	wire [4-1:0] node45248;
	wire [4-1:0] node45251;
	wire [4-1:0] node45252;
	wire [4-1:0] node45253;
	wire [4-1:0] node45254;
	wire [4-1:0] node45257;
	wire [4-1:0] node45260;
	wire [4-1:0] node45261;
	wire [4-1:0] node45264;
	wire [4-1:0] node45267;
	wire [4-1:0] node45268;
	wire [4-1:0] node45270;
	wire [4-1:0] node45273;
	wire [4-1:0] node45274;
	wire [4-1:0] node45277;
	wire [4-1:0] node45280;
	wire [4-1:0] node45281;
	wire [4-1:0] node45282;
	wire [4-1:0] node45283;
	wire [4-1:0] node45284;
	wire [4-1:0] node45285;
	wire [4-1:0] node45288;
	wire [4-1:0] node45291;
	wire [4-1:0] node45293;
	wire [4-1:0] node45294;
	wire [4-1:0] node45297;
	wire [4-1:0] node45300;
	wire [4-1:0] node45301;
	wire [4-1:0] node45302;
	wire [4-1:0] node45305;
	wire [4-1:0] node45308;
	wire [4-1:0] node45311;
	wire [4-1:0] node45312;
	wire [4-1:0] node45313;
	wire [4-1:0] node45316;
	wire [4-1:0] node45317;
	wire [4-1:0] node45320;
	wire [4-1:0] node45323;
	wire [4-1:0] node45324;
	wire [4-1:0] node45325;
	wire [4-1:0] node45326;
	wire [4-1:0] node45330;
	wire [4-1:0] node45331;
	wire [4-1:0] node45334;
	wire [4-1:0] node45337;
	wire [4-1:0] node45338;
	wire [4-1:0] node45341;
	wire [4-1:0] node45344;
	wire [4-1:0] node45345;
	wire [4-1:0] node45346;
	wire [4-1:0] node45347;
	wire [4-1:0] node45349;
	wire [4-1:0] node45352;
	wire [4-1:0] node45354;
	wire [4-1:0] node45357;
	wire [4-1:0] node45358;
	wire [4-1:0] node45359;
	wire [4-1:0] node45362;
	wire [4-1:0] node45365;
	wire [4-1:0] node45366;
	wire [4-1:0] node45370;
	wire [4-1:0] node45371;
	wire [4-1:0] node45372;
	wire [4-1:0] node45374;
	wire [4-1:0] node45377;
	wire [4-1:0] node45378;
	wire [4-1:0] node45381;
	wire [4-1:0] node45384;
	wire [4-1:0] node45385;
	wire [4-1:0] node45387;
	wire [4-1:0] node45390;
	wire [4-1:0] node45391;
	wire [4-1:0] node45394;
	wire [4-1:0] node45397;
	wire [4-1:0] node45398;
	wire [4-1:0] node45399;
	wire [4-1:0] node45400;
	wire [4-1:0] node45401;
	wire [4-1:0] node45404;
	wire [4-1:0] node45407;
	wire [4-1:0] node45408;
	wire [4-1:0] node45409;
	wire [4-1:0] node45410;
	wire [4-1:0] node45411;
	wire [4-1:0] node45414;
	wire [4-1:0] node45417;
	wire [4-1:0] node45418;
	wire [4-1:0] node45421;
	wire [4-1:0] node45424;
	wire [4-1:0] node45425;
	wire [4-1:0] node45426;
	wire [4-1:0] node45429;
	wire [4-1:0] node45432;
	wire [4-1:0] node45433;
	wire [4-1:0] node45436;
	wire [4-1:0] node45439;
	wire [4-1:0] node45440;
	wire [4-1:0] node45443;
	wire [4-1:0] node45446;
	wire [4-1:0] node45447;
	wire [4-1:0] node45448;
	wire [4-1:0] node45449;
	wire [4-1:0] node45450;
	wire [4-1:0] node45452;
	wire [4-1:0] node45453;
	wire [4-1:0] node45456;
	wire [4-1:0] node45459;
	wire [4-1:0] node45460;
	wire [4-1:0] node45462;
	wire [4-1:0] node45465;
	wire [4-1:0] node45467;
	wire [4-1:0] node45470;
	wire [4-1:0] node45471;
	wire [4-1:0] node45473;
	wire [4-1:0] node45474;
	wire [4-1:0] node45477;
	wire [4-1:0] node45480;
	wire [4-1:0] node45481;
	wire [4-1:0] node45484;
	wire [4-1:0] node45487;
	wire [4-1:0] node45488;
	wire [4-1:0] node45491;
	wire [4-1:0] node45494;
	wire [4-1:0] node45495;
	wire [4-1:0] node45496;
	wire [4-1:0] node45497;
	wire [4-1:0] node45499;
	wire [4-1:0] node45502;
	wire [4-1:0] node45503;
	wire [4-1:0] node45504;
	wire [4-1:0] node45507;
	wire [4-1:0] node45510;
	wire [4-1:0] node45511;
	wire [4-1:0] node45514;
	wire [4-1:0] node45517;
	wire [4-1:0] node45518;
	wire [4-1:0] node45519;
	wire [4-1:0] node45522;
	wire [4-1:0] node45525;
	wire [4-1:0] node45526;
	wire [4-1:0] node45529;
	wire [4-1:0] node45532;
	wire [4-1:0] node45533;
	wire [4-1:0] node45534;
	wire [4-1:0] node45536;
	wire [4-1:0] node45538;
	wire [4-1:0] node45541;
	wire [4-1:0] node45542;
	wire [4-1:0] node45545;
	wire [4-1:0] node45548;
	wire [4-1:0] node45549;
	wire [4-1:0] node45550;
	wire [4-1:0] node45553;
	wire [4-1:0] node45556;
	wire [4-1:0] node45557;
	wire [4-1:0] node45560;
	wire [4-1:0] node45563;
	wire [4-1:0] node45564;
	wire [4-1:0] node45565;
	wire [4-1:0] node45566;
	wire [4-1:0] node45567;
	wire [4-1:0] node45568;
	wire [4-1:0] node45569;
	wire [4-1:0] node45572;
	wire [4-1:0] node45575;
	wire [4-1:0] node45576;
	wire [4-1:0] node45580;
	wire [4-1:0] node45581;
	wire [4-1:0] node45584;
	wire [4-1:0] node45587;
	wire [4-1:0] node45588;
	wire [4-1:0] node45591;
	wire [4-1:0] node45594;
	wire [4-1:0] node45595;
	wire [4-1:0] node45596;
	wire [4-1:0] node45597;
	wire [4-1:0] node45598;
	wire [4-1:0] node45601;
	wire [4-1:0] node45602;
	wire [4-1:0] node45606;
	wire [4-1:0] node45608;
	wire [4-1:0] node45611;
	wire [4-1:0] node45612;
	wire [4-1:0] node45614;
	wire [4-1:0] node45617;
	wire [4-1:0] node45618;
	wire [4-1:0] node45621;
	wire [4-1:0] node45624;
	wire [4-1:0] node45625;
	wire [4-1:0] node45626;
	wire [4-1:0] node45627;
	wire [4-1:0] node45630;
	wire [4-1:0] node45633;
	wire [4-1:0] node45634;
	wire [4-1:0] node45637;
	wire [4-1:0] node45640;
	wire [4-1:0] node45641;
	wire [4-1:0] node45644;
	wire [4-1:0] node45647;
	wire [4-1:0] node45648;
	wire [4-1:0] node45649;
	wire [4-1:0] node45650;
	wire [4-1:0] node45651;
	wire [4-1:0] node45654;
	wire [4-1:0] node45657;
	wire [4-1:0] node45658;
	wire [4-1:0] node45660;
	wire [4-1:0] node45663;
	wire [4-1:0] node45664;
	wire [4-1:0] node45667;
	wire [4-1:0] node45670;
	wire [4-1:0] node45671;
	wire [4-1:0] node45672;
	wire [4-1:0] node45674;
	wire [4-1:0] node45676;
	wire [4-1:0] node45679;
	wire [4-1:0] node45680;
	wire [4-1:0] node45683;
	wire [4-1:0] node45686;
	wire [4-1:0] node45687;
	wire [4-1:0] node45688;
	wire [4-1:0] node45691;
	wire [4-1:0] node45694;
	wire [4-1:0] node45695;
	wire [4-1:0] node45698;
	wire [4-1:0] node45701;
	wire [4-1:0] node45702;
	wire [4-1:0] node45703;
	wire [4-1:0] node45706;
	wire [4-1:0] node45709;
	wire [4-1:0] node45710;
	wire [4-1:0] node45713;
	wire [4-1:0] node45716;
	wire [4-1:0] node45717;
	wire [4-1:0] node45718;
	wire [4-1:0] node45719;
	wire [4-1:0] node45720;
	wire [4-1:0] node45721;
	wire [4-1:0] node45722;
	wire [4-1:0] node45723;
	wire [4-1:0] node45726;
	wire [4-1:0] node45729;
	wire [4-1:0] node45730;
	wire [4-1:0] node45731;
	wire [4-1:0] node45735;
	wire [4-1:0] node45736;
	wire [4-1:0] node45739;
	wire [4-1:0] node45742;
	wire [4-1:0] node45743;
	wire [4-1:0] node45744;
	wire [4-1:0] node45746;
	wire [4-1:0] node45749;
	wire [4-1:0] node45750;
	wire [4-1:0] node45753;
	wire [4-1:0] node45756;
	wire [4-1:0] node45757;
	wire [4-1:0] node45760;
	wire [4-1:0] node45763;
	wire [4-1:0] node45764;
	wire [4-1:0] node45765;
	wire [4-1:0] node45766;
	wire [4-1:0] node45769;
	wire [4-1:0] node45772;
	wire [4-1:0] node45773;
	wire [4-1:0] node45775;
	wire [4-1:0] node45776;
	wire [4-1:0] node45779;
	wire [4-1:0] node45782;
	wire [4-1:0] node45783;
	wire [4-1:0] node45786;
	wire [4-1:0] node45789;
	wire [4-1:0] node45791;
	wire [4-1:0] node45792;
	wire [4-1:0] node45793;
	wire [4-1:0] node45796;
	wire [4-1:0] node45799;
	wire [4-1:0] node45800;
	wire [4-1:0] node45804;
	wire [4-1:0] node45805;
	wire [4-1:0] node45806;
	wire [4-1:0] node45807;
	wire [4-1:0] node45808;
	wire [4-1:0] node45810;
	wire [4-1:0] node45813;
	wire [4-1:0] node45814;
	wire [4-1:0] node45817;
	wire [4-1:0] node45818;
	wire [4-1:0] node45822;
	wire [4-1:0] node45824;
	wire [4-1:0] node45825;
	wire [4-1:0] node45828;
	wire [4-1:0] node45831;
	wire [4-1:0] node45832;
	wire [4-1:0] node45833;
	wire [4-1:0] node45836;
	wire [4-1:0] node45839;
	wire [4-1:0] node45840;
	wire [4-1:0] node45841;
	wire [4-1:0] node45842;
	wire [4-1:0] node45845;
	wire [4-1:0] node45848;
	wire [4-1:0] node45849;
	wire [4-1:0] node45853;
	wire [4-1:0] node45854;
	wire [4-1:0] node45858;
	wire [4-1:0] node45859;
	wire [4-1:0] node45860;
	wire [4-1:0] node45861;
	wire [4-1:0] node45863;
	wire [4-1:0] node45867;
	wire [4-1:0] node45868;
	wire [4-1:0] node45870;
	wire [4-1:0] node45873;
	wire [4-1:0] node45875;
	wire [4-1:0] node45878;
	wire [4-1:0] node45879;
	wire [4-1:0] node45880;
	wire [4-1:0] node45883;
	wire [4-1:0] node45886;
	wire [4-1:0] node45887;
	wire [4-1:0] node45888;
	wire [4-1:0] node45889;
	wire [4-1:0] node45892;
	wire [4-1:0] node45896;
	wire [4-1:0] node45898;
	wire [4-1:0] node45901;
	wire [4-1:0] node45902;
	wire [4-1:0] node45903;
	wire [4-1:0] node45904;
	wire [4-1:0] node45905;
	wire [4-1:0] node45906;
	wire [4-1:0] node45909;
	wire [4-1:0] node45912;
	wire [4-1:0] node45913;
	wire [4-1:0] node45914;
	wire [4-1:0] node45917;
	wire [4-1:0] node45920;
	wire [4-1:0] node45922;
	wire [4-1:0] node45926;
	wire [4-1:0] node45927;
	wire [4-1:0] node45928;
	wire [4-1:0] node45929;
	wire [4-1:0] node45930;
	wire [4-1:0] node45931;
	wire [4-1:0] node45934;
	wire [4-1:0] node45938;
	wire [4-1:0] node45940;
	wire [4-1:0] node45941;
	wire [4-1:0] node45944;
	wire [4-1:0] node45947;
	wire [4-1:0] node45949;
	wire [4-1:0] node45950;
	wire [4-1:0] node45953;
	wire [4-1:0] node45957;
	wire [4-1:0] node45958;
	wire [4-1:0] node45959;
	wire [4-1:0] node45960;
	wire [4-1:0] node45961;
	wire [4-1:0] node45964;
	wire [4-1:0] node45967;
	wire [4-1:0] node45968;
	wire [4-1:0] node45969;
	wire [4-1:0] node45970;
	wire [4-1:0] node45973;
	wire [4-1:0] node45977;
	wire [4-1:0] node45978;
	wire [4-1:0] node45979;
	wire [4-1:0] node45982;
	wire [4-1:0] node45985;
	wire [4-1:0] node45986;
	wire [4-1:0] node45991;
	wire [4-1:0] node45992;
	wire [4-1:0] node45993;
	wire [4-1:0] node45996;
	wire [4-1:0] node46000;
	wire [4-1:0] node46001;
	wire [4-1:0] node46002;
	wire [4-1:0] node46003;
	wire [4-1:0] node46004;
	wire [4-1:0] node46005;
	wire [4-1:0] node46007;
	wire [4-1:0] node46010;
	wire [4-1:0] node46011;
	wire [4-1:0] node46014;
	wire [4-1:0] node46018;
	wire [4-1:0] node46019;
	wire [4-1:0] node46020;
	wire [4-1:0] node46021;
	wire [4-1:0] node46022;
	wire [4-1:0] node46026;
	wire [4-1:0] node46027;
	wire [4-1:0] node46031;
	wire [4-1:0] node46032;
	wire [4-1:0] node46033;
	wire [4-1:0] node46036;
	wire [4-1:0] node46041;
	wire [4-1:0] node46042;
	wire [4-1:0] node46043;
	wire [4-1:0] node46044;
	wire [4-1:0] node46047;
	wire [4-1:0] node46051;
	wire [4-1:0] node46052;
	wire [4-1:0] node46053;
	wire [4-1:0] node46056;
	wire [4-1:0] node46060;
	wire [4-1:0] node46061;
	wire [4-1:0] node46062;
	wire [4-1:0] node46063;
	wire [4-1:0] node46064;
	wire [4-1:0] node46065;
	wire [4-1:0] node46066;
	wire [4-1:0] node46069;
	wire [4-1:0] node46073;
	wire [4-1:0] node46074;
	wire [4-1:0] node46075;
	wire [4-1:0] node46078;
	wire [4-1:0] node46082;
	wire [4-1:0] node46083;
	wire [4-1:0] node46084;
	wire [4-1:0] node46085;
	wire [4-1:0] node46090;
	wire [4-1:0] node46091;
	wire [4-1:0] node46092;
	wire [4-1:0] node46095;
	wire [4-1:0] node46099;
	wire [4-1:0] node46100;
	wire [4-1:0] node46101;
	wire [4-1:0] node46102;
	wire [4-1:0] node46104;
	wire [4-1:0] node46107;
	wire [4-1:0] node46108;
	wire [4-1:0] node46112;
	wire [4-1:0] node46113;
	wire [4-1:0] node46115;
	wire [4-1:0] node46118;
	wire [4-1:0] node46119;
	wire [4-1:0] node46123;
	wire [4-1:0] node46124;
	wire [4-1:0] node46125;
	wire [4-1:0] node46126;
	wire [4-1:0] node46130;
	wire [4-1:0] node46131;
	wire [4-1:0] node46135;
	wire [4-1:0] node46136;
	wire [4-1:0] node46137;
	wire [4-1:0] node46141;
	wire [4-1:0] node46142;
	wire [4-1:0] node46146;
	wire [4-1:0] node46147;
	wire [4-1:0] node46148;
	wire [4-1:0] node46149;
	wire [4-1:0] node46150;
	wire [4-1:0] node46153;
	wire [4-1:0] node46156;
	wire [4-1:0] node46157;
	wire [4-1:0] node46158;
	wire [4-1:0] node46159;
	wire [4-1:0] node46162;
	wire [4-1:0] node46165;
	wire [4-1:0] node46166;
	wire [4-1:0] node46169;
	wire [4-1:0] node46172;
	wire [4-1:0] node46173;
	wire [4-1:0] node46174;
	wire [4-1:0] node46178;
	wire [4-1:0] node46179;
	wire [4-1:0] node46182;
	wire [4-1:0] node46185;
	wire [4-1:0] node46186;
	wire [4-1:0] node46187;
	wire [4-1:0] node46188;
	wire [4-1:0] node46189;
	wire [4-1:0] node46193;
	wire [4-1:0] node46194;
	wire [4-1:0] node46197;
	wire [4-1:0] node46200;
	wire [4-1:0] node46201;
	wire [4-1:0] node46202;
	wire [4-1:0] node46205;
	wire [4-1:0] node46208;
	wire [4-1:0] node46209;
	wire [4-1:0] node46212;
	wire [4-1:0] node46215;
	wire [4-1:0] node46216;
	wire [4-1:0] node46217;
	wire [4-1:0] node46220;
	wire [4-1:0] node46223;
	wire [4-1:0] node46224;
	wire [4-1:0] node46227;
	wire [4-1:0] node46230;
	wire [4-1:0] node46231;
	wire [4-1:0] node46232;
	wire [4-1:0] node46233;
	wire [4-1:0] node46234;
	wire [4-1:0] node46238;
	wire [4-1:0] node46239;
	wire [4-1:0] node46243;
	wire [4-1:0] node46244;
	wire [4-1:0] node46245;
	wire [4-1:0] node46246;
	wire [4-1:0] node46249;
	wire [4-1:0] node46254;
	wire [4-1:0] node46255;
	wire [4-1:0] node46256;
	wire [4-1:0] node46257;
	wire [4-1:0] node46261;
	wire [4-1:0] node46262;
	wire [4-1:0] node46266;
	wire [4-1:0] node46267;
	wire [4-1:0] node46268;
	wire [4-1:0] node46272;
	wire [4-1:0] node46273;
	wire [4-1:0] node46277;
	wire [4-1:0] node46278;
	wire [4-1:0] node46279;
	wire [4-1:0] node46280;
	wire [4-1:0] node46281;
	wire [4-1:0] node46282;
	wire [4-1:0] node46283;
	wire [4-1:0] node46284;
	wire [4-1:0] node46285;
	wire [4-1:0] node46288;
	wire [4-1:0] node46291;
	wire [4-1:0] node46292;
	wire [4-1:0] node46295;
	wire [4-1:0] node46298;
	wire [4-1:0] node46299;
	wire [4-1:0] node46300;
	wire [4-1:0] node46301;
	wire [4-1:0] node46304;
	wire [4-1:0] node46307;
	wire [4-1:0] node46308;
	wire [4-1:0] node46311;
	wire [4-1:0] node46314;
	wire [4-1:0] node46315;
	wire [4-1:0] node46316;
	wire [4-1:0] node46318;
	wire [4-1:0] node46321;
	wire [4-1:0] node46322;
	wire [4-1:0] node46325;
	wire [4-1:0] node46328;
	wire [4-1:0] node46329;
	wire [4-1:0] node46330;
	wire [4-1:0] node46333;
	wire [4-1:0] node46337;
	wire [4-1:0] node46338;
	wire [4-1:0] node46339;
	wire [4-1:0] node46340;
	wire [4-1:0] node46343;
	wire [4-1:0] node46346;
	wire [4-1:0] node46347;
	wire [4-1:0] node46348;
	wire [4-1:0] node46349;
	wire [4-1:0] node46352;
	wire [4-1:0] node46356;
	wire [4-1:0] node46357;
	wire [4-1:0] node46359;
	wire [4-1:0] node46362;
	wire [4-1:0] node46363;
	wire [4-1:0] node46367;
	wire [4-1:0] node46368;
	wire [4-1:0] node46369;
	wire [4-1:0] node46371;
	wire [4-1:0] node46372;
	wire [4-1:0] node46375;
	wire [4-1:0] node46378;
	wire [4-1:0] node46379;
	wire [4-1:0] node46382;
	wire [4-1:0] node46385;
	wire [4-1:0] node46386;
	wire [4-1:0] node46388;
	wire [4-1:0] node46391;
	wire [4-1:0] node46392;
	wire [4-1:0] node46395;
	wire [4-1:0] node46398;
	wire [4-1:0] node46399;
	wire [4-1:0] node46400;
	wire [4-1:0] node46403;
	wire [4-1:0] node46406;
	wire [4-1:0] node46407;
	wire [4-1:0] node46408;
	wire [4-1:0] node46409;
	wire [4-1:0] node46412;
	wire [4-1:0] node46415;
	wire [4-1:0] node46416;
	wire [4-1:0] node46417;
	wire [4-1:0] node46420;
	wire [4-1:0] node46423;
	wire [4-1:0] node46424;
	wire [4-1:0] node46427;
	wire [4-1:0] node46430;
	wire [4-1:0] node46431;
	wire [4-1:0] node46432;
	wire [4-1:0] node46433;
	wire [4-1:0] node46436;
	wire [4-1:0] node46439;
	wire [4-1:0] node46440;
	wire [4-1:0] node46443;
	wire [4-1:0] node46446;
	wire [4-1:0] node46447;
	wire [4-1:0] node46448;
	wire [4-1:0] node46451;
	wire [4-1:0] node46454;
	wire [4-1:0] node46455;
	wire [4-1:0] node46456;
	wire [4-1:0] node46459;
	wire [4-1:0] node46462;
	wire [4-1:0] node46463;
	wire [4-1:0] node46467;
	wire [4-1:0] node46468;
	wire [4-1:0] node46471;
	wire [4-1:0] node46474;
	wire [4-1:0] node46475;
	wire [4-1:0] node46476;
	wire [4-1:0] node46477;
	wire [4-1:0] node46478;
	wire [4-1:0] node46479;
	wire [4-1:0] node46480;
	wire [4-1:0] node46481;
	wire [4-1:0] node46485;
	wire [4-1:0] node46486;
	wire [4-1:0] node46487;
	wire [4-1:0] node46491;
	wire [4-1:0] node46492;
	wire [4-1:0] node46495;
	wire [4-1:0] node46498;
	wire [4-1:0] node46499;
	wire [4-1:0] node46500;
	wire [4-1:0] node46503;
	wire [4-1:0] node46506;
	wire [4-1:0] node46507;
	wire [4-1:0] node46508;
	wire [4-1:0] node46513;
	wire [4-1:0] node46514;
	wire [4-1:0] node46515;
	wire [4-1:0] node46516;
	wire [4-1:0] node46519;
	wire [4-1:0] node46522;
	wire [4-1:0] node46523;
	wire [4-1:0] node46524;
	wire [4-1:0] node46527;
	wire [4-1:0] node46530;
	wire [4-1:0] node46531;
	wire [4-1:0] node46534;
	wire [4-1:0] node46537;
	wire [4-1:0] node46538;
	wire [4-1:0] node46540;
	wire [4-1:0] node46543;
	wire [4-1:0] node46544;
	wire [4-1:0] node46545;
	wire [4-1:0] node46548;
	wire [4-1:0] node46551;
	wire [4-1:0] node46552;
	wire [4-1:0] node46555;
	wire [4-1:0] node46559;
	wire [4-1:0] node46560;
	wire [4-1:0] node46561;
	wire [4-1:0] node46562;
	wire [4-1:0] node46563;
	wire [4-1:0] node46564;
	wire [4-1:0] node46567;
	wire [4-1:0] node46570;
	wire [4-1:0] node46571;
	wire [4-1:0] node46574;
	wire [4-1:0] node46577;
	wire [4-1:0] node46578;
	wire [4-1:0] node46579;
	wire [4-1:0] node46582;
	wire [4-1:0] node46585;
	wire [4-1:0] node46586;
	wire [4-1:0] node46589;
	wire [4-1:0] node46592;
	wire [4-1:0] node46593;
	wire [4-1:0] node46596;
	wire [4-1:0] node46600;
	wire [4-1:0] node46601;
	wire [4-1:0] node46602;
	wire [4-1:0] node46606;
	wire [4-1:0] node46607;
	wire [4-1:0] node46611;
	wire [4-1:0] node46612;
	wire [4-1:0] node46613;
	wire [4-1:0] node46614;
	wire [4-1:0] node46615;
	wire [4-1:0] node46616;
	wire [4-1:0] node46619;
	wire [4-1:0] node46622;
	wire [4-1:0] node46623;
	wire [4-1:0] node46626;
	wire [4-1:0] node46629;
	wire [4-1:0] node46630;
	wire [4-1:0] node46631;
	wire [4-1:0] node46632;
	wire [4-1:0] node46635;
	wire [4-1:0] node46638;
	wire [4-1:0] node46639;
	wire [4-1:0] node46640;
	wire [4-1:0] node46643;
	wire [4-1:0] node46646;
	wire [4-1:0] node46647;
	wire [4-1:0] node46650;
	wire [4-1:0] node46653;
	wire [4-1:0] node46654;
	wire [4-1:0] node46655;
	wire [4-1:0] node46656;
	wire [4-1:0] node46657;
	wire [4-1:0] node46660;
	wire [4-1:0] node46663;
	wire [4-1:0] node46664;
	wire [4-1:0] node46667;
	wire [4-1:0] node46670;
	wire [4-1:0] node46671;
	wire [4-1:0] node46674;
	wire [4-1:0] node46677;
	wire [4-1:0] node46678;
	wire [4-1:0] node46679;
	wire [4-1:0] node46680;
	wire [4-1:0] node46683;
	wire [4-1:0] node46686;
	wire [4-1:0] node46687;
	wire [4-1:0] node46689;
	wire [4-1:0] node46692;
	wire [4-1:0] node46693;
	wire [4-1:0] node46696;
	wire [4-1:0] node46699;
	wire [4-1:0] node46701;
	wire [4-1:0] node46704;
	wire [4-1:0] node46705;
	wire [4-1:0] node46706;
	wire [4-1:0] node46709;
	wire [4-1:0] node46712;
	wire [4-1:0] node46713;
	wire [4-1:0] node46714;
	wire [4-1:0] node46717;
	wire [4-1:0] node46720;
	wire [4-1:0] node46721;
	wire [4-1:0] node46722;
	wire [4-1:0] node46723;
	wire [4-1:0] node46724;
	wire [4-1:0] node46725;
	wire [4-1:0] node46729;
	wire [4-1:0] node46730;
	wire [4-1:0] node46734;
	wire [4-1:0] node46735;
	wire [4-1:0] node46736;
	wire [4-1:0] node46739;
	wire [4-1:0] node46742;
	wire [4-1:0] node46743;
	wire [4-1:0] node46746;
	wire [4-1:0] node46749;
	wire [4-1:0] node46750;
	wire [4-1:0] node46751;
	wire [4-1:0] node46754;
	wire [4-1:0] node46757;
	wire [4-1:0] node46758;
	wire [4-1:0] node46761;
	wire [4-1:0] node46764;
	wire [4-1:0] node46765;
	wire [4-1:0] node46768;
	wire [4-1:0] node46771;
	wire [4-1:0] node46772;
	wire [4-1:0] node46773;
	wire [4-1:0] node46777;
	wire [4-1:0] node46778;
	wire [4-1:0] node46782;
	wire [4-1:0] node46783;
	wire [4-1:0] node46784;
	wire [4-1:0] node46785;
	wire [4-1:0] node46786;
	wire [4-1:0] node46787;
	wire [4-1:0] node46788;
	wire [4-1:0] node46789;
	wire [4-1:0] node46790;
	wire [4-1:0] node46791;
	wire [4-1:0] node46795;
	wire [4-1:0] node46796;
	wire [4-1:0] node46800;
	wire [4-1:0] node46801;
	wire [4-1:0] node46802;
	wire [4-1:0] node46806;
	wire [4-1:0] node46807;
	wire [4-1:0] node46811;
	wire [4-1:0] node46812;
	wire [4-1:0] node46813;
	wire [4-1:0] node46816;
	wire [4-1:0] node46819;
	wire [4-1:0] node46820;
	wire [4-1:0] node46821;
	wire [4-1:0] node46822;
	wire [4-1:0] node46825;
	wire [4-1:0] node46828;
	wire [4-1:0] node46829;
	wire [4-1:0] node46832;
	wire [4-1:0] node46835;
	wire [4-1:0] node46837;
	wire [4-1:0] node46838;
	wire [4-1:0] node46841;
	wire [4-1:0] node46844;
	wire [4-1:0] node46845;
	wire [4-1:0] node46846;
	wire [4-1:0] node46847;
	wire [4-1:0] node46849;
	wire [4-1:0] node46850;
	wire [4-1:0] node46853;
	wire [4-1:0] node46856;
	wire [4-1:0] node46857;
	wire [4-1:0] node46860;
	wire [4-1:0] node46863;
	wire [4-1:0] node46864;
	wire [4-1:0] node46865;
	wire [4-1:0] node46867;
	wire [4-1:0] node46868;
	wire [4-1:0] node46872;
	wire [4-1:0] node46873;
	wire [4-1:0] node46876;
	wire [4-1:0] node46879;
	wire [4-1:0] node46880;
	wire [4-1:0] node46881;
	wire [4-1:0] node46883;
	wire [4-1:0] node46886;
	wire [4-1:0] node46887;
	wire [4-1:0] node46890;
	wire [4-1:0] node46893;
	wire [4-1:0] node46895;
	wire [4-1:0] node46896;
	wire [4-1:0] node46899;
	wire [4-1:0] node46902;
	wire [4-1:0] node46903;
	wire [4-1:0] node46904;
	wire [4-1:0] node46905;
	wire [4-1:0] node46906;
	wire [4-1:0] node46907;
	wire [4-1:0] node46910;
	wire [4-1:0] node46913;
	wire [4-1:0] node46914;
	wire [4-1:0] node46918;
	wire [4-1:0] node46919;
	wire [4-1:0] node46920;
	wire [4-1:0] node46923;
	wire [4-1:0] node46926;
	wire [4-1:0] node46928;
	wire [4-1:0] node46931;
	wire [4-1:0] node46932;
	wire [4-1:0] node46933;
	wire [4-1:0] node46936;
	wire [4-1:0] node46939;
	wire [4-1:0] node46940;
	wire [4-1:0] node46941;
	wire [4-1:0] node46945;
	wire [4-1:0] node46946;
	wire [4-1:0] node46949;
	wire [4-1:0] node46952;
	wire [4-1:0] node46953;
	wire [4-1:0] node46954;
	wire [4-1:0] node46958;
	wire [4-1:0] node46959;
	wire [4-1:0] node46961;
	wire [4-1:0] node46962;
	wire [4-1:0] node46965;
	wire [4-1:0] node46968;
	wire [4-1:0] node46969;
	wire [4-1:0] node46972;
	wire [4-1:0] node46975;
	wire [4-1:0] node46976;
	wire [4-1:0] node46977;
	wire [4-1:0] node46978;
	wire [4-1:0] node46979;
	wire [4-1:0] node46980;
	wire [4-1:0] node46981;
	wire [4-1:0] node46985;
	wire [4-1:0] node46988;
	wire [4-1:0] node46989;
	wire [4-1:0] node46990;
	wire [4-1:0] node46994;
	wire [4-1:0] node46995;
	wire [4-1:0] node46999;
	wire [4-1:0] node47000;
	wire [4-1:0] node47001;
	wire [4-1:0] node47002;
	wire [4-1:0] node47003;
	wire [4-1:0] node47006;
	wire [4-1:0] node47009;
	wire [4-1:0] node47010;
	wire [4-1:0] node47013;
	wire [4-1:0] node47016;
	wire [4-1:0] node47017;
	wire [4-1:0] node47021;
	wire [4-1:0] node47022;
	wire [4-1:0] node47023;
	wire [4-1:0] node47026;
	wire [4-1:0] node47029;
	wire [4-1:0] node47030;
	wire [4-1:0] node47033;
	wire [4-1:0] node47036;
	wire [4-1:0] node47037;
	wire [4-1:0] node47038;
	wire [4-1:0] node47039;
	wire [4-1:0] node47043;
	wire [4-1:0] node47044;
	wire [4-1:0] node47045;
	wire [4-1:0] node47049;
	wire [4-1:0] node47050;
	wire [4-1:0] node47054;
	wire [4-1:0] node47055;
	wire [4-1:0] node47056;
	wire [4-1:0] node47057;
	wire [4-1:0] node47060;
	wire [4-1:0] node47063;
	wire [4-1:0] node47064;
	wire [4-1:0] node47065;
	wire [4-1:0] node47068;
	wire [4-1:0] node47071;
	wire [4-1:0] node47072;
	wire [4-1:0] node47075;
	wire [4-1:0] node47078;
	wire [4-1:0] node47079;
	wire [4-1:0] node47082;
	wire [4-1:0] node47085;
	wire [4-1:0] node47086;
	wire [4-1:0] node47087;
	wire [4-1:0] node47088;
	wire [4-1:0] node47089;
	wire [4-1:0] node47090;
	wire [4-1:0] node47092;
	wire [4-1:0] node47095;
	wire [4-1:0] node47096;
	wire [4-1:0] node47100;
	wire [4-1:0] node47101;
	wire [4-1:0] node47104;
	wire [4-1:0] node47107;
	wire [4-1:0] node47108;
	wire [4-1:0] node47111;
	wire [4-1:0] node47114;
	wire [4-1:0] node47115;
	wire [4-1:0] node47116;
	wire [4-1:0] node47117;
	wire [4-1:0] node47118;
	wire [4-1:0] node47122;
	wire [4-1:0] node47123;
	wire [4-1:0] node47127;
	wire [4-1:0] node47129;
	wire [4-1:0] node47130;
	wire [4-1:0] node47134;
	wire [4-1:0] node47135;
	wire [4-1:0] node47136;
	wire [4-1:0] node47137;
	wire [4-1:0] node47142;
	wire [4-1:0] node47143;
	wire [4-1:0] node47144;
	wire [4-1:0] node47149;
	wire [4-1:0] node47150;
	wire [4-1:0] node47151;
	wire [4-1:0] node47152;
	wire [4-1:0] node47156;
	wire [4-1:0] node47157;
	wire [4-1:0] node47161;
	wire [4-1:0] node47162;
	wire [4-1:0] node47163;
	wire [4-1:0] node47167;
	wire [4-1:0] node47168;
	wire [4-1:0] node47172;
	wire [4-1:0] node47173;
	wire [4-1:0] node47174;
	wire [4-1:0] node47175;
	wire [4-1:0] node47177;
	wire [4-1:0] node47180;
	wire [4-1:0] node47182;
	wire [4-1:0] node47185;
	wire [4-1:0] node47186;
	wire [4-1:0] node47188;
	wire [4-1:0] node47191;
	wire [4-1:0] node47193;
	wire [4-1:0] node47196;
	wire [4-1:0] node47197;
	wire [4-1:0] node47198;
	wire [4-1:0] node47199;
	wire [4-1:0] node47200;
	wire [4-1:0] node47201;
	wire [4-1:0] node47202;
	wire [4-1:0] node47205;
	wire [4-1:0] node47207;
	wire [4-1:0] node47210;
	wire [4-1:0] node47211;
	wire [4-1:0] node47213;
	wire [4-1:0] node47216;
	wire [4-1:0] node47218;
	wire [4-1:0] node47221;
	wire [4-1:0] node47222;
	wire [4-1:0] node47223;
	wire [4-1:0] node47226;
	wire [4-1:0] node47229;
	wire [4-1:0] node47231;
	wire [4-1:0] node47234;
	wire [4-1:0] node47235;
	wire [4-1:0] node47236;
	wire [4-1:0] node47239;
	wire [4-1:0] node47242;
	wire [4-1:0] node47243;
	wire [4-1:0] node47246;
	wire [4-1:0] node47249;
	wire [4-1:0] node47250;
	wire [4-1:0] node47253;
	wire [4-1:0] node47256;
	wire [4-1:0] node47257;
	wire [4-1:0] node47258;
	wire [4-1:0] node47259;
	wire [4-1:0] node47263;
	wire [4-1:0] node47264;
	wire [4-1:0] node47268;
	wire [4-1:0] node47269;
	wire [4-1:0] node47270;
	wire [4-1:0] node47274;
	wire [4-1:0] node47275;
	wire [4-1:0] node47279;
	wire [4-1:0] node47280;
	wire [4-1:0] node47281;
	wire [4-1:0] node47282;
	wire [4-1:0] node47283;
	wire [4-1:0] node47284;
	wire [4-1:0] node47285;
	wire [4-1:0] node47286;
	wire [4-1:0] node47287;
	wire [4-1:0] node47292;
	wire [4-1:0] node47293;
	wire [4-1:0] node47294;
	wire [4-1:0] node47298;
	wire [4-1:0] node47299;
	wire [4-1:0] node47303;
	wire [4-1:0] node47304;
	wire [4-1:0] node47305;
	wire [4-1:0] node47306;
	wire [4-1:0] node47310;
	wire [4-1:0] node47311;
	wire [4-1:0] node47315;
	wire [4-1:0] node47316;
	wire [4-1:0] node47319;
	wire [4-1:0] node47320;
	wire [4-1:0] node47324;
	wire [4-1:0] node47325;
	wire [4-1:0] node47326;
	wire [4-1:0] node47327;
	wire [4-1:0] node47328;
	wire [4-1:0] node47332;
	wire [4-1:0] node47333;
	wire [4-1:0] node47337;
	wire [4-1:0] node47338;
	wire [4-1:0] node47339;
	wire [4-1:0] node47344;
	wire [4-1:0] node47345;
	wire [4-1:0] node47346;
	wire [4-1:0] node47347;
	wire [4-1:0] node47348;
	wire [4-1:0] node47353;
	wire [4-1:0] node47356;
	wire [4-1:0] node47357;
	wire [4-1:0] node47358;
	wire [4-1:0] node47360;
	wire [4-1:0] node47363;
	wire [4-1:0] node47364;
	wire [4-1:0] node47367;
	wire [4-1:0] node47370;
	wire [4-1:0] node47371;
	wire [4-1:0] node47374;
	wire [4-1:0] node47377;
	wire [4-1:0] node47378;
	wire [4-1:0] node47379;
	wire [4-1:0] node47380;
	wire [4-1:0] node47381;
	wire [4-1:0] node47382;
	wire [4-1:0] node47386;
	wire [4-1:0] node47387;
	wire [4-1:0] node47391;
	wire [4-1:0] node47392;
	wire [4-1:0] node47393;
	wire [4-1:0] node47397;
	wire [4-1:0] node47398;
	wire [4-1:0] node47402;
	wire [4-1:0] node47403;
	wire [4-1:0] node47404;
	wire [4-1:0] node47405;
	wire [4-1:0] node47406;
	wire [4-1:0] node47410;
	wire [4-1:0] node47411;
	wire [4-1:0] node47415;
	wire [4-1:0] node47416;
	wire [4-1:0] node47419;
	wire [4-1:0] node47420;
	wire [4-1:0] node47424;
	wire [4-1:0] node47425;
	wire [4-1:0] node47426;
	wire [4-1:0] node47427;
	wire [4-1:0] node47431;
	wire [4-1:0] node47432;
	wire [4-1:0] node47436;
	wire [4-1:0] node47437;
	wire [4-1:0] node47440;
	wire [4-1:0] node47441;
	wire [4-1:0] node47445;
	wire [4-1:0] node47446;
	wire [4-1:0] node47447;
	wire [4-1:0] node47448;
	wire [4-1:0] node47451;
	wire [4-1:0] node47454;
	wire [4-1:0] node47455;
	wire [4-1:0] node47456;
	wire [4-1:0] node47459;
	wire [4-1:0] node47462;
	wire [4-1:0] node47463;
	wire [4-1:0] node47466;
	wire [4-1:0] node47469;
	wire [4-1:0] node47470;
	wire [4-1:0] node47471;
	wire [4-1:0] node47474;
	wire [4-1:0] node47477;
	wire [4-1:0] node47478;
	wire [4-1:0] node47479;
	wire [4-1:0] node47482;
	wire [4-1:0] node47485;
	wire [4-1:0] node47486;
	wire [4-1:0] node47487;
	wire [4-1:0] node47490;
	wire [4-1:0] node47493;
	wire [4-1:0] node47494;
	wire [4-1:0] node47497;
	wire [4-1:0] node47500;
	wire [4-1:0] node47501;
	wire [4-1:0] node47502;
	wire [4-1:0] node47503;
	wire [4-1:0] node47504;
	wire [4-1:0] node47507;
	wire [4-1:0] node47510;
	wire [4-1:0] node47511;
	wire [4-1:0] node47512;
	wire [4-1:0] node47514;
	wire [4-1:0] node47517;
	wire [4-1:0] node47518;
	wire [4-1:0] node47519;
	wire [4-1:0] node47522;
	wire [4-1:0] node47526;
	wire [4-1:0] node47527;
	wire [4-1:0] node47528;
	wire [4-1:0] node47532;
	wire [4-1:0] node47533;
	wire [4-1:0] node47536;
	wire [4-1:0] node47539;
	wire [4-1:0] node47540;
	wire [4-1:0] node47541;
	wire [4-1:0] node47542;
	wire [4-1:0] node47543;
	wire [4-1:0] node47544;
	wire [4-1:0] node47547;
	wire [4-1:0] node47550;
	wire [4-1:0] node47551;
	wire [4-1:0] node47555;
	wire [4-1:0] node47556;
	wire [4-1:0] node47557;
	wire [4-1:0] node47560;
	wire [4-1:0] node47563;
	wire [4-1:0] node47564;
	wire [4-1:0] node47567;
	wire [4-1:0] node47570;
	wire [4-1:0] node47571;
	wire [4-1:0] node47572;
	wire [4-1:0] node47574;
	wire [4-1:0] node47577;
	wire [4-1:0] node47578;
	wire [4-1:0] node47581;
	wire [4-1:0] node47584;
	wire [4-1:0] node47585;
	wire [4-1:0] node47588;
	wire [4-1:0] node47591;
	wire [4-1:0] node47592;
	wire [4-1:0] node47593;
	wire [4-1:0] node47594;
	wire [4-1:0] node47595;
	wire [4-1:0] node47600;
	wire [4-1:0] node47601;
	wire [4-1:0] node47605;
	wire [4-1:0] node47606;
	wire [4-1:0] node47607;
	wire [4-1:0] node47608;
	wire [4-1:0] node47611;
	wire [4-1:0] node47615;
	wire [4-1:0] node47616;
	wire [4-1:0] node47617;
	wire [4-1:0] node47621;
	wire [4-1:0] node47622;
	wire [4-1:0] node47626;
	wire [4-1:0] node47627;
	wire [4-1:0] node47628;
	wire [4-1:0] node47629;
	wire [4-1:0] node47630;
	wire [4-1:0] node47631;
	wire [4-1:0] node47633;
	wire [4-1:0] node47636;
	wire [4-1:0] node47637;
	wire [4-1:0] node47640;
	wire [4-1:0] node47643;
	wire [4-1:0] node47644;
	wire [4-1:0] node47645;
	wire [4-1:0] node47648;
	wire [4-1:0] node47651;
	wire [4-1:0] node47652;
	wire [4-1:0] node47655;
	wire [4-1:0] node47658;
	wire [4-1:0] node47659;
	wire [4-1:0] node47662;
	wire [4-1:0] node47665;
	wire [4-1:0] node47666;
	wire [4-1:0] node47667;
	wire [4-1:0] node47669;
	wire [4-1:0] node47670;
	wire [4-1:0] node47673;
	wire [4-1:0] node47676;
	wire [4-1:0] node47677;
	wire [4-1:0] node47679;
	wire [4-1:0] node47682;
	wire [4-1:0] node47685;
	wire [4-1:0] node47686;
	wire [4-1:0] node47687;
	wire [4-1:0] node47689;
	wire [4-1:0] node47692;
	wire [4-1:0] node47693;
	wire [4-1:0] node47696;
	wire [4-1:0] node47699;
	wire [4-1:0] node47700;
	wire [4-1:0] node47704;
	wire [4-1:0] node47705;
	wire [4-1:0] node47706;
	wire [4-1:0] node47707;
	wire [4-1:0] node47711;
	wire [4-1:0] node47712;
	wire [4-1:0] node47716;
	wire [4-1:0] node47717;
	wire [4-1:0] node47718;
	wire [4-1:0] node47722;
	wire [4-1:0] node47723;
	wire [4-1:0] node47727;
	wire [4-1:0] node47728;
	wire [4-1:0] node47729;
	wire [4-1:0] node47730;
	wire [4-1:0] node47731;
	wire [4-1:0] node47735;
	wire [4-1:0] node47736;
	wire [4-1:0] node47741;
	wire [4-1:0] node47742;
	wire [4-1:0] node47743;
	wire [4-1:0] node47744;
	wire [4-1:0] node47748;
	wire [4-1:0] node47749;
	wire [4-1:0] node47754;
	wire [4-1:0] node47755;
	wire [4-1:0] node47756;
	wire [4-1:0] node47757;
	wire [4-1:0] node47758;
	wire [4-1:0] node47759;
	wire [4-1:0] node47760;
	wire [4-1:0] node47761;
	wire [4-1:0] node47764;
	wire [4-1:0] node47767;
	wire [4-1:0] node47768;
	wire [4-1:0] node47769;
	wire [4-1:0] node47772;
	wire [4-1:0] node47775;
	wire [4-1:0] node47776;
	wire [4-1:0] node47779;
	wire [4-1:0] node47783;
	wire [4-1:0] node47784;
	wire [4-1:0] node47788;
	wire [4-1:0] node47789;
	wire [4-1:0] node47790;
	wire [4-1:0] node47791;
	wire [4-1:0] node47792;
	wire [4-1:0] node47795;
	wire [4-1:0] node47798;
	wire [4-1:0] node47799;
	wire [4-1:0] node47800;
	wire [4-1:0] node47803;
	wire [4-1:0] node47806;
	wire [4-1:0] node47807;
	wire [4-1:0] node47810;
	wire [4-1:0] node47814;
	wire [4-1:0] node47815;
	wire [4-1:0] node47819;
	wire [4-1:0] node47820;
	wire [4-1:0] node47821;
	wire [4-1:0] node47825;
	wire [4-1:0] node47826;
	wire [4-1:0] node47830;
	wire [4-1:0] node47831;
	wire [4-1:0] node47832;
	wire [4-1:0] node47833;
	wire [4-1:0] node47834;
	wire [4-1:0] node47835;
	wire [4-1:0] node47839;
	wire [4-1:0] node47840;
	wire [4-1:0] node47845;
	wire [4-1:0] node47846;
	wire [4-1:0] node47850;
	wire [4-1:0] node47851;
	wire [4-1:0] node47852;
	wire [4-1:0] node47853;
	wire [4-1:0] node47854;
	wire [4-1:0] node47859;
	wire [4-1:0] node47860;
	wire [4-1:0] node47861;

	assign outp = (inp[3]) ? node26504 : node1;
		assign node1 = (inp[6]) ? node16561 : node2;
			assign node2 = (inp[8]) ? node9624 : node3;
				assign node3 = (inp[14]) ? node4739 : node4;
					assign node4 = (inp[12]) ? node2204 : node5;
						assign node5 = (inp[7]) ? node1217 : node6;
							assign node6 = (inp[4]) ? node584 : node7;
								assign node7 = (inp[15]) ? node303 : node8;
									assign node8 = (inp[0]) ? node142 : node9;
										assign node9 = (inp[2]) ? node73 : node10;
											assign node10 = (inp[13]) ? node40 : node11;
												assign node11 = (inp[1]) ? node29 : node12;
													assign node12 = (inp[5]) ? node22 : node13;
														assign node13 = (inp[11]) ? node15 : 4'b0001;
															assign node15 = (inp[9]) ? node19 : node16;
																assign node16 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node19 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node22 = (inp[10]) ? node26 : node23;
															assign node23 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node26 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node29 = (inp[5]) ? node35 : node30;
														assign node30 = (inp[10]) ? node32 : 4'b0000;
															assign node32 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node35 = (inp[9]) ? 4'b0101 : node36;
															assign node36 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node40 = (inp[5]) ? node62 : node41;
													assign node41 = (inp[1]) ? node49 : node42;
														assign node42 = (inp[9]) ? node46 : node43;
															assign node43 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node46 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node49 = (inp[11]) ? node57 : node50;
															assign node50 = (inp[9]) ? node54 : node51;
																assign node51 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node54 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node57 = (inp[9]) ? node59 : 4'b0100;
																assign node59 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node62 = (inp[1]) ? node70 : node63;
														assign node63 = (inp[9]) ? node67 : node64;
															assign node64 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node67 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node70 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node73 = (inp[13]) ? node105 : node74;
												assign node74 = (inp[5]) ? node80 : node75;
													assign node75 = (inp[10]) ? 4'b0100 : node76;
														assign node76 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node80 = (inp[1]) ? node92 : node81;
														assign node81 = (inp[11]) ? node87 : node82;
															assign node82 = (inp[9]) ? node84 : 4'b0101;
																assign node84 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node87 = (inp[9]) ? 4'b0100 : node88;
																assign node88 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node92 = (inp[9]) ? node98 : node93;
															assign node93 = (inp[10]) ? 4'b0001 : node94;
																assign node94 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node98 = (inp[11]) ? node102 : node99;
																assign node99 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node102 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node105 = (inp[1]) ? node123 : node106;
													assign node106 = (inp[11]) ? node116 : node107;
														assign node107 = (inp[5]) ? node109 : 4'b0000;
															assign node109 = (inp[10]) ? node113 : node110;
																assign node110 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node113 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node116 = (inp[10]) ? node120 : node117;
															assign node117 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node120 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node123 = (inp[5]) ? node133 : node124;
														assign node124 = (inp[9]) ? 4'b0000 : node125;
															assign node125 = (inp[11]) ? node129 : node126;
																assign node126 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node129 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node133 = (inp[11]) ? node135 : 4'b0100;
															assign node135 = (inp[10]) ? node139 : node136;
																assign node136 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node139 = (inp[9]) ? 4'b0101 : 4'b0100;
										assign node142 = (inp[10]) ? node224 : node143;
											assign node143 = (inp[9]) ? node189 : node144;
												assign node144 = (inp[11]) ? node168 : node145;
													assign node145 = (inp[13]) ? node157 : node146;
														assign node146 = (inp[2]) ? node152 : node147;
															assign node147 = (inp[1]) ? node149 : 4'b0000;
																assign node149 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node152 = (inp[1]) ? node154 : 4'b0100;
																assign node154 = (inp[5]) ? 4'b0001 : 4'b0100;
														assign node157 = (inp[2]) ? node163 : node158;
															assign node158 = (inp[1]) ? node160 : 4'b0100;
																assign node160 = (inp[5]) ? 4'b0001 : 4'b0100;
															assign node163 = (inp[5]) ? node165 : 4'b0001;
																assign node165 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node168 = (inp[1]) ? node180 : node169;
														assign node169 = (inp[5]) ? node175 : node170;
															assign node170 = (inp[2]) ? node172 : 4'b0101;
																assign node172 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node175 = (inp[2]) ? 4'b0001 : node176;
																assign node176 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node180 = (inp[2]) ? node182 : 4'b0001;
															assign node182 = (inp[13]) ? node186 : node183;
																assign node183 = (inp[5]) ? 4'b0001 : 4'b0101;
																assign node186 = (inp[5]) ? 4'b0101 : 4'b0001;
												assign node189 = (inp[11]) ? node207 : node190;
													assign node190 = (inp[13]) ? node198 : node191;
														assign node191 = (inp[2]) ? 4'b0101 : node192;
															assign node192 = (inp[5]) ? node194 : 4'b0001;
																assign node194 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node198 = (inp[2]) ? node202 : node199;
															assign node199 = (inp[5]) ? 4'b0000 : 4'b0101;
															assign node202 = (inp[5]) ? node204 : 4'b0000;
																assign node204 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node207 = (inp[1]) ? node215 : node208;
														assign node208 = (inp[13]) ? node212 : node209;
															assign node209 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node212 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node215 = (inp[2]) ? node217 : 4'b0000;
															assign node217 = (inp[13]) ? node221 : node218;
																assign node218 = (inp[5]) ? 4'b0000 : 4'b0100;
																assign node221 = (inp[5]) ? 4'b0100 : 4'b0000;
											assign node224 = (inp[9]) ? node266 : node225;
												assign node225 = (inp[11]) ? node245 : node226;
													assign node226 = (inp[2]) ? node238 : node227;
														assign node227 = (inp[13]) ? node233 : node228;
															assign node228 = (inp[5]) ? node230 : 4'b0001;
																assign node230 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node233 = (inp[5]) ? node235 : 4'b0101;
																assign node235 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node238 = (inp[13]) ? node242 : node239;
															assign node239 = (inp[5]) ? 4'b0000 : 4'b0101;
															assign node242 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node245 = (inp[2]) ? node257 : node246;
														assign node246 = (inp[13]) ? node252 : node247;
															assign node247 = (inp[1]) ? node249 : 4'b0000;
																assign node249 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node252 = (inp[5]) ? node254 : 4'b0100;
																assign node254 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node257 = (inp[13]) ? node263 : node258;
															assign node258 = (inp[5]) ? node260 : 4'b0100;
																assign node260 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node263 = (inp[5]) ? 4'b0100 : 4'b0000;
												assign node266 = (inp[11]) ? node282 : node267;
													assign node267 = (inp[2]) ? node273 : node268;
														assign node268 = (inp[13]) ? 4'b0100 : node269;
															assign node269 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node273 = (inp[13]) ? node279 : node274;
															assign node274 = (inp[5]) ? node276 : 4'b0100;
																assign node276 = (inp[1]) ? 4'b0001 : 4'b0100;
															assign node279 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node282 = (inp[13]) ? node292 : node283;
														assign node283 = (inp[2]) ? node287 : node284;
															assign node284 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node287 = (inp[5]) ? node289 : 4'b0101;
																assign node289 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node292 = (inp[2]) ? node298 : node293;
															assign node293 = (inp[5]) ? node295 : 4'b0101;
																assign node295 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node298 = (inp[1]) ? node300 : 4'b0001;
																assign node300 = (inp[5]) ? 4'b0101 : 4'b0001;
									assign node303 = (inp[13]) ? node439 : node304;
										assign node304 = (inp[2]) ? node374 : node305;
											assign node305 = (inp[1]) ? node329 : node306;
												assign node306 = (inp[9]) ? node318 : node307;
													assign node307 = (inp[10]) ? node313 : node308;
														assign node308 = (inp[11]) ? node310 : 4'b0000;
															assign node310 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node313 = (inp[0]) ? node315 : 4'b0001;
															assign node315 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node318 = (inp[10]) ? node324 : node319;
														assign node319 = (inp[0]) ? node321 : 4'b0001;
															assign node321 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node324 = (inp[11]) ? node326 : 4'b0000;
															assign node326 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node329 = (inp[5]) ? node347 : node330;
													assign node330 = (inp[0]) ? node340 : node331;
														assign node331 = (inp[11]) ? node333 : 4'b0001;
															assign node333 = (inp[10]) ? node337 : node334;
																assign node334 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node337 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node340 = (inp[10]) ? node344 : node341;
															assign node341 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node344 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node347 = (inp[0]) ? node363 : node348;
														assign node348 = (inp[9]) ? node356 : node349;
															assign node349 = (inp[11]) ? node353 : node350;
																assign node350 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node353 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node356 = (inp[11]) ? node360 : node357;
																assign node357 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node360 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node363 = (inp[11]) ? node369 : node364;
															assign node364 = (inp[9]) ? 4'b0101 : node365;
																assign node365 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node369 = (inp[9]) ? node371 : 4'b0101;
																assign node371 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node374 = (inp[5]) ? node412 : node375;
												assign node375 = (inp[10]) ? node391 : node376;
													assign node376 = (inp[9]) ? node384 : node377;
														assign node377 = (inp[1]) ? node379 : 4'b0100;
															assign node379 = (inp[0]) ? 4'b0101 : node380;
																assign node380 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node384 = (inp[1]) ? 4'b0100 : node385;
															assign node385 = (inp[0]) ? node387 : 4'b0101;
																assign node387 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node391 = (inp[0]) ? node401 : node392;
														assign node392 = (inp[9]) ? node398 : node393;
															assign node393 = (inp[1]) ? node395 : 4'b0101;
																assign node395 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node398 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node401 = (inp[9]) ? node407 : node402;
															assign node402 = (inp[11]) ? 4'b0100 : node403;
																assign node403 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node407 = (inp[11]) ? 4'b0101 : node408;
																assign node408 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node412 = (inp[1]) ? node424 : node413;
													assign node413 = (inp[9]) ? node419 : node414;
														assign node414 = (inp[10]) ? node416 : 4'b0100;
															assign node416 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node419 = (inp[10]) ? node421 : 4'b0101;
															assign node421 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node424 = (inp[11]) ? node430 : node425;
														assign node425 = (inp[0]) ? node427 : 4'b0000;
															assign node427 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node430 = (inp[10]) ? 4'b0001 : node431;
															assign node431 = (inp[0]) ? node435 : node432;
																assign node432 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node435 = (inp[9]) ? 4'b0001 : 4'b0000;
										assign node439 = (inp[2]) ? node513 : node440;
											assign node440 = (inp[1]) ? node478 : node441;
												assign node441 = (inp[11]) ? node453 : node442;
													assign node442 = (inp[0]) ? node448 : node443;
														assign node443 = (inp[10]) ? node445 : 4'b0101;
															assign node445 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node448 = (inp[5]) ? node450 : 4'b0100;
															assign node450 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node453 = (inp[5]) ? node463 : node454;
														assign node454 = (inp[10]) ? node456 : 4'b0100;
															assign node456 = (inp[9]) ? node460 : node457;
																assign node457 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node460 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node463 = (inp[9]) ? node471 : node464;
															assign node464 = (inp[10]) ? node468 : node465;
																assign node465 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node468 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node471 = (inp[0]) ? node475 : node472;
																assign node472 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node475 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node478 = (inp[5]) ? node492 : node479;
													assign node479 = (inp[0]) ? node487 : node480;
														assign node480 = (inp[11]) ? 4'b0100 : node481;
															assign node481 = (inp[9]) ? node483 : 4'b0101;
																assign node483 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node487 = (inp[9]) ? node489 : 4'b0100;
															assign node489 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node492 = (inp[0]) ? node500 : node493;
														assign node493 = (inp[9]) ? node497 : node494;
															assign node494 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node497 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node500 = (inp[10]) ? node506 : node501;
															assign node501 = (inp[11]) ? node503 : 4'b0001;
																assign node503 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node506 = (inp[11]) ? node510 : node507;
																assign node507 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node510 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node513 = (inp[5]) ? node549 : node514;
												assign node514 = (inp[9]) ? node536 : node515;
													assign node515 = (inp[10]) ? node527 : node516;
														assign node516 = (inp[0]) ? node522 : node517;
															assign node517 = (inp[11]) ? 4'b0000 : node518;
																assign node518 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node522 = (inp[1]) ? node524 : 4'b0000;
																assign node524 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node527 = (inp[0]) ? node533 : node528;
															assign node528 = (inp[1]) ? 4'b0001 : node529;
																assign node529 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node533 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node536 = (inp[10]) ? node544 : node537;
														assign node537 = (inp[11]) ? 4'b0001 : node538;
															assign node538 = (inp[0]) ? 4'b0001 : node539;
																assign node539 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node544 = (inp[0]) ? 4'b0000 : node545;
															assign node545 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node549 = (inp[1]) ? node569 : node550;
													assign node550 = (inp[0]) ? node564 : node551;
														assign node551 = (inp[10]) ? node559 : node552;
															assign node552 = (inp[11]) ? node556 : node553;
																assign node553 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node556 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node559 = (inp[9]) ? 4'b0000 : node560;
																assign node560 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node564 = (inp[10]) ? 4'b0000 : node565;
															assign node565 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node569 = (inp[10]) ? node579 : node570;
														assign node570 = (inp[9]) ? node576 : node571;
															assign node571 = (inp[0]) ? node573 : 4'b0100;
																assign node573 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node576 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node579 = (inp[9]) ? node581 : 4'b0101;
															assign node581 = (inp[0]) ? 4'b0101 : 4'b0100;
								assign node584 = (inp[15]) ? node898 : node585;
									assign node585 = (inp[11]) ? node707 : node586;
										assign node586 = (inp[10]) ? node648 : node587;
											assign node587 = (inp[9]) ? node617 : node588;
												assign node588 = (inp[5]) ? node598 : node589;
													assign node589 = (inp[2]) ? node593 : node590;
														assign node590 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node593 = (inp[13]) ? node595 : 4'b0101;
															assign node595 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node598 = (inp[2]) ? node612 : node599;
														assign node599 = (inp[0]) ? node607 : node600;
															assign node600 = (inp[13]) ? node604 : node601;
																assign node601 = (inp[1]) ? 4'b0100 : 4'b0000;
																assign node604 = (inp[1]) ? 4'b0001 : 4'b0100;
															assign node607 = (inp[13]) ? 4'b0001 : node608;
																assign node608 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node612 = (inp[13]) ? node614 : 4'b0000;
															assign node614 = (inp[1]) ? 4'b0100 : 4'b0000;
												assign node617 = (inp[13]) ? node635 : node618;
													assign node618 = (inp[2]) ? node628 : node619;
														assign node619 = (inp[5]) ? node621 : 4'b0001;
															assign node621 = (inp[0]) ? node625 : node622;
																assign node622 = (inp[1]) ? 4'b0101 : 4'b0001;
																assign node625 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node628 = (inp[5]) ? node630 : 4'b0100;
															assign node630 = (inp[1]) ? 4'b0001 : node631;
																assign node631 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node635 = (inp[2]) ? node641 : node636;
														assign node636 = (inp[5]) ? node638 : 4'b0101;
															assign node638 = (inp[1]) ? 4'b0000 : 4'b0101;
														assign node641 = (inp[1]) ? node645 : node642;
															assign node642 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node645 = (inp[5]) ? 4'b0101 : 4'b0001;
											assign node648 = (inp[9]) ? node678 : node649;
												assign node649 = (inp[13]) ? node665 : node650;
													assign node650 = (inp[2]) ? node658 : node651;
														assign node651 = (inp[5]) ? node653 : 4'b0001;
															assign node653 = (inp[0]) ? node655 : 4'b0001;
																assign node655 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node658 = (inp[5]) ? node660 : 4'b0100;
															assign node660 = (inp[1]) ? 4'b0001 : node661;
																assign node661 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node665 = (inp[5]) ? node671 : node666;
														assign node666 = (inp[2]) ? node668 : 4'b0101;
															assign node668 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node671 = (inp[2]) ? 4'b0101 : node672;
															assign node672 = (inp[1]) ? 4'b0000 : node673;
																assign node673 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node678 = (inp[5]) ? node688 : node679;
													assign node679 = (inp[2]) ? node683 : node680;
														assign node680 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node683 = (inp[0]) ? 4'b0000 : node684;
															assign node684 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node688 = (inp[2]) ? node698 : node689;
														assign node689 = (inp[0]) ? node693 : node690;
															assign node690 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node693 = (inp[13]) ? 4'b0101 : node694;
																assign node694 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node698 = (inp[13]) ? node704 : node699;
															assign node699 = (inp[1]) ? 4'b0000 : node700;
																assign node700 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node704 = (inp[1]) ? 4'b0100 : 4'b0000;
										assign node707 = (inp[5]) ? node817 : node708;
											assign node708 = (inp[1]) ? node768 : node709;
												assign node709 = (inp[9]) ? node739 : node710;
													assign node710 = (inp[10]) ? node724 : node711;
														assign node711 = (inp[0]) ? node717 : node712;
															assign node712 = (inp[13]) ? node714 : 4'b0000;
																assign node714 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node717 = (inp[2]) ? node721 : node718;
																assign node718 = (inp[13]) ? 4'b0101 : 4'b0001;
																assign node721 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node724 = (inp[0]) ? node732 : node725;
															assign node725 = (inp[13]) ? node729 : node726;
																assign node726 = (inp[2]) ? 4'b0100 : 4'b0001;
																assign node729 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node732 = (inp[2]) ? node736 : node733;
																assign node733 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node736 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node739 = (inp[10]) ? node753 : node740;
														assign node740 = (inp[2]) ? node748 : node741;
															assign node741 = (inp[0]) ? node745 : node742;
																assign node742 = (inp[13]) ? 4'b0101 : 4'b0001;
																assign node745 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node748 = (inp[13]) ? 4'b0001 : node749;
																assign node749 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node753 = (inp[0]) ? node761 : node754;
															assign node754 = (inp[2]) ? node758 : node755;
																assign node755 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node758 = (inp[13]) ? 4'b0000 : 4'b0101;
															assign node761 = (inp[2]) ? node765 : node762;
																assign node762 = (inp[13]) ? 4'b0101 : 4'b0001;
																assign node765 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node768 = (inp[9]) ? node792 : node769;
													assign node769 = (inp[10]) ? node779 : node770;
														assign node770 = (inp[13]) ? node774 : node771;
															assign node771 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node774 = (inp[2]) ? 4'b0000 : node775;
																assign node775 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node779 = (inp[13]) ? node787 : node780;
															assign node780 = (inp[2]) ? node784 : node781;
																assign node781 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node784 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node787 = (inp[2]) ? 4'b0001 : node788;
																assign node788 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node792 = (inp[0]) ? node804 : node793;
														assign node793 = (inp[13]) ? node801 : node794;
															assign node794 = (inp[2]) ? node798 : node795;
																assign node795 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node798 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node801 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node804 = (inp[10]) ? node812 : node805;
															assign node805 = (inp[2]) ? node809 : node806;
																assign node806 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node809 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node812 = (inp[2]) ? 4'b0000 : node813;
																assign node813 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node817 = (inp[10]) ? node849 : node818;
												assign node818 = (inp[9]) ? node838 : node819;
													assign node819 = (inp[2]) ? node829 : node820;
														assign node820 = (inp[1]) ? node824 : node821;
															assign node821 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node824 = (inp[13]) ? node826 : 4'b0101;
																assign node826 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node829 = (inp[0]) ? node831 : 4'b0100;
															assign node831 = (inp[13]) ? node835 : node832;
																assign node832 = (inp[1]) ? 4'b0001 : 4'b0100;
																assign node835 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node838 = (inp[2]) ? node844 : node839;
														assign node839 = (inp[1]) ? node841 : 4'b0100;
															assign node841 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node844 = (inp[13]) ? 4'b0101 : node845;
															assign node845 = (inp[1]) ? 4'b0000 : 4'b0101;
												assign node849 = (inp[9]) ? node877 : node850;
													assign node850 = (inp[2]) ? node864 : node851;
														assign node851 = (inp[0]) ? node859 : node852;
															assign node852 = (inp[13]) ? node856 : node853;
																assign node853 = (inp[1]) ? 4'b0100 : 4'b0000;
																assign node856 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node859 = (inp[13]) ? node861 : 4'b0100;
																assign node861 = (inp[1]) ? 4'b0001 : 4'b0100;
														assign node864 = (inp[0]) ? node872 : node865;
															assign node865 = (inp[1]) ? node869 : node866;
																assign node866 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node869 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node872 = (inp[13]) ? node874 : 4'b0000;
																assign node874 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node877 = (inp[2]) ? node885 : node878;
														assign node878 = (inp[0]) ? 4'b0101 : node879;
															assign node879 = (inp[1]) ? 4'b0001 : node880;
																assign node880 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node885 = (inp[0]) ? node891 : node886;
															assign node886 = (inp[1]) ? 4'b0000 : node887;
																assign node887 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node891 = (inp[1]) ? node895 : node892;
																assign node892 = (inp[13]) ? 4'b0001 : 4'b0100;
																assign node895 = (inp[13]) ? 4'b0101 : 4'b0001;
									assign node898 = (inp[0]) ? node1064 : node899;
										assign node899 = (inp[5]) ? node985 : node900;
											assign node900 = (inp[11]) ? node944 : node901;
												assign node901 = (inp[10]) ? node923 : node902;
													assign node902 = (inp[9]) ? node910 : node903;
														assign node903 = (inp[2]) ? 4'b0111 : node904;
															assign node904 = (inp[1]) ? node906 : 4'b0111;
																assign node906 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node910 = (inp[13]) ? node918 : node911;
															assign node911 = (inp[1]) ? node915 : node912;
																assign node912 = (inp[2]) ? 4'b0110 : 4'b0011;
																assign node915 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node918 = (inp[1]) ? 4'b0110 : node919;
																assign node919 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node923 = (inp[1]) ? node937 : node924;
														assign node924 = (inp[2]) ? node932 : node925;
															assign node925 = (inp[13]) ? node929 : node926;
																assign node926 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node929 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node932 = (inp[13]) ? node934 : 4'b0111;
																assign node934 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node937 = (inp[9]) ? 4'b0111 : node938;
															assign node938 = (inp[2]) ? 4'b0011 : node939;
																assign node939 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node944 = (inp[9]) ? node960 : node945;
													assign node945 = (inp[10]) ? node951 : node946;
														assign node946 = (inp[1]) ? 4'b0111 : node947;
															assign node947 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node951 = (inp[2]) ? node953 : 4'b0110;
															assign node953 = (inp[1]) ? node957 : node954;
																assign node954 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node957 = (inp[13]) ? 4'b0110 : 4'b0011;
													assign node960 = (inp[1]) ? node972 : node961;
														assign node961 = (inp[2]) ? node969 : node962;
															assign node962 = (inp[13]) ? node966 : node963;
																assign node963 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node966 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node969 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node972 = (inp[2]) ? node980 : node973;
															assign node973 = (inp[13]) ? node977 : node974;
																assign node974 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node977 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node980 = (inp[13]) ? 4'b0110 : node981;
																assign node981 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node985 = (inp[1]) ? node1021 : node986;
												assign node986 = (inp[10]) ? node1004 : node987;
													assign node987 = (inp[11]) ? node997 : node988;
														assign node988 = (inp[13]) ? node992 : node989;
															assign node989 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node992 = (inp[2]) ? node994 : 4'b0010;
																assign node994 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node997 = (inp[2]) ? node1001 : node998;
															assign node998 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node1001 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node1004 = (inp[2]) ? node1016 : node1005;
														assign node1005 = (inp[13]) ? node1013 : node1006;
															assign node1006 = (inp[9]) ? node1010 : node1007;
																assign node1007 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node1010 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node1013 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node1016 = (inp[13]) ? node1018 : 4'b0010;
															assign node1018 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node1021 = (inp[2]) ? node1043 : node1022;
													assign node1022 = (inp[13]) ? node1028 : node1023;
														assign node1023 = (inp[9]) ? node1025 : 4'b0111;
															assign node1025 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node1028 = (inp[11]) ? node1036 : node1029;
															assign node1029 = (inp[9]) ? node1033 : node1030;
																assign node1030 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node1033 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node1036 = (inp[9]) ? node1040 : node1037;
																assign node1037 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node1040 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node1043 = (inp[13]) ? node1057 : node1044;
														assign node1044 = (inp[10]) ? node1052 : node1045;
															assign node1045 = (inp[11]) ? node1049 : node1046;
																assign node1046 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node1049 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node1052 = (inp[11]) ? node1054 : 4'b0011;
																assign node1054 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node1057 = (inp[10]) ? node1059 : 4'b0111;
															assign node1059 = (inp[9]) ? 4'b0111 : node1060;
																assign node1060 = (inp[11]) ? 4'b0111 : 4'b0110;
										assign node1064 = (inp[13]) ? node1136 : node1065;
											assign node1065 = (inp[2]) ? node1105 : node1066;
												assign node1066 = (inp[5]) ? node1084 : node1067;
													assign node1067 = (inp[1]) ? node1077 : node1068;
														assign node1068 = (inp[11]) ? node1070 : 4'b0011;
															assign node1070 = (inp[10]) ? node1074 : node1071;
																assign node1071 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node1074 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node1077 = (inp[9]) ? node1081 : node1078;
															assign node1078 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node1081 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node1084 = (inp[11]) ? node1092 : node1085;
														assign node1085 = (inp[9]) ? node1089 : node1086;
															assign node1086 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node1089 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node1092 = (inp[1]) ? node1100 : node1093;
															assign node1093 = (inp[10]) ? node1097 : node1094;
																assign node1094 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node1097 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node1100 = (inp[9]) ? 4'b0111 : node1101;
																assign node1101 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node1105 = (inp[1]) ? node1123 : node1106;
													assign node1106 = (inp[5]) ? node1116 : node1107;
														assign node1107 = (inp[9]) ? 4'b0110 : node1108;
															assign node1108 = (inp[10]) ? node1112 : node1109;
																assign node1109 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node1112 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node1116 = (inp[11]) ? 4'b0010 : node1117;
															assign node1117 = (inp[9]) ? node1119 : 4'b0011;
																assign node1119 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node1123 = (inp[9]) ? node1129 : node1124;
														assign node1124 = (inp[10]) ? node1126 : 4'b0011;
															assign node1126 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node1129 = (inp[11]) ? 4'b0011 : node1130;
															assign node1130 = (inp[10]) ? node1132 : 4'b0010;
																assign node1132 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node1136 = (inp[2]) ? node1176 : node1137;
												assign node1137 = (inp[5]) ? node1157 : node1138;
													assign node1138 = (inp[1]) ? node1150 : node1139;
														assign node1139 = (inp[11]) ? node1145 : node1140;
															assign node1140 = (inp[10]) ? node1142 : 4'b0111;
																assign node1142 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node1145 = (inp[9]) ? node1147 : 4'b0110;
																assign node1147 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node1150 = (inp[9]) ? node1152 : 4'b0010;
															assign node1152 = (inp[11]) ? 4'b0011 : node1153;
																assign node1153 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node1157 = (inp[9]) ? node1169 : node1158;
														assign node1158 = (inp[10]) ? node1164 : node1159;
															assign node1159 = (inp[1]) ? 4'b0011 : node1160;
																assign node1160 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node1164 = (inp[1]) ? 4'b0010 : node1165;
																assign node1165 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node1169 = (inp[10]) ? 4'b0011 : node1170;
															assign node1170 = (inp[1]) ? 4'b0010 : node1171;
																assign node1171 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node1176 = (inp[5]) ? node1196 : node1177;
													assign node1177 = (inp[1]) ? node1185 : node1178;
														assign node1178 = (inp[10]) ? node1182 : node1179;
															assign node1179 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node1182 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node1185 = (inp[9]) ? node1191 : node1186;
															assign node1186 = (inp[10]) ? node1188 : 4'b0111;
																assign node1188 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node1191 = (inp[10]) ? node1193 : 4'b0110;
																assign node1193 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node1196 = (inp[10]) ? node1206 : node1197;
														assign node1197 = (inp[9]) ? node1203 : node1198;
															assign node1198 = (inp[1]) ? 4'b0110 : node1199;
																assign node1199 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node1203 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node1206 = (inp[9]) ? node1212 : node1207;
															assign node1207 = (inp[1]) ? 4'b0111 : node1208;
																assign node1208 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node1212 = (inp[11]) ? 4'b0110 : node1213;
																assign node1213 = (inp[1]) ? 4'b0110 : 4'b0111;
							assign node1217 = (inp[15]) ? node1643 : node1218;
								assign node1218 = (inp[10]) ? node1426 : node1219;
									assign node1219 = (inp[9]) ? node1327 : node1220;
										assign node1220 = (inp[2]) ? node1274 : node1221;
											assign node1221 = (inp[13]) ? node1253 : node1222;
												assign node1222 = (inp[1]) ? node1240 : node1223;
													assign node1223 = (inp[4]) ? node1233 : node1224;
														assign node1224 = (inp[5]) ? node1228 : node1225;
															assign node1225 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node1228 = (inp[11]) ? node1230 : 4'b0011;
																assign node1230 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node1233 = (inp[0]) ? node1235 : 4'b0010;
															assign node1235 = (inp[11]) ? node1237 : 4'b0010;
																assign node1237 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node1240 = (inp[5]) ? node1246 : node1241;
														assign node1241 = (inp[11]) ? node1243 : 4'b0010;
															assign node1243 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1246 = (inp[11]) ? 4'b0110 : node1247;
															assign node1247 = (inp[4]) ? node1249 : 4'b0111;
																assign node1249 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node1253 = (inp[5]) ? node1259 : node1254;
													assign node1254 = (inp[11]) ? node1256 : 4'b0110;
														assign node1256 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node1259 = (inp[1]) ? node1263 : node1260;
														assign node1260 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node1263 = (inp[11]) ? node1269 : node1264;
															assign node1264 = (inp[4]) ? 4'b0010 : node1265;
																assign node1265 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node1269 = (inp[4]) ? node1271 : 4'b0010;
																assign node1271 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node1274 = (inp[13]) ? node1300 : node1275;
												assign node1275 = (inp[5]) ? node1287 : node1276;
													assign node1276 = (inp[4]) ? node1282 : node1277;
														assign node1277 = (inp[11]) ? node1279 : 4'b0110;
															assign node1279 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node1282 = (inp[0]) ? node1284 : 4'b0111;
															assign node1284 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node1287 = (inp[1]) ? node1293 : node1288;
														assign node1288 = (inp[4]) ? 4'b0111 : node1289;
															assign node1289 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node1293 = (inp[0]) ? node1295 : 4'b0011;
															assign node1295 = (inp[11]) ? 4'b0010 : node1296;
																assign node1296 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node1300 = (inp[5]) ? node1312 : node1301;
													assign node1301 = (inp[4]) ? node1307 : node1302;
														assign node1302 = (inp[0]) ? 4'b0011 : node1303;
															assign node1303 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node1307 = (inp[0]) ? 4'b0010 : node1308;
															assign node1308 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1312 = (inp[1]) ? node1320 : node1313;
														assign node1313 = (inp[4]) ? 4'b0011 : node1314;
															assign node1314 = (inp[0]) ? 4'b0010 : node1315;
																assign node1315 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node1320 = (inp[4]) ? node1322 : 4'b0110;
															assign node1322 = (inp[0]) ? node1324 : 4'b0111;
																assign node1324 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node1327 = (inp[2]) ? node1371 : node1328;
											assign node1328 = (inp[13]) ? node1346 : node1329;
												assign node1329 = (inp[5]) ? node1335 : node1330;
													assign node1330 = (inp[0]) ? node1332 : 4'b0011;
														assign node1332 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1335 = (inp[1]) ? node1341 : node1336;
														assign node1336 = (inp[11]) ? 4'b0011 : node1337;
															assign node1337 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1341 = (inp[11]) ? 4'b0111 : node1342;
															assign node1342 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node1346 = (inp[1]) ? node1360 : node1347;
													assign node1347 = (inp[11]) ? node1355 : node1348;
														assign node1348 = (inp[5]) ? node1350 : 4'b0111;
															assign node1350 = (inp[0]) ? node1352 : 4'b0110;
																assign node1352 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node1355 = (inp[0]) ? node1357 : 4'b0111;
															assign node1357 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node1360 = (inp[5]) ? node1366 : node1361;
														assign node1361 = (inp[11]) ? node1363 : 4'b0111;
															assign node1363 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node1366 = (inp[11]) ? 4'b0011 : node1367;
															assign node1367 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node1371 = (inp[13]) ? node1389 : node1372;
												assign node1372 = (inp[4]) ? node1380 : node1373;
													assign node1373 = (inp[5]) ? node1375 : 4'b0111;
														assign node1375 = (inp[1]) ? 4'b0010 : node1376;
															assign node1376 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node1380 = (inp[1]) ? node1386 : node1381;
														assign node1381 = (inp[11]) ? 4'b0110 : node1382;
															assign node1382 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node1386 = (inp[5]) ? 4'b0010 : 4'b0110;
												assign node1389 = (inp[1]) ? node1409 : node1390;
													assign node1390 = (inp[0]) ? node1400 : node1391;
														assign node1391 = (inp[5]) ? 4'b0010 : node1392;
															assign node1392 = (inp[4]) ? node1396 : node1393;
																assign node1393 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node1396 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node1400 = (inp[5]) ? node1404 : node1401;
															assign node1401 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node1404 = (inp[4]) ? node1406 : 4'b0011;
																assign node1406 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node1409 = (inp[5]) ? node1415 : node1410;
														assign node1410 = (inp[4]) ? 4'b0011 : node1411;
															assign node1411 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node1415 = (inp[4]) ? node1421 : node1416;
															assign node1416 = (inp[11]) ? 4'b0111 : node1417;
																assign node1417 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node1421 = (inp[0]) ? node1423 : 4'b0110;
																assign node1423 = (inp[11]) ? 4'b0111 : 4'b0110;
									assign node1426 = (inp[9]) ? node1536 : node1427;
										assign node1427 = (inp[2]) ? node1483 : node1428;
											assign node1428 = (inp[13]) ? node1450 : node1429;
												assign node1429 = (inp[5]) ? node1435 : node1430;
													assign node1430 = (inp[11]) ? node1432 : 4'b0011;
														assign node1432 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node1435 = (inp[1]) ? node1443 : node1436;
														assign node1436 = (inp[11]) ? node1438 : 4'b0010;
															assign node1438 = (inp[4]) ? 4'b0011 : node1439;
																assign node1439 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1443 = (inp[11]) ? node1445 : 4'b0110;
															assign node1445 = (inp[4]) ? 4'b0111 : node1446;
																assign node1446 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node1450 = (inp[1]) ? node1472 : node1451;
													assign node1451 = (inp[4]) ? node1463 : node1452;
														assign node1452 = (inp[5]) ? node1458 : node1453;
															assign node1453 = (inp[0]) ? node1455 : 4'b0111;
																assign node1455 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node1458 = (inp[11]) ? node1460 : 4'b0110;
																assign node1460 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node1463 = (inp[11]) ? node1467 : node1464;
															assign node1464 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node1467 = (inp[5]) ? 4'b0111 : node1468;
																assign node1468 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node1472 = (inp[5]) ? node1474 : 4'b0111;
														assign node1474 = (inp[11]) ? node1480 : node1475;
															assign node1475 = (inp[0]) ? 4'b0011 : node1476;
																assign node1476 = (inp[4]) ? 4'b0011 : 4'b0010;
															assign node1480 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node1483 = (inp[13]) ? node1513 : node1484;
												assign node1484 = (inp[1]) ? node1496 : node1485;
													assign node1485 = (inp[4]) ? node1487 : 4'b0110;
														assign node1487 = (inp[5]) ? node1491 : node1488;
															assign node1488 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node1491 = (inp[0]) ? 4'b0110 : node1492;
																assign node1492 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node1496 = (inp[5]) ? node1506 : node1497;
														assign node1497 = (inp[4]) ? node1503 : node1498;
															assign node1498 = (inp[0]) ? node1500 : 4'b0111;
																assign node1500 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node1503 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node1506 = (inp[11]) ? 4'b0011 : node1507;
															assign node1507 = (inp[0]) ? node1509 : 4'b0010;
																assign node1509 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node1513 = (inp[5]) ? node1525 : node1514;
													assign node1514 = (inp[4]) ? node1520 : node1515;
														assign node1515 = (inp[0]) ? 4'b0010 : node1516;
															assign node1516 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node1520 = (inp[11]) ? 4'b0011 : node1521;
															assign node1521 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node1525 = (inp[1]) ? node1533 : node1526;
														assign node1526 = (inp[4]) ? node1528 : 4'b0011;
															assign node1528 = (inp[11]) ? node1530 : 4'b0010;
																assign node1530 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1533 = (inp[11]) ? 4'b0111 : 4'b0110;
										assign node1536 = (inp[2]) ? node1582 : node1537;
											assign node1537 = (inp[13]) ? node1563 : node1538;
												assign node1538 = (inp[1]) ? node1558 : node1539;
													assign node1539 = (inp[11]) ? node1545 : node1540;
														assign node1540 = (inp[5]) ? node1542 : 4'b0010;
															assign node1542 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node1545 = (inp[4]) ? node1553 : node1546;
															assign node1546 = (inp[0]) ? node1550 : node1547;
																assign node1547 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node1550 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node1553 = (inp[0]) ? node1555 : 4'b0010;
																assign node1555 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node1558 = (inp[5]) ? node1560 : 4'b0010;
														assign node1560 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node1563 = (inp[5]) ? node1569 : node1564;
													assign node1564 = (inp[11]) ? node1566 : 4'b0110;
														assign node1566 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node1569 = (inp[1]) ? node1577 : node1570;
														assign node1570 = (inp[11]) ? node1572 : 4'b0111;
															assign node1572 = (inp[4]) ? 4'b0110 : node1573;
																assign node1573 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node1577 = (inp[4]) ? 4'b0011 : node1578;
															assign node1578 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node1582 = (inp[13]) ? node1616 : node1583;
												assign node1583 = (inp[1]) ? node1599 : node1584;
													assign node1584 = (inp[5]) ? node1592 : node1585;
														assign node1585 = (inp[4]) ? node1589 : node1586;
															assign node1586 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node1589 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node1592 = (inp[4]) ? 4'b0111 : node1593;
															assign node1593 = (inp[11]) ? node1595 : 4'b0111;
																assign node1595 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node1599 = (inp[5]) ? node1609 : node1600;
														assign node1600 = (inp[4]) ? node1604 : node1601;
															assign node1601 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node1604 = (inp[0]) ? node1606 : 4'b0111;
																assign node1606 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node1609 = (inp[4]) ? node1611 : 4'b0010;
															assign node1611 = (inp[11]) ? node1613 : 4'b0011;
																assign node1613 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node1616 = (inp[1]) ? node1630 : node1617;
													assign node1617 = (inp[11]) ? node1625 : node1618;
														assign node1618 = (inp[0]) ? node1620 : 4'b0011;
															assign node1620 = (inp[4]) ? node1622 : 4'b0010;
																assign node1622 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node1625 = (inp[5]) ? 4'b0010 : node1626;
															assign node1626 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node1630 = (inp[5]) ? node1636 : node1631;
														assign node1631 = (inp[4]) ? 4'b0010 : node1632;
															assign node1632 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1636 = (inp[11]) ? 4'b0110 : node1637;
															assign node1637 = (inp[0]) ? node1639 : 4'b0111;
																assign node1639 = (inp[4]) ? 4'b0111 : 4'b0110;
								assign node1643 = (inp[4]) ? node1903 : node1644;
									assign node1644 = (inp[9]) ? node1774 : node1645;
										assign node1645 = (inp[10]) ? node1709 : node1646;
											assign node1646 = (inp[2]) ? node1680 : node1647;
												assign node1647 = (inp[13]) ? node1663 : node1648;
													assign node1648 = (inp[5]) ? node1656 : node1649;
														assign node1649 = (inp[1]) ? node1651 : 4'b0110;
															assign node1651 = (inp[0]) ? 4'b0111 : node1652;
																assign node1652 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node1656 = (inp[1]) ? node1660 : node1657;
															assign node1657 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node1660 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node1663 = (inp[1]) ? node1671 : node1664;
														assign node1664 = (inp[11]) ? 4'b0010 : node1665;
															assign node1665 = (inp[0]) ? 4'b0011 : node1666;
																assign node1666 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node1671 = (inp[5]) ? node1675 : node1672;
															assign node1672 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1675 = (inp[0]) ? node1677 : 4'b0111;
																assign node1677 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node1680 = (inp[13]) ? node1694 : node1681;
													assign node1681 = (inp[1]) ? node1687 : node1682;
														assign node1682 = (inp[5]) ? 4'b0010 : node1683;
															assign node1683 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1687 = (inp[5]) ? node1691 : node1688;
															assign node1688 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node1691 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node1694 = (inp[1]) ? node1702 : node1695;
														assign node1695 = (inp[5]) ? node1697 : 4'b0110;
															assign node1697 = (inp[0]) ? 4'b0111 : node1698;
																assign node1698 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node1702 = (inp[5]) ? 4'b0010 : node1703;
															assign node1703 = (inp[0]) ? node1705 : 4'b0110;
																assign node1705 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node1709 = (inp[2]) ? node1747 : node1710;
												assign node1710 = (inp[13]) ? node1726 : node1711;
													assign node1711 = (inp[5]) ? node1719 : node1712;
														assign node1712 = (inp[11]) ? 4'b0110 : node1713;
															assign node1713 = (inp[1]) ? node1715 : 4'b0111;
																assign node1715 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node1719 = (inp[1]) ? node1723 : node1720;
															assign node1720 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node1723 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1726 = (inp[5]) ? node1738 : node1727;
														assign node1727 = (inp[1]) ? node1733 : node1728;
															assign node1728 = (inp[11]) ? 4'b0011 : node1729;
																assign node1729 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1733 = (inp[11]) ? node1735 : 4'b0011;
																assign node1735 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node1738 = (inp[1]) ? node1742 : node1739;
															assign node1739 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node1742 = (inp[0]) ? node1744 : 4'b0110;
																assign node1744 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node1747 = (inp[13]) ? node1761 : node1748;
													assign node1748 = (inp[5]) ? node1752 : node1749;
														assign node1749 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node1752 = (inp[1]) ? node1756 : node1753;
															assign node1753 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node1756 = (inp[0]) ? node1758 : 4'b0111;
																assign node1758 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node1761 = (inp[5]) ? node1769 : node1762;
														assign node1762 = (inp[11]) ? node1766 : node1763;
															assign node1763 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node1766 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node1769 = (inp[11]) ? 4'b0110 : node1770;
															assign node1770 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node1774 = (inp[2]) ? node1838 : node1775;
											assign node1775 = (inp[13]) ? node1805 : node1776;
												assign node1776 = (inp[1]) ? node1792 : node1777;
													assign node1777 = (inp[11]) ? node1785 : node1778;
														assign node1778 = (inp[10]) ? node1782 : node1779;
															assign node1779 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node1782 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node1785 = (inp[10]) ? node1787 : 4'b0110;
															assign node1787 = (inp[0]) ? 4'b0110 : node1788;
																assign node1788 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node1792 = (inp[5]) ? node1796 : node1793;
														assign node1793 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node1796 = (inp[10]) ? node1800 : node1797;
															assign node1797 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node1800 = (inp[11]) ? node1802 : 4'b0010;
																assign node1802 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node1805 = (inp[1]) ? node1823 : node1806;
													assign node1806 = (inp[10]) ? node1816 : node1807;
														assign node1807 = (inp[5]) ? node1813 : node1808;
															assign node1808 = (inp[11]) ? 4'b0011 : node1809;
																assign node1809 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node1813 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node1816 = (inp[5]) ? node1818 : 4'b0010;
															assign node1818 = (inp[0]) ? 4'b0011 : node1819;
																assign node1819 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node1823 = (inp[5]) ? node1829 : node1824;
														assign node1824 = (inp[10]) ? node1826 : 4'b0011;
															assign node1826 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node1829 = (inp[10]) ? node1833 : node1830;
															assign node1830 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node1833 = (inp[0]) ? node1835 : 4'b0111;
																assign node1835 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node1838 = (inp[13]) ? node1866 : node1839;
												assign node1839 = (inp[1]) ? node1851 : node1840;
													assign node1840 = (inp[10]) ? node1846 : node1841;
														assign node1841 = (inp[5]) ? node1843 : 4'b0010;
															assign node1843 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node1846 = (inp[5]) ? node1848 : 4'b0011;
															assign node1848 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node1851 = (inp[5]) ? node1855 : node1852;
														assign node1852 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node1855 = (inp[10]) ? node1861 : node1856;
															assign node1856 = (inp[0]) ? node1858 : 4'b0111;
																assign node1858 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node1861 = (inp[0]) ? node1863 : 4'b0110;
																assign node1863 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node1866 = (inp[1]) ? node1886 : node1867;
													assign node1867 = (inp[0]) ? node1881 : node1868;
														assign node1868 = (inp[10]) ? node1876 : node1869;
															assign node1869 = (inp[5]) ? node1873 : node1870;
																assign node1870 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node1873 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node1876 = (inp[11]) ? node1878 : 4'b0111;
																assign node1878 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node1881 = (inp[10]) ? 4'b0110 : node1882;
															assign node1882 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node1886 = (inp[5]) ? node1894 : node1887;
														assign node1887 = (inp[10]) ? node1889 : 4'b0111;
															assign node1889 = (inp[11]) ? node1891 : 4'b0110;
																assign node1891 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node1894 = (inp[11]) ? 4'b0010 : node1895;
															assign node1895 = (inp[10]) ? node1899 : node1896;
																assign node1896 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node1899 = (inp[0]) ? 4'b0010 : 4'b0011;
									assign node1903 = (inp[5]) ? node2057 : node1904;
										assign node1904 = (inp[2]) ? node1986 : node1905;
											assign node1905 = (inp[13]) ? node1945 : node1906;
												assign node1906 = (inp[11]) ? node1924 : node1907;
													assign node1907 = (inp[9]) ? node1917 : node1908;
														assign node1908 = (inp[10]) ? node1912 : node1909;
															assign node1909 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node1912 = (inp[0]) ? 4'b0000 : node1913;
																assign node1913 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node1917 = (inp[10]) ? 4'b0001 : node1918;
															assign node1918 = (inp[0]) ? 4'b0000 : node1919;
																assign node1919 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node1924 = (inp[10]) ? node1936 : node1925;
														assign node1925 = (inp[9]) ? node1931 : node1926;
															assign node1926 = (inp[1]) ? node1928 : 4'b0001;
																assign node1928 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node1931 = (inp[1]) ? node1933 : 4'b0000;
																assign node1933 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node1936 = (inp[9]) ? node1942 : node1937;
															assign node1937 = (inp[1]) ? node1939 : 4'b0000;
																assign node1939 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node1942 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node1945 = (inp[1]) ? node1965 : node1946;
													assign node1946 = (inp[11]) ? node1956 : node1947;
														assign node1947 = (inp[9]) ? node1949 : 4'b0100;
															assign node1949 = (inp[10]) ? node1953 : node1950;
																assign node1950 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node1953 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node1956 = (inp[0]) ? 4'b0101 : node1957;
															assign node1957 = (inp[10]) ? node1961 : node1958;
																assign node1958 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node1961 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node1965 = (inp[11]) ? node1979 : node1966;
														assign node1966 = (inp[0]) ? node1972 : node1967;
															assign node1967 = (inp[9]) ? 4'b0101 : node1968;
																assign node1968 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node1972 = (inp[10]) ? node1976 : node1973;
																assign node1973 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node1976 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node1979 = (inp[0]) ? 4'b0100 : node1980;
															assign node1980 = (inp[9]) ? 4'b0100 : node1981;
																assign node1981 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node1986 = (inp[13]) ? node2020 : node1987;
												assign node1987 = (inp[9]) ? node2005 : node1988;
													assign node1988 = (inp[10]) ? node1994 : node1989;
														assign node1989 = (inp[0]) ? 4'b0101 : node1990;
															assign node1990 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node1994 = (inp[0]) ? node2000 : node1995;
															assign node1995 = (inp[11]) ? 4'b0101 : node1996;
																assign node1996 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node2000 = (inp[1]) ? node2002 : 4'b0101;
																assign node2002 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node2005 = (inp[10]) ? node2015 : node2006;
														assign node2006 = (inp[1]) ? node2010 : node2007;
															assign node2007 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node2010 = (inp[11]) ? node2012 : 4'b0101;
																assign node2012 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node2015 = (inp[11]) ? node2017 : 4'b0100;
															assign node2017 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node2020 = (inp[11]) ? node2038 : node2021;
													assign node2021 = (inp[10]) ? node2027 : node2022;
														assign node2022 = (inp[9]) ? 4'b0000 : node2023;
															assign node2023 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node2027 = (inp[9]) ? node2033 : node2028;
															assign node2028 = (inp[1]) ? node2030 : 4'b0000;
																assign node2030 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node2033 = (inp[0]) ? node2035 : 4'b0001;
																assign node2035 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node2038 = (inp[10]) ? node2050 : node2039;
														assign node2039 = (inp[9]) ? node2045 : node2040;
															assign node2040 = (inp[1]) ? 4'b0000 : node2041;
																assign node2041 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node2045 = (inp[1]) ? 4'b0001 : node2046;
																assign node2046 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node2050 = (inp[9]) ? node2052 : 4'b0001;
															assign node2052 = (inp[1]) ? 4'b0000 : node2053;
																assign node2053 = (inp[0]) ? 4'b0000 : 4'b0001;
										assign node2057 = (inp[1]) ? node2133 : node2058;
											assign node2058 = (inp[13]) ? node2098 : node2059;
												assign node2059 = (inp[2]) ? node2075 : node2060;
													assign node2060 = (inp[11]) ? node2064 : node2061;
														assign node2061 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node2064 = (inp[10]) ? node2070 : node2065;
															assign node2065 = (inp[0]) ? 4'b0000 : node2066;
																assign node2066 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node2070 = (inp[9]) ? 4'b0001 : node2071;
																assign node2071 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node2075 = (inp[11]) ? node2083 : node2076;
														assign node2076 = (inp[10]) ? node2080 : node2077;
															assign node2077 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node2080 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node2083 = (inp[9]) ? node2091 : node2084;
															assign node2084 = (inp[0]) ? node2088 : node2085;
																assign node2085 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node2088 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node2091 = (inp[0]) ? node2095 : node2092;
																assign node2092 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node2095 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node2098 = (inp[2]) ? node2114 : node2099;
													assign node2099 = (inp[9]) ? node2109 : node2100;
														assign node2100 = (inp[10]) ? node2106 : node2101;
															assign node2101 = (inp[11]) ? node2103 : 4'b0101;
																assign node2103 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node2106 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node2109 = (inp[10]) ? 4'b0101 : node2110;
															assign node2110 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node2114 = (inp[0]) ? node2124 : node2115;
														assign node2115 = (inp[9]) ? 4'b0001 : node2116;
															assign node2116 = (inp[11]) ? node2120 : node2117;
																assign node2117 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node2120 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node2124 = (inp[11]) ? 4'b0000 : node2125;
															assign node2125 = (inp[10]) ? node2129 : node2126;
																assign node2126 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node2129 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node2133 = (inp[10]) ? node2169 : node2134;
												assign node2134 = (inp[13]) ? node2154 : node2135;
													assign node2135 = (inp[2]) ? node2145 : node2136;
														assign node2136 = (inp[9]) ? node2142 : node2137;
															assign node2137 = (inp[11]) ? 4'b0101 : node2138;
																assign node2138 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node2142 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node2145 = (inp[11]) ? node2149 : node2146;
															assign node2146 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node2149 = (inp[0]) ? node2151 : 4'b0001;
																assign node2151 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node2154 = (inp[2]) ? node2162 : node2155;
														assign node2155 = (inp[9]) ? node2157 : 4'b0000;
															assign node2157 = (inp[11]) ? node2159 : 4'b0001;
																assign node2159 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node2162 = (inp[9]) ? node2164 : 4'b0101;
															assign node2164 = (inp[0]) ? node2166 : 4'b0100;
																assign node2166 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node2169 = (inp[11]) ? node2189 : node2170;
													assign node2170 = (inp[9]) ? node2180 : node2171;
														assign node2171 = (inp[0]) ? 4'b0100 : node2172;
															assign node2172 = (inp[13]) ? node2176 : node2173;
																assign node2173 = (inp[2]) ? 4'b0001 : 4'b0101;
																assign node2176 = (inp[2]) ? 4'b0100 : 4'b0001;
														assign node2180 = (inp[2]) ? node2186 : node2181;
															assign node2181 = (inp[13]) ? 4'b0000 : node2182;
																assign node2182 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node2186 = (inp[13]) ? 4'b0101 : 4'b0000;
													assign node2189 = (inp[0]) ? node2201 : node2190;
														assign node2190 = (inp[13]) ? node2196 : node2191;
															assign node2191 = (inp[2]) ? node2193 : 4'b0101;
																assign node2193 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node2196 = (inp[2]) ? node2198 : 4'b0000;
																assign node2198 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node2201 = (inp[9]) ? 4'b0001 : 4'b0000;
						assign node2204 = (inp[7]) ? node3464 : node2205;
							assign node2205 = (inp[15]) ? node2863 : node2206;
								assign node2206 = (inp[4]) ? node2518 : node2207;
									assign node2207 = (inp[9]) ? node2357 : node2208;
										assign node2208 = (inp[10]) ? node2274 : node2209;
											assign node2209 = (inp[1]) ? node2233 : node2210;
												assign node2210 = (inp[11]) ? node2220 : node2211;
													assign node2211 = (inp[13]) ? node2215 : node2212;
														assign node2212 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node2215 = (inp[2]) ? node2217 : 4'b0110;
															assign node2217 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node2220 = (inp[0]) ? node2228 : node2221;
														assign node2221 = (inp[2]) ? node2225 : node2222;
															assign node2222 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node2225 = (inp[13]) ? 4'b0011 : 4'b0110;
														assign node2228 = (inp[2]) ? node2230 : 4'b0011;
															assign node2230 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node2233 = (inp[11]) ? node2257 : node2234;
													assign node2234 = (inp[0]) ? node2248 : node2235;
														assign node2235 = (inp[13]) ? node2243 : node2236;
															assign node2236 = (inp[2]) ? node2240 : node2237;
																assign node2237 = (inp[5]) ? 4'b0111 : 4'b0011;
																assign node2240 = (inp[5]) ? 4'b0011 : 4'b0111;
															assign node2243 = (inp[2]) ? node2245 : 4'b0111;
																assign node2245 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node2248 = (inp[13]) ? 4'b0010 : node2249;
															assign node2249 = (inp[5]) ? node2253 : node2250;
																assign node2250 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node2253 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node2257 = (inp[2]) ? node2267 : node2258;
														assign node2258 = (inp[0]) ? 4'b0010 : node2259;
															assign node2259 = (inp[5]) ? node2263 : node2260;
																assign node2260 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node2263 = (inp[13]) ? 4'b0010 : 4'b0111;
														assign node2267 = (inp[13]) ? node2271 : node2268;
															assign node2268 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node2271 = (inp[5]) ? 4'b0110 : 4'b0010;
											assign node2274 = (inp[1]) ? node2300 : node2275;
												assign node2275 = (inp[0]) ? node2285 : node2276;
													assign node2276 = (inp[13]) ? node2280 : node2277;
														assign node2277 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node2280 = (inp[2]) ? node2282 : 4'b0111;
															assign node2282 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node2285 = (inp[11]) ? node2291 : node2286;
														assign node2286 = (inp[2]) ? 4'b0010 : node2287;
															assign node2287 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node2291 = (inp[5]) ? node2293 : 4'b0110;
															assign node2293 = (inp[2]) ? node2297 : node2294;
																assign node2294 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node2297 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node2300 = (inp[0]) ? node2332 : node2301;
													assign node2301 = (inp[11]) ? node2317 : node2302;
														assign node2302 = (inp[2]) ? node2310 : node2303;
															assign node2303 = (inp[13]) ? node2307 : node2304;
																assign node2304 = (inp[5]) ? 4'b0110 : 4'b0010;
																assign node2307 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node2310 = (inp[13]) ? node2314 : node2311;
																assign node2311 = (inp[5]) ? 4'b0010 : 4'b0110;
																assign node2314 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node2317 = (inp[5]) ? node2325 : node2318;
															assign node2318 = (inp[2]) ? node2322 : node2319;
																assign node2319 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node2322 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node2325 = (inp[2]) ? node2329 : node2326;
																assign node2326 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node2329 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node2332 = (inp[11]) ? node2348 : node2333;
														assign node2333 = (inp[2]) ? node2341 : node2334;
															assign node2334 = (inp[5]) ? node2338 : node2335;
																assign node2335 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node2338 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node2341 = (inp[5]) ? node2345 : node2342;
																assign node2342 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node2345 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node2348 = (inp[2]) ? node2350 : 4'b0011;
															assign node2350 = (inp[13]) ? node2354 : node2351;
																assign node2351 = (inp[5]) ? 4'b0011 : 4'b0111;
																assign node2354 = (inp[5]) ? 4'b0111 : 4'b0011;
										assign node2357 = (inp[10]) ? node2431 : node2358;
											assign node2358 = (inp[0]) ? node2394 : node2359;
												assign node2359 = (inp[1]) ? node2375 : node2360;
													assign node2360 = (inp[11]) ? node2368 : node2361;
														assign node2361 = (inp[2]) ? node2365 : node2362;
															assign node2362 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node2365 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node2368 = (inp[13]) ? node2372 : node2369;
															assign node2369 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node2372 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node2375 = (inp[11]) ? node2383 : node2376;
														assign node2376 = (inp[2]) ? 4'b0010 : node2377;
															assign node2377 = (inp[13]) ? node2379 : 4'b0110;
																assign node2379 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node2383 = (inp[13]) ? node2389 : node2384;
															assign node2384 = (inp[5]) ? node2386 : 4'b0110;
																assign node2386 = (inp[2]) ? 4'b0011 : 4'b0110;
															assign node2389 = (inp[5]) ? node2391 : 4'b0011;
																assign node2391 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node2394 = (inp[1]) ? node2410 : node2395;
													assign node2395 = (inp[11]) ? node2403 : node2396;
														assign node2396 = (inp[2]) ? node2400 : node2397;
															assign node2397 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node2400 = (inp[13]) ? 4'b0010 : 4'b0111;
														assign node2403 = (inp[2]) ? node2407 : node2404;
															assign node2404 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node2407 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node2410 = (inp[11]) ? node2418 : node2411;
														assign node2411 = (inp[13]) ? 4'b0011 : node2412;
															assign node2412 = (inp[2]) ? 4'b0011 : node2413;
																assign node2413 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node2418 = (inp[13]) ? node2424 : node2419;
															assign node2419 = (inp[5]) ? node2421 : 4'b0111;
																assign node2421 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node2424 = (inp[5]) ? node2428 : node2425;
																assign node2425 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node2428 = (inp[2]) ? 4'b0111 : 4'b0011;
											assign node2431 = (inp[5]) ? node2477 : node2432;
												assign node2432 = (inp[11]) ? node2448 : node2433;
													assign node2433 = (inp[1]) ? node2439 : node2434;
														assign node2434 = (inp[13]) ? 4'b0011 : node2435;
															assign node2435 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node2439 = (inp[2]) ? node2443 : node2440;
															assign node2440 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node2443 = (inp[13]) ? node2445 : 4'b0111;
																assign node2445 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node2448 = (inp[1]) ? node2464 : node2449;
														assign node2449 = (inp[0]) ? node2457 : node2450;
															assign node2450 = (inp[2]) ? node2454 : node2451;
																assign node2451 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node2454 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node2457 = (inp[13]) ? node2461 : node2458;
																assign node2458 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node2461 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node2464 = (inp[0]) ? node2470 : node2465;
															assign node2465 = (inp[13]) ? 4'b0010 : node2466;
																assign node2466 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node2470 = (inp[2]) ? node2474 : node2471;
																assign node2471 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node2474 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node2477 = (inp[11]) ? node2495 : node2478;
													assign node2478 = (inp[2]) ? node2486 : node2479;
														assign node2479 = (inp[13]) ? node2483 : node2480;
															assign node2480 = (inp[1]) ? 4'b0111 : 4'b0010;
															assign node2483 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node2486 = (inp[13]) ? node2492 : node2487;
															assign node2487 = (inp[1]) ? node2489 : 4'b0110;
																assign node2489 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node2492 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node2495 = (inp[1]) ? node2511 : node2496;
														assign node2496 = (inp[0]) ? node2504 : node2497;
															assign node2497 = (inp[2]) ? node2501 : node2498;
																assign node2498 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node2501 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node2504 = (inp[2]) ? node2508 : node2505;
																assign node2505 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node2508 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node2511 = (inp[13]) ? node2515 : node2512;
															assign node2512 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node2515 = (inp[2]) ? 4'b0110 : 4'b0010;
									assign node2518 = (inp[10]) ? node2688 : node2519;
										assign node2519 = (inp[0]) ? node2599 : node2520;
											assign node2520 = (inp[5]) ? node2558 : node2521;
												assign node2521 = (inp[2]) ? node2539 : node2522;
													assign node2522 = (inp[13]) ? node2530 : node2523;
														assign node2523 = (inp[1]) ? node2527 : node2524;
															assign node2524 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node2527 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node2530 = (inp[9]) ? 4'b0011 : node2531;
															assign node2531 = (inp[1]) ? node2535 : node2532;
																assign node2532 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node2535 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node2539 = (inp[13]) ? node2545 : node2540;
														assign node2540 = (inp[9]) ? node2542 : 4'b0011;
															assign node2542 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node2545 = (inp[11]) ? node2553 : node2546;
															assign node2546 = (inp[1]) ? node2550 : node2547;
																assign node2547 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node2550 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node2553 = (inp[1]) ? node2555 : 4'b0110;
																assign node2555 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node2558 = (inp[9]) ? node2580 : node2559;
													assign node2559 = (inp[13]) ? node2567 : node2560;
														assign node2560 = (inp[1]) ? node2564 : node2561;
															assign node2561 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node2564 = (inp[2]) ? 4'b0111 : 4'b0010;
														assign node2567 = (inp[11]) ? node2575 : node2568;
															assign node2568 = (inp[2]) ? node2572 : node2569;
																assign node2569 = (inp[1]) ? 4'b0110 : 4'b0011;
																assign node2572 = (inp[1]) ? 4'b0011 : 4'b0110;
															assign node2575 = (inp[1]) ? node2577 : 4'b0110;
																assign node2577 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node2580 = (inp[2]) ? node2590 : node2581;
														assign node2581 = (inp[1]) ? node2587 : node2582;
															assign node2582 = (inp[13]) ? 4'b0010 : node2583;
																assign node2583 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node2587 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node2590 = (inp[1]) ? node2594 : node2591;
															assign node2591 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node2594 = (inp[13]) ? node2596 : 4'b0110;
																assign node2596 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node2599 = (inp[9]) ? node2643 : node2600;
												assign node2600 = (inp[11]) ? node2620 : node2601;
													assign node2601 = (inp[13]) ? node2613 : node2602;
														assign node2602 = (inp[1]) ? node2606 : node2603;
															assign node2603 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node2606 = (inp[5]) ? node2610 : node2607;
																assign node2607 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node2610 = (inp[2]) ? 4'b0111 : 4'b0010;
														assign node2613 = (inp[1]) ? node2615 : 4'b0110;
															assign node2615 = (inp[5]) ? node2617 : 4'b0010;
																assign node2617 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node2620 = (inp[5]) ? node2636 : node2621;
														assign node2621 = (inp[1]) ? node2629 : node2622;
															assign node2622 = (inp[2]) ? node2626 : node2623;
																assign node2623 = (inp[13]) ? 4'b0011 : 4'b0111;
																assign node2626 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node2629 = (inp[2]) ? node2633 : node2630;
																assign node2630 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node2633 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node2636 = (inp[1]) ? node2638 : 4'b0111;
															assign node2638 = (inp[2]) ? node2640 : 4'b0111;
																assign node2640 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node2643 = (inp[11]) ? node2667 : node2644;
													assign node2644 = (inp[1]) ? node2654 : node2645;
														assign node2645 = (inp[2]) ? node2651 : node2646;
															assign node2646 = (inp[13]) ? 4'b0010 : node2647;
																assign node2647 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node2651 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node2654 = (inp[2]) ? node2662 : node2655;
															assign node2655 = (inp[5]) ? node2659 : node2656;
																assign node2656 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node2659 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node2662 = (inp[5]) ? 4'b0110 : node2663;
																assign node2663 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node2667 = (inp[13]) ? node2677 : node2668;
														assign node2668 = (inp[2]) ? node2672 : node2669;
															assign node2669 = (inp[1]) ? 4'b0010 : 4'b0110;
															assign node2672 = (inp[1]) ? 4'b0010 : node2673;
																assign node2673 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node2677 = (inp[5]) ? node2681 : node2678;
															assign node2678 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node2681 = (inp[1]) ? node2685 : node2682;
																assign node2682 = (inp[2]) ? 4'b0110 : 4'b0011;
																assign node2685 = (inp[2]) ? 4'b0011 : 4'b0110;
										assign node2688 = (inp[0]) ? node2772 : node2689;
											assign node2689 = (inp[11]) ? node2735 : node2690;
												assign node2690 = (inp[5]) ? node2714 : node2691;
													assign node2691 = (inp[1]) ? node2699 : node2692;
														assign node2692 = (inp[9]) ? 4'b0110 : node2693;
															assign node2693 = (inp[2]) ? node2695 : 4'b0011;
																assign node2695 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node2699 = (inp[2]) ? node2707 : node2700;
															assign node2700 = (inp[13]) ? node2704 : node2701;
																assign node2701 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node2704 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node2707 = (inp[9]) ? node2711 : node2708;
																assign node2708 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node2711 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node2714 = (inp[1]) ? node2722 : node2715;
														assign node2715 = (inp[9]) ? 4'b0011 : node2716;
															assign node2716 = (inp[2]) ? node2718 : 4'b0111;
																assign node2718 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node2722 = (inp[9]) ? node2730 : node2723;
															assign node2723 = (inp[2]) ? node2727 : node2724;
																assign node2724 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node2727 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node2730 = (inp[2]) ? node2732 : 4'b0010;
																assign node2732 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node2735 = (inp[1]) ? node2757 : node2736;
													assign node2736 = (inp[5]) ? node2748 : node2737;
														assign node2737 = (inp[9]) ? node2741 : node2738;
															assign node2738 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node2741 = (inp[2]) ? node2745 : node2742;
																assign node2742 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node2745 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node2748 = (inp[2]) ? node2754 : node2749;
															assign node2749 = (inp[9]) ? 4'b0111 : node2750;
																assign node2750 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node2754 = (inp[13]) ? 4'b0111 : 4'b0010;
													assign node2757 = (inp[2]) ? node2761 : node2758;
														assign node2758 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node2761 = (inp[13]) ? node2765 : node2762;
															assign node2762 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node2765 = (inp[5]) ? node2769 : node2766;
																assign node2766 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node2769 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node2772 = (inp[1]) ? node2820 : node2773;
												assign node2773 = (inp[5]) ? node2791 : node2774;
													assign node2774 = (inp[9]) ? node2784 : node2775;
														assign node2775 = (inp[2]) ? node2781 : node2776;
															assign node2776 = (inp[13]) ? 4'b0010 : node2777;
																assign node2777 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node2781 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node2784 = (inp[2]) ? node2788 : node2785;
															assign node2785 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node2788 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node2791 = (inp[9]) ? node2807 : node2792;
														assign node2792 = (inp[11]) ? node2800 : node2793;
															assign node2793 = (inp[2]) ? node2797 : node2794;
																assign node2794 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node2797 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node2800 = (inp[13]) ? node2804 : node2801;
																assign node2801 = (inp[2]) ? 4'b0010 : 4'b0110;
																assign node2804 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node2807 = (inp[11]) ? node2815 : node2808;
															assign node2808 = (inp[2]) ? node2812 : node2809;
																assign node2809 = (inp[13]) ? 4'b0011 : 4'b0111;
																assign node2812 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node2815 = (inp[2]) ? node2817 : 4'b0010;
																assign node2817 = (inp[13]) ? 4'b0111 : 4'b0011;
												assign node2820 = (inp[13]) ? node2848 : node2821;
													assign node2821 = (inp[9]) ? node2835 : node2822;
														assign node2822 = (inp[11]) ? node2830 : node2823;
															assign node2823 = (inp[2]) ? node2827 : node2824;
																assign node2824 = (inp[5]) ? 4'b0011 : 4'b0110;
																assign node2827 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node2830 = (inp[5]) ? 4'b0111 : node2831;
																assign node2831 = (inp[2]) ? 4'b0010 : 4'b0111;
														assign node2835 = (inp[11]) ? node2841 : node2836;
															assign node2836 = (inp[2]) ? node2838 : 4'b0111;
																assign node2838 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node2841 = (inp[2]) ? node2845 : node2842;
																assign node2842 = (inp[5]) ? 4'b0011 : 4'b0110;
																assign node2845 = (inp[5]) ? 4'b0110 : 4'b0011;
													assign node2848 = (inp[9]) ? node2854 : node2849;
														assign node2849 = (inp[5]) ? 4'b0011 : node2850;
															assign node2850 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node2854 = (inp[11]) ? node2858 : node2855;
															assign node2855 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node2858 = (inp[5]) ? node2860 : 4'b0111;
																assign node2860 = (inp[2]) ? 4'b0010 : 4'b0111;
								assign node2863 = (inp[4]) ? node3161 : node2864;
									assign node2864 = (inp[5]) ? node3018 : node2865;
										assign node2865 = (inp[13]) ? node2939 : node2866;
											assign node2866 = (inp[2]) ? node2904 : node2867;
												assign node2867 = (inp[0]) ? node2883 : node2868;
													assign node2868 = (inp[10]) ? node2878 : node2869;
														assign node2869 = (inp[11]) ? node2875 : node2870;
															assign node2870 = (inp[1]) ? node2872 : 4'b0010;
																assign node2872 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node2875 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node2878 = (inp[9]) ? node2880 : 4'b0011;
															assign node2880 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node2883 = (inp[11]) ? node2891 : node2884;
														assign node2884 = (inp[9]) ? node2888 : node2885;
															assign node2885 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node2888 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node2891 = (inp[9]) ? node2897 : node2892;
															assign node2892 = (inp[1]) ? 4'b0011 : node2893;
																assign node2893 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node2897 = (inp[1]) ? node2901 : node2898;
																assign node2898 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node2901 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node2904 = (inp[0]) ? node2924 : node2905;
													assign node2905 = (inp[9]) ? node2915 : node2906;
														assign node2906 = (inp[10]) ? node2912 : node2907;
															assign node2907 = (inp[11]) ? 4'b0110 : node2908;
																assign node2908 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node2912 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node2915 = (inp[11]) ? 4'b0111 : node2916;
															assign node2916 = (inp[10]) ? node2920 : node2917;
																assign node2917 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node2920 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node2924 = (inp[1]) ? node2926 : 4'b0111;
														assign node2926 = (inp[11]) ? node2932 : node2927;
															assign node2927 = (inp[9]) ? 4'b0111 : node2928;
																assign node2928 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node2932 = (inp[9]) ? node2936 : node2933;
																assign node2933 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node2936 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node2939 = (inp[2]) ? node2989 : node2940;
												assign node2940 = (inp[1]) ? node2970 : node2941;
													assign node2941 = (inp[0]) ? node2957 : node2942;
														assign node2942 = (inp[11]) ? node2950 : node2943;
															assign node2943 = (inp[10]) ? node2947 : node2944;
																assign node2944 = (inp[9]) ? 4'b0110 : 4'b0111;
																assign node2947 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node2950 = (inp[9]) ? node2954 : node2951;
																assign node2951 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node2954 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node2957 = (inp[9]) ? node2963 : node2958;
															assign node2958 = (inp[10]) ? 4'b0111 : node2959;
																assign node2959 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node2963 = (inp[11]) ? node2967 : node2964;
																assign node2964 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node2967 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node2970 = (inp[11]) ? node2982 : node2971;
														assign node2971 = (inp[10]) ? node2977 : node2972;
															assign node2972 = (inp[9]) ? node2974 : 4'b0111;
																assign node2974 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node2977 = (inp[9]) ? node2979 : 4'b0110;
																assign node2979 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node2982 = (inp[10]) ? node2986 : node2983;
															assign node2983 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node2986 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node2989 = (inp[0]) ? node3001 : node2990;
													assign node2990 = (inp[9]) ? node2992 : 4'b0010;
														assign node2992 = (inp[11]) ? node2994 : 4'b0010;
															assign node2994 = (inp[10]) ? node2998 : node2995;
																assign node2995 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node2998 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node3001 = (inp[9]) ? node3011 : node3002;
														assign node3002 = (inp[10]) ? node3006 : node3003;
															assign node3003 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node3006 = (inp[11]) ? 4'b0011 : node3007;
																assign node3007 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node3011 = (inp[1]) ? node3013 : 4'b0010;
															assign node3013 = (inp[11]) ? 4'b0010 : node3014;
																assign node3014 = (inp[10]) ? 4'b0011 : 4'b0010;
										assign node3018 = (inp[9]) ? node3080 : node3019;
											assign node3019 = (inp[2]) ? node3047 : node3020;
												assign node3020 = (inp[11]) ? node3036 : node3021;
													assign node3021 = (inp[13]) ? node3031 : node3022;
														assign node3022 = (inp[1]) ? node3026 : node3023;
															assign node3023 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node3026 = (inp[10]) ? 4'b0110 : node3027;
																assign node3027 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node3031 = (inp[1]) ? node3033 : 4'b0110;
															assign node3033 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node3036 = (inp[1]) ? node3040 : node3037;
														assign node3037 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node3040 = (inp[13]) ? node3042 : 4'b0110;
															assign node3042 = (inp[0]) ? 4'b0010 : node3043;
																assign node3043 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node3047 = (inp[10]) ? node3067 : node3048;
													assign node3048 = (inp[1]) ? node3056 : node3049;
														assign node3049 = (inp[13]) ? node3051 : 4'b0110;
															assign node3051 = (inp[0]) ? 4'b0010 : node3052;
																assign node3052 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node3056 = (inp[13]) ? node3062 : node3057;
															assign node3057 = (inp[11]) ? node3059 : 4'b0010;
																assign node3059 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node3062 = (inp[0]) ? node3064 : 4'b0111;
																assign node3064 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node3067 = (inp[1]) ? node3071 : node3068;
														assign node3068 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node3071 = (inp[13]) ? node3075 : node3072;
															assign node3072 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node3075 = (inp[0]) ? node3077 : 4'b0110;
																assign node3077 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node3080 = (inp[10]) ? node3122 : node3081;
												assign node3081 = (inp[13]) ? node3101 : node3082;
													assign node3082 = (inp[11]) ? node3088 : node3083;
														assign node3083 = (inp[1]) ? node3085 : 4'b0111;
															assign node3085 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node3088 = (inp[0]) ? node3094 : node3089;
															assign node3089 = (inp[1]) ? 4'b0111 : node3090;
																assign node3090 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node3094 = (inp[1]) ? node3098 : node3095;
																assign node3095 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node3098 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node3101 = (inp[0]) ? node3113 : node3102;
														assign node3102 = (inp[11]) ? node3108 : node3103;
															assign node3103 = (inp[2]) ? 4'b0010 : node3104;
																assign node3104 = (inp[1]) ? 4'b0010 : 4'b0110;
															assign node3108 = (inp[2]) ? 4'b0110 : node3109;
																assign node3109 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node3113 = (inp[11]) ? node3115 : 4'b0110;
															assign node3115 = (inp[1]) ? node3119 : node3116;
																assign node3116 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node3119 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node3122 = (inp[13]) ? node3142 : node3123;
													assign node3123 = (inp[11]) ? node3131 : node3124;
														assign node3124 = (inp[2]) ? node3128 : node3125;
															assign node3125 = (inp[1]) ? 4'b0110 : 4'b0010;
															assign node3128 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node3131 = (inp[0]) ? node3137 : node3132;
															assign node3132 = (inp[1]) ? node3134 : 4'b0010;
																assign node3134 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node3137 = (inp[1]) ? node3139 : 4'b0011;
																assign node3139 = (inp[2]) ? 4'b0011 : 4'b0110;
													assign node3142 = (inp[0]) ? node3152 : node3143;
														assign node3143 = (inp[2]) ? node3147 : node3144;
															assign node3144 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node3147 = (inp[1]) ? 4'b0111 : node3148;
																assign node3148 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node3152 = (inp[11]) ? node3156 : node3153;
															assign node3153 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node3156 = (inp[2]) ? node3158 : 4'b0110;
																assign node3158 = (inp[1]) ? 4'b0110 : 4'b0010;
									assign node3161 = (inp[0]) ? node3307 : node3162;
										assign node3162 = (inp[5]) ? node3228 : node3163;
											assign node3163 = (inp[9]) ? node3199 : node3164;
												assign node3164 = (inp[10]) ? node3186 : node3165;
													assign node3165 = (inp[2]) ? node3175 : node3166;
														assign node3166 = (inp[13]) ? node3172 : node3167;
															assign node3167 = (inp[1]) ? 4'b0000 : node3168;
																assign node3168 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node3172 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node3175 = (inp[13]) ? node3181 : node3176;
															assign node3176 = (inp[1]) ? 4'b0101 : node3177;
																assign node3177 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node3181 = (inp[11]) ? 4'b0001 : node3182;
																assign node3182 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node3186 = (inp[13]) ? node3192 : node3187;
														assign node3187 = (inp[2]) ? node3189 : 4'b0001;
															assign node3189 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node3192 = (inp[2]) ? node3194 : 4'b0100;
															assign node3194 = (inp[11]) ? 4'b0000 : node3195;
																assign node3195 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node3199 = (inp[10]) ? node3211 : node3200;
													assign node3200 = (inp[2]) ? node3208 : node3201;
														assign node3201 = (inp[13]) ? 4'b0100 : node3202;
															assign node3202 = (inp[1]) ? 4'b0001 : node3203;
																assign node3203 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node3208 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node3211 = (inp[2]) ? node3223 : node3212;
														assign node3212 = (inp[13]) ? node3218 : node3213;
															assign node3213 = (inp[1]) ? 4'b0000 : node3214;
																assign node3214 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node3218 = (inp[11]) ? node3220 : 4'b0101;
																assign node3220 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node3223 = (inp[13]) ? node3225 : 4'b0101;
															assign node3225 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node3228 = (inp[9]) ? node3268 : node3229;
												assign node3229 = (inp[10]) ? node3243 : node3230;
													assign node3230 = (inp[13]) ? node3238 : node3231;
														assign node3231 = (inp[2]) ? node3235 : node3232;
															assign node3232 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node3235 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node3238 = (inp[2]) ? node3240 : 4'b0000;
															assign node3240 = (inp[11]) ? 4'b0101 : 4'b0001;
													assign node3243 = (inp[11]) ? node3259 : node3244;
														assign node3244 = (inp[2]) ? node3252 : node3245;
															assign node3245 = (inp[1]) ? node3249 : node3246;
																assign node3246 = (inp[13]) ? 4'b0101 : 4'b0000;
																assign node3249 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node3252 = (inp[13]) ? node3256 : node3253;
																assign node3253 = (inp[1]) ? 4'b0001 : 4'b0101;
																assign node3256 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node3259 = (inp[13]) ? node3263 : node3260;
															assign node3260 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node3263 = (inp[2]) ? node3265 : 4'b0001;
																assign node3265 = (inp[1]) ? 4'b0100 : 4'b0001;
												assign node3268 = (inp[10]) ? node3286 : node3269;
													assign node3269 = (inp[13]) ? node3279 : node3270;
														assign node3270 = (inp[2]) ? node3276 : node3271;
															assign node3271 = (inp[1]) ? node3273 : 4'b0000;
																assign node3273 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node3276 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node3279 = (inp[2]) ? node3283 : node3280;
															assign node3280 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node3283 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node3286 = (inp[1]) ? node3294 : node3287;
														assign node3287 = (inp[2]) ? node3291 : node3288;
															assign node3288 = (inp[13]) ? 4'b0100 : 4'b0001;
															assign node3291 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node3294 = (inp[11]) ? node3302 : node3295;
															assign node3295 = (inp[13]) ? node3299 : node3296;
																assign node3296 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node3299 = (inp[2]) ? 4'b0101 : 4'b0000;
															assign node3302 = (inp[2]) ? 4'b0101 : node3303;
																assign node3303 = (inp[13]) ? 4'b0000 : 4'b0101;
										assign node3307 = (inp[10]) ? node3389 : node3308;
											assign node3308 = (inp[11]) ? node3356 : node3309;
												assign node3309 = (inp[2]) ? node3329 : node3310;
													assign node3310 = (inp[13]) ? node3318 : node3311;
														assign node3311 = (inp[9]) ? node3315 : node3312;
															assign node3312 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node3315 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node3318 = (inp[1]) ? node3322 : node3319;
															assign node3319 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node3322 = (inp[5]) ? node3326 : node3323;
																assign node3323 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node3326 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node3329 = (inp[13]) ? node3345 : node3330;
														assign node3330 = (inp[5]) ? node3338 : node3331;
															assign node3331 = (inp[9]) ? node3335 : node3332;
																assign node3332 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node3335 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node3338 = (inp[1]) ? node3342 : node3339;
																assign node3339 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node3342 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node3345 = (inp[5]) ? node3349 : node3346;
															assign node3346 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node3349 = (inp[1]) ? node3353 : node3350;
																assign node3350 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node3353 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node3356 = (inp[9]) ? node3376 : node3357;
													assign node3357 = (inp[13]) ? node3367 : node3358;
														assign node3358 = (inp[5]) ? node3362 : node3359;
															assign node3359 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node3362 = (inp[2]) ? node3364 : 4'b0101;
																assign node3364 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node3367 = (inp[2]) ? node3371 : node3368;
															assign node3368 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node3371 = (inp[5]) ? node3373 : 4'b0001;
																assign node3373 = (inp[1]) ? 4'b0100 : 4'b0000;
													assign node3376 = (inp[13]) ? node3380 : node3377;
														assign node3377 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node3380 = (inp[2]) ? node3384 : node3381;
															assign node3381 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node3384 = (inp[1]) ? node3386 : 4'b0001;
																assign node3386 = (inp[5]) ? 4'b0101 : 4'b0000;
											assign node3389 = (inp[13]) ? node3425 : node3390;
												assign node3390 = (inp[2]) ? node3410 : node3391;
													assign node3391 = (inp[9]) ? node3401 : node3392;
														assign node3392 = (inp[1]) ? node3398 : node3393;
															assign node3393 = (inp[11]) ? node3395 : 4'b0000;
																assign node3395 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node3398 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node3401 = (inp[5]) ? node3405 : node3402;
															assign node3402 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node3405 = (inp[1]) ? 4'b0101 : node3406;
																assign node3406 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node3410 = (inp[5]) ? node3420 : node3411;
														assign node3411 = (inp[9]) ? node3415 : node3412;
															assign node3412 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node3415 = (inp[11]) ? 4'b0100 : node3416;
																assign node3416 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node3420 = (inp[1]) ? node3422 : 4'b0100;
															assign node3422 = (inp[9]) ? 4'b0001 : 4'b0000;
												assign node3425 = (inp[2]) ? node3449 : node3426;
													assign node3426 = (inp[1]) ? node3438 : node3427;
														assign node3427 = (inp[9]) ? node3433 : node3428;
															assign node3428 = (inp[5]) ? node3430 : 4'b0101;
																assign node3430 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node3433 = (inp[11]) ? node3435 : 4'b0100;
																assign node3435 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node3438 = (inp[5]) ? node3442 : node3439;
															assign node3439 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node3442 = (inp[11]) ? node3446 : node3443;
																assign node3443 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node3446 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node3449 = (inp[5]) ? node3455 : node3450;
														assign node3450 = (inp[9]) ? 4'b0001 : node3451;
															assign node3451 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node3455 = (inp[1]) ? node3459 : node3456;
															assign node3456 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node3459 = (inp[9]) ? node3461 : 4'b0101;
																assign node3461 = (inp[11]) ? 4'b0100 : 4'b0101;
							assign node3464 = (inp[4]) ? node4116 : node3465;
								assign node3465 = (inp[9]) ? node3781 : node3466;
									assign node3466 = (inp[13]) ? node3618 : node3467;
										assign node3467 = (inp[15]) ? node3543 : node3468;
											assign node3468 = (inp[2]) ? node3502 : node3469;
												assign node3469 = (inp[1]) ? node3485 : node3470;
													assign node3470 = (inp[5]) ? node3482 : node3471;
														assign node3471 = (inp[10]) ? node3477 : node3472;
															assign node3472 = (inp[11]) ? 4'b0001 : node3473;
																assign node3473 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node3477 = (inp[0]) ? 4'b0000 : node3478;
																assign node3478 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node3482 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node3485 = (inp[11]) ? node3497 : node3486;
														assign node3486 = (inp[0]) ? node3492 : node3487;
															assign node3487 = (inp[5]) ? node3489 : 4'b0100;
																assign node3489 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node3492 = (inp[5]) ? node3494 : 4'b0101;
																assign node3494 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node3497 = (inp[0]) ? node3499 : 4'b0101;
															assign node3499 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node3502 = (inp[5]) ? node3520 : node3503;
													assign node3503 = (inp[1]) ? node3511 : node3504;
														assign node3504 = (inp[10]) ? node3506 : 4'b0101;
															assign node3506 = (inp[11]) ? 4'b0100 : node3507;
																assign node3507 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node3511 = (inp[10]) ? node3517 : node3512;
															assign node3512 = (inp[0]) ? node3514 : 4'b0000;
																assign node3514 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node3517 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node3520 = (inp[1]) ? node3532 : node3521;
														assign node3521 = (inp[10]) ? node3527 : node3522;
															assign node3522 = (inp[11]) ? node3524 : 4'b0000;
																assign node3524 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node3527 = (inp[0]) ? node3529 : 4'b0001;
																assign node3529 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node3532 = (inp[10]) ? node3538 : node3533;
															assign node3533 = (inp[11]) ? node3535 : 4'b0001;
																assign node3535 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node3538 = (inp[0]) ? node3540 : 4'b0000;
																assign node3540 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node3543 = (inp[2]) ? node3573 : node3544;
												assign node3544 = (inp[5]) ? node3556 : node3545;
													assign node3545 = (inp[1]) ? node3551 : node3546;
														assign node3546 = (inp[10]) ? 4'b0100 : node3547;
															assign node3547 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node3551 = (inp[10]) ? 4'b0000 : node3552;
															assign node3552 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node3556 = (inp[10]) ? node3564 : node3557;
														assign node3557 = (inp[0]) ? 4'b0001 : node3558;
															assign node3558 = (inp[1]) ? node3560 : 4'b0000;
																assign node3560 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node3564 = (inp[0]) ? node3570 : node3565;
															assign node3565 = (inp[1]) ? node3567 : 4'b0001;
																assign node3567 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node3570 = (inp[1]) ? 4'b0001 : 4'b0000;
												assign node3573 = (inp[1]) ? node3591 : node3574;
													assign node3574 = (inp[5]) ? node3586 : node3575;
														assign node3575 = (inp[10]) ? node3581 : node3576;
															assign node3576 = (inp[0]) ? node3578 : 4'b0001;
																assign node3578 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node3581 = (inp[0]) ? node3583 : 4'b0000;
																assign node3583 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node3586 = (inp[10]) ? node3588 : 4'b0100;
															assign node3588 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node3591 = (inp[11]) ? node3605 : node3592;
														assign node3592 = (inp[5]) ? node3598 : node3593;
															assign node3593 = (inp[10]) ? 4'b0101 : node3594;
																assign node3594 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node3598 = (inp[10]) ? node3602 : node3599;
																assign node3599 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node3602 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node3605 = (inp[0]) ? node3613 : node3606;
															assign node3606 = (inp[10]) ? node3610 : node3607;
																assign node3607 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node3610 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node3613 = (inp[10]) ? 4'b0100 : node3614;
																assign node3614 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node3618 = (inp[1]) ? node3686 : node3619;
											assign node3619 = (inp[15]) ? node3653 : node3620;
												assign node3620 = (inp[10]) ? node3638 : node3621;
													assign node3621 = (inp[0]) ? node3629 : node3622;
														assign node3622 = (inp[5]) ? node3626 : node3623;
															assign node3623 = (inp[2]) ? 4'b0001 : 4'b0100;
															assign node3626 = (inp[11]) ? 4'b0100 : 4'b0000;
														assign node3629 = (inp[2]) ? node3633 : node3630;
															assign node3630 = (inp[5]) ? 4'b0001 : 4'b0101;
															assign node3633 = (inp[5]) ? node3635 : 4'b0000;
																assign node3635 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node3638 = (inp[11]) ? node3646 : node3639;
														assign node3639 = (inp[0]) ? 4'b0001 : node3640;
															assign node3640 = (inp[2]) ? node3642 : 4'b0101;
																assign node3642 = (inp[5]) ? 4'b0101 : 4'b0000;
														assign node3646 = (inp[5]) ? node3648 : 4'b0100;
															assign node3648 = (inp[2]) ? 4'b0100 : node3649;
																assign node3649 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node3653 = (inp[5]) ? node3669 : node3654;
													assign node3654 = (inp[2]) ? node3664 : node3655;
														assign node3655 = (inp[10]) ? node3659 : node3656;
															assign node3656 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node3659 = (inp[11]) ? node3661 : 4'b0001;
																assign node3661 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node3664 = (inp[10]) ? 4'b0101 : node3665;
															assign node3665 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node3669 = (inp[2]) ? node3677 : node3670;
														assign node3670 = (inp[10]) ? 4'b0100 : node3671;
															assign node3671 = (inp[0]) ? node3673 : 4'b0101;
																assign node3673 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node3677 = (inp[11]) ? 4'b0001 : node3678;
															assign node3678 = (inp[10]) ? node3682 : node3679;
																assign node3679 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node3682 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node3686 = (inp[10]) ? node3732 : node3687;
												assign node3687 = (inp[5]) ? node3705 : node3688;
													assign node3688 = (inp[0]) ? node3696 : node3689;
														assign node3689 = (inp[15]) ? node3691 : 4'b0000;
															assign node3691 = (inp[2]) ? 4'b0000 : node3692;
																assign node3692 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node3696 = (inp[11]) ? node3698 : 4'b0000;
															assign node3698 = (inp[2]) ? node3702 : node3699;
																assign node3699 = (inp[15]) ? 4'b0100 : 4'b0001;
																assign node3702 = (inp[15]) ? 4'b0001 : 4'b0101;
													assign node3705 = (inp[0]) ? node3719 : node3706;
														assign node3706 = (inp[11]) ? node3712 : node3707;
															assign node3707 = (inp[2]) ? node3709 : 4'b0001;
																assign node3709 = (inp[15]) ? 4'b0001 : 4'b0101;
															assign node3712 = (inp[2]) ? node3716 : node3713;
																assign node3713 = (inp[15]) ? 4'b0101 : 4'b0001;
																assign node3716 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node3719 = (inp[11]) ? node3725 : node3720;
															assign node3720 = (inp[15]) ? 4'b0001 : node3721;
																assign node3721 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node3725 = (inp[2]) ? node3729 : node3726;
																assign node3726 = (inp[15]) ? 4'b0101 : 4'b0000;
																assign node3729 = (inp[15]) ? 4'b0000 : 4'b0100;
												assign node3732 = (inp[5]) ? node3760 : node3733;
													assign node3733 = (inp[0]) ? node3747 : node3734;
														assign node3734 = (inp[11]) ? node3740 : node3735;
															assign node3735 = (inp[2]) ? 4'b0001 : node3736;
																assign node3736 = (inp[15]) ? 4'b0100 : 4'b0001;
															assign node3740 = (inp[2]) ? node3744 : node3741;
																assign node3741 = (inp[15]) ? 4'b0101 : 4'b0001;
																assign node3744 = (inp[15]) ? 4'b0001 : 4'b0101;
														assign node3747 = (inp[11]) ? node3753 : node3748;
															assign node3748 = (inp[15]) ? node3750 : 4'b0001;
																assign node3750 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node3753 = (inp[2]) ? node3757 : node3754;
																assign node3754 = (inp[15]) ? 4'b0101 : 4'b0000;
																assign node3757 = (inp[15]) ? 4'b0000 : 4'b0100;
													assign node3760 = (inp[11]) ? node3774 : node3761;
														assign node3761 = (inp[0]) ? node3767 : node3762;
															assign node3762 = (inp[15]) ? 4'b0101 : node3763;
																assign node3763 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node3767 = (inp[15]) ? node3771 : node3768;
																assign node3768 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node3771 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node3774 = (inp[0]) ? 4'b0001 : node3775;
															assign node3775 = (inp[15]) ? 4'b0000 : node3776;
																assign node3776 = (inp[2]) ? 4'b0100 : 4'b0000;
									assign node3781 = (inp[0]) ? node3955 : node3782;
										assign node3782 = (inp[10]) ? node3874 : node3783;
											assign node3783 = (inp[1]) ? node3835 : node3784;
												assign node3784 = (inp[5]) ? node3816 : node3785;
													assign node3785 = (inp[11]) ? node3801 : node3786;
														assign node3786 = (inp[2]) ? node3794 : node3787;
															assign node3787 = (inp[15]) ? node3791 : node3788;
																assign node3788 = (inp[13]) ? 4'b0101 : 4'b0001;
																assign node3791 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node3794 = (inp[13]) ? node3798 : node3795;
																assign node3795 = (inp[15]) ? 4'b0000 : 4'b0101;
																assign node3798 = (inp[15]) ? 4'b0101 : 4'b0000;
														assign node3801 = (inp[13]) ? node3809 : node3802;
															assign node3802 = (inp[2]) ? node3806 : node3803;
																assign node3803 = (inp[15]) ? 4'b0100 : 4'b0000;
																assign node3806 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node3809 = (inp[15]) ? node3813 : node3810;
																assign node3810 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node3813 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node3816 = (inp[2]) ? node3824 : node3817;
														assign node3817 = (inp[11]) ? node3819 : 4'b0100;
															assign node3819 = (inp[15]) ? 4'b0100 : node3820;
																assign node3820 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node3824 = (inp[11]) ? node3830 : node3825;
															assign node3825 = (inp[15]) ? 4'b0000 : node3826;
																assign node3826 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node3830 = (inp[13]) ? node3832 : 4'b0101;
																assign node3832 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node3835 = (inp[5]) ? node3853 : node3836;
													assign node3836 = (inp[15]) ? node3846 : node3837;
														assign node3837 = (inp[2]) ? node3843 : node3838;
															assign node3838 = (inp[13]) ? 4'b0001 : node3839;
																assign node3839 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node3843 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node3846 = (inp[13]) ? node3850 : node3847;
															assign node3847 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node3850 = (inp[2]) ? 4'b0001 : 4'b0100;
													assign node3853 = (inp[15]) ? node3863 : node3854;
														assign node3854 = (inp[13]) ? node3860 : node3855;
															assign node3855 = (inp[2]) ? 4'b0000 : node3856;
																assign node3856 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node3860 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node3863 = (inp[13]) ? node3869 : node3864;
															assign node3864 = (inp[11]) ? node3866 : 4'b0000;
																assign node3866 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node3869 = (inp[2]) ? 4'b0000 : node3870;
																assign node3870 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node3874 = (inp[11]) ? node3910 : node3875;
												assign node3875 = (inp[5]) ? node3895 : node3876;
													assign node3876 = (inp[2]) ? node3884 : node3877;
														assign node3877 = (inp[1]) ? 4'b0101 : node3878;
															assign node3878 = (inp[13]) ? node3880 : 4'b0100;
																assign node3880 = (inp[15]) ? 4'b0000 : 4'b0100;
														assign node3884 = (inp[1]) ? node3888 : node3885;
															assign node3885 = (inp[15]) ? 4'b0001 : 4'b0100;
															assign node3888 = (inp[15]) ? node3892 : node3889;
																assign node3889 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node3892 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node3895 = (inp[1]) ? node3907 : node3896;
														assign node3896 = (inp[15]) ? node3900 : node3897;
															assign node3897 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node3900 = (inp[13]) ? node3904 : node3901;
																assign node3901 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node3904 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node3907 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node3910 = (inp[5]) ? node3936 : node3911;
													assign node3911 = (inp[1]) ? node3923 : node3912;
														assign node3912 = (inp[13]) ? node3918 : node3913;
															assign node3913 = (inp[2]) ? node3915 : 4'b0001;
																assign node3915 = (inp[15]) ? 4'b0001 : 4'b0101;
															assign node3918 = (inp[15]) ? node3920 : 4'b0001;
																assign node3920 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node3923 = (inp[13]) ? node3929 : node3924;
															assign node3924 = (inp[15]) ? 4'b0001 : node3925;
																assign node3925 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node3929 = (inp[15]) ? node3933 : node3930;
																assign node3930 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node3933 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node3936 = (inp[13]) ? node3944 : node3937;
														assign node3937 = (inp[2]) ? node3941 : node3938;
															assign node3938 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node3941 = (inp[15]) ? 4'b0100 : 4'b0000;
														assign node3944 = (inp[1]) ? node3952 : node3945;
															assign node3945 = (inp[2]) ? node3949 : node3946;
																assign node3946 = (inp[15]) ? 4'b0101 : 4'b0000;
																assign node3949 = (inp[15]) ? 4'b0000 : 4'b0100;
															assign node3952 = (inp[15]) ? 4'b0001 : 4'b0101;
										assign node3955 = (inp[13]) ? node4043 : node3956;
											assign node3956 = (inp[15]) ? node3996 : node3957;
												assign node3957 = (inp[2]) ? node3977 : node3958;
													assign node3958 = (inp[5]) ? node3966 : node3959;
														assign node3959 = (inp[1]) ? node3963 : node3960;
															assign node3960 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node3963 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node3966 = (inp[11]) ? node3972 : node3967;
															assign node3967 = (inp[1]) ? 4'b0100 : node3968;
																assign node3968 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node3972 = (inp[1]) ? node3974 : 4'b0101;
																assign node3974 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node3977 = (inp[1]) ? node3987 : node3978;
														assign node3978 = (inp[5]) ? node3982 : node3979;
															assign node3979 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node3982 = (inp[10]) ? node3984 : 4'b0001;
																assign node3984 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node3987 = (inp[5]) ? 4'b0001 : node3988;
															assign node3988 = (inp[10]) ? node3992 : node3989;
																assign node3989 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node3992 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node3996 = (inp[2]) ? node4012 : node3997;
													assign node3997 = (inp[5]) ? node4005 : node3998;
														assign node3998 = (inp[10]) ? node4002 : node3999;
															assign node3999 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node4002 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node4005 = (inp[10]) ? 4'b0000 : node4006;
															assign node4006 = (inp[11]) ? node4008 : 4'b0001;
																assign node4008 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node4012 = (inp[1]) ? node4028 : node4013;
														assign node4013 = (inp[5]) ? node4021 : node4014;
															assign node4014 = (inp[11]) ? node4018 : node4015;
																assign node4015 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node4018 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node4021 = (inp[11]) ? node4025 : node4022;
																assign node4022 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node4025 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node4028 = (inp[11]) ? node4036 : node4029;
															assign node4029 = (inp[10]) ? node4033 : node4030;
																assign node4030 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node4033 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node4036 = (inp[10]) ? node4040 : node4037;
																assign node4037 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node4040 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node4043 = (inp[5]) ? node4083 : node4044;
												assign node4044 = (inp[2]) ? node4066 : node4045;
													assign node4045 = (inp[11]) ? node4057 : node4046;
														assign node4046 = (inp[10]) ? node4050 : node4047;
															assign node4047 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node4050 = (inp[15]) ? node4054 : node4051;
																assign node4051 = (inp[1]) ? 4'b0000 : 4'b0101;
																assign node4054 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node4057 = (inp[10]) ? 4'b0001 : node4058;
															assign node4058 = (inp[1]) ? node4062 : node4059;
																assign node4059 = (inp[15]) ? 4'b0000 : 4'b0100;
																assign node4062 = (inp[15]) ? 4'b0101 : 4'b0000;
													assign node4066 = (inp[15]) ? node4074 : node4067;
														assign node4067 = (inp[1]) ? node4069 : 4'b0001;
															assign node4069 = (inp[11]) ? node4071 : 4'b0101;
																assign node4071 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node4074 = (inp[1]) ? node4078 : node4075;
															assign node4075 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node4078 = (inp[11]) ? 4'b0000 : node4079;
																assign node4079 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node4083 = (inp[11]) ? node4105 : node4084;
													assign node4084 = (inp[15]) ? node4094 : node4085;
														assign node4085 = (inp[2]) ? 4'b0100 : node4086;
															assign node4086 = (inp[1]) ? node4090 : node4087;
																assign node4087 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node4090 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node4094 = (inp[2]) ? node4098 : node4095;
															assign node4095 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node4098 = (inp[1]) ? node4102 : node4099;
																assign node4099 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node4102 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node4105 = (inp[15]) ? node4111 : node4106;
														assign node4106 = (inp[2]) ? 4'b0100 : node4107;
															assign node4107 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node4111 = (inp[2]) ? node4113 : 4'b0100;
															assign node4113 = (inp[10]) ? 4'b0000 : 4'b0001;
								assign node4116 = (inp[15]) ? node4420 : node4117;
									assign node4117 = (inp[10]) ? node4285 : node4118;
										assign node4118 = (inp[5]) ? node4190 : node4119;
											assign node4119 = (inp[2]) ? node4147 : node4120;
												assign node4120 = (inp[1]) ? node4130 : node4121;
													assign node4121 = (inp[13]) ? 4'b0000 : node4122;
														assign node4122 = (inp[9]) ? node4124 : 4'b0101;
															assign node4124 = (inp[0]) ? 4'b0100 : node4125;
																assign node4125 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node4130 = (inp[13]) ? node4138 : node4131;
														assign node4131 = (inp[9]) ? node4133 : 4'b0000;
															assign node4133 = (inp[11]) ? node4135 : 4'b0001;
																assign node4135 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node4138 = (inp[9]) ? node4142 : node4139;
															assign node4139 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node4142 = (inp[11]) ? node4144 : 4'b0101;
																assign node4144 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node4147 = (inp[11]) ? node4165 : node4148;
													assign node4148 = (inp[9]) ? node4158 : node4149;
														assign node4149 = (inp[1]) ? node4153 : node4150;
															assign node4150 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node4153 = (inp[13]) ? node4155 : 4'b0101;
																assign node4155 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node4158 = (inp[1]) ? node4162 : node4159;
															assign node4159 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node4162 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node4165 = (inp[9]) ? node4177 : node4166;
														assign node4166 = (inp[13]) ? node4172 : node4167;
															assign node4167 = (inp[1]) ? node4169 : 4'b0001;
																assign node4169 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node4172 = (inp[1]) ? 4'b0000 : node4173;
																assign node4173 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node4177 = (inp[1]) ? node4185 : node4178;
															assign node4178 = (inp[13]) ? node4182 : node4179;
																assign node4179 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node4182 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node4185 = (inp[13]) ? 4'b0001 : node4186;
																assign node4186 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node4190 = (inp[9]) ? node4238 : node4191;
												assign node4191 = (inp[11]) ? node4217 : node4192;
													assign node4192 = (inp[1]) ? node4206 : node4193;
														assign node4193 = (inp[2]) ? node4201 : node4194;
															assign node4194 = (inp[13]) ? node4198 : node4195;
																assign node4195 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node4198 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node4201 = (inp[0]) ? node4203 : 4'b0101;
																assign node4203 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node4206 = (inp[0]) ? node4210 : node4207;
															assign node4207 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node4210 = (inp[2]) ? node4214 : node4211;
																assign node4211 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node4214 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node4217 = (inp[0]) ? node4229 : node4218;
														assign node4218 = (inp[1]) ? node4224 : node4219;
															assign node4219 = (inp[2]) ? 4'b0100 : node4220;
																assign node4220 = (inp[13]) ? 4'b0101 : 4'b0001;
															assign node4224 = (inp[2]) ? node4226 : 4'b0100;
																assign node4226 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node4229 = (inp[1]) ? node4235 : node4230;
															assign node4230 = (inp[13]) ? node4232 : 4'b0001;
																assign node4232 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node4235 = (inp[13]) ? 4'b0000 : 4'b0101;
												assign node4238 = (inp[11]) ? node4260 : node4239;
													assign node4239 = (inp[0]) ? node4247 : node4240;
														assign node4240 = (inp[1]) ? node4242 : 4'b0001;
															assign node4242 = (inp[2]) ? node4244 : 4'b0000;
																assign node4244 = (inp[13]) ? 4'b0000 : 4'b0101;
														assign node4247 = (inp[13]) ? node4255 : node4248;
															assign node4248 = (inp[2]) ? node4252 : node4249;
																assign node4249 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node4252 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node4255 = (inp[2]) ? 4'b0001 : node4256;
																assign node4256 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node4260 = (inp[0]) ? node4276 : node4261;
														assign node4261 = (inp[13]) ? node4269 : node4262;
															assign node4262 = (inp[2]) ? node4266 : node4263;
																assign node4263 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node4266 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node4269 = (inp[2]) ? node4273 : node4270;
																assign node4270 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node4273 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node4276 = (inp[1]) ? node4282 : node4277;
															assign node4277 = (inp[2]) ? 4'b0000 : node4278;
																assign node4278 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node4282 = (inp[13]) ? 4'b0001 : 4'b0100;
										assign node4285 = (inp[2]) ? node4347 : node4286;
											assign node4286 = (inp[13]) ? node4318 : node4287;
												assign node4287 = (inp[1]) ? node4305 : node4288;
													assign node4288 = (inp[5]) ? node4298 : node4289;
														assign node4289 = (inp[0]) ? 4'b0101 : node4290;
															assign node4290 = (inp[11]) ? node4294 : node4291;
																assign node4291 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node4294 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node4298 = (inp[11]) ? 4'b0000 : node4299;
															assign node4299 = (inp[0]) ? node4301 : 4'b0001;
																assign node4301 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node4305 = (inp[11]) ? node4307 : 4'b0001;
														assign node4307 = (inp[9]) ? node4313 : node4308;
															assign node4308 = (inp[5]) ? 4'b0001 : node4309;
																assign node4309 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node4313 = (inp[5]) ? 4'b0000 : node4314;
																assign node4314 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node4318 = (inp[1]) ? node4332 : node4319;
													assign node4319 = (inp[5]) ? node4325 : node4320;
														assign node4320 = (inp[9]) ? 4'b0001 : node4321;
															assign node4321 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node4325 = (inp[11]) ? 4'b0101 : node4326;
															assign node4326 = (inp[9]) ? 4'b0100 : node4327;
																assign node4327 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node4332 = (inp[9]) ? node4338 : node4333;
														assign node4333 = (inp[0]) ? node4335 : 4'b0101;
															assign node4335 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node4338 = (inp[0]) ? node4344 : node4339;
															assign node4339 = (inp[11]) ? 4'b0100 : node4340;
																assign node4340 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node4344 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node4347 = (inp[13]) ? node4383 : node4348;
												assign node4348 = (inp[5]) ? node4366 : node4349;
													assign node4349 = (inp[1]) ? node4361 : node4350;
														assign node4350 = (inp[9]) ? node4356 : node4351;
															assign node4351 = (inp[11]) ? node4353 : 4'b0001;
																assign node4353 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node4356 = (inp[11]) ? node4358 : 4'b0000;
																assign node4358 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node4361 = (inp[9]) ? 4'b0101 : node4362;
															assign node4362 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node4366 = (inp[11]) ? node4378 : node4367;
														assign node4367 = (inp[9]) ? node4373 : node4368;
															assign node4368 = (inp[1]) ? 4'b0101 : node4369;
																assign node4369 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node4373 = (inp[0]) ? node4375 : 4'b0100;
																assign node4375 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node4378 = (inp[9]) ? 4'b0101 : node4379;
															assign node4379 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node4383 = (inp[1]) ? node4403 : node4384;
													assign node4384 = (inp[5]) ? node4392 : node4385;
														assign node4385 = (inp[11]) ? node4387 : 4'b0101;
															assign node4387 = (inp[0]) ? node4389 : 4'b0101;
																assign node4389 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node4392 = (inp[9]) ? node4398 : node4393;
															assign node4393 = (inp[0]) ? node4395 : 4'b0001;
																assign node4395 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node4398 = (inp[11]) ? node4400 : 4'b0000;
																assign node4400 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node4403 = (inp[5]) ? node4415 : node4404;
														assign node4404 = (inp[9]) ? node4410 : node4405;
															assign node4405 = (inp[0]) ? 4'b0001 : node4406;
																assign node4406 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node4410 = (inp[0]) ? 4'b0000 : node4411;
																assign node4411 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node4415 = (inp[9]) ? node4417 : 4'b0000;
															assign node4417 = (inp[0]) ? 4'b0000 : 4'b0001;
									assign node4420 = (inp[10]) ? node4574 : node4421;
										assign node4421 = (inp[11]) ? node4491 : node4422;
											assign node4422 = (inp[5]) ? node4456 : node4423;
												assign node4423 = (inp[0]) ? node4433 : node4424;
													assign node4424 = (inp[13]) ? node4428 : node4425;
														assign node4425 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node4428 = (inp[2]) ? 4'b0111 : node4429;
															assign node4429 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node4433 = (inp[13]) ? node4445 : node4434;
														assign node4434 = (inp[2]) ? node4438 : node4435;
															assign node4435 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node4438 = (inp[9]) ? node4442 : node4439;
																assign node4439 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node4442 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node4445 = (inp[2]) ? node4451 : node4446;
															assign node4446 = (inp[9]) ? node4448 : 4'b0010;
																assign node4448 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node4451 = (inp[9]) ? 4'b0110 : node4452;
																assign node4452 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node4456 = (inp[13]) ? node4478 : node4457;
													assign node4457 = (inp[9]) ? node4469 : node4458;
														assign node4458 = (inp[1]) ? node4464 : node4459;
															assign node4459 = (inp[2]) ? 4'b0010 : node4460;
																assign node4460 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node4464 = (inp[2]) ? node4466 : 4'b0011;
																assign node4466 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node4469 = (inp[2]) ? node4475 : node4470;
															assign node4470 = (inp[0]) ? 4'b0010 : node4471;
																assign node4471 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node4475 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node4478 = (inp[9]) ? node4482 : node4479;
														assign node4479 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node4482 = (inp[2]) ? node4488 : node4483;
															assign node4483 = (inp[1]) ? node4485 : 4'b0011;
																assign node4485 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node4488 = (inp[1]) ? 4'b0010 : 4'b0110;
											assign node4491 = (inp[9]) ? node4535 : node4492;
												assign node4492 = (inp[5]) ? node4514 : node4493;
													assign node4493 = (inp[1]) ? node4501 : node4494;
														assign node4494 = (inp[13]) ? 4'b0011 : node4495;
															assign node4495 = (inp[2]) ? 4'b0011 : node4496;
																assign node4496 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node4501 = (inp[13]) ? node4507 : node4502;
															assign node4502 = (inp[2]) ? node4504 : 4'b0111;
																assign node4504 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node4507 = (inp[2]) ? node4511 : node4508;
																assign node4508 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node4511 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node4514 = (inp[2]) ? node4522 : node4515;
														assign node4515 = (inp[0]) ? node4517 : 4'b0010;
															assign node4517 = (inp[1]) ? node4519 : 4'b0011;
																assign node4519 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node4522 = (inp[0]) ? node4530 : node4523;
															assign node4523 = (inp[13]) ? node4527 : node4524;
																assign node4524 = (inp[1]) ? 4'b0110 : 4'b0010;
																assign node4527 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node4530 = (inp[13]) ? node4532 : 4'b0011;
																assign node4532 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node4535 = (inp[13]) ? node4553 : node4536;
													assign node4536 = (inp[2]) ? node4546 : node4537;
														assign node4537 = (inp[5]) ? node4543 : node4538;
															assign node4538 = (inp[0]) ? node4540 : 4'b0110;
																assign node4540 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node4543 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node4546 = (inp[0]) ? 4'b0010 : node4547;
															assign node4547 = (inp[1]) ? 4'b0011 : node4548;
																assign node4548 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node4553 = (inp[2]) ? node4565 : node4554;
														assign node4554 = (inp[5]) ? node4560 : node4555;
															assign node4555 = (inp[1]) ? node4557 : 4'b0010;
																assign node4557 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node4560 = (inp[1]) ? 4'b0111 : node4561;
																assign node4561 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node4565 = (inp[5]) ? node4567 : 4'b0111;
															assign node4567 = (inp[0]) ? node4571 : node4568;
																assign node4568 = (inp[1]) ? 4'b0010 : 4'b0110;
																assign node4571 = (inp[1]) ? 4'b0011 : 4'b0111;
										assign node4574 = (inp[11]) ? node4656 : node4575;
											assign node4575 = (inp[0]) ? node4615 : node4576;
												assign node4576 = (inp[9]) ? node4594 : node4577;
													assign node4577 = (inp[1]) ? node4585 : node4578;
														assign node4578 = (inp[2]) ? node4582 : node4579;
															assign node4579 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node4582 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node4585 = (inp[5]) ? node4587 : 4'b0011;
															assign node4587 = (inp[2]) ? node4591 : node4588;
																assign node4588 = (inp[13]) ? 4'b0110 : 4'b0011;
																assign node4591 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node4594 = (inp[13]) ? node4606 : node4595;
														assign node4595 = (inp[2]) ? node4601 : node4596;
															assign node4596 = (inp[1]) ? node4598 : 4'b0111;
																assign node4598 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node4601 = (inp[5]) ? node4603 : 4'b0010;
																assign node4603 = (inp[1]) ? 4'b0111 : 4'b0010;
														assign node4606 = (inp[2]) ? node4612 : node4607;
															assign node4607 = (inp[1]) ? node4609 : 4'b0010;
																assign node4609 = (inp[5]) ? 4'b0111 : 4'b0010;
															assign node4612 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node4615 = (inp[9]) ? node4635 : node4616;
													assign node4616 = (inp[2]) ? node4624 : node4617;
														assign node4617 = (inp[13]) ? node4619 : 4'b0110;
															assign node4619 = (inp[5]) ? node4621 : 4'b0011;
																assign node4621 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node4624 = (inp[13]) ? node4630 : node4625;
															assign node4625 = (inp[5]) ? 4'b0011 : node4626;
																assign node4626 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node4630 = (inp[5]) ? node4632 : 4'b0110;
																assign node4632 = (inp[1]) ? 4'b0010 : 4'b0110;
													assign node4635 = (inp[2]) ? node4643 : node4636;
														assign node4636 = (inp[13]) ? node4640 : node4637;
															assign node4637 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node4640 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node4643 = (inp[13]) ? node4649 : node4644;
															assign node4644 = (inp[1]) ? node4646 : 4'b0011;
																assign node4646 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node4649 = (inp[5]) ? node4653 : node4650;
																assign node4650 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node4653 = (inp[1]) ? 4'b0011 : 4'b0111;
											assign node4656 = (inp[5]) ? node4696 : node4657;
												assign node4657 = (inp[9]) ? node4677 : node4658;
													assign node4658 = (inp[2]) ? node4668 : node4659;
														assign node4659 = (inp[13]) ? node4665 : node4660;
															assign node4660 = (inp[1]) ? 4'b0110 : node4661;
																assign node4661 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node4665 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node4668 = (inp[13]) ? node4674 : node4669;
															assign node4669 = (inp[1]) ? node4671 : 4'b0010;
																assign node4671 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node4674 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node4677 = (inp[13]) ? node4687 : node4678;
														assign node4678 = (inp[2]) ? node4684 : node4679;
															assign node4679 = (inp[0]) ? node4681 : 4'b0111;
																assign node4681 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node4684 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node4687 = (inp[2]) ? node4691 : node4688;
															assign node4688 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node4691 = (inp[1]) ? node4693 : 4'b0110;
																assign node4693 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node4696 = (inp[13]) ? node4714 : node4697;
													assign node4697 = (inp[9]) ? node4707 : node4698;
														assign node4698 = (inp[0]) ? node4702 : node4699;
															assign node4699 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node4702 = (inp[2]) ? 4'b0010 : node4703;
																assign node4703 = (inp[1]) ? 4'b0010 : 4'b0110;
														assign node4707 = (inp[2]) ? node4709 : 4'b0011;
															assign node4709 = (inp[1]) ? 4'b0110 : node4710;
																assign node4710 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node4714 = (inp[9]) ? node4728 : node4715;
														assign node4715 = (inp[0]) ? node4721 : node4716;
															assign node4716 = (inp[2]) ? 4'b0010 : node4717;
																assign node4717 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node4721 = (inp[1]) ? node4725 : node4722;
																assign node4722 = (inp[2]) ? 4'b0111 : 4'b0010;
																assign node4725 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node4728 = (inp[1]) ? node4734 : node4729;
															assign node4729 = (inp[2]) ? 4'b0111 : node4730;
																assign node4730 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node4734 = (inp[2]) ? node4736 : 4'b0110;
																assign node4736 = (inp[0]) ? 4'b0010 : 4'b0011;
					assign node4739 = (inp[10]) ? node7171 : node4740;
						assign node4740 = (inp[9]) ? node5912 : node4741;
							assign node4741 = (inp[11]) ? node5289 : node4742;
								assign node4742 = (inp[1]) ? node5046 : node4743;
									assign node4743 = (inp[12]) ? node4889 : node4744;
										assign node4744 = (inp[7]) ? node4806 : node4745;
											assign node4745 = (inp[15]) ? node4765 : node4746;
												assign node4746 = (inp[2]) ? node4756 : node4747;
													assign node4747 = (inp[5]) ? node4751 : node4748;
														assign node4748 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node4751 = (inp[0]) ? node4753 : 4'b1100;
															assign node4753 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node4756 = (inp[13]) ? node4762 : node4757;
														assign node4757 = (inp[4]) ? 4'b1101 : node4758;
															assign node4758 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node4762 = (inp[5]) ? 4'b1101 : 4'b1001;
												assign node4765 = (inp[4]) ? node4787 : node4766;
													assign node4766 = (inp[0]) ? node4782 : node4767;
														assign node4767 = (inp[13]) ? node4775 : node4768;
															assign node4768 = (inp[2]) ? node4772 : node4769;
																assign node4769 = (inp[5]) ? 4'b1110 : 4'b1010;
																assign node4772 = (inp[5]) ? 4'b1011 : 4'b1110;
															assign node4775 = (inp[2]) ? node4779 : node4776;
																assign node4776 = (inp[5]) ? 4'b1011 : 4'b1111;
																assign node4779 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node4782 = (inp[2]) ? node4784 : 4'b1010;
															assign node4784 = (inp[13]) ? 4'b1010 : 4'b1111;
													assign node4787 = (inp[13]) ? node4797 : node4788;
														assign node4788 = (inp[0]) ? node4794 : node4789;
															assign node4789 = (inp[2]) ? node4791 : 4'b1100;
																assign node4791 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node4794 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node4797 = (inp[5]) ? node4803 : node4798;
															assign node4798 = (inp[2]) ? 4'b1101 : node4799;
																assign node4799 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node4803 = (inp[2]) ? 4'b1000 : 4'b1100;
											assign node4806 = (inp[4]) ? node4844 : node4807;
												assign node4807 = (inp[15]) ? node4825 : node4808;
													assign node4808 = (inp[0]) ? node4818 : node4809;
														assign node4809 = (inp[13]) ? node4811 : 4'b1110;
															assign node4811 = (inp[5]) ? node4815 : node4812;
																assign node4812 = (inp[2]) ? 4'b1011 : 4'b1110;
																assign node4815 = (inp[2]) ? 4'b1110 : 4'b1011;
														assign node4818 = (inp[13]) ? node4820 : 4'b1010;
															assign node4820 = (inp[5]) ? node4822 : 4'b1110;
																assign node4822 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node4825 = (inp[0]) ? node4835 : node4826;
														assign node4826 = (inp[13]) ? 4'b1001 : node4827;
															assign node4827 = (inp[2]) ? node4831 : node4828;
																assign node4828 = (inp[5]) ? 4'b1101 : 4'b1100;
																assign node4831 = (inp[5]) ? 4'b1000 : 4'b1001;
														assign node4835 = (inp[13]) ? node4839 : node4836;
															assign node4836 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node4839 = (inp[2]) ? 4'b1100 : node4840;
																assign node4840 = (inp[5]) ? 4'b1001 : 4'b1000;
												assign node4844 = (inp[0]) ? node4868 : node4845;
													assign node4845 = (inp[2]) ? node4857 : node4846;
														assign node4846 = (inp[15]) ? node4852 : node4847;
															assign node4847 = (inp[13]) ? node4849 : 4'b1010;
																assign node4849 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node4852 = (inp[13]) ? node4854 : 4'b1110;
																assign node4854 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node4857 = (inp[15]) ? node4861 : node4858;
															assign node4858 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node4861 = (inp[13]) ? node4865 : node4862;
																assign node4862 = (inp[5]) ? 4'b1010 : 4'b1110;
																assign node4865 = (inp[5]) ? 4'b1111 : 4'b1011;
													assign node4868 = (inp[15]) ? node4876 : node4869;
														assign node4869 = (inp[5]) ? 4'b1110 : node4870;
															assign node4870 = (inp[2]) ? node4872 : 4'b1010;
																assign node4872 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node4876 = (inp[2]) ? node4884 : node4877;
															assign node4877 = (inp[5]) ? node4881 : node4878;
																assign node4878 = (inp[13]) ? 4'b1110 : 4'b1011;
																assign node4881 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node4884 = (inp[13]) ? node4886 : 4'b1010;
																assign node4886 = (inp[5]) ? 4'b1111 : 4'b1010;
										assign node4889 = (inp[7]) ? node4971 : node4890;
											assign node4890 = (inp[15]) ? node4930 : node4891;
												assign node4891 = (inp[5]) ? node4909 : node4892;
													assign node4892 = (inp[4]) ? node4902 : node4893;
														assign node4893 = (inp[2]) ? node4897 : node4894;
															assign node4894 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node4897 = (inp[13]) ? 4'b1011 : node4898;
																assign node4898 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node4902 = (inp[2]) ? node4906 : node4903;
															assign node4903 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node4906 = (inp[13]) ? 4'b1110 : 4'b1010;
													assign node4909 = (inp[4]) ? node4923 : node4910;
														assign node4910 = (inp[0]) ? node4916 : node4911;
															assign node4911 = (inp[2]) ? 4'b1011 : node4912;
																assign node4912 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node4916 = (inp[13]) ? node4920 : node4917;
																assign node4917 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node4920 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node4923 = (inp[13]) ? node4927 : node4924;
															assign node4924 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node4927 = (inp[2]) ? 4'b1111 : 4'b1011;
												assign node4930 = (inp[4]) ? node4956 : node4931;
													assign node4931 = (inp[5]) ? node4941 : node4932;
														assign node4932 = (inp[13]) ? node4936 : node4933;
															assign node4933 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node4936 = (inp[2]) ? 4'b1100 : node4937;
																assign node4937 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node4941 = (inp[0]) ? node4949 : node4942;
															assign node4942 = (inp[13]) ? node4946 : node4943;
																assign node4943 = (inp[2]) ? 4'b1101 : 4'b1000;
																assign node4946 = (inp[2]) ? 4'b1000 : 4'b1101;
															assign node4949 = (inp[13]) ? node4953 : node4950;
																assign node4950 = (inp[2]) ? 4'b1101 : 4'b1001;
																assign node4953 = (inp[2]) ? 4'b1001 : 4'b1100;
													assign node4956 = (inp[13]) ? node4962 : node4957;
														assign node4957 = (inp[2]) ? node4959 : 4'b1010;
															assign node4959 = (inp[5]) ? 4'b1111 : 4'b1110;
														assign node4962 = (inp[2]) ? node4964 : 4'b1111;
															assign node4964 = (inp[5]) ? node4968 : node4965;
																assign node4965 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node4968 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node4971 = (inp[4]) ? node5009 : node4972;
												assign node4972 = (inp[15]) ? node4990 : node4973;
													assign node4973 = (inp[13]) ? node4981 : node4974;
														assign node4974 = (inp[0]) ? 4'b1101 : node4975;
															assign node4975 = (inp[5]) ? node4977 : 4'b1100;
																assign node4977 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node4981 = (inp[2]) ? node4985 : node4982;
															assign node4982 = (inp[5]) ? 4'b1100 : 4'b1001;
															assign node4985 = (inp[5]) ? 4'b1001 : node4986;
																assign node4986 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node4990 = (inp[5]) ? node5000 : node4991;
														assign node4991 = (inp[2]) ? node4995 : node4992;
															assign node4992 = (inp[13]) ? 4'b1110 : 4'b1011;
															assign node4995 = (inp[13]) ? 4'b1011 : node4996;
																assign node4996 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node5000 = (inp[0]) ? node5002 : 4'b1110;
															assign node5002 = (inp[13]) ? node5006 : node5003;
																assign node5003 = (inp[2]) ? 4'b1011 : 4'b1110;
																assign node5006 = (inp[2]) ? 4'b1110 : 4'b1010;
												assign node5009 = (inp[0]) ? node5033 : node5010;
													assign node5010 = (inp[13]) ? node5022 : node5011;
														assign node5011 = (inp[15]) ? node5015 : node5012;
															assign node5012 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node5015 = (inp[5]) ? node5019 : node5016;
																assign node5016 = (inp[2]) ? 4'b1101 : 4'b1001;
																assign node5019 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node5022 = (inp[15]) ? node5030 : node5023;
															assign node5023 = (inp[5]) ? node5027 : node5024;
																assign node5024 = (inp[2]) ? 4'b1001 : 4'b1101;
																assign node5027 = (inp[2]) ? 4'b1100 : 4'b1001;
															assign node5030 = (inp[2]) ? 4'b1000 : 4'b1100;
													assign node5033 = (inp[15]) ? 4'b1001 : node5034;
														assign node5034 = (inp[2]) ? node5040 : node5035;
															assign node5035 = (inp[13]) ? 4'b1101 : node5036;
																assign node5036 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node5040 = (inp[13]) ? 4'b1001 : node5041;
																assign node5041 = (inp[5]) ? 4'b1001 : 4'b1101;
									assign node5046 = (inp[13]) ? node5182 : node5047;
										assign node5047 = (inp[2]) ? node5111 : node5048;
											assign node5048 = (inp[15]) ? node5082 : node5049;
												assign node5049 = (inp[12]) ? node5063 : node5050;
													assign node5050 = (inp[7]) ? node5058 : node5051;
														assign node5051 = (inp[5]) ? node5053 : 4'b1000;
															assign node5053 = (inp[0]) ? 4'b1001 : node5054;
																assign node5054 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node5058 = (inp[0]) ? 4'b1010 : node5059;
															assign node5059 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node5063 = (inp[7]) ? node5077 : node5064;
														assign node5064 = (inp[0]) ? node5070 : node5065;
															assign node5065 = (inp[4]) ? 4'b1011 : node5066;
																assign node5066 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node5070 = (inp[4]) ? node5074 : node5071;
																assign node5071 = (inp[5]) ? 4'b1010 : 4'b1111;
																assign node5074 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node5077 = (inp[4]) ? 4'b1000 : node5078;
															assign node5078 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node5082 = (inp[4]) ? node5098 : node5083;
													assign node5083 = (inp[5]) ? node5093 : node5084;
														assign node5084 = (inp[12]) ? node5090 : node5085;
															assign node5085 = (inp[7]) ? 4'b1001 : node5086;
																assign node5086 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node5090 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node5093 = (inp[12]) ? node5095 : 4'b1100;
															assign node5095 = (inp[7]) ? 4'b1010 : 4'b1100;
													assign node5098 = (inp[7]) ? node5108 : node5099;
														assign node5099 = (inp[12]) ? node5105 : node5100;
															assign node5100 = (inp[0]) ? 4'b1101 : node5101;
																assign node5101 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node5105 = (inp[5]) ? 4'b1011 : 4'b1110;
														assign node5108 = (inp[12]) ? 4'b1001 : 4'b1011;
											assign node5111 = (inp[7]) ? node5149 : node5112;
												assign node5112 = (inp[12]) ? node5134 : node5113;
													assign node5113 = (inp[4]) ? node5125 : node5114;
														assign node5114 = (inp[15]) ? node5120 : node5115;
															assign node5115 = (inp[0]) ? 4'b1101 : node5116;
																assign node5116 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node5120 = (inp[5]) ? node5122 : 4'b1111;
																assign node5122 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node5125 = (inp[15]) ? node5127 : 4'b1100;
															assign node5127 = (inp[0]) ? node5131 : node5128;
																assign node5128 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node5131 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node5134 = (inp[15]) ? node5142 : node5135;
														assign node5135 = (inp[5]) ? node5139 : node5136;
															assign node5136 = (inp[4]) ? 4'b1111 : 4'b1010;
															assign node5139 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node5142 = (inp[4]) ? node5146 : node5143;
															assign node5143 = (inp[5]) ? 4'b1001 : 4'b1000;
															assign node5146 = (inp[0]) ? 4'b1010 : 4'b1110;
												assign node5149 = (inp[12]) ? node5171 : node5150;
													assign node5150 = (inp[4]) ? node5158 : node5151;
														assign node5151 = (inp[15]) ? node5153 : 4'b1110;
															assign node5153 = (inp[5]) ? 4'b1001 : node5154;
																assign node5154 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node5158 = (inp[5]) ? node5166 : node5159;
															assign node5159 = (inp[0]) ? node5163 : node5160;
																assign node5160 = (inp[15]) ? 4'b1110 : 4'b1111;
																assign node5163 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node5166 = (inp[0]) ? node5168 : 4'b1110;
																assign node5168 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node5171 = (inp[15]) ? node5177 : node5172;
														assign node5172 = (inp[4]) ? node5174 : 4'b1000;
															assign node5174 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node5177 = (inp[4]) ? node5179 : 4'b1111;
															assign node5179 = (inp[5]) ? 4'b1101 : 4'b1100;
										assign node5182 = (inp[2]) ? node5230 : node5183;
											assign node5183 = (inp[7]) ? node5215 : node5184;
												assign node5184 = (inp[12]) ? node5198 : node5185;
													assign node5185 = (inp[4]) ? node5191 : node5186;
														assign node5186 = (inp[15]) ? node5188 : 4'b1100;
															assign node5188 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node5191 = (inp[15]) ? node5195 : node5192;
															assign node5192 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node5195 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node5198 = (inp[4]) ? node5204 : node5199;
														assign node5199 = (inp[15]) ? 4'b1001 : node5200;
															assign node5200 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node5204 = (inp[5]) ? node5210 : node5205;
															assign node5205 = (inp[0]) ? 4'b1010 : node5206;
																assign node5206 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node5210 = (inp[15]) ? 4'b1110 : node5211;
																assign node5211 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node5215 = (inp[4]) ? node5227 : node5216;
													assign node5216 = (inp[15]) ? node5220 : node5217;
														assign node5217 = (inp[12]) ? 4'b1000 : 4'b1110;
														assign node5220 = (inp[12]) ? 4'b1111 : node5221;
															assign node5221 = (inp[5]) ? node5223 : 4'b1100;
																assign node5223 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node5227 = (inp[12]) ? 4'b1100 : 4'b1110;
											assign node5230 = (inp[4]) ? node5272 : node5231;
												assign node5231 = (inp[12]) ? node5251 : node5232;
													assign node5232 = (inp[5]) ? node5246 : node5233;
														assign node5233 = (inp[0]) ? node5239 : node5234;
															assign node5234 = (inp[15]) ? node5236 : 4'b1001;
																assign node5236 = (inp[7]) ? 4'b1001 : 4'b1010;
															assign node5239 = (inp[7]) ? node5243 : node5240;
																assign node5240 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node5243 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node5246 = (inp[15]) ? 4'b1100 : node5247;
															assign node5247 = (inp[7]) ? 4'b1011 : 4'b1000;
													assign node5251 = (inp[0]) ? node5263 : node5252;
														assign node5252 = (inp[15]) ? node5258 : node5253;
															assign node5253 = (inp[7]) ? 4'b1100 : node5254;
																assign node5254 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node5258 = (inp[7]) ? 4'b1010 : node5259;
																assign node5259 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node5263 = (inp[7]) ? node5267 : node5264;
															assign node5264 = (inp[15]) ? 4'b1100 : 4'b1011;
															assign node5267 = (inp[15]) ? 4'b1011 : node5268;
																assign node5268 = (inp[5]) ? 4'b1100 : 4'b1101;
												assign node5272 = (inp[7]) ? node5286 : node5273;
													assign node5273 = (inp[12]) ? node5279 : node5274;
														assign node5274 = (inp[15]) ? 4'b1100 : node5275;
															assign node5275 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node5279 = (inp[5]) ? node5283 : node5280;
															assign node5280 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node5283 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node5286 = (inp[12]) ? 4'b1000 : 4'b1010;
								assign node5289 = (inp[0]) ? node5603 : node5290;
									assign node5290 = (inp[13]) ? node5444 : node5291;
										assign node5291 = (inp[2]) ? node5373 : node5292;
											assign node5292 = (inp[1]) ? node5334 : node5293;
												assign node5293 = (inp[5]) ? node5311 : node5294;
													assign node5294 = (inp[7]) ? node5306 : node5295;
														assign node5295 = (inp[15]) ? node5299 : node5296;
															assign node5296 = (inp[4]) ? 4'b1001 : 4'b1011;
															assign node5299 = (inp[4]) ? node5303 : node5300;
																assign node5300 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node5303 = (inp[12]) ? 4'b1010 : 4'b1101;
														assign node5306 = (inp[12]) ? 4'b1100 : node5307;
															assign node5307 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node5311 = (inp[7]) ? node5325 : node5312;
														assign node5312 = (inp[12]) ? node5318 : node5313;
															assign node5313 = (inp[15]) ? 4'b1000 : node5314;
																assign node5314 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node5318 = (inp[15]) ? node5322 : node5319;
																assign node5319 = (inp[4]) ? 4'b1110 : 4'b1010;
																assign node5322 = (inp[4]) ? 4'b1011 : 4'b1000;
														assign node5325 = (inp[12]) ? node5329 : node5326;
															assign node5326 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node5329 = (inp[4]) ? 4'b1100 : node5330;
																assign node5330 = (inp[15]) ? 4'b1111 : 4'b1001;
												assign node5334 = (inp[7]) ? node5358 : node5335;
													assign node5335 = (inp[12]) ? node5345 : node5336;
														assign node5336 = (inp[5]) ? node5338 : 4'b1001;
															assign node5338 = (inp[4]) ? node5342 : node5339;
																assign node5339 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node5342 = (inp[15]) ? 4'b1101 : 4'b1000;
														assign node5345 = (inp[4]) ? node5351 : node5346;
															assign node5346 = (inp[15]) ? 4'b1101 : node5347;
																assign node5347 = (inp[5]) ? 4'b1011 : 4'b1110;
															assign node5351 = (inp[5]) ? node5355 : node5352;
																assign node5352 = (inp[15]) ? 4'b1111 : 4'b1011;
																assign node5355 = (inp[15]) ? 4'b1010 : 4'b1111;
													assign node5358 = (inp[15]) ? node5364 : node5359;
														assign node5359 = (inp[12]) ? node5361 : 4'b1011;
															assign node5361 = (inp[4]) ? 4'b1001 : 4'b1100;
														assign node5364 = (inp[4]) ? node5370 : node5365;
															assign node5365 = (inp[5]) ? 4'b1011 : node5366;
																assign node5366 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node5370 = (inp[12]) ? 4'b1000 : 4'b1010;
											assign node5373 = (inp[4]) ? node5413 : node5374;
												assign node5374 = (inp[7]) ? node5392 : node5375;
													assign node5375 = (inp[15]) ? node5385 : node5376;
														assign node5376 = (inp[12]) ? node5382 : node5377;
															assign node5377 = (inp[1]) ? 4'b1100 : node5378;
																assign node5378 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node5382 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node5385 = (inp[12]) ? node5389 : node5386;
															assign node5386 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node5389 = (inp[5]) ? 4'b1100 : 4'b1000;
													assign node5392 = (inp[15]) ? node5404 : node5393;
														assign node5393 = (inp[12]) ? node5399 : node5394;
															assign node5394 = (inp[5]) ? node5396 : 4'b1110;
																assign node5396 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node5399 = (inp[1]) ? node5401 : 4'b1100;
																assign node5401 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node5404 = (inp[12]) ? node5410 : node5405;
															assign node5405 = (inp[1]) ? node5407 : 4'b1000;
																assign node5407 = (inp[5]) ? 4'b1000 : 4'b1101;
															assign node5410 = (inp[5]) ? 4'b1110 : 4'b1111;
												assign node5413 = (inp[5]) ? node5429 : node5414;
													assign node5414 = (inp[7]) ? node5422 : node5415;
														assign node5415 = (inp[15]) ? node5417 : 4'b1101;
															assign node5417 = (inp[12]) ? 4'b1011 : node5418;
																assign node5418 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node5422 = (inp[12]) ? 4'b1101 : node5423;
															assign node5423 = (inp[1]) ? node5425 : 4'b1111;
																assign node5425 = (inp[15]) ? 4'b1110 : 4'b1111;
													assign node5429 = (inp[1]) ? node5435 : node5430;
														assign node5430 = (inp[12]) ? node5432 : 4'b1011;
															assign node5432 = (inp[7]) ? 4'b1000 : 4'b1010;
														assign node5435 = (inp[15]) ? node5439 : node5436;
															assign node5436 = (inp[12]) ? 4'b1101 : 4'b1100;
															assign node5439 = (inp[7]) ? 4'b1110 : node5440;
																assign node5440 = (inp[12]) ? 4'b1110 : 4'b1001;
										assign node5444 = (inp[2]) ? node5520 : node5445;
											assign node5445 = (inp[1]) ? node5487 : node5446;
												assign node5446 = (inp[5]) ? node5466 : node5447;
													assign node5447 = (inp[12]) ? node5459 : node5448;
														assign node5448 = (inp[15]) ? node5452 : node5449;
															assign node5449 = (inp[7]) ? 4'b1111 : 4'b1101;
															assign node5452 = (inp[4]) ? node5456 : node5453;
																assign node5453 = (inp[7]) ? 4'b1001 : 4'b1110;
																assign node5456 = (inp[7]) ? 4'b1111 : 4'b1001;
														assign node5459 = (inp[7]) ? node5463 : node5460;
															assign node5460 = (inp[4]) ? 4'b1010 : 4'b1111;
															assign node5463 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node5466 = (inp[12]) ? node5476 : node5467;
														assign node5467 = (inp[7]) ? node5473 : node5468;
															assign node5468 = (inp[15]) ? node5470 : 4'b1000;
																assign node5470 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node5473 = (inp[4]) ? 4'b1011 : 4'b1000;
														assign node5476 = (inp[4]) ? node5482 : node5477;
															assign node5477 = (inp[7]) ? node5479 : 4'b1101;
																assign node5479 = (inp[15]) ? 4'b1011 : 4'b1101;
															assign node5482 = (inp[15]) ? node5484 : 4'b1011;
																assign node5484 = (inp[7]) ? 4'b1000 : 4'b1110;
												assign node5487 = (inp[15]) ? node5499 : node5488;
													assign node5488 = (inp[7]) ? node5494 : node5489;
														assign node5489 = (inp[12]) ? 4'b1111 : node5490;
															assign node5490 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node5494 = (inp[12]) ? node5496 : 4'b1111;
															assign node5496 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node5499 = (inp[7]) ? node5511 : node5500;
														assign node5500 = (inp[12]) ? node5506 : node5501;
															assign node5501 = (inp[4]) ? node5503 : 4'b1111;
																assign node5503 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node5506 = (inp[4]) ? 4'b1011 : node5507;
																assign node5507 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node5511 = (inp[4]) ? node5517 : node5512;
															assign node5512 = (inp[12]) ? 4'b1110 : node5513;
																assign node5513 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node5517 = (inp[12]) ? 4'b1101 : 4'b1111;
											assign node5520 = (inp[1]) ? node5564 : node5521;
												assign node5521 = (inp[5]) ? node5541 : node5522;
													assign node5522 = (inp[7]) ? node5534 : node5523;
														assign node5523 = (inp[12]) ? node5529 : node5524;
															assign node5524 = (inp[4]) ? node5526 : 4'b1011;
																assign node5526 = (inp[15]) ? 4'b1100 : 4'b1001;
															assign node5529 = (inp[4]) ? node5531 : 4'b1101;
																assign node5531 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node5534 = (inp[12]) ? node5538 : node5535;
															assign node5535 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node5538 = (inp[4]) ? 4'b1000 : 4'b1010;
													assign node5541 = (inp[7]) ? node5551 : node5542;
														assign node5542 = (inp[15]) ? node5546 : node5543;
															assign node5543 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node5546 = (inp[4]) ? node5548 : 4'b1111;
																assign node5548 = (inp[12]) ? 4'b1010 : 4'b1001;
														assign node5551 = (inp[4]) ? node5557 : node5552;
															assign node5552 = (inp[15]) ? node5554 : 4'b1111;
																assign node5554 = (inp[12]) ? 4'b1111 : 4'b1101;
															assign node5557 = (inp[12]) ? node5561 : node5558;
																assign node5558 = (inp[15]) ? 4'b1110 : 4'b1111;
																assign node5561 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node5564 = (inp[4]) ? node5590 : node5565;
													assign node5565 = (inp[5]) ? node5577 : node5566;
														assign node5566 = (inp[12]) ? node5572 : node5567;
															assign node5567 = (inp[15]) ? node5569 : 4'b1000;
																assign node5569 = (inp[7]) ? 4'b1000 : 4'b1010;
															assign node5572 = (inp[7]) ? node5574 : 4'b1101;
																assign node5574 = (inp[15]) ? 4'b1010 : 4'b1100;
														assign node5577 = (inp[7]) ? node5585 : node5578;
															assign node5578 = (inp[15]) ? node5582 : node5579;
																assign node5579 = (inp[12]) ? 4'b1010 : 4'b1001;
																assign node5582 = (inp[12]) ? 4'b1101 : 4'b1010;
															assign node5585 = (inp[15]) ? node5587 : 4'b1101;
																assign node5587 = (inp[12]) ? 4'b1011 : 4'b1101;
													assign node5590 = (inp[7]) ? node5600 : node5591;
														assign node5591 = (inp[12]) ? node5595 : node5592;
															assign node5592 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node5595 = (inp[15]) ? node5597 : 4'b1011;
																assign node5597 = (inp[5]) ? 4'b1011 : 4'b1110;
														assign node5600 = (inp[12]) ? 4'b1001 : 4'b1011;
									assign node5603 = (inp[4]) ? node5751 : node5604;
										assign node5604 = (inp[13]) ? node5674 : node5605;
											assign node5605 = (inp[1]) ? node5639 : node5606;
												assign node5606 = (inp[2]) ? node5624 : node5607;
													assign node5607 = (inp[12]) ? node5617 : node5608;
														assign node5608 = (inp[7]) ? node5614 : node5609;
															assign node5609 = (inp[5]) ? node5611 : 4'b1010;
																assign node5611 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node5614 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node5617 = (inp[5]) ? node5619 : 4'b1011;
															assign node5619 = (inp[7]) ? 4'b1000 : node5620;
																assign node5620 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node5624 = (inp[12]) ? node5632 : node5625;
														assign node5625 = (inp[5]) ? node5627 : 4'b1100;
															assign node5627 = (inp[7]) ? node5629 : 4'b1001;
																assign node5629 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node5632 = (inp[5]) ? node5636 : node5633;
															assign node5633 = (inp[15]) ? 4'b1111 : 4'b1001;
															assign node5636 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node5639 = (inp[2]) ? node5659 : node5640;
													assign node5640 = (inp[12]) ? node5650 : node5641;
														assign node5641 = (inp[5]) ? node5645 : node5642;
															assign node5642 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node5645 = (inp[15]) ? node5647 : 4'b1011;
																assign node5647 = (inp[7]) ? 4'b1100 : 4'b1011;
														assign node5650 = (inp[15]) ? node5656 : node5651;
															assign node5651 = (inp[7]) ? 4'b1101 : node5652;
																assign node5652 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node5656 = (inp[7]) ? 4'b1010 : 4'b1101;
													assign node5659 = (inp[12]) ? node5667 : node5660;
														assign node5660 = (inp[15]) ? node5664 : node5661;
															assign node5661 = (inp[7]) ? 4'b1110 : 4'b1101;
															assign node5664 = (inp[7]) ? 4'b1001 : 4'b1111;
														assign node5667 = (inp[15]) ? 4'b1110 : node5668;
															assign node5668 = (inp[7]) ? 4'b1000 : node5669;
																assign node5669 = (inp[5]) ? 4'b1110 : 4'b1010;
											assign node5674 = (inp[2]) ? node5708 : node5675;
												assign node5675 = (inp[15]) ? node5687 : node5676;
													assign node5676 = (inp[7]) ? node5680 : node5677;
														assign node5677 = (inp[12]) ? 4'b1110 : 4'b1100;
														assign node5680 = (inp[12]) ? node5684 : node5681;
															assign node5681 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node5684 = (inp[1]) ? 4'b1001 : 4'b1100;
													assign node5687 = (inp[7]) ? node5699 : node5688;
														assign node5688 = (inp[12]) ? node5694 : node5689;
															assign node5689 = (inp[5]) ? node5691 : 4'b1111;
																assign node5691 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node5694 = (inp[5]) ? node5696 : 4'b1001;
																assign node5696 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node5699 = (inp[12]) ? node5705 : node5700;
															assign node5700 = (inp[5]) ? 4'b1001 : node5701;
																assign node5701 = (inp[1]) ? 4'b1100 : 4'b1001;
															assign node5705 = (inp[1]) ? 4'b1111 : 4'b1110;
												assign node5708 = (inp[1]) ? node5732 : node5709;
													assign node5709 = (inp[15]) ? node5723 : node5710;
														assign node5710 = (inp[5]) ? node5718 : node5711;
															assign node5711 = (inp[7]) ? node5715 : node5712;
																assign node5712 = (inp[12]) ? 4'b1011 : 4'b1001;
																assign node5715 = (inp[12]) ? 4'b1101 : 4'b1011;
															assign node5718 = (inp[12]) ? node5720 : 4'b1101;
																assign node5720 = (inp[7]) ? 4'b1001 : 4'b1011;
														assign node5723 = (inp[7]) ? node5729 : node5724;
															assign node5724 = (inp[12]) ? 4'b1000 : node5725;
																assign node5725 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node5729 = (inp[5]) ? 4'b1101 : 4'b1011;
													assign node5732 = (inp[12]) ? node5740 : node5733;
														assign node5733 = (inp[7]) ? node5737 : node5734;
															assign node5734 = (inp[5]) ? 4'b1011 : 4'b1010;
															assign node5737 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node5740 = (inp[15]) ? node5746 : node5741;
															assign node5741 = (inp[7]) ? 4'b1100 : node5742;
																assign node5742 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node5746 = (inp[7]) ? 4'b1010 : node5747;
																assign node5747 = (inp[5]) ? 4'b1100 : 4'b1101;
										assign node5751 = (inp[13]) ? node5837 : node5752;
											assign node5752 = (inp[12]) ? node5796 : node5753;
												assign node5753 = (inp[7]) ? node5779 : node5754;
													assign node5754 = (inp[1]) ? node5766 : node5755;
														assign node5755 = (inp[15]) ? node5761 : node5756;
															assign node5756 = (inp[5]) ? node5758 : 4'b1000;
																assign node5758 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node5761 = (inp[5]) ? 4'b1100 : node5762;
																assign node5762 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node5766 = (inp[5]) ? node5774 : node5767;
															assign node5767 = (inp[2]) ? node5771 : node5768;
																assign node5768 = (inp[15]) ? 4'b1100 : 4'b1000;
																assign node5771 = (inp[15]) ? 4'b1000 : 4'b1101;
															assign node5774 = (inp[15]) ? 4'b1001 : node5775;
																assign node5775 = (inp[2]) ? 4'b1100 : 4'b1001;
													assign node5779 = (inp[15]) ? node5787 : node5780;
														assign node5780 = (inp[2]) ? node5784 : node5781;
															assign node5781 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node5784 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node5787 = (inp[1]) ? node5793 : node5788;
															assign node5788 = (inp[2]) ? 4'b1010 : node5789;
																assign node5789 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node5793 = (inp[2]) ? 4'b1110 : 4'b1011;
												assign node5796 = (inp[7]) ? node5816 : node5797;
													assign node5797 = (inp[1]) ? node5809 : node5798;
														assign node5798 = (inp[5]) ? node5802 : node5799;
															assign node5799 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node5802 = (inp[15]) ? node5806 : node5803;
																assign node5803 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node5806 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node5809 = (inp[5]) ? node5813 : node5810;
															assign node5810 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node5813 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node5816 = (inp[2]) ? node5828 : node5817;
														assign node5817 = (inp[15]) ? node5823 : node5818;
															assign node5818 = (inp[5]) ? 4'b1100 : node5819;
																assign node5819 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node5823 = (inp[1]) ? 4'b1001 : node5824;
																assign node5824 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node5828 = (inp[1]) ? node5834 : node5829;
															assign node5829 = (inp[15]) ? node5831 : 4'b1000;
																assign node5831 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node5834 = (inp[15]) ? 4'b1100 : 4'b1101;
											assign node5837 = (inp[2]) ? node5881 : node5838;
												assign node5838 = (inp[5]) ? node5858 : node5839;
													assign node5839 = (inp[12]) ? node5849 : node5840;
														assign node5840 = (inp[7]) ? node5844 : node5841;
															assign node5841 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node5844 = (inp[15]) ? node5846 : 4'b1110;
																assign node5846 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node5849 = (inp[7]) ? node5855 : node5850;
															assign node5850 = (inp[1]) ? node5852 : 4'b1111;
																assign node5852 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node5855 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node5858 = (inp[12]) ? node5872 : node5859;
														assign node5859 = (inp[7]) ? node5867 : node5860;
															assign node5860 = (inp[15]) ? node5864 : node5861;
																assign node5861 = (inp[1]) ? 4'b1101 : 4'b1001;
																assign node5864 = (inp[1]) ? 4'b1001 : 4'b1100;
															assign node5867 = (inp[1]) ? 4'b1110 : node5868;
																assign node5868 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node5872 = (inp[7]) ? node5878 : node5873;
															assign node5873 = (inp[15]) ? 4'b1110 : node5874;
																assign node5874 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node5878 = (inp[15]) ? 4'b1000 : 4'b1100;
												assign node5881 = (inp[1]) ? node5897 : node5882;
													assign node5882 = (inp[5]) ? node5888 : node5883;
														assign node5883 = (inp[15]) ? 4'b1011 : node5884;
															assign node5884 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node5888 = (inp[7]) ? node5894 : node5889;
															assign node5889 = (inp[12]) ? 4'b1010 : node5890;
																assign node5890 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node5894 = (inp[12]) ? 4'b1100 : 4'b1111;
													assign node5897 = (inp[7]) ? node5909 : node5898;
														assign node5898 = (inp[12]) ? node5902 : node5899;
															assign node5899 = (inp[5]) ? 4'b1001 : 4'b1000;
															assign node5902 = (inp[5]) ? node5906 : node5903;
																assign node5903 = (inp[15]) ? 4'b1111 : 4'b1011;
																assign node5906 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node5909 = (inp[12]) ? 4'b1000 : 4'b1010;
							assign node5912 = (inp[11]) ? node6536 : node5913;
								assign node5913 = (inp[5]) ? node6181 : node5914;
									assign node5914 = (inp[2]) ? node6030 : node5915;
										assign node5915 = (inp[13]) ? node5969 : node5916;
											assign node5916 = (inp[7]) ? node5938 : node5917;
												assign node5917 = (inp[12]) ? node5923 : node5918;
													assign node5918 = (inp[15]) ? node5920 : 4'b1001;
														assign node5920 = (inp[4]) ? 4'b1101 : 4'b1011;
													assign node5923 = (inp[15]) ? node5933 : node5924;
														assign node5924 = (inp[1]) ? node5928 : node5925;
															assign node5925 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node5928 = (inp[4]) ? node5930 : 4'b1110;
																assign node5930 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node5933 = (inp[4]) ? node5935 : 4'b1101;
															assign node5935 = (inp[0]) ? 4'b1111 : 4'b1011;
												assign node5938 = (inp[12]) ? node5950 : node5939;
													assign node5939 = (inp[15]) ? node5941 : 4'b1011;
														assign node5941 = (inp[4]) ? node5945 : node5942;
															assign node5942 = (inp[1]) ? 4'b1000 : 4'b1101;
															assign node5945 = (inp[1]) ? 4'b1010 : node5946;
																assign node5946 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node5950 = (inp[15]) ? node5960 : node5951;
														assign node5951 = (inp[4]) ? node5957 : node5952;
															assign node5952 = (inp[1]) ? node5954 : 4'b1101;
																assign node5954 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node5957 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node5960 = (inp[4]) ? node5966 : node5961;
															assign node5961 = (inp[1]) ? node5963 : 4'b1010;
																assign node5963 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node5966 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node5969 = (inp[12]) ? node5989 : node5970;
												assign node5970 = (inp[15]) ? node5974 : node5971;
													assign node5971 = (inp[7]) ? 4'b1111 : 4'b1101;
													assign node5974 = (inp[1]) ? node5980 : node5975;
														assign node5975 = (inp[0]) ? 4'b1001 : node5976;
															assign node5976 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node5980 = (inp[7]) ? node5986 : node5981;
															assign node5981 = (inp[4]) ? 4'b1001 : node5982;
																assign node5982 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node5986 = (inp[4]) ? 4'b1111 : 4'b1101;
												assign node5989 = (inp[7]) ? node6013 : node5990;
													assign node5990 = (inp[4]) ? node6000 : node5991;
														assign node5991 = (inp[15]) ? node5995 : node5992;
															assign node5992 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node5995 = (inp[1]) ? 4'b1000 : node5996;
																assign node5996 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node6000 = (inp[0]) ? node6006 : node6001;
															assign node6001 = (inp[15]) ? node6003 : 4'b1011;
																assign node6003 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node6006 = (inp[1]) ? node6010 : node6007;
																assign node6007 = (inp[15]) ? 4'b1111 : 4'b1010;
																assign node6010 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node6013 = (inp[4]) ? node6023 : node6014;
														assign node6014 = (inp[15]) ? node6018 : node6015;
															assign node6015 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node6018 = (inp[1]) ? node6020 : 4'b1111;
																assign node6020 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node6023 = (inp[1]) ? 4'b1101 : node6024;
															assign node6024 = (inp[0]) ? 4'b1100 : node6025;
																assign node6025 = (inp[15]) ? 4'b1101 : 4'b1100;
										assign node6030 = (inp[13]) ? node6112 : node6031;
											assign node6031 = (inp[7]) ? node6069 : node6032;
												assign node6032 = (inp[12]) ? node6050 : node6033;
													assign node6033 = (inp[4]) ? node6043 : node6034;
														assign node6034 = (inp[15]) ? node6038 : node6035;
															assign node6035 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node6038 = (inp[0]) ? 4'b1110 : node6039;
																assign node6039 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node6043 = (inp[15]) ? node6045 : 4'b1100;
															assign node6045 = (inp[1]) ? node6047 : 4'b1001;
																assign node6047 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node6050 = (inp[4]) ? node6062 : node6051;
														assign node6051 = (inp[15]) ? node6057 : node6052;
															assign node6052 = (inp[1]) ? 4'b1011 : node6053;
																assign node6053 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node6057 = (inp[0]) ? 4'b1000 : node6058;
																assign node6058 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node6062 = (inp[1]) ? node6066 : node6063;
															assign node6063 = (inp[15]) ? 4'b1111 : 4'b1011;
															assign node6066 = (inp[15]) ? 4'b1011 : 4'b1110;
												assign node6069 = (inp[12]) ? node6091 : node6070;
													assign node6070 = (inp[15]) ? node6082 : node6071;
														assign node6071 = (inp[1]) ? node6077 : node6072;
															assign node6072 = (inp[0]) ? 4'b1111 : node6073;
																assign node6073 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node6077 = (inp[0]) ? node6079 : 4'b1111;
																assign node6079 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node6082 = (inp[4]) ? node6088 : node6083;
															assign node6083 = (inp[1]) ? node6085 : 4'b1000;
																assign node6085 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node6088 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node6091 = (inp[15]) ? node6103 : node6092;
														assign node6092 = (inp[4]) ? node6100 : node6093;
															assign node6093 = (inp[0]) ? node6097 : node6094;
																assign node6094 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node6097 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node6100 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node6103 = (inp[4]) ? node6107 : node6104;
															assign node6104 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node6107 = (inp[0]) ? 4'b1100 : node6108;
																assign node6108 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node6112 = (inp[7]) ? node6154 : node6113;
												assign node6113 = (inp[12]) ? node6129 : node6114;
													assign node6114 = (inp[4]) ? node6122 : node6115;
														assign node6115 = (inp[15]) ? node6117 : 4'b1000;
															assign node6117 = (inp[0]) ? node6119 : 4'b1011;
																assign node6119 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node6122 = (inp[15]) ? node6124 : 4'b1001;
															assign node6124 = (inp[1]) ? node6126 : 4'b1100;
																assign node6126 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node6129 = (inp[4]) ? node6139 : node6130;
														assign node6130 = (inp[15]) ? node6134 : node6131;
															assign node6131 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node6134 = (inp[1]) ? node6136 : 4'b1101;
																assign node6136 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node6139 = (inp[0]) ? node6147 : node6140;
															assign node6140 = (inp[1]) ? node6144 : node6141;
																assign node6141 = (inp[15]) ? 4'b1010 : 4'b1111;
																assign node6144 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node6147 = (inp[1]) ? node6151 : node6148;
																assign node6148 = (inp[15]) ? 4'b1011 : 4'b1111;
																assign node6151 = (inp[15]) ? 4'b1110 : 4'b1011;
												assign node6154 = (inp[4]) ? node6172 : node6155;
													assign node6155 = (inp[12]) ? node6161 : node6156;
														assign node6156 = (inp[15]) ? node6158 : 4'b1010;
															assign node6158 = (inp[1]) ? 4'b1000 : 4'b1101;
														assign node6161 = (inp[15]) ? node6167 : node6162;
															assign node6162 = (inp[1]) ? node6164 : 4'b1101;
																assign node6164 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node6167 = (inp[1]) ? node6169 : 4'b1010;
																assign node6169 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node6172 = (inp[12]) ? node6174 : 4'b1011;
														assign node6174 = (inp[1]) ? 4'b1001 : node6175;
															assign node6175 = (inp[15]) ? node6177 : 4'b1000;
																assign node6177 = (inp[0]) ? 4'b1000 : 4'b1001;
									assign node6181 = (inp[7]) ? node6367 : node6182;
										assign node6182 = (inp[12]) ? node6280 : node6183;
											assign node6183 = (inp[15]) ? node6241 : node6184;
												assign node6184 = (inp[0]) ? node6212 : node6185;
													assign node6185 = (inp[2]) ? node6199 : node6186;
														assign node6186 = (inp[4]) ? node6192 : node6187;
															assign node6187 = (inp[1]) ? node6189 : 4'b1101;
																assign node6189 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node6192 = (inp[1]) ? node6196 : node6193;
																assign node6193 = (inp[13]) ? 4'b1000 : 4'b1101;
																assign node6196 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node6199 = (inp[4]) ? node6207 : node6200;
															assign node6200 = (inp[13]) ? node6204 : node6201;
																assign node6201 = (inp[1]) ? 4'b1100 : 4'b1000;
																assign node6204 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node6207 = (inp[1]) ? node6209 : 4'b1101;
																assign node6209 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node6212 = (inp[4]) ? node6226 : node6213;
														assign node6213 = (inp[13]) ? node6221 : node6214;
															assign node6214 = (inp[2]) ? node6218 : node6215;
																assign node6215 = (inp[1]) ? 4'b1000 : 4'b1101;
																assign node6218 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node6221 = (inp[2]) ? 4'b1001 : node6222;
																assign node6222 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node6226 = (inp[2]) ? node6234 : node6227;
															assign node6227 = (inp[13]) ? node6231 : node6228;
																assign node6228 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node6231 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node6234 = (inp[1]) ? node6238 : node6235;
																assign node6235 = (inp[13]) ? 4'b1100 : 4'b1000;
																assign node6238 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node6241 = (inp[4]) ? node6261 : node6242;
													assign node6242 = (inp[0]) ? node6250 : node6243;
														assign node6243 = (inp[13]) ? 4'b1010 : node6244;
															assign node6244 = (inp[1]) ? node6246 : 4'b1111;
																assign node6246 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node6250 = (inp[13]) ? node6258 : node6251;
															assign node6251 = (inp[1]) ? node6255 : node6252;
																assign node6252 = (inp[2]) ? 4'b1010 : 4'b1111;
																assign node6255 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node6258 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node6261 = (inp[13]) ? node6271 : node6262;
														assign node6262 = (inp[0]) ? node6268 : node6263;
															assign node6263 = (inp[2]) ? 4'b1000 : node6264;
																assign node6264 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node6268 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node6271 = (inp[1]) ? node6275 : node6272;
															assign node6272 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node6275 = (inp[2]) ? node6277 : 4'b1000;
																assign node6277 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node6280 = (inp[4]) ? node6324 : node6281;
												assign node6281 = (inp[15]) ? node6305 : node6282;
													assign node6282 = (inp[13]) ? node6292 : node6283;
														assign node6283 = (inp[2]) ? node6289 : node6284;
															assign node6284 = (inp[1]) ? node6286 : 4'b1011;
																assign node6286 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node6289 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node6292 = (inp[2]) ? node6298 : node6293;
															assign node6293 = (inp[0]) ? 4'b1111 : node6294;
																assign node6294 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node6298 = (inp[1]) ? node6302 : node6299;
																assign node6299 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node6302 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node6305 = (inp[13]) ? node6315 : node6306;
														assign node6306 = (inp[2]) ? node6312 : node6307;
															assign node6307 = (inp[0]) ? 4'b1000 : node6308;
																assign node6308 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node6312 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node6315 = (inp[0]) ? node6319 : node6316;
															assign node6316 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node6319 = (inp[1]) ? node6321 : 4'b1101;
																assign node6321 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node6324 = (inp[1]) ? node6348 : node6325;
													assign node6325 = (inp[2]) ? node6335 : node6326;
														assign node6326 = (inp[15]) ? node6330 : node6327;
															assign node6327 = (inp[13]) ? 4'b1010 : 4'b1110;
															assign node6330 = (inp[13]) ? 4'b1111 : node6331;
																assign node6331 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6335 = (inp[0]) ? node6341 : node6336;
															assign node6336 = (inp[15]) ? 4'b1110 : node6337;
																assign node6337 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node6341 = (inp[13]) ? node6345 : node6342;
																assign node6342 = (inp[15]) ? 4'b1110 : 4'b1010;
																assign node6345 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node6348 = (inp[2]) ? node6358 : node6349;
														assign node6349 = (inp[15]) ? node6355 : node6350;
															assign node6350 = (inp[13]) ? node6352 : 4'b1111;
																assign node6352 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node6355 = (inp[13]) ? 4'b1111 : 4'b1010;
														assign node6358 = (inp[13]) ? node6364 : node6359;
															assign node6359 = (inp[15]) ? node6361 : 4'b1011;
																assign node6361 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node6364 = (inp[15]) ? 4'b1011 : 4'b1111;
										assign node6367 = (inp[12]) ? node6443 : node6368;
											assign node6368 = (inp[4]) ? node6402 : node6369;
												assign node6369 = (inp[15]) ? node6389 : node6370;
													assign node6370 = (inp[2]) ? node6378 : node6371;
														assign node6371 = (inp[0]) ? 4'b1011 : node6372;
															assign node6372 = (inp[13]) ? 4'b1010 : node6373;
																assign node6373 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node6378 = (inp[0]) ? node6384 : node6379;
															assign node6379 = (inp[13]) ? node6381 : 4'b1111;
																assign node6381 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node6384 = (inp[13]) ? 4'b1010 : node6385;
																assign node6385 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node6389 = (inp[13]) ? node6391 : 4'b1101;
														assign node6391 = (inp[2]) ? node6397 : node6392;
															assign node6392 = (inp[1]) ? node6394 : 4'b1000;
																assign node6394 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node6397 = (inp[1]) ? 4'b1101 : node6398;
																assign node6398 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node6402 = (inp[0]) ? node6424 : node6403;
													assign node6403 = (inp[1]) ? node6415 : node6404;
														assign node6404 = (inp[13]) ? node6410 : node6405;
															assign node6405 = (inp[15]) ? node6407 : 4'b1110;
																assign node6407 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node6410 = (inp[2]) ? 4'b1110 : node6411;
																assign node6411 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node6415 = (inp[2]) ? node6421 : node6416;
															assign node6416 = (inp[13]) ? 4'b1111 : node6417;
																assign node6417 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node6421 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node6424 = (inp[15]) ? node6436 : node6425;
														assign node6425 = (inp[13]) ? node6431 : node6426;
															assign node6426 = (inp[1]) ? 4'b1111 : node6427;
																assign node6427 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node6431 = (inp[2]) ? node6433 : 4'b1011;
																assign node6433 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node6436 = (inp[13]) ? node6438 : 4'b1010;
															assign node6438 = (inp[2]) ? 4'b1011 : node6439;
																assign node6439 = (inp[1]) ? 4'b1111 : 4'b1011;
											assign node6443 = (inp[15]) ? node6499 : node6444;
												assign node6444 = (inp[1]) ? node6474 : node6445;
													assign node6445 = (inp[0]) ? node6459 : node6446;
														assign node6446 = (inp[13]) ? node6454 : node6447;
															assign node6447 = (inp[2]) ? node6451 : node6448;
																assign node6448 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node6451 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node6454 = (inp[4]) ? node6456 : 4'b1101;
																assign node6456 = (inp[2]) ? 4'b1101 : 4'b1000;
														assign node6459 = (inp[4]) ? node6467 : node6460;
															assign node6460 = (inp[2]) ? node6464 : node6461;
																assign node6461 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node6464 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node6467 = (inp[2]) ? node6471 : node6468;
																assign node6468 = (inp[13]) ? 4'b1000 : 4'b1100;
																assign node6471 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node6474 = (inp[0]) ? node6488 : node6475;
														assign node6475 = (inp[13]) ? node6481 : node6476;
															assign node6476 = (inp[2]) ? node6478 : 4'b1100;
																assign node6478 = (inp[4]) ? 4'b1100 : 4'b1001;
															assign node6481 = (inp[2]) ? node6485 : node6482;
																assign node6482 = (inp[4]) ? 4'b1101 : 4'b1000;
																assign node6485 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node6488 = (inp[13]) ? node6494 : node6489;
															assign node6489 = (inp[2]) ? node6491 : 4'b1001;
																assign node6491 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node6494 = (inp[2]) ? node6496 : 4'b1101;
																assign node6496 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node6499 = (inp[4]) ? node6517 : node6500;
													assign node6500 = (inp[2]) ? node6510 : node6501;
														assign node6501 = (inp[13]) ? node6505 : node6502;
															assign node6502 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node6505 = (inp[1]) ? 4'b1110 : node6506;
																assign node6506 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node6510 = (inp[13]) ? node6514 : node6511;
															assign node6511 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node6514 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node6517 = (inp[13]) ? node6527 : node6518;
														assign node6518 = (inp[1]) ? node6522 : node6519;
															assign node6519 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node6522 = (inp[2]) ? node6524 : 4'b1000;
																assign node6524 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node6527 = (inp[0]) ? node6533 : node6528;
															assign node6528 = (inp[2]) ? node6530 : 4'b1001;
																assign node6530 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node6533 = (inp[1]) ? 4'b1101 : 4'b1000;
								assign node6536 = (inp[0]) ? node6844 : node6537;
									assign node6537 = (inp[13]) ? node6689 : node6538;
										assign node6538 = (inp[2]) ? node6616 : node6539;
											assign node6539 = (inp[5]) ? node6577 : node6540;
												assign node6540 = (inp[7]) ? node6558 : node6541;
													assign node6541 = (inp[12]) ? node6549 : node6542;
														assign node6542 = (inp[15]) ? node6544 : 4'b1000;
															assign node6544 = (inp[4]) ? 4'b1101 : node6545;
																assign node6545 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node6549 = (inp[4]) ? node6553 : node6550;
															assign node6550 = (inp[15]) ? 4'b1100 : 4'b1111;
															assign node6553 = (inp[1]) ? node6555 : 4'b1110;
																assign node6555 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node6558 = (inp[12]) ? node6566 : node6559;
														assign node6559 = (inp[4]) ? node6563 : node6560;
															assign node6560 = (inp[15]) ? 4'b1100 : 4'b1010;
															assign node6563 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node6566 = (inp[15]) ? node6572 : node6567;
															assign node6567 = (inp[1]) ? 4'b1100 : node6568;
																assign node6568 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node6572 = (inp[4]) ? node6574 : 4'b1011;
																assign node6574 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node6577 = (inp[4]) ? node6601 : node6578;
													assign node6578 = (inp[1]) ? node6588 : node6579;
														assign node6579 = (inp[15]) ? node6583 : node6580;
															assign node6580 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node6583 = (inp[12]) ? 4'b1110 : node6584;
																assign node6584 = (inp[7]) ? 4'b1100 : 4'b1110;
														assign node6588 = (inp[12]) ? node6594 : node6589;
															assign node6589 = (inp[7]) ? 4'b1010 : node6590;
																assign node6590 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node6594 = (inp[15]) ? node6598 : node6595;
																assign node6595 = (inp[7]) ? 4'b1101 : 4'b1010;
																assign node6598 = (inp[7]) ? 4'b1010 : 4'b1100;
													assign node6601 = (inp[1]) ? node6611 : node6602;
														assign node6602 = (inp[7]) ? node6608 : node6603;
															assign node6603 = (inp[12]) ? 4'b1111 : node6604;
																assign node6604 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node6608 = (inp[12]) ? 4'b1101 : 4'b1110;
														assign node6611 = (inp[12]) ? node6613 : 4'b1100;
															assign node6613 = (inp[15]) ? 4'b1001 : 4'b1000;
											assign node6616 = (inp[15]) ? node6652 : node6617;
												assign node6617 = (inp[7]) ? node6635 : node6618;
													assign node6618 = (inp[12]) ? node6624 : node6619;
														assign node6619 = (inp[4]) ? node6621 : 4'b1101;
															assign node6621 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node6624 = (inp[4]) ? node6628 : node6625;
															assign node6625 = (inp[1]) ? 4'b1010 : 4'b1111;
															assign node6628 = (inp[1]) ? node6632 : node6629;
																assign node6629 = (inp[5]) ? 4'b1011 : 4'b1010;
																assign node6632 = (inp[5]) ? 4'b1010 : 4'b1111;
													assign node6635 = (inp[12]) ? node6645 : node6636;
														assign node6636 = (inp[1]) ? node6640 : node6637;
															assign node6637 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node6640 = (inp[5]) ? 4'b1110 : node6641;
																assign node6641 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node6645 = (inp[4]) ? 4'b1100 : node6646;
															assign node6646 = (inp[1]) ? 4'b1000 : node6647;
																assign node6647 = (inp[5]) ? 4'b1101 : 4'b1000;
												assign node6652 = (inp[12]) ? node6676 : node6653;
													assign node6653 = (inp[1]) ? node6667 : node6654;
														assign node6654 = (inp[4]) ? node6660 : node6655;
															assign node6655 = (inp[7]) ? 4'b1001 : node6656;
																assign node6656 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node6660 = (inp[7]) ? node6664 : node6661;
																assign node6661 = (inp[5]) ? 4'b1101 : 4'b1000;
																assign node6664 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node6667 = (inp[4]) ? node6671 : node6668;
															assign node6668 = (inp[7]) ? 4'b1100 : 4'b1110;
															assign node6671 = (inp[7]) ? 4'b1111 : node6672;
																assign node6672 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node6676 = (inp[4]) ? node6682 : node6677;
														assign node6677 = (inp[7]) ? node6679 : 4'b1001;
															assign node6679 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node6682 = (inp[7]) ? node6684 : 4'b1111;
															assign node6684 = (inp[5]) ? node6686 : 4'b1101;
																assign node6686 = (inp[1]) ? 4'b1101 : 4'b1001;
										assign node6689 = (inp[2]) ? node6763 : node6690;
											assign node6690 = (inp[5]) ? node6728 : node6691;
												assign node6691 = (inp[12]) ? node6709 : node6692;
													assign node6692 = (inp[15]) ? node6696 : node6693;
														assign node6693 = (inp[7]) ? 4'b1110 : 4'b1100;
														assign node6696 = (inp[1]) ? node6704 : node6697;
															assign node6697 = (inp[7]) ? node6701 : node6698;
																assign node6698 = (inp[4]) ? 4'b1000 : 4'b1111;
																assign node6701 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node6704 = (inp[4]) ? 4'b1110 : node6705;
																assign node6705 = (inp[7]) ? 4'b1100 : 4'b1110;
													assign node6709 = (inp[7]) ? node6719 : node6710;
														assign node6710 = (inp[15]) ? node6714 : node6711;
															assign node6711 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node6714 = (inp[4]) ? 4'b1010 : node6715;
																assign node6715 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node6719 = (inp[15]) ? node6725 : node6720;
															assign node6720 = (inp[4]) ? 4'b1100 : node6721;
																assign node6721 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node6725 = (inp[4]) ? 4'b1101 : 4'b1110;
												assign node6728 = (inp[1]) ? node6746 : node6729;
													assign node6729 = (inp[12]) ? node6735 : node6730;
														assign node6730 = (inp[7]) ? 4'b1010 : node6731;
															assign node6731 = (inp[15]) ? 4'b1100 : 4'b1001;
														assign node6735 = (inp[7]) ? node6743 : node6736;
															assign node6736 = (inp[4]) ? node6740 : node6737;
																assign node6737 = (inp[15]) ? 4'b1100 : 4'b1111;
																assign node6740 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node6743 = (inp[4]) ? 4'b1001 : 4'b1100;
													assign node6746 = (inp[15]) ? node6754 : node6747;
														assign node6747 = (inp[12]) ? node6751 : node6748;
															assign node6748 = (inp[7]) ? 4'b1110 : 4'b1101;
															assign node6751 = (inp[7]) ? 4'b1100 : 4'b1110;
														assign node6754 = (inp[4]) ? 4'b1100 : node6755;
															assign node6755 = (inp[12]) ? node6759 : node6756;
																assign node6756 = (inp[7]) ? 4'b1000 : 4'b1110;
																assign node6759 = (inp[7]) ? 4'b1111 : 4'b1000;
											assign node6763 = (inp[7]) ? node6809 : node6764;
												assign node6764 = (inp[12]) ? node6786 : node6765;
													assign node6765 = (inp[4]) ? node6773 : node6766;
														assign node6766 = (inp[15]) ? 4'b1011 : node6767;
															assign node6767 = (inp[5]) ? node6769 : 4'b1001;
																assign node6769 = (inp[1]) ? 4'b1000 : 4'b1101;
														assign node6773 = (inp[15]) ? node6779 : node6774;
															assign node6774 = (inp[5]) ? node6776 : 4'b1000;
																assign node6776 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node6779 = (inp[1]) ? node6783 : node6780;
																assign node6780 = (inp[5]) ? 4'b1000 : 4'b1101;
																assign node6783 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node6786 = (inp[1]) ? node6798 : node6787;
														assign node6787 = (inp[4]) ? node6795 : node6788;
															assign node6788 = (inp[15]) ? node6792 : node6789;
																assign node6789 = (inp[5]) ? 4'b1010 : 4'b1011;
																assign node6792 = (inp[5]) ? 4'b1001 : 4'b1100;
															assign node6795 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node6798 = (inp[4]) ? node6802 : node6799;
															assign node6799 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node6802 = (inp[5]) ? node6806 : node6803;
																assign node6803 = (inp[15]) ? 4'b1111 : 4'b1010;
																assign node6806 = (inp[15]) ? 4'b1010 : 4'b1110;
												assign node6809 = (inp[12]) ? node6827 : node6810;
													assign node6810 = (inp[4]) ? node6822 : node6811;
														assign node6811 = (inp[15]) ? node6817 : node6812;
															assign node6812 = (inp[1]) ? 4'b1011 : node6813;
																assign node6813 = (inp[5]) ? 4'b1110 : 4'b1011;
															assign node6817 = (inp[1]) ? node6819 : 4'b1100;
																assign node6819 = (inp[5]) ? 4'b1100 : 4'b1001;
														assign node6822 = (inp[5]) ? node6824 : 4'b1010;
															assign node6824 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node6827 = (inp[1]) ? node6837 : node6828;
														assign node6828 = (inp[5]) ? node6834 : node6829;
															assign node6829 = (inp[15]) ? 4'b1011 : node6830;
																assign node6830 = (inp[4]) ? 4'b1001 : 4'b1100;
															assign node6834 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node6837 = (inp[4]) ? 4'b1000 : node6838;
															assign node6838 = (inp[15]) ? node6840 : 4'b1100;
																assign node6840 = (inp[5]) ? 4'b1010 : 4'b1011;
									assign node6844 = (inp[15]) ? node7000 : node6845;
										assign node6845 = (inp[13]) ? node6931 : node6846;
											assign node6846 = (inp[2]) ? node6882 : node6847;
												assign node6847 = (inp[5]) ? node6859 : node6848;
													assign node6848 = (inp[7]) ? node6854 : node6849;
														assign node6849 = (inp[12]) ? node6851 : 4'b1001;
															assign node6851 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node6854 = (inp[12]) ? node6856 : 4'b1011;
															assign node6856 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node6859 = (inp[1]) ? node6869 : node6860;
														assign node6860 = (inp[12]) ? node6864 : node6861;
															assign node6861 = (inp[7]) ? 4'b1110 : 4'b1101;
															assign node6864 = (inp[4]) ? 4'b1110 : node6865;
																assign node6865 = (inp[7]) ? 4'b1001 : 4'b1011;
														assign node6869 = (inp[4]) ? node6877 : node6870;
															assign node6870 = (inp[12]) ? node6874 : node6871;
																assign node6871 = (inp[7]) ? 4'b1010 : 4'b1001;
																assign node6874 = (inp[7]) ? 4'b1100 : 4'b1010;
															assign node6877 = (inp[7]) ? node6879 : 4'b1111;
																assign node6879 = (inp[12]) ? 4'b1001 : 4'b1011;
												assign node6882 = (inp[12]) ? node6904 : node6883;
													assign node6883 = (inp[7]) ? node6897 : node6884;
														assign node6884 = (inp[1]) ? node6890 : node6885;
															assign node6885 = (inp[5]) ? 4'b1000 : node6886;
																assign node6886 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node6890 = (inp[4]) ? node6894 : node6891;
																assign node6891 = (inp[5]) ? 4'b1100 : 4'b1101;
																assign node6894 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node6897 = (inp[4]) ? node6901 : node6898;
															assign node6898 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node6901 = (inp[5]) ? 4'b1010 : 4'b1110;
													assign node6904 = (inp[7]) ? node6918 : node6905;
														assign node6905 = (inp[4]) ? node6913 : node6906;
															assign node6906 = (inp[1]) ? node6910 : node6907;
																assign node6907 = (inp[5]) ? 4'b1110 : 4'b1111;
																assign node6910 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node6913 = (inp[1]) ? 4'b1011 : node6914;
																assign node6914 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node6918 = (inp[5]) ? node6926 : node6919;
															assign node6919 = (inp[4]) ? node6923 : node6920;
																assign node6920 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node6923 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node6926 = (inp[4]) ? 4'b1001 : node6927;
																assign node6927 = (inp[1]) ? 4'b1001 : 4'b1101;
											assign node6931 = (inp[2]) ? node6965 : node6932;
												assign node6932 = (inp[5]) ? node6946 : node6933;
													assign node6933 = (inp[12]) ? node6937 : node6934;
														assign node6934 = (inp[7]) ? 4'b1111 : 4'b1101;
														assign node6937 = (inp[7]) ? node6943 : node6938;
															assign node6938 = (inp[1]) ? 4'b1010 : node6939;
																assign node6939 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node6943 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node6946 = (inp[1]) ? node6954 : node6947;
														assign node6947 = (inp[4]) ? node6949 : 4'b1101;
															assign node6949 = (inp[12]) ? node6951 : 4'b1000;
																assign node6951 = (inp[7]) ? 4'b1000 : 4'b1010;
														assign node6954 = (inp[12]) ? node6962 : node6955;
															assign node6955 = (inp[7]) ? node6959 : node6956;
																assign node6956 = (inp[4]) ? 4'b1100 : 4'b1101;
																assign node6959 = (inp[4]) ? 4'b1111 : 4'b1110;
															assign node6962 = (inp[7]) ? 4'b1000 : 4'b1110;
												assign node6965 = (inp[7]) ? node6983 : node6966;
													assign node6966 = (inp[12]) ? node6976 : node6967;
														assign node6967 = (inp[1]) ? 4'b1000 : node6968;
															assign node6968 = (inp[5]) ? node6972 : node6969;
																assign node6969 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node6972 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node6976 = (inp[5]) ? node6978 : 4'b1010;
															assign node6978 = (inp[4]) ? node6980 : 4'b1010;
																assign node6980 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node6983 = (inp[12]) ? node6993 : node6984;
														assign node6984 = (inp[1]) ? 4'b1011 : node6985;
															assign node6985 = (inp[5]) ? node6989 : node6986;
																assign node6986 = (inp[4]) ? 4'b1011 : 4'b1010;
																assign node6989 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node6993 = (inp[4]) ? 4'b1101 : node6994;
															assign node6994 = (inp[5]) ? 4'b1000 : node6995;
																assign node6995 = (inp[1]) ? 4'b1101 : 4'b1100;
										assign node7000 = (inp[4]) ? node7086 : node7001;
											assign node7001 = (inp[12]) ? node7043 : node7002;
												assign node7002 = (inp[7]) ? node7020 : node7003;
													assign node7003 = (inp[5]) ? node7011 : node7004;
														assign node7004 = (inp[13]) ? node7008 : node7005;
															assign node7005 = (inp[2]) ? 4'b1110 : 4'b1011;
															assign node7008 = (inp[2]) ? 4'b1011 : 4'b1110;
														assign node7011 = (inp[1]) ? node7013 : 4'b1010;
															assign node7013 = (inp[13]) ? node7017 : node7014;
																assign node7014 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node7017 = (inp[2]) ? 4'b1010 : 4'b1111;
													assign node7020 = (inp[5]) ? node7036 : node7021;
														assign node7021 = (inp[13]) ? node7029 : node7022;
															assign node7022 = (inp[1]) ? node7026 : node7023;
																assign node7023 = (inp[2]) ? 4'b1000 : 4'b1101;
																assign node7026 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node7029 = (inp[2]) ? node7033 : node7030;
																assign node7030 = (inp[1]) ? 4'b1101 : 4'b1000;
																assign node7033 = (inp[1]) ? 4'b1000 : 4'b1101;
														assign node7036 = (inp[2]) ? node7040 : node7037;
															assign node7037 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node7040 = (inp[1]) ? 4'b1000 : 4'b1001;
												assign node7043 = (inp[7]) ? node7067 : node7044;
													assign node7044 = (inp[2]) ? node7056 : node7045;
														assign node7045 = (inp[13]) ? node7051 : node7046;
															assign node7046 = (inp[5]) ? node7048 : 4'b1100;
																assign node7048 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node7051 = (inp[5]) ? node7053 : 4'b1000;
																assign node7053 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node7056 = (inp[13]) ? node7060 : node7057;
															assign node7057 = (inp[1]) ? 4'b1001 : 4'b1100;
															assign node7060 = (inp[1]) ? node7064 : node7061;
																assign node7061 = (inp[5]) ? 4'b1001 : 4'b1101;
																assign node7064 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node7067 = (inp[2]) ? node7079 : node7068;
														assign node7068 = (inp[13]) ? node7074 : node7069;
															assign node7069 = (inp[5]) ? 4'b1111 : node7070;
																assign node7070 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node7074 = (inp[1]) ? 4'b1110 : node7075;
																assign node7075 = (inp[5]) ? 4'b1010 : 4'b1111;
														assign node7079 = (inp[13]) ? node7083 : node7080;
															assign node7080 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node7083 = (inp[5]) ? 4'b1011 : 4'b1010;
											assign node7086 = (inp[2]) ? node7130 : node7087;
												assign node7087 = (inp[13]) ? node7107 : node7088;
													assign node7088 = (inp[5]) ? node7096 : node7089;
														assign node7089 = (inp[7]) ? node7093 : node7090;
															assign node7090 = (inp[12]) ? 4'b1111 : 4'b1101;
															assign node7093 = (inp[1]) ? 4'b1010 : 4'b1000;
														assign node7096 = (inp[12]) ? node7102 : node7097;
															assign node7097 = (inp[7]) ? 4'b1010 : node7098;
																assign node7098 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node7102 = (inp[7]) ? node7104 : 4'b1010;
																assign node7104 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node7107 = (inp[5]) ? node7121 : node7108;
														assign node7108 = (inp[7]) ? node7116 : node7109;
															assign node7109 = (inp[12]) ? node7113 : node7110;
																assign node7110 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node7113 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node7116 = (inp[12]) ? 4'b1101 : node7117;
																assign node7117 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node7121 = (inp[7]) ? node7125 : node7122;
															assign node7122 = (inp[12]) ? 4'b1111 : 4'b1101;
															assign node7125 = (inp[1]) ? node7127 : 4'b1010;
																assign node7127 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node7130 = (inp[1]) ? node7150 : node7131;
													assign node7131 = (inp[5]) ? node7143 : node7132;
														assign node7132 = (inp[13]) ? node7140 : node7133;
															assign node7133 = (inp[12]) ? node7137 : node7134;
																assign node7134 = (inp[7]) ? 4'b1111 : 4'b1001;
																assign node7137 = (inp[7]) ? 4'b1100 : 4'b1111;
															assign node7140 = (inp[7]) ? 4'b1001 : 4'b1010;
														assign node7143 = (inp[13]) ? node7147 : node7144;
															assign node7144 = (inp[12]) ? 4'b1110 : 4'b1101;
															assign node7147 = (inp[12]) ? 4'b1101 : 4'b1110;
													assign node7150 = (inp[7]) ? node7166 : node7151;
														assign node7151 = (inp[12]) ? node7159 : node7152;
															assign node7152 = (inp[13]) ? node7156 : node7153;
																assign node7153 = (inp[5]) ? 4'b1000 : 4'b1001;
																assign node7156 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node7159 = (inp[5]) ? node7163 : node7160;
																assign node7160 = (inp[13]) ? 4'b1110 : 4'b1011;
																assign node7163 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node7166 = (inp[12]) ? node7168 : 4'b1011;
															assign node7168 = (inp[13]) ? 4'b1001 : 4'b1101;
						assign node7171 = (inp[9]) ? node8411 : node7172;
							assign node7172 = (inp[11]) ? node7800 : node7173;
								assign node7173 = (inp[15]) ? node7479 : node7174;
									assign node7174 = (inp[5]) ? node7288 : node7175;
										assign node7175 = (inp[2]) ? node7223 : node7176;
											assign node7176 = (inp[13]) ? node7196 : node7177;
												assign node7177 = (inp[12]) ? node7181 : node7178;
													assign node7178 = (inp[7]) ? 4'b1011 : 4'b1001;
													assign node7181 = (inp[7]) ? node7189 : node7182;
														assign node7182 = (inp[1]) ? node7186 : node7183;
															assign node7183 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node7186 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node7189 = (inp[4]) ? 4'b1001 : node7190;
															assign node7190 = (inp[1]) ? 4'b1100 : node7191;
																assign node7191 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node7196 = (inp[12]) ? node7200 : node7197;
													assign node7197 = (inp[7]) ? 4'b1111 : 4'b1101;
													assign node7200 = (inp[7]) ? node7216 : node7201;
														assign node7201 = (inp[0]) ? node7209 : node7202;
															assign node7202 = (inp[1]) ? node7206 : node7203;
																assign node7203 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node7206 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node7209 = (inp[4]) ? node7213 : node7210;
																assign node7210 = (inp[1]) ? 4'b1011 : 4'b1111;
																assign node7213 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node7216 = (inp[4]) ? node7220 : node7217;
															assign node7217 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node7220 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node7223 = (inp[13]) ? node7261 : node7224;
												assign node7224 = (inp[12]) ? node7244 : node7225;
													assign node7225 = (inp[7]) ? node7237 : node7226;
														assign node7226 = (inp[1]) ? node7232 : node7227;
															assign node7227 = (inp[4]) ? 4'b1101 : node7228;
																assign node7228 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node7232 = (inp[4]) ? node7234 : 4'b1100;
																assign node7234 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node7237 = (inp[0]) ? node7241 : node7238;
															assign node7238 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node7241 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node7244 = (inp[7]) ? node7252 : node7245;
														assign node7245 = (inp[1]) ? node7249 : node7246;
															assign node7246 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node7249 = (inp[4]) ? 4'b1110 : 4'b1011;
														assign node7252 = (inp[4]) ? node7256 : node7253;
															assign node7253 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node7256 = (inp[0]) ? node7258 : 4'b1101;
																assign node7258 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node7261 = (inp[4]) ? node7275 : node7262;
													assign node7262 = (inp[12]) ? node7266 : node7263;
														assign node7263 = (inp[7]) ? 4'b1010 : 4'b1000;
														assign node7266 = (inp[7]) ? node7270 : node7267;
															assign node7267 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node7270 = (inp[0]) ? 4'b1100 : node7271;
																assign node7271 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node7275 = (inp[12]) ? node7279 : node7276;
														assign node7276 = (inp[7]) ? 4'b1011 : 4'b1001;
														assign node7279 = (inp[7]) ? node7285 : node7280;
															assign node7280 = (inp[1]) ? node7282 : 4'b1111;
																assign node7282 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node7285 = (inp[1]) ? 4'b1001 : 4'b1000;
										assign node7288 = (inp[7]) ? node7380 : node7289;
											assign node7289 = (inp[12]) ? node7337 : node7290;
												assign node7290 = (inp[0]) ? node7320 : node7291;
													assign node7291 = (inp[2]) ? node7307 : node7292;
														assign node7292 = (inp[4]) ? node7300 : node7293;
															assign node7293 = (inp[13]) ? node7297 : node7294;
																assign node7294 = (inp[1]) ? 4'b1001 : 4'b1101;
																assign node7297 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node7300 = (inp[1]) ? node7304 : node7301;
																assign node7301 = (inp[13]) ? 4'b1000 : 4'b1101;
																assign node7304 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node7307 = (inp[4]) ? node7315 : node7308;
															assign node7308 = (inp[13]) ? node7312 : node7309;
																assign node7309 = (inp[1]) ? 4'b1100 : 4'b1000;
																assign node7312 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node7315 = (inp[1]) ? 4'b1101 : node7316;
																assign node7316 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node7320 = (inp[1]) ? node7330 : node7321;
														assign node7321 = (inp[4]) ? node7323 : 4'b1000;
															assign node7323 = (inp[2]) ? node7327 : node7324;
																assign node7324 = (inp[13]) ? 4'b1000 : 4'b1100;
																assign node7327 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node7330 = (inp[2]) ? node7332 : 4'b1100;
															assign node7332 = (inp[13]) ? node7334 : 4'b1100;
																assign node7334 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node7337 = (inp[1]) ? node7355 : node7338;
													assign node7338 = (inp[13]) ? node7344 : node7339;
														assign node7339 = (inp[4]) ? node7341 : 4'b1110;
															assign node7341 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node7344 = (inp[2]) ? node7350 : node7345;
															assign node7345 = (inp[4]) ? 4'b1011 : node7346;
																assign node7346 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node7350 = (inp[4]) ? 4'b1110 : node7351;
																assign node7351 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node7355 = (inp[4]) ? node7367 : node7356;
														assign node7356 = (inp[0]) ? node7362 : node7357;
															assign node7357 = (inp[2]) ? 4'b1111 : node7358;
																assign node7358 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node7362 = (inp[2]) ? 4'b1010 : node7363;
																assign node7363 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node7367 = (inp[0]) ? node7375 : node7368;
															assign node7368 = (inp[13]) ? node7372 : node7369;
																assign node7369 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node7372 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node7375 = (inp[2]) ? node7377 : 4'b1010;
																assign node7377 = (inp[13]) ? 4'b1111 : 4'b1011;
											assign node7380 = (inp[12]) ? node7432 : node7381;
												assign node7381 = (inp[0]) ? node7413 : node7382;
													assign node7382 = (inp[2]) ? node7398 : node7383;
														assign node7383 = (inp[4]) ? node7391 : node7384;
															assign node7384 = (inp[1]) ? node7388 : node7385;
																assign node7385 = (inp[13]) ? 4'b1010 : 4'b1110;
																assign node7388 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node7391 = (inp[1]) ? node7395 : node7392;
																assign node7392 = (inp[13]) ? 4'b1011 : 4'b1110;
																assign node7395 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node7398 = (inp[4]) ? node7406 : node7399;
															assign node7399 = (inp[13]) ? node7403 : node7400;
																assign node7400 = (inp[1]) ? 4'b1111 : 4'b1011;
																assign node7403 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node7406 = (inp[1]) ? node7410 : node7407;
																assign node7407 = (inp[13]) ? 4'b1110 : 4'b1010;
																assign node7410 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node7413 = (inp[4]) ? node7425 : node7414;
														assign node7414 = (inp[2]) ? node7420 : node7415;
															assign node7415 = (inp[1]) ? node7417 : 4'b1011;
																assign node7417 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node7420 = (inp[13]) ? node7422 : 4'b1111;
																assign node7422 = (inp[1]) ? 4'b1010 : 4'b1111;
														assign node7425 = (inp[2]) ? node7427 : 4'b1011;
															assign node7427 = (inp[13]) ? node7429 : 4'b1011;
																assign node7429 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node7432 = (inp[0]) ? node7450 : node7433;
													assign node7433 = (inp[13]) ? node7443 : node7434;
														assign node7434 = (inp[1]) ? 4'b1001 : node7435;
															assign node7435 = (inp[4]) ? node7439 : node7436;
																assign node7436 = (inp[2]) ? 4'b1101 : 4'b1001;
																assign node7439 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node7443 = (inp[1]) ? node7445 : 4'b1101;
															assign node7445 = (inp[4]) ? node7447 : 4'b1101;
																assign node7447 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node7450 = (inp[1]) ? node7466 : node7451;
														assign node7451 = (inp[4]) ? node7459 : node7452;
															assign node7452 = (inp[2]) ? node7456 : node7453;
																assign node7453 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node7456 = (inp[13]) ? 4'b1000 : 4'b1100;
															assign node7459 = (inp[13]) ? node7463 : node7460;
																assign node7460 = (inp[2]) ? 4'b1000 : 4'b1100;
																assign node7463 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node7466 = (inp[2]) ? node7472 : node7467;
															assign node7467 = (inp[13]) ? node7469 : 4'b1100;
																assign node7469 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node7472 = (inp[13]) ? node7476 : node7473;
																assign node7473 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node7476 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node7479 = (inp[13]) ? node7649 : node7480;
										assign node7480 = (inp[0]) ? node7560 : node7481;
											assign node7481 = (inp[5]) ? node7521 : node7482;
												assign node7482 = (inp[7]) ? node7506 : node7483;
													assign node7483 = (inp[4]) ? node7495 : node7484;
														assign node7484 = (inp[12]) ? node7488 : node7485;
															assign node7485 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node7488 = (inp[2]) ? node7492 : node7489;
																assign node7489 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node7492 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node7495 = (inp[12]) ? node7499 : node7496;
															assign node7496 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node7499 = (inp[1]) ? node7503 : node7500;
																assign node7500 = (inp[2]) ? 4'b1111 : 4'b1011;
																assign node7503 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node7506 = (inp[2]) ? node7514 : node7507;
														assign node7507 = (inp[4]) ? 4'b1000 : node7508;
															assign node7508 = (inp[12]) ? node7510 : 4'b1000;
																assign node7510 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node7514 = (inp[4]) ? 4'b1101 : node7515;
															assign node7515 = (inp[12]) ? 4'b1110 : node7516;
																assign node7516 = (inp[1]) ? 4'b1100 : 4'b1000;
												assign node7521 = (inp[7]) ? node7547 : node7522;
													assign node7522 = (inp[2]) ? node7534 : node7523;
														assign node7523 = (inp[4]) ? node7531 : node7524;
															assign node7524 = (inp[12]) ? node7528 : node7525;
																assign node7525 = (inp[1]) ? 4'b1010 : 4'b1111;
																assign node7528 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node7531 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node7534 = (inp[4]) ? node7542 : node7535;
															assign node7535 = (inp[12]) ? node7539 : node7536;
																assign node7536 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node7539 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node7542 = (inp[12]) ? node7544 : 4'b1101;
																assign node7544 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node7547 = (inp[12]) ? node7557 : node7548;
														assign node7548 = (inp[2]) ? node7554 : node7549;
															assign node7549 = (inp[4]) ? 4'b1111 : node7550;
																assign node7550 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node7554 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node7557 = (inp[4]) ? 4'b1101 : 4'b1111;
											assign node7560 = (inp[2]) ? node7606 : node7561;
												assign node7561 = (inp[1]) ? node7585 : node7562;
													assign node7562 = (inp[4]) ? node7574 : node7563;
														assign node7563 = (inp[5]) ? node7569 : node7564;
															assign node7564 = (inp[12]) ? 4'b1010 : node7565;
																assign node7565 = (inp[7]) ? 4'b1101 : 4'b1011;
															assign node7569 = (inp[12]) ? 4'b1111 : node7570;
																assign node7570 = (inp[7]) ? 4'b1101 : 4'b1111;
														assign node7574 = (inp[7]) ? node7580 : node7575;
															assign node7575 = (inp[12]) ? 4'b1011 : node7576;
																assign node7576 = (inp[5]) ? 4'b1000 : 4'b1101;
															assign node7580 = (inp[12]) ? 4'b1100 : node7581;
																assign node7581 = (inp[5]) ? 4'b1111 : 4'b1010;
													assign node7585 = (inp[7]) ? node7595 : node7586;
														assign node7586 = (inp[4]) ? node7590 : node7587;
															assign node7587 = (inp[12]) ? 4'b1101 : 4'b1010;
															assign node7590 = (inp[12]) ? 4'b1010 : node7591;
																assign node7591 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node7595 = (inp[4]) ? node7603 : node7596;
															assign node7596 = (inp[12]) ? node7600 : node7597;
																assign node7597 = (inp[5]) ? 4'b1101 : 4'b1000;
																assign node7600 = (inp[5]) ? 4'b1011 : 4'b1010;
															assign node7603 = (inp[12]) ? 4'b1000 : 4'b1010;
												assign node7606 = (inp[4]) ? node7628 : node7607;
													assign node7607 = (inp[12]) ? node7621 : node7608;
														assign node7608 = (inp[7]) ? node7616 : node7609;
															assign node7609 = (inp[1]) ? node7613 : node7610;
																assign node7610 = (inp[5]) ? 4'b1010 : 4'b1110;
																assign node7613 = (inp[5]) ? 4'b1111 : 4'b1110;
															assign node7616 = (inp[5]) ? 4'b1000 : node7617;
																assign node7617 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node7621 = (inp[7]) ? 4'b1110 : node7622;
															assign node7622 = (inp[5]) ? node7624 : 4'b1000;
																assign node7624 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node7628 = (inp[5]) ? node7638 : node7629;
														assign node7629 = (inp[7]) ? node7633 : node7630;
															assign node7630 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node7633 = (inp[12]) ? 4'b1100 : node7634;
																assign node7634 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node7638 = (inp[1]) ? node7644 : node7639;
															assign node7639 = (inp[7]) ? 4'b1000 : node7640;
																assign node7640 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node7644 = (inp[12]) ? node7646 : 4'b1110;
																assign node7646 = (inp[7]) ? 4'b1100 : 4'b1110;
										assign node7649 = (inp[1]) ? node7739 : node7650;
											assign node7650 = (inp[12]) ? node7696 : node7651;
												assign node7651 = (inp[0]) ? node7673 : node7652;
													assign node7652 = (inp[2]) ? node7660 : node7653;
														assign node7653 = (inp[4]) ? node7657 : node7654;
															assign node7654 = (inp[7]) ? 4'b1000 : 4'b1010;
															assign node7657 = (inp[7]) ? 4'b1110 : 4'b1000;
														assign node7660 = (inp[4]) ? node7668 : node7661;
															assign node7661 = (inp[7]) ? node7665 : node7662;
																assign node7662 = (inp[5]) ? 4'b1111 : 4'b1011;
																assign node7665 = (inp[5]) ? 4'b1100 : 4'b1101;
															assign node7668 = (inp[7]) ? node7670 : 4'b1100;
																assign node7670 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node7673 = (inp[2]) ? node7687 : node7674;
														assign node7674 = (inp[4]) ? node7682 : node7675;
															assign node7675 = (inp[7]) ? node7679 : node7676;
																assign node7676 = (inp[5]) ? 4'b1011 : 4'b1110;
																assign node7679 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node7682 = (inp[7]) ? node7684 : 4'b1101;
																assign node7684 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node7687 = (inp[5]) ? node7689 : 4'b1100;
															assign node7689 = (inp[7]) ? node7693 : node7690;
																assign node7690 = (inp[4]) ? 4'b1001 : 4'b1111;
																assign node7693 = (inp[4]) ? 4'b1110 : 4'b1101;
												assign node7696 = (inp[0]) ? node7718 : node7697;
													assign node7697 = (inp[4]) ? node7709 : node7698;
														assign node7698 = (inp[7]) ? node7704 : node7699;
															assign node7699 = (inp[2]) ? 4'b1101 : node7700;
																assign node7700 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node7704 = (inp[5]) ? 4'b1111 : node7705;
																assign node7705 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node7709 = (inp[7]) ? node7713 : node7710;
															assign node7710 = (inp[2]) ? 4'b1011 : 4'b1111;
															assign node7713 = (inp[5]) ? node7715 : 4'b1101;
																assign node7715 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node7718 = (inp[4]) ? node7732 : node7719;
														assign node7719 = (inp[7]) ? node7727 : node7720;
															assign node7720 = (inp[5]) ? node7724 : node7721;
																assign node7721 = (inp[2]) ? 4'b1101 : 4'b1001;
																assign node7724 = (inp[2]) ? 4'b1000 : 4'b1101;
															assign node7727 = (inp[2]) ? node7729 : 4'b1111;
																assign node7729 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node7732 = (inp[2]) ? node7736 : node7733;
															assign node7733 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node7736 = (inp[5]) ? 4'b1101 : 4'b1000;
											assign node7739 = (inp[4]) ? node7773 : node7740;
												assign node7740 = (inp[2]) ? node7756 : node7741;
													assign node7741 = (inp[12]) ? node7749 : node7742;
														assign node7742 = (inp[7]) ? node7746 : node7743;
															assign node7743 = (inp[5]) ? 4'b1111 : 4'b1110;
															assign node7746 = (inp[5]) ? 4'b1001 : 4'b1101;
														assign node7749 = (inp[7]) ? 4'b1110 : node7750;
															assign node7750 = (inp[5]) ? node7752 : 4'b1000;
																assign node7752 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node7756 = (inp[12]) ? node7766 : node7757;
														assign node7757 = (inp[7]) ? node7763 : node7758;
															assign node7758 = (inp[0]) ? 4'b1010 : node7759;
																assign node7759 = (inp[5]) ? 4'b1010 : 4'b1011;
															assign node7763 = (inp[5]) ? 4'b1101 : 4'b1000;
														assign node7766 = (inp[7]) ? 4'b1011 : node7767;
															assign node7767 = (inp[5]) ? 4'b1101 : node7768;
																assign node7768 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node7773 = (inp[7]) ? node7793 : node7774;
													assign node7774 = (inp[12]) ? node7786 : node7775;
														assign node7775 = (inp[2]) ? node7779 : node7776;
															assign node7776 = (inp[5]) ? 4'b1000 : 4'b1001;
															assign node7779 = (inp[0]) ? node7783 : node7780;
																assign node7780 = (inp[5]) ? 4'b1101 : 4'b1100;
																assign node7783 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node7786 = (inp[5]) ? node7790 : node7787;
															assign node7787 = (inp[0]) ? 4'b1110 : 4'b1010;
															assign node7790 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node7793 = (inp[12]) ? node7797 : node7794;
														assign node7794 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node7797 = (inp[2]) ? 4'b1001 : 4'b1101;
								assign node7800 = (inp[0]) ? node8088 : node7801;
									assign node7801 = (inp[2]) ? node7939 : node7802;
										assign node7802 = (inp[13]) ? node7878 : node7803;
											assign node7803 = (inp[5]) ? node7831 : node7804;
												assign node7804 = (inp[7]) ? node7816 : node7805;
													assign node7805 = (inp[12]) ? node7809 : node7806;
														assign node7806 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node7809 = (inp[4]) ? node7811 : 4'b1100;
															assign node7811 = (inp[15]) ? node7813 : 4'b1110;
																assign node7813 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node7816 = (inp[12]) ? node7822 : node7817;
														assign node7817 = (inp[15]) ? node7819 : 4'b1010;
															assign node7819 = (inp[4]) ? 4'b1011 : 4'b1100;
														assign node7822 = (inp[15]) ? node7826 : node7823;
															assign node7823 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node7826 = (inp[4]) ? node7828 : 4'b1011;
																assign node7828 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node7831 = (inp[7]) ? node7857 : node7832;
													assign node7832 = (inp[12]) ? node7846 : node7833;
														assign node7833 = (inp[1]) ? node7839 : node7834;
															assign node7834 = (inp[15]) ? 4'b1001 : node7835;
																assign node7835 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node7839 = (inp[4]) ? node7843 : node7840;
																assign node7840 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node7843 = (inp[15]) ? 4'b1100 : 4'b1001;
														assign node7846 = (inp[15]) ? node7850 : node7847;
															assign node7847 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node7850 = (inp[4]) ? node7854 : node7851;
																assign node7851 = (inp[1]) ? 4'b1100 : 4'b1001;
																assign node7854 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node7857 = (inp[12]) ? node7869 : node7858;
														assign node7858 = (inp[1]) ? node7864 : node7859;
															assign node7859 = (inp[15]) ? node7861 : 4'b1111;
																assign node7861 = (inp[4]) ? 4'b1110 : 4'b1100;
															assign node7864 = (inp[15]) ? node7866 : 4'b1010;
																assign node7866 = (inp[4]) ? 4'b1011 : 4'b1100;
														assign node7869 = (inp[15]) ? 4'b1010 : node7870;
															assign node7870 = (inp[1]) ? node7874 : node7871;
																assign node7871 = (inp[4]) ? 4'b1101 : 4'b1000;
																assign node7874 = (inp[4]) ? 4'b1000 : 4'b1101;
											assign node7878 = (inp[7]) ? node7918 : node7879;
												assign node7879 = (inp[12]) ? node7897 : node7880;
													assign node7880 = (inp[4]) ? node7888 : node7881;
														assign node7881 = (inp[15]) ? node7883 : 4'b1101;
															assign node7883 = (inp[5]) ? 4'b1010 : node7884;
																assign node7884 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node7888 = (inp[5]) ? node7892 : node7889;
															assign node7889 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node7892 = (inp[15]) ? node7894 : 4'b1001;
																assign node7894 = (inp[1]) ? 4'b1001 : 4'b1100;
													assign node7897 = (inp[4]) ? node7905 : node7898;
														assign node7898 = (inp[15]) ? node7900 : 4'b1110;
															assign node7900 = (inp[1]) ? 4'b1001 : node7901;
																assign node7901 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node7905 = (inp[15]) ? node7913 : node7906;
															assign node7906 = (inp[1]) ? node7910 : node7907;
																assign node7907 = (inp[5]) ? 4'b1010 : 4'b1011;
																assign node7910 = (inp[5]) ? 4'b1011 : 4'b1110;
															assign node7913 = (inp[1]) ? 4'b1110 : node7914;
																assign node7914 = (inp[5]) ? 4'b1111 : 4'b1110;
												assign node7918 = (inp[12]) ? node7924 : node7919;
													assign node7919 = (inp[5]) ? node7921 : 4'b1110;
														assign node7921 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node7924 = (inp[1]) ? node7932 : node7925;
														assign node7925 = (inp[4]) ? node7929 : node7926;
															assign node7926 = (inp[15]) ? 4'b1110 : 4'b1001;
															assign node7929 = (inp[5]) ? 4'b1001 : 4'b1101;
														assign node7932 = (inp[4]) ? 4'b1100 : node7933;
															assign node7933 = (inp[15]) ? node7935 : 4'b1000;
																assign node7935 = (inp[5]) ? 4'b1111 : 4'b1110;
										assign node7939 = (inp[13]) ? node8009 : node7940;
											assign node7940 = (inp[4]) ? node7972 : node7941;
												assign node7941 = (inp[15]) ? node7961 : node7942;
													assign node7942 = (inp[5]) ? node7948 : node7943;
														assign node7943 = (inp[1]) ? node7945 : 4'b1111;
															assign node7945 = (inp[7]) ? 4'b1111 : 4'b1101;
														assign node7948 = (inp[1]) ? node7956 : node7949;
															assign node7949 = (inp[12]) ? node7953 : node7950;
																assign node7950 = (inp[7]) ? 4'b1010 : 4'b1001;
																assign node7953 = (inp[7]) ? 4'b1101 : 4'b1111;
															assign node7956 = (inp[12]) ? node7958 : 4'b1110;
																assign node7958 = (inp[7]) ? 4'b1000 : 4'b1110;
													assign node7961 = (inp[7]) ? node7969 : node7962;
														assign node7962 = (inp[12]) ? node7966 : node7963;
															assign node7963 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node7966 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node7969 = (inp[12]) ? 4'b1111 : 4'b1001;
												assign node7972 = (inp[12]) ? node7990 : node7973;
													assign node7973 = (inp[7]) ? node7983 : node7974;
														assign node7974 = (inp[15]) ? node7978 : node7975;
															assign node7975 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node7978 = (inp[5]) ? 4'b1000 : node7979;
																assign node7979 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node7983 = (inp[1]) ? node7987 : node7984;
															assign node7984 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node7987 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node7990 = (inp[7]) ? node8002 : node7991;
														assign node7991 = (inp[5]) ? node7997 : node7992;
															assign node7992 = (inp[15]) ? node7994 : 4'b1111;
																assign node7994 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node7997 = (inp[15]) ? 4'b1111 : node7998;
																assign node7998 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node8002 = (inp[1]) ? node8006 : node8003;
															assign node8003 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node8006 = (inp[15]) ? 4'b1101 : 4'b1100;
											assign node8009 = (inp[1]) ? node8051 : node8010;
												assign node8010 = (inp[5]) ? node8030 : node8011;
													assign node8011 = (inp[4]) ? node8019 : node8012;
														assign node8012 = (inp[15]) ? 4'b1100 : node8013;
															assign node8013 = (inp[7]) ? 4'b1100 : node8014;
																assign node8014 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node8019 = (inp[7]) ? node8027 : node8020;
															assign node8020 = (inp[12]) ? node8024 : node8021;
																assign node8021 = (inp[15]) ? 4'b1101 : 4'b1000;
																assign node8024 = (inp[15]) ? 4'b1010 : 4'b1110;
															assign node8027 = (inp[12]) ? 4'b1001 : 4'b1010;
													assign node8030 = (inp[7]) ? node8040 : node8031;
														assign node8031 = (inp[12]) ? node8033 : 4'b1101;
															assign node8033 = (inp[15]) ? node8037 : node8034;
																assign node8034 = (inp[4]) ? 4'b1111 : 4'b1010;
																assign node8037 = (inp[4]) ? 4'b1011 : 4'b1001;
														assign node8040 = (inp[4]) ? node8044 : node8041;
															assign node8041 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node8044 = (inp[12]) ? node8048 : node8045;
																assign node8045 = (inp[15]) ? 4'b1111 : 4'b1110;
																assign node8048 = (inp[15]) ? 4'b1100 : 4'b1101;
												assign node8051 = (inp[4]) ? node8071 : node8052;
													assign node8052 = (inp[5]) ? node8062 : node8053;
														assign node8053 = (inp[12]) ? 4'b1011 : node8054;
															assign node8054 = (inp[15]) ? node8058 : node8055;
																assign node8055 = (inp[7]) ? 4'b1011 : 4'b1001;
																assign node8058 = (inp[7]) ? 4'b1001 : 4'b1011;
														assign node8062 = (inp[7]) ? node8068 : node8063;
															assign node8063 = (inp[15]) ? 4'b1011 : node8064;
																assign node8064 = (inp[12]) ? 4'b1011 : 4'b1000;
															assign node8068 = (inp[15]) ? 4'b1010 : 4'b1100;
													assign node8071 = (inp[7]) ? node8085 : node8072;
														assign node8072 = (inp[12]) ? node8080 : node8073;
															assign node8073 = (inp[15]) ? node8077 : node8074;
																assign node8074 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node8077 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node8080 = (inp[5]) ? node8082 : 4'b1010;
																assign node8082 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node8085 = (inp[12]) ? 4'b1000 : 4'b1010;
									assign node8088 = (inp[13]) ? node8240 : node8089;
										assign node8089 = (inp[2]) ? node8163 : node8090;
											assign node8090 = (inp[15]) ? node8128 : node8091;
												assign node8091 = (inp[1]) ? node8111 : node8092;
													assign node8092 = (inp[5]) ? node8104 : node8093;
														assign node8093 = (inp[12]) ? node8097 : node8094;
															assign node8094 = (inp[7]) ? 4'b1011 : 4'b1001;
															assign node8097 = (inp[7]) ? node8101 : node8098;
																assign node8098 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node8101 = (inp[4]) ? 4'b1000 : 4'b1101;
														assign node8104 = (inp[12]) ? node8106 : 4'b1101;
															assign node8106 = (inp[7]) ? node8108 : 4'b1011;
																assign node8108 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node8111 = (inp[12]) ? node8119 : node8112;
														assign node8112 = (inp[7]) ? 4'b1011 : node8113;
															assign node8113 = (inp[4]) ? node8115 : 4'b1001;
																assign node8115 = (inp[5]) ? 4'b1000 : 4'b1001;
														assign node8119 = (inp[7]) ? node8125 : node8120;
															assign node8120 = (inp[5]) ? node8122 : 4'b1010;
																assign node8122 = (inp[4]) ? 4'b1111 : 4'b1010;
															assign node8125 = (inp[4]) ? 4'b1001 : 4'b1100;
												assign node8128 = (inp[12]) ? node8148 : node8129;
													assign node8129 = (inp[5]) ? node8139 : node8130;
														assign node8130 = (inp[4]) ? node8136 : node8131;
															assign node8131 = (inp[7]) ? node8133 : 4'b1011;
																assign node8133 = (inp[1]) ? 4'b1000 : 4'b1101;
															assign node8136 = (inp[7]) ? 4'b1011 : 4'b1101;
														assign node8139 = (inp[4]) ? node8143 : node8140;
															assign node8140 = (inp[7]) ? 4'b1101 : 4'b1111;
															assign node8143 = (inp[7]) ? 4'b1010 : node8144;
																assign node8144 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node8148 = (inp[1]) ? node8158 : node8149;
														assign node8149 = (inp[7]) ? node8155 : node8150;
															assign node8150 = (inp[4]) ? node8152 : 4'b1001;
																assign node8152 = (inp[5]) ? 4'b1010 : 4'b1011;
															assign node8155 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node8158 = (inp[4]) ? node8160 : 4'b1100;
															assign node8160 = (inp[7]) ? 4'b1000 : 4'b1010;
											assign node8163 = (inp[5]) ? node8195 : node8164;
												assign node8164 = (inp[12]) ? node8182 : node8165;
													assign node8165 = (inp[7]) ? node8173 : node8166;
														assign node8166 = (inp[15]) ? node8170 : node8167;
															assign node8167 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node8170 = (inp[4]) ? 4'b1001 : 4'b1111;
														assign node8173 = (inp[1]) ? node8175 : 4'b1111;
															assign node8175 = (inp[4]) ? node8179 : node8176;
																assign node8176 = (inp[15]) ? 4'b1100 : 4'b1111;
																assign node8179 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node8182 = (inp[4]) ? node8186 : node8183;
														assign node8183 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node8186 = (inp[7]) ? node8190 : node8187;
															assign node8187 = (inp[15]) ? 4'b1111 : 4'b1011;
															assign node8190 = (inp[15]) ? 4'b1100 : node8191;
																assign node8191 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node8195 = (inp[1]) ? node8219 : node8196;
													assign node8196 = (inp[12]) ? node8208 : node8197;
														assign node8197 = (inp[7]) ? node8203 : node8198;
															assign node8198 = (inp[15]) ? 4'b1101 : node8199;
																assign node8199 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node8203 = (inp[4]) ? node8205 : 4'b1001;
																assign node8205 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node8208 = (inp[7]) ? node8214 : node8209;
															assign node8209 = (inp[15]) ? 4'b1110 : node8210;
																assign node8210 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node8214 = (inp[15]) ? node8216 : 4'b1101;
																assign node8216 = (inp[4]) ? 4'b1000 : 4'b1010;
													assign node8219 = (inp[4]) ? node8227 : node8220;
														assign node8220 = (inp[15]) ? 4'b1000 : node8221;
															assign node8221 = (inp[7]) ? node8223 : 4'b1100;
																assign node8223 = (inp[12]) ? 4'b1001 : 4'b1111;
														assign node8227 = (inp[15]) ? node8233 : node8228;
															assign node8228 = (inp[7]) ? node8230 : 4'b1101;
																assign node8230 = (inp[12]) ? 4'b1100 : 4'b1110;
															assign node8233 = (inp[7]) ? node8237 : node8234;
																assign node8234 = (inp[12]) ? 4'b1111 : 4'b1000;
																assign node8237 = (inp[12]) ? 4'b1101 : 4'b1111;
										assign node8240 = (inp[2]) ? node8330 : node8241;
											assign node8241 = (inp[15]) ? node8285 : node8242;
												assign node8242 = (inp[5]) ? node8262 : node8243;
													assign node8243 = (inp[12]) ? node8247 : node8244;
														assign node8244 = (inp[7]) ? 4'b1111 : 4'b1101;
														assign node8247 = (inp[7]) ? node8255 : node8248;
															assign node8248 = (inp[1]) ? node8252 : node8249;
																assign node8249 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node8252 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node8255 = (inp[4]) ? node8259 : node8256;
																assign node8256 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node8259 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node8262 = (inp[1]) ? node8276 : node8263;
														assign node8263 = (inp[4]) ? node8269 : node8264;
															assign node8264 = (inp[12]) ? node8266 : 4'b1010;
																assign node8266 = (inp[7]) ? 4'b1101 : 4'b1111;
															assign node8269 = (inp[7]) ? node8273 : node8270;
																assign node8270 = (inp[12]) ? 4'b1010 : 4'b1000;
																assign node8273 = (inp[12]) ? 4'b1000 : 4'b1011;
														assign node8276 = (inp[4]) ? node8278 : 4'b1110;
															assign node8278 = (inp[7]) ? node8282 : node8279;
																assign node8279 = (inp[12]) ? 4'b1011 : 4'b1100;
																assign node8282 = (inp[12]) ? 4'b1101 : 4'b1111;
												assign node8285 = (inp[4]) ? node8309 : node8286;
													assign node8286 = (inp[5]) ? node8298 : node8287;
														assign node8287 = (inp[7]) ? node8291 : node8288;
															assign node8288 = (inp[12]) ? 4'b1000 : 4'b1110;
															assign node8291 = (inp[12]) ? node8295 : node8292;
																assign node8292 = (inp[1]) ? 4'b1101 : 4'b1000;
																assign node8295 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node8298 = (inp[1]) ? node8302 : node8299;
															assign node8299 = (inp[7]) ? 4'b1000 : 4'b1100;
															assign node8302 = (inp[12]) ? node8306 : node8303;
																assign node8303 = (inp[7]) ? 4'b1000 : 4'b1111;
																assign node8306 = (inp[7]) ? 4'b1110 : 4'b1000;
													assign node8309 = (inp[5]) ? node8323 : node8310;
														assign node8310 = (inp[7]) ? node8318 : node8311;
															assign node8311 = (inp[12]) ? node8315 : node8312;
																assign node8312 = (inp[1]) ? 4'b1001 : 4'b1000;
																assign node8315 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node8318 = (inp[12]) ? 4'b1101 : node8319;
																assign node8319 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node8323 = (inp[7]) ? node8327 : node8324;
															assign node8324 = (inp[12]) ? 4'b1111 : 4'b1101;
															assign node8327 = (inp[12]) ? 4'b1001 : 4'b1010;
											assign node8330 = (inp[1]) ? node8374 : node8331;
												assign node8331 = (inp[12]) ? node8359 : node8332;
													assign node8332 = (inp[5]) ? node8346 : node8333;
														assign node8333 = (inp[15]) ? node8339 : node8334;
															assign node8334 = (inp[4]) ? node8336 : 4'b1000;
																assign node8336 = (inp[7]) ? 4'b1011 : 4'b1001;
															assign node8339 = (inp[4]) ? node8343 : node8340;
																assign node8340 = (inp[7]) ? 4'b1101 : 4'b1011;
																assign node8343 = (inp[7]) ? 4'b1010 : 4'b1100;
														assign node8346 = (inp[7]) ? node8354 : node8347;
															assign node8347 = (inp[4]) ? node8351 : node8348;
																assign node8348 = (inp[15]) ? 4'b1111 : 4'b1100;
																assign node8351 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node8354 = (inp[15]) ? 4'b1100 : node8355;
																assign node8355 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node8359 = (inp[4]) ? node8369 : node8360;
														assign node8360 = (inp[15]) ? node8366 : node8361;
															assign node8361 = (inp[7]) ? node8363 : 4'b1010;
																assign node8363 = (inp[5]) ? 4'b1000 : 4'b1100;
															assign node8366 = (inp[7]) ? 4'b1111 : 4'b1101;
														assign node8369 = (inp[15]) ? node8371 : 4'b1111;
															assign node8371 = (inp[5]) ? 4'b1011 : 4'b1010;
												assign node8374 = (inp[7]) ? node8398 : node8375;
													assign node8375 = (inp[12]) ? node8387 : node8376;
														assign node8376 = (inp[15]) ? node8382 : node8377;
															assign node8377 = (inp[5]) ? 4'b1000 : node8378;
																assign node8378 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node8382 = (inp[4]) ? 4'b1101 : node8383;
																assign node8383 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node8387 = (inp[5]) ? node8393 : node8388;
															assign node8388 = (inp[4]) ? 4'b1010 : node8389;
																assign node8389 = (inp[15]) ? 4'b1100 : 4'b1111;
															assign node8393 = (inp[4]) ? node8395 : 4'b1011;
																assign node8395 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node8398 = (inp[12]) ? node8406 : node8399;
														assign node8399 = (inp[4]) ? 4'b1011 : node8400;
															assign node8400 = (inp[15]) ? 4'b1101 : node8401;
																assign node8401 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node8406 = (inp[15]) ? 4'b1011 : node8407;
															assign node8407 = (inp[4]) ? 4'b1001 : 4'b1101;
							assign node8411 = (inp[11]) ? node8979 : node8412;
								assign node8412 = (inp[4]) ? node8718 : node8413;
									assign node8413 = (inp[15]) ? node8553 : node8414;
										assign node8414 = (inp[2]) ? node8480 : node8415;
											assign node8415 = (inp[12]) ? node8439 : node8416;
												assign node8416 = (inp[7]) ? node8432 : node8417;
													assign node8417 = (inp[13]) ? node8423 : node8418;
														assign node8418 = (inp[5]) ? node8420 : 4'b1000;
															assign node8420 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node8423 = (inp[5]) ? node8425 : 4'b1100;
															assign node8425 = (inp[1]) ? node8429 : node8426;
																assign node8426 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node8429 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node8432 = (inp[13]) ? node8434 : 4'b1010;
														assign node8434 = (inp[5]) ? node8436 : 4'b1110;
															assign node8436 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node8439 = (inp[7]) ? node8461 : node8440;
													assign node8440 = (inp[13]) ? node8450 : node8441;
														assign node8441 = (inp[1]) ? node8445 : node8442;
															assign node8442 = (inp[5]) ? 4'b1011 : 4'b1010;
															assign node8445 = (inp[5]) ? node8447 : 4'b1111;
																assign node8447 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node8450 = (inp[5]) ? node8456 : node8451;
															assign node8451 = (inp[1]) ? node8453 : 4'b1110;
																assign node8453 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node8456 = (inp[1]) ? node8458 : 4'b1110;
																assign node8458 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node8461 = (inp[13]) ? node8471 : node8462;
														assign node8462 = (inp[5]) ? 4'b1101 : node8463;
															assign node8463 = (inp[1]) ? node8467 : node8464;
																assign node8464 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node8467 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node8471 = (inp[1]) ? node8475 : node8472;
															assign node8472 = (inp[5]) ? 4'b1100 : 4'b1001;
															assign node8475 = (inp[5]) ? node8477 : 4'b1000;
																assign node8477 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node8480 = (inp[13]) ? node8518 : node8481;
												assign node8481 = (inp[7]) ? node8497 : node8482;
													assign node8482 = (inp[12]) ? node8488 : node8483;
														assign node8483 = (inp[0]) ? 4'b1101 : node8484;
															assign node8484 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node8488 = (inp[1]) ? node8494 : node8489;
															assign node8489 = (inp[5]) ? 4'b1111 : node8490;
																assign node8490 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node8494 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node8497 = (inp[12]) ? node8505 : node8498;
														assign node8498 = (inp[5]) ? node8502 : node8499;
															assign node8499 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node8502 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node8505 = (inp[5]) ? node8513 : node8506;
															assign node8506 = (inp[0]) ? node8510 : node8507;
																assign node8507 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node8510 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node8513 = (inp[1]) ? 4'b1000 : node8514;
																assign node8514 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node8518 = (inp[7]) ? node8536 : node8519;
													assign node8519 = (inp[12]) ? node8525 : node8520;
														assign node8520 = (inp[5]) ? node8522 : 4'b1001;
															assign node8522 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node8525 = (inp[1]) ? node8531 : node8526;
															assign node8526 = (inp[5]) ? node8528 : 4'b1011;
																assign node8528 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node8531 = (inp[5]) ? node8533 : 4'b1110;
																assign node8533 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node8536 = (inp[12]) ? node8544 : node8537;
														assign node8537 = (inp[5]) ? node8539 : 4'b1011;
															assign node8539 = (inp[1]) ? node8541 : 4'b1110;
																assign node8541 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node8544 = (inp[1]) ? node8548 : node8545;
															assign node8545 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node8548 = (inp[5]) ? 4'b1100 : node8549;
																assign node8549 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node8553 = (inp[0]) ? node8653 : node8554;
											assign node8554 = (inp[1]) ? node8606 : node8555;
												assign node8555 = (inp[12]) ? node8579 : node8556;
													assign node8556 = (inp[7]) ? node8566 : node8557;
														assign node8557 = (inp[13]) ? node8563 : node8558;
															assign node8558 = (inp[5]) ? node8560 : 4'b1110;
																assign node8560 = (inp[2]) ? 4'b1011 : 4'b1110;
															assign node8563 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node8566 = (inp[5]) ? node8572 : node8567;
															assign node8567 = (inp[13]) ? 4'b1100 : node8568;
																assign node8568 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node8572 = (inp[13]) ? node8576 : node8573;
																assign node8573 = (inp[2]) ? 4'b1000 : 4'b1101;
																assign node8576 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node8579 = (inp[7]) ? node8595 : node8580;
														assign node8580 = (inp[13]) ? node8588 : node8581;
															assign node8581 = (inp[2]) ? node8585 : node8582;
																assign node8582 = (inp[5]) ? 4'b1000 : 4'b1100;
																assign node8585 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node8588 = (inp[2]) ? node8592 : node8589;
																assign node8589 = (inp[5]) ? 4'b1101 : 4'b1001;
																assign node8592 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node8595 = (inp[5]) ? node8601 : node8596;
															assign node8596 = (inp[2]) ? 4'b1011 : node8597;
																assign node8597 = (inp[13]) ? 4'b1110 : 4'b1011;
															assign node8601 = (inp[13]) ? node8603 : 4'b1110;
																assign node8603 = (inp[2]) ? 4'b1110 : 4'b1011;
												assign node8606 = (inp[12]) ? node8628 : node8607;
													assign node8607 = (inp[7]) ? node8621 : node8608;
														assign node8608 = (inp[2]) ? node8616 : node8609;
															assign node8609 = (inp[13]) ? node8613 : node8610;
																assign node8610 = (inp[5]) ? 4'b1011 : 4'b1010;
																assign node8613 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node8616 = (inp[13]) ? node8618 : 4'b1111;
																assign node8618 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node8621 = (inp[5]) ? node8625 : node8622;
															assign node8622 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node8625 = (inp[2]) ? 4'b1001 : 4'b1100;
													assign node8628 = (inp[7]) ? node8642 : node8629;
														assign node8629 = (inp[2]) ? node8635 : node8630;
															assign node8630 = (inp[13]) ? 4'b1001 : node8631;
																assign node8631 = (inp[5]) ? 4'b1100 : 4'b1101;
															assign node8635 = (inp[13]) ? node8639 : node8636;
																assign node8636 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node8639 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node8642 = (inp[5]) ? node8650 : node8643;
															assign node8643 = (inp[2]) ? node8647 : node8644;
																assign node8644 = (inp[13]) ? 4'b1111 : 4'b1010;
																assign node8647 = (inp[13]) ? 4'b1010 : 4'b1111;
															assign node8650 = (inp[13]) ? 4'b1111 : 4'b1110;
											assign node8653 = (inp[13]) ? node8685 : node8654;
												assign node8654 = (inp[2]) ? node8668 : node8655;
													assign node8655 = (inp[1]) ? node8663 : node8656;
														assign node8656 = (inp[5]) ? 4'b1110 : node8657;
															assign node8657 = (inp[12]) ? 4'b1011 : node8658;
																assign node8658 = (inp[7]) ? 4'b1100 : 4'b1010;
														assign node8663 = (inp[7]) ? node8665 : 4'b1011;
															assign node8665 = (inp[5]) ? 4'b1010 : 4'b1011;
													assign node8668 = (inp[1]) ? node8678 : node8669;
														assign node8669 = (inp[7]) ? node8675 : node8670;
															assign node8670 = (inp[12]) ? 4'b1101 : node8671;
																assign node8671 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node8675 = (inp[12]) ? 4'b1011 : 4'b1001;
														assign node8678 = (inp[12]) ? node8682 : node8679;
															assign node8679 = (inp[7]) ? 4'b1100 : 4'b1111;
															assign node8682 = (inp[7]) ? 4'b1111 : 4'b1001;
												assign node8685 = (inp[5]) ? node8699 : node8686;
													assign node8686 = (inp[7]) ? node8694 : node8687;
														assign node8687 = (inp[12]) ? 4'b1100 : node8688;
															assign node8688 = (inp[2]) ? node8690 : 4'b1111;
																assign node8690 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node8694 = (inp[12]) ? 4'b1011 : node8695;
															assign node8695 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node8699 = (inp[2]) ? node8707 : node8700;
														assign node8700 = (inp[12]) ? 4'b1100 : node8701;
															assign node8701 = (inp[7]) ? node8703 : 4'b1010;
																assign node8703 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node8707 = (inp[7]) ? node8713 : node8708;
															assign node8708 = (inp[12]) ? 4'b1001 : node8709;
																assign node8709 = (inp[1]) ? 4'b1011 : 4'b1110;
															assign node8713 = (inp[12]) ? node8715 : 4'b1100;
																assign node8715 = (inp[1]) ? 4'b1010 : 4'b1110;
									assign node8718 = (inp[13]) ? node8860 : node8719;
										assign node8719 = (inp[2]) ? node8787 : node8720;
											assign node8720 = (inp[5]) ? node8754 : node8721;
												assign node8721 = (inp[7]) ? node8739 : node8722;
													assign node8722 = (inp[12]) ? node8728 : node8723;
														assign node8723 = (inp[15]) ? node8725 : 4'b1000;
															assign node8725 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node8728 = (inp[15]) ? node8734 : node8729;
															assign node8729 = (inp[1]) ? node8731 : 4'b1110;
																assign node8731 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node8734 = (inp[1]) ? 4'b1110 : node8735;
																assign node8735 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node8739 = (inp[12]) ? node8747 : node8740;
														assign node8740 = (inp[15]) ? node8742 : 4'b1010;
															assign node8742 = (inp[1]) ? 4'b1011 : node8743;
																assign node8743 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node8747 = (inp[1]) ? node8751 : node8748;
															assign node8748 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node8751 = (inp[15]) ? 4'b1001 : 4'b1000;
												assign node8754 = (inp[1]) ? node8770 : node8755;
													assign node8755 = (inp[7]) ? node8765 : node8756;
														assign node8756 = (inp[15]) ? node8760 : node8757;
															assign node8757 = (inp[12]) ? 4'b1111 : 4'b1100;
															assign node8760 = (inp[12]) ? node8762 : 4'b1001;
																assign node8762 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node8765 = (inp[12]) ? node8767 : 4'b1110;
															assign node8767 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node8770 = (inp[7]) ? node8780 : node8771;
														assign node8771 = (inp[12]) ? node8777 : node8772;
															assign node8772 = (inp[15]) ? node8774 : 4'b1001;
																assign node8774 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8777 = (inp[15]) ? 4'b1011 : 4'b1110;
														assign node8780 = (inp[15]) ? node8784 : node8781;
															assign node8781 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node8784 = (inp[12]) ? 4'b1001 : 4'b1011;
											assign node8787 = (inp[7]) ? node8829 : node8788;
												assign node8788 = (inp[12]) ? node8816 : node8789;
													assign node8789 = (inp[15]) ? node8803 : node8790;
														assign node8790 = (inp[1]) ? node8796 : node8791;
															assign node8791 = (inp[5]) ? 4'b1000 : node8792;
																assign node8792 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node8796 = (inp[0]) ? node8800 : node8797;
																assign node8797 = (inp[5]) ? 4'b1100 : 4'b1101;
																assign node8800 = (inp[5]) ? 4'b1101 : 4'b1100;
														assign node8803 = (inp[1]) ? node8809 : node8804;
															assign node8804 = (inp[5]) ? node8806 : 4'b1000;
																assign node8806 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node8809 = (inp[0]) ? node8813 : node8810;
																assign node8810 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node8813 = (inp[5]) ? 4'b1000 : 4'b1001;
													assign node8816 = (inp[15]) ? node8824 : node8817;
														assign node8817 = (inp[5]) ? node8821 : node8818;
															assign node8818 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node8821 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node8824 = (inp[5]) ? 4'b1111 : node8825;
															assign node8825 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node8829 = (inp[12]) ? node8849 : node8830;
													assign node8830 = (inp[1]) ? node8842 : node8831;
														assign node8831 = (inp[5]) ? node8837 : node8832;
															assign node8832 = (inp[0]) ? 4'b1110 : node8833;
																assign node8833 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node8837 = (inp[0]) ? 4'b1010 : node8838;
																assign node8838 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node8842 = (inp[0]) ? node8846 : node8843;
															assign node8843 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node8846 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node8849 = (inp[15]) ? node8851 : 4'b1100;
														assign node8851 = (inp[0]) ? node8855 : node8852;
															assign node8852 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node8855 = (inp[1]) ? 4'b1101 : node8856;
																assign node8856 = (inp[5]) ? 4'b1001 : 4'b1101;
										assign node8860 = (inp[2]) ? node8924 : node8861;
											assign node8861 = (inp[1]) ? node8901 : node8862;
												assign node8862 = (inp[12]) ? node8884 : node8863;
													assign node8863 = (inp[7]) ? node8875 : node8864;
														assign node8864 = (inp[0]) ? node8872 : node8865;
															assign node8865 = (inp[15]) ? node8869 : node8866;
																assign node8866 = (inp[5]) ? 4'b1001 : 4'b1100;
																assign node8869 = (inp[5]) ? 4'b1100 : 4'b1001;
															assign node8872 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node8875 = (inp[5]) ? node8881 : node8876;
															assign node8876 = (inp[15]) ? node8878 : 4'b1110;
																assign node8878 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node8881 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node8884 = (inp[7]) ? node8898 : node8885;
														assign node8885 = (inp[15]) ? node8891 : node8886;
															assign node8886 = (inp[0]) ? node8888 : 4'b1010;
																assign node8888 = (inp[5]) ? 4'b1010 : 4'b1011;
															assign node8891 = (inp[5]) ? node8895 : node8892;
																assign node8892 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node8895 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node8898 = (inp[5]) ? 4'b1001 : 4'b1101;
												assign node8901 = (inp[7]) ? node8921 : node8902;
													assign node8902 = (inp[12]) ? node8910 : node8903;
														assign node8903 = (inp[5]) ? node8907 : node8904;
															assign node8904 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node8907 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node8910 = (inp[15]) ? node8918 : node8911;
															assign node8911 = (inp[5]) ? node8915 : node8912;
																assign node8912 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node8915 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node8918 = (inp[5]) ? 4'b1110 : 4'b1010;
													assign node8921 = (inp[12]) ? 4'b1100 : 4'b1110;
											assign node8924 = (inp[1]) ? node8964 : node8925;
												assign node8925 = (inp[5]) ? node8945 : node8926;
													assign node8926 = (inp[0]) ? node8936 : node8927;
														assign node8927 = (inp[15]) ? node8929 : 4'b1000;
															assign node8929 = (inp[7]) ? node8933 : node8930;
																assign node8930 = (inp[12]) ? 4'b1011 : 4'b1101;
																assign node8933 = (inp[12]) ? 4'b1000 : 4'b1011;
														assign node8936 = (inp[15]) ? 4'b1010 : node8937;
															assign node8937 = (inp[12]) ? node8941 : node8938;
																assign node8938 = (inp[7]) ? 4'b1010 : 4'b1000;
																assign node8941 = (inp[7]) ? 4'b1001 : 4'b1110;
													assign node8945 = (inp[7]) ? node8955 : node8946;
														assign node8946 = (inp[15]) ? node8950 : node8947;
															assign node8947 = (inp[12]) ? 4'b1111 : 4'b1101;
															assign node8950 = (inp[12]) ? node8952 : 4'b1000;
																assign node8952 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node8955 = (inp[12]) ? node8961 : node8956;
															assign node8956 = (inp[0]) ? node8958 : 4'b1111;
																assign node8958 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node8961 = (inp[15]) ? 4'b1100 : 4'b1101;
												assign node8964 = (inp[7]) ? node8976 : node8965;
													assign node8965 = (inp[12]) ? node8971 : node8966;
														assign node8966 = (inp[15]) ? 4'b1100 : node8967;
															assign node8967 = (inp[5]) ? 4'b1001 : 4'b1000;
														assign node8971 = (inp[5]) ? node8973 : 4'b1111;
															assign node8973 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node8976 = (inp[12]) ? 4'b1000 : 4'b1010;
								assign node8979 = (inp[0]) ? node9289 : node8980;
									assign node8980 = (inp[2]) ? node9140 : node8981;
										assign node8981 = (inp[13]) ? node9071 : node8982;
											assign node8982 = (inp[15]) ? node9020 : node8983;
												assign node8983 = (inp[1]) ? node9003 : node8984;
													assign node8984 = (inp[12]) ? node8994 : node8985;
														assign node8985 = (inp[5]) ? node8989 : node8986;
															assign node8986 = (inp[7]) ? 4'b1011 : 4'b1001;
															assign node8989 = (inp[7]) ? 4'b1111 : node8990;
																assign node8990 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node8994 = (inp[7]) ? node9000 : node8995;
															assign node8995 = (inp[5]) ? node8997 : 4'b1111;
																assign node8997 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node9000 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node9003 = (inp[12]) ? node9009 : node9004;
														assign node9004 = (inp[7]) ? 4'b1011 : node9005;
															assign node9005 = (inp[5]) ? 4'b1000 : 4'b1001;
														assign node9009 = (inp[7]) ? node9015 : node9010;
															assign node9010 = (inp[5]) ? node9012 : 4'b1011;
																assign node9012 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node9015 = (inp[5]) ? 4'b1100 : node9016;
																assign node9016 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node9020 = (inp[7]) ? node9046 : node9021;
													assign node9021 = (inp[5]) ? node9033 : node9022;
														assign node9022 = (inp[12]) ? node9028 : node9023;
															assign node9023 = (inp[4]) ? node9025 : 4'b1010;
																assign node9025 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node9028 = (inp[4]) ? node9030 : 4'b1101;
																assign node9030 = (inp[1]) ? 4'b1111 : 4'b1010;
														assign node9033 = (inp[1]) ? node9039 : node9034;
															assign node9034 = (inp[4]) ? 4'b1000 : node9035;
																assign node9035 = (inp[12]) ? 4'b1000 : 4'b1111;
															assign node9039 = (inp[12]) ? node9043 : node9040;
																assign node9040 = (inp[4]) ? 4'b1101 : 4'b1010;
																assign node9043 = (inp[4]) ? 4'b1010 : 4'b1101;
													assign node9046 = (inp[1]) ? node9060 : node9047;
														assign node9047 = (inp[5]) ? node9055 : node9048;
															assign node9048 = (inp[4]) ? node9052 : node9049;
																assign node9049 = (inp[12]) ? 4'b1010 : 4'b1101;
																assign node9052 = (inp[12]) ? 4'b1001 : 4'b1010;
															assign node9055 = (inp[4]) ? node9057 : 4'b1111;
																assign node9057 = (inp[12]) ? 4'b1100 : 4'b1111;
														assign node9060 = (inp[5]) ? node9066 : node9061;
															assign node9061 = (inp[12]) ? node9063 : 4'b1000;
																assign node9063 = (inp[4]) ? 4'b1000 : 4'b1010;
															assign node9066 = (inp[4]) ? node9068 : 4'b1101;
																assign node9068 = (inp[12]) ? 4'b1000 : 4'b1010;
											assign node9071 = (inp[1]) ? node9115 : node9072;
												assign node9072 = (inp[5]) ? node9094 : node9073;
													assign node9073 = (inp[4]) ? node9087 : node9074;
														assign node9074 = (inp[12]) ? node9080 : node9075;
															assign node9075 = (inp[7]) ? node9077 : 4'b1110;
																assign node9077 = (inp[15]) ? 4'b1001 : 4'b1111;
															assign node9080 = (inp[15]) ? node9084 : node9081;
																assign node9081 = (inp[7]) ? 4'b1000 : 4'b1111;
																assign node9084 = (inp[7]) ? 4'b1111 : 4'b1001;
														assign node9087 = (inp[12]) ? 4'b1100 : node9088;
															assign node9088 = (inp[7]) ? 4'b1111 : node9089;
																assign node9089 = (inp[15]) ? 4'b1001 : 4'b1101;
													assign node9094 = (inp[7]) ? node9106 : node9095;
														assign node9095 = (inp[15]) ? node9101 : node9096;
															assign node9096 = (inp[4]) ? 4'b1011 : node9097;
																assign node9097 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node9101 = (inp[4]) ? node9103 : 4'b1101;
																assign node9103 = (inp[12]) ? 4'b1110 : 4'b1101;
														assign node9106 = (inp[12]) ? node9110 : node9107;
															assign node9107 = (inp[4]) ? 4'b1011 : 4'b1000;
															assign node9110 = (inp[15]) ? 4'b1011 : node9111;
																assign node9111 = (inp[4]) ? 4'b1000 : 4'b1101;
												assign node9115 = (inp[7]) ? node9131 : node9116;
													assign node9116 = (inp[12]) ? node9122 : node9117;
														assign node9117 = (inp[15]) ? 4'b1111 : node9118;
															assign node9118 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node9122 = (inp[15]) ? node9128 : node9123;
															assign node9123 = (inp[5]) ? 4'b1111 : node9124;
																assign node9124 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node9128 = (inp[4]) ? 4'b1011 : 4'b1000;
													assign node9131 = (inp[12]) ? 4'b1101 : node9132;
														assign node9132 = (inp[4]) ? 4'b1111 : node9133;
															assign node9133 = (inp[15]) ? node9135 : 4'b1111;
																assign node9135 = (inp[5]) ? 4'b1001 : 4'b1101;
										assign node9140 = (inp[4]) ? node9216 : node9141;
											assign node9141 = (inp[13]) ? node9177 : node9142;
												assign node9142 = (inp[5]) ? node9160 : node9143;
													assign node9143 = (inp[12]) ? node9151 : node9144;
														assign node9144 = (inp[7]) ? node9148 : node9145;
															assign node9145 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node9148 = (inp[15]) ? 4'b1101 : 4'b1110;
														assign node9151 = (inp[7]) ? node9155 : node9152;
															assign node9152 = (inp[15]) ? 4'b1000 : 4'b1011;
															assign node9155 = (inp[15]) ? node9157 : 4'b1000;
																assign node9157 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node9160 = (inp[15]) ? node9166 : node9161;
														assign node9161 = (inp[7]) ? 4'b1011 : node9162;
															assign node9162 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node9166 = (inp[7]) ? node9174 : node9167;
															assign node9167 = (inp[12]) ? node9171 : node9168;
																assign node9168 = (inp[1]) ? 4'b1111 : 4'b1010;
																assign node9171 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node9174 = (inp[12]) ? 4'b1010 : 4'b1000;
												assign node9177 = (inp[1]) ? node9201 : node9178;
													assign node9178 = (inp[15]) ? node9194 : node9179;
														assign node9179 = (inp[7]) ? node9187 : node9180;
															assign node9180 = (inp[12]) ? node9184 : node9181;
																assign node9181 = (inp[5]) ? 4'b1100 : 4'b1000;
																assign node9184 = (inp[5]) ? 4'b1011 : 4'b1010;
															assign node9187 = (inp[12]) ? node9191 : node9188;
																assign node9188 = (inp[5]) ? 4'b1111 : 4'b1010;
																assign node9191 = (inp[5]) ? 4'b1000 : 4'b1101;
														assign node9194 = (inp[12]) ? node9198 : node9195;
															assign node9195 = (inp[7]) ? 4'b1101 : 4'b1111;
															assign node9198 = (inp[7]) ? 4'b1010 : 4'b1101;
													assign node9201 = (inp[12]) ? node9203 : 4'b1010;
														assign node9203 = (inp[15]) ? node9211 : node9204;
															assign node9204 = (inp[7]) ? node9208 : node9205;
																assign node9205 = (inp[5]) ? 4'b1010 : 4'b1111;
																assign node9208 = (inp[5]) ? 4'b1101 : 4'b1100;
															assign node9211 = (inp[7]) ? node9213 : 4'b1101;
																assign node9213 = (inp[5]) ? 4'b1011 : 4'b1010;
											assign node9216 = (inp[13]) ? node9260 : node9217;
												assign node9217 = (inp[5]) ? node9239 : node9218;
													assign node9218 = (inp[7]) ? node9232 : node9219;
														assign node9219 = (inp[12]) ? node9225 : node9220;
															assign node9220 = (inp[15]) ? node9222 : 4'b1101;
																assign node9222 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node9225 = (inp[15]) ? node9229 : node9226;
																assign node9226 = (inp[1]) ? 4'b1110 : 4'b1011;
																assign node9229 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node9232 = (inp[12]) ? node9236 : node9233;
															assign node9233 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node9236 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node9239 = (inp[1]) ? node9249 : node9240;
														assign node9240 = (inp[15]) ? node9246 : node9241;
															assign node9241 = (inp[12]) ? node9243 : 4'b1011;
																assign node9243 = (inp[7]) ? 4'b1000 : 4'b1010;
															assign node9246 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node9249 = (inp[7]) ? node9255 : node9250;
															assign node9250 = (inp[12]) ? 4'b1011 : node9251;
																assign node9251 = (inp[15]) ? 4'b1001 : 4'b1100;
															assign node9255 = (inp[15]) ? node9257 : 4'b1101;
																assign node9257 = (inp[12]) ? 4'b1100 : 4'b1110;
												assign node9260 = (inp[1]) ? node9280 : node9261;
													assign node9261 = (inp[5]) ? node9267 : node9262;
														assign node9262 = (inp[7]) ? node9264 : 4'b1111;
															assign node9264 = (inp[12]) ? 4'b1000 : 4'b1011;
														assign node9267 = (inp[15]) ? node9275 : node9268;
															assign node9268 = (inp[12]) ? node9272 : node9269;
																assign node9269 = (inp[7]) ? 4'b1111 : 4'b1100;
																assign node9272 = (inp[7]) ? 4'b1100 : 4'b1110;
															assign node9275 = (inp[7]) ? 4'b1101 : node9276;
																assign node9276 = (inp[12]) ? 4'b1010 : 4'b1001;
													assign node9280 = (inp[12]) ? node9286 : node9281;
														assign node9281 = (inp[7]) ? 4'b1011 : node9282;
															assign node9282 = (inp[5]) ? 4'b1100 : 4'b1001;
														assign node9286 = (inp[7]) ? 4'b1001 : 4'b1011;
									assign node9289 = (inp[4]) ? node9467 : node9290;
										assign node9290 = (inp[15]) ? node9378 : node9291;
											assign node9291 = (inp[7]) ? node9337 : node9292;
												assign node9292 = (inp[12]) ? node9312 : node9293;
													assign node9293 = (inp[2]) ? node9301 : node9294;
														assign node9294 = (inp[1]) ? 4'b1100 : node9295;
															assign node9295 = (inp[13]) ? node9297 : 4'b1100;
																assign node9297 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node9301 = (inp[13]) ? node9307 : node9302;
															assign node9302 = (inp[5]) ? node9304 : 4'b1100;
																assign node9304 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node9307 = (inp[1]) ? 4'b1001 : node9308;
																assign node9308 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node9312 = (inp[2]) ? node9324 : node9313;
														assign node9313 = (inp[1]) ? node9317 : node9314;
															assign node9314 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node9317 = (inp[13]) ? node9321 : node9318;
																assign node9318 = (inp[5]) ? 4'b1011 : 4'b1111;
																assign node9321 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node9324 = (inp[1]) ? node9330 : node9325;
															assign node9325 = (inp[13]) ? 4'b1011 : node9326;
																assign node9326 = (inp[5]) ? 4'b1111 : 4'b1110;
															assign node9330 = (inp[13]) ? node9334 : node9331;
																assign node9331 = (inp[5]) ? 4'b1110 : 4'b1010;
																assign node9334 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node9337 = (inp[12]) ? node9355 : node9338;
													assign node9338 = (inp[13]) ? node9346 : node9339;
														assign node9339 = (inp[2]) ? node9343 : node9340;
															assign node9340 = (inp[5]) ? 4'b1011 : 4'b1010;
															assign node9343 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node9346 = (inp[2]) ? node9350 : node9347;
															assign node9347 = (inp[5]) ? 4'b1111 : 4'b1110;
															assign node9350 = (inp[5]) ? node9352 : 4'b1011;
																assign node9352 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node9355 = (inp[2]) ? node9369 : node9356;
														assign node9356 = (inp[1]) ? node9364 : node9357;
															assign node9357 = (inp[5]) ? node9361 : node9358;
																assign node9358 = (inp[13]) ? 4'b1001 : 4'b1100;
																assign node9361 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node9364 = (inp[5]) ? node9366 : 4'b1000;
																assign node9366 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node9369 = (inp[13]) ? 4'b1100 : node9370;
															assign node9370 = (inp[5]) ? node9374 : node9371;
																assign node9371 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node9374 = (inp[1]) ? 4'b1000 : 4'b1100;
											assign node9378 = (inp[1]) ? node9430 : node9379;
												assign node9379 = (inp[7]) ? node9403 : node9380;
													assign node9380 = (inp[12]) ? node9392 : node9381;
														assign node9381 = (inp[2]) ? node9387 : node9382;
															assign node9382 = (inp[13]) ? node9384 : 4'b1110;
																assign node9384 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node9387 = (inp[13]) ? node9389 : 4'b1110;
																assign node9389 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node9392 = (inp[13]) ? node9398 : node9393;
															assign node9393 = (inp[2]) ? node9395 : 4'b1000;
																assign node9395 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node9398 = (inp[2]) ? node9400 : 4'b1101;
																assign node9400 = (inp[5]) ? 4'b1000 : 4'b1100;
													assign node9403 = (inp[12]) ? node9419 : node9404;
														assign node9404 = (inp[5]) ? node9412 : node9405;
															assign node9405 = (inp[2]) ? node9409 : node9406;
																assign node9406 = (inp[13]) ? 4'b1001 : 4'b1100;
																assign node9409 = (inp[13]) ? 4'b1100 : 4'b1001;
															assign node9412 = (inp[2]) ? node9416 : node9413;
																assign node9413 = (inp[13]) ? 4'b1001 : 4'b1101;
																assign node9416 = (inp[13]) ? 4'b1101 : 4'b1000;
														assign node9419 = (inp[2]) ? node9425 : node9420;
															assign node9420 = (inp[13]) ? 4'b1110 : node9421;
																assign node9421 = (inp[5]) ? 4'b1110 : 4'b1011;
															assign node9425 = (inp[5]) ? node9427 : 4'b1011;
																assign node9427 = (inp[13]) ? 4'b1110 : 4'b1011;
												assign node9430 = (inp[5]) ? node9452 : node9431;
													assign node9431 = (inp[13]) ? node9441 : node9432;
														assign node9432 = (inp[2]) ? node9434 : 4'b1001;
															assign node9434 = (inp[7]) ? node9438 : node9435;
																assign node9435 = (inp[12]) ? 4'b1000 : 4'b1111;
																assign node9438 = (inp[12]) ? 4'b1111 : 4'b1101;
														assign node9441 = (inp[2]) ? node9447 : node9442;
															assign node9442 = (inp[7]) ? node9444 : 4'b1111;
																assign node9444 = (inp[12]) ? 4'b1111 : 4'b1100;
															assign node9447 = (inp[7]) ? 4'b1010 : node9448;
																assign node9448 = (inp[12]) ? 4'b1101 : 4'b1010;
													assign node9452 = (inp[7]) ? node9460 : node9453;
														assign node9453 = (inp[12]) ? 4'b1001 : node9454;
															assign node9454 = (inp[13]) ? 4'b1011 : node9455;
																assign node9455 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node9460 = (inp[12]) ? node9462 : 4'b1001;
															assign node9462 = (inp[13]) ? 4'b1111 : node9463;
																assign node9463 = (inp[2]) ? 4'b1110 : 4'b1010;
										assign node9467 = (inp[13]) ? node9547 : node9468;
											assign node9468 = (inp[2]) ? node9498 : node9469;
												assign node9469 = (inp[7]) ? node9487 : node9470;
													assign node9470 = (inp[12]) ? node9478 : node9471;
														assign node9471 = (inp[5]) ? node9475 : node9472;
															assign node9472 = (inp[15]) ? 4'b1100 : 4'b1000;
															assign node9475 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node9478 = (inp[15]) ? node9484 : node9479;
															assign node9479 = (inp[1]) ? node9481 : 4'b1110;
																assign node9481 = (inp[5]) ? 4'b1110 : 4'b1011;
															assign node9484 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node9487 = (inp[12]) ? node9493 : node9488;
														assign node9488 = (inp[1]) ? node9490 : 4'b1111;
															assign node9490 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node9493 = (inp[5]) ? node9495 : 4'b1001;
															assign node9495 = (inp[15]) ? 4'b1101 : 4'b1000;
												assign node9498 = (inp[15]) ? node9524 : node9499;
													assign node9499 = (inp[1]) ? node9513 : node9500;
														assign node9500 = (inp[5]) ? node9506 : node9501;
															assign node9501 = (inp[7]) ? node9503 : 4'b1010;
																assign node9503 = (inp[12]) ? 4'b1100 : 4'b1111;
															assign node9506 = (inp[12]) ? node9510 : node9507;
																assign node9507 = (inp[7]) ? 4'b1011 : 4'b1000;
																assign node9510 = (inp[7]) ? 4'b1000 : 4'b1011;
														assign node9513 = (inp[5]) ? node9521 : node9514;
															assign node9514 = (inp[12]) ? node9518 : node9515;
																assign node9515 = (inp[7]) ? 4'b1111 : 4'b1101;
																assign node9518 = (inp[7]) ? 4'b1101 : 4'b1111;
															assign node9521 = (inp[12]) ? 4'b1101 : 4'b1100;
													assign node9524 = (inp[5]) ? node9534 : node9525;
														assign node9525 = (inp[7]) ? node9531 : node9526;
															assign node9526 = (inp[12]) ? node9528 : 4'b1000;
																assign node9528 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node9531 = (inp[12]) ? 4'b1100 : 4'b1110;
														assign node9534 = (inp[7]) ? node9540 : node9535;
															assign node9535 = (inp[1]) ? 4'b1001 : node9536;
																assign node9536 = (inp[12]) ? 4'b1111 : 4'b1100;
															assign node9540 = (inp[12]) ? node9544 : node9541;
																assign node9541 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node9544 = (inp[1]) ? 4'b1100 : 4'b1001;
											assign node9547 = (inp[2]) ? node9583 : node9548;
												assign node9548 = (inp[7]) ? node9570 : node9549;
													assign node9549 = (inp[12]) ? node9561 : node9550;
														assign node9550 = (inp[5]) ? node9554 : node9551;
															assign node9551 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node9554 = (inp[15]) ? node9558 : node9555;
																assign node9555 = (inp[1]) ? 4'b1101 : 4'b1001;
																assign node9558 = (inp[1]) ? 4'b1001 : 4'b1100;
														assign node9561 = (inp[5]) ? node9567 : node9562;
															assign node9562 = (inp[1]) ? node9564 : 4'b1010;
																assign node9564 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node9567 = (inp[15]) ? 4'b1110 : 4'b1010;
													assign node9570 = (inp[12]) ? node9578 : node9571;
														assign node9571 = (inp[1]) ? 4'b1110 : node9572;
															assign node9572 = (inp[5]) ? 4'b1011 : node9573;
																assign node9573 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node9578 = (inp[1]) ? 4'b1100 : node9579;
															assign node9579 = (inp[15]) ? 4'b1000 : 4'b1101;
												assign node9583 = (inp[1]) ? node9607 : node9584;
													assign node9584 = (inp[5]) ? node9596 : node9585;
														assign node9585 = (inp[7]) ? node9589 : node9586;
															assign node9586 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node9589 = (inp[12]) ? node9593 : node9590;
																assign node9590 = (inp[15]) ? 4'b1011 : 4'b1010;
																assign node9593 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node9596 = (inp[7]) ? node9604 : node9597;
															assign node9597 = (inp[15]) ? node9601 : node9598;
																assign node9598 = (inp[12]) ? 4'b1111 : 4'b1100;
																assign node9601 = (inp[12]) ? 4'b1010 : 4'b1000;
															assign node9604 = (inp[12]) ? 4'b1100 : 4'b1111;
													assign node9607 = (inp[7]) ? node9621 : node9608;
														assign node9608 = (inp[12]) ? node9616 : node9609;
															assign node9609 = (inp[15]) ? node9613 : node9610;
																assign node9610 = (inp[5]) ? 4'b1001 : 4'b1000;
																assign node9613 = (inp[5]) ? 4'b1100 : 4'b1101;
															assign node9616 = (inp[5]) ? 4'b1010 : node9617;
																assign node9617 = (inp[15]) ? 4'b1111 : 4'b1011;
														assign node9621 = (inp[12]) ? 4'b1000 : 4'b1010;
				assign node9624 = (inp[7]) ? node12438 : node9625;
					assign node9625 = (inp[10]) ? node11001 : node9626;
						assign node9626 = (inp[0]) ? node10328 : node9627;
							assign node9627 = (inp[13]) ? node9939 : node9628;
								assign node9628 = (inp[1]) ? node9760 : node9629;
									assign node9629 = (inp[2]) ? node9687 : node9630;
										assign node9630 = (inp[4]) ? node9652 : node9631;
											assign node9631 = (inp[12]) ? node9641 : node9632;
												assign node9632 = (inp[11]) ? node9634 : 4'b1000;
													assign node9634 = (inp[14]) ? node9636 : 4'b1000;
														assign node9636 = (inp[5]) ? node9638 : 4'b1001;
															assign node9638 = (inp[15]) ? 4'b1000 : 4'b1101;
												assign node9641 = (inp[14]) ? node9643 : 4'b1010;
													assign node9643 = (inp[5]) ? 4'b1010 : node9644;
														assign node9644 = (inp[15]) ? node9648 : node9645;
															assign node9645 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node9648 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node9652 = (inp[12]) ? node9672 : node9653;
												assign node9653 = (inp[5]) ? node9663 : node9654;
													assign node9654 = (inp[14]) ? node9656 : 4'b1010;
														assign node9656 = (inp[11]) ? node9660 : node9657;
															assign node9657 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node9660 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node9663 = (inp[14]) ? node9669 : node9664;
														assign node9664 = (inp[15]) ? node9666 : 4'b1011;
															assign node9666 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node9669 = (inp[15]) ? 4'b1011 : 4'b1110;
												assign node9672 = (inp[5]) ? node9680 : node9673;
													assign node9673 = (inp[15]) ? node9677 : node9674;
														assign node9674 = (inp[14]) ? 4'b1000 : 4'b1100;
														assign node9677 = (inp[14]) ? 4'b1100 : 4'b1001;
													assign node9680 = (inp[14]) ? node9682 : 4'b1001;
														assign node9682 = (inp[15]) ? 4'b1001 : node9683;
															assign node9683 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node9687 = (inp[4]) ? node9715 : node9688;
											assign node9688 = (inp[12]) ? node9702 : node9689;
												assign node9689 = (inp[14]) ? node9691 : 4'b1100;
													assign node9691 = (inp[15]) ? node9697 : node9692;
														assign node9692 = (inp[5]) ? node9694 : 4'b1100;
															assign node9694 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node9697 = (inp[11]) ? 4'b1100 : node9698;
															assign node9698 = (inp[5]) ? 4'b1101 : 4'b1100;
												assign node9702 = (inp[14]) ? node9704 : 4'b1110;
													assign node9704 = (inp[11]) ? node9710 : node9705;
														assign node9705 = (inp[5]) ? 4'b1111 : node9706;
															assign node9706 = (inp[15]) ? 4'b1011 : 4'b1110;
														assign node9710 = (inp[5]) ? 4'b1110 : node9711;
															assign node9711 = (inp[15]) ? 4'b1010 : 4'b1110;
											assign node9715 = (inp[12]) ? node9733 : node9716;
												assign node9716 = (inp[5]) ? node9724 : node9717;
													assign node9717 = (inp[15]) ? node9719 : 4'b1111;
														assign node9719 = (inp[14]) ? node9721 : 4'b1111;
															assign node9721 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node9724 = (inp[15]) ? node9730 : node9725;
														assign node9725 = (inp[14]) ? 4'b1010 : node9726;
															assign node9726 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node9730 = (inp[14]) ? 4'b1110 : 4'b1010;
												assign node9733 = (inp[11]) ? node9749 : node9734;
													assign node9734 = (inp[15]) ? node9740 : node9735;
														assign node9735 = (inp[14]) ? node9737 : 4'b1001;
															assign node9737 = (inp[5]) ? 4'b1001 : 4'b1100;
														assign node9740 = (inp[9]) ? node9742 : 4'b1101;
															assign node9742 = (inp[14]) ? node9746 : node9743;
																assign node9743 = (inp[5]) ? 4'b1100 : 4'b1101;
																assign node9746 = (inp[5]) ? 4'b1101 : 4'b1000;
													assign node9749 = (inp[5]) ? node9755 : node9750;
														assign node9750 = (inp[15]) ? node9752 : 4'b1101;
															assign node9752 = (inp[14]) ? 4'b1000 : 4'b1100;
														assign node9755 = (inp[15]) ? 4'b1100 : node9756;
															assign node9756 = (inp[14]) ? 4'b1000 : 4'b1100;
									assign node9760 = (inp[2]) ? node9840 : node9761;
										assign node9761 = (inp[4]) ? node9797 : node9762;
											assign node9762 = (inp[12]) ? node9778 : node9763;
												assign node9763 = (inp[15]) ? node9771 : node9764;
													assign node9764 = (inp[14]) ? node9766 : 4'b1100;
														assign node9766 = (inp[5]) ? 4'b1000 : node9767;
															assign node9767 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node9771 = (inp[14]) ? node9773 : 4'b1101;
														assign node9773 = (inp[11]) ? 4'b1100 : node9774;
															assign node9774 = (inp[5]) ? 4'b1101 : 4'b1100;
												assign node9778 = (inp[5]) ? node9790 : node9779;
													assign node9779 = (inp[11]) ? node9785 : node9780;
														assign node9780 = (inp[14]) ? node9782 : 4'b1111;
															assign node9782 = (inp[9]) ? 4'b1111 : 4'b1010;
														assign node9785 = (inp[15]) ? node9787 : 4'b1110;
															assign node9787 = (inp[14]) ? 4'b1011 : 4'b1110;
													assign node9790 = (inp[15]) ? node9792 : 4'b1111;
														assign node9792 = (inp[11]) ? node9794 : 4'b1111;
															assign node9794 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node9797 = (inp[12]) ? node9817 : node9798;
												assign node9798 = (inp[14]) ? node9810 : node9799;
													assign node9799 = (inp[15]) ? node9805 : node9800;
														assign node9800 = (inp[11]) ? node9802 : 4'b1110;
															assign node9802 = (inp[5]) ? 4'b1111 : 4'b1110;
														assign node9805 = (inp[5]) ? node9807 : 4'b1111;
															assign node9807 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node9810 = (inp[5]) ? node9814 : node9811;
														assign node9811 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node9814 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node9817 = (inp[5]) ? node9827 : node9818;
													assign node9818 = (inp[15]) ? node9824 : node9819;
														assign node9819 = (inp[14]) ? 4'b1101 : node9820;
															assign node9820 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node9824 = (inp[14]) ? 4'b1000 : 4'b1100;
													assign node9827 = (inp[15]) ? node9831 : node9828;
														assign node9828 = (inp[14]) ? 4'b1000 : 4'b1100;
														assign node9831 = (inp[9]) ? node9833 : 4'b1101;
															assign node9833 = (inp[14]) ? node9837 : node9834;
																assign node9834 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node9837 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node9840 = (inp[4]) ? node9882 : node9841;
											assign node9841 = (inp[12]) ? node9859 : node9842;
												assign node9842 = (inp[15]) ? node9852 : node9843;
													assign node9843 = (inp[14]) ? node9847 : node9844;
														assign node9844 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node9847 = (inp[5]) ? 4'b1100 : node9848;
															assign node9848 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node9852 = (inp[11]) ? 4'b1001 : node9853;
														assign node9853 = (inp[14]) ? node9855 : 4'b1001;
															assign node9855 = (inp[5]) ? 4'b1000 : 4'b1001;
												assign node9859 = (inp[15]) ? node9875 : node9860;
													assign node9860 = (inp[5]) ? node9868 : node9861;
														assign node9861 = (inp[11]) ? node9865 : node9862;
															assign node9862 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node9865 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node9868 = (inp[9]) ? node9870 : 4'b1010;
															assign node9870 = (inp[14]) ? 4'b1010 : node9871;
																assign node9871 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node9875 = (inp[14]) ? node9877 : 4'b1010;
														assign node9877 = (inp[5]) ? node9879 : 4'b1110;
															assign node9879 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node9882 = (inp[12]) ? node9904 : node9883;
												assign node9883 = (inp[15]) ? node9895 : node9884;
													assign node9884 = (inp[5]) ? node9892 : node9885;
														assign node9885 = (inp[11]) ? node9889 : node9886;
															assign node9886 = (inp[14]) ? 4'b1010 : 4'b1011;
															assign node9889 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node9892 = (inp[14]) ? 4'b1110 : 4'b1010;
													assign node9895 = (inp[5]) ? node9899 : node9896;
														assign node9896 = (inp[14]) ? 4'b1110 : 4'b1010;
														assign node9899 = (inp[14]) ? 4'b1011 : node9900;
															assign node9900 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node9904 = (inp[15]) ? node9926 : node9905;
													assign node9905 = (inp[11]) ? node9919 : node9906;
														assign node9906 = (inp[9]) ? node9914 : node9907;
															assign node9907 = (inp[5]) ? node9911 : node9908;
																assign node9908 = (inp[14]) ? 4'b1001 : 4'b1100;
																assign node9911 = (inp[14]) ? 4'b1100 : 4'b1001;
															assign node9914 = (inp[14]) ? 4'b1100 : node9915;
																assign node9915 = (inp[5]) ? 4'b1001 : 4'b1100;
														assign node9919 = (inp[14]) ? node9923 : node9920;
															assign node9920 = (inp[5]) ? 4'b1000 : 4'b1101;
															assign node9923 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node9926 = (inp[5]) ? node9934 : node9927;
														assign node9927 = (inp[14]) ? node9931 : node9928;
															assign node9928 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node9931 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node9934 = (inp[14]) ? node9936 : 4'b1000;
															assign node9936 = (inp[11]) ? 4'b1000 : 4'b1001;
								assign node9939 = (inp[4]) ? node10103 : node9940;
									assign node9940 = (inp[12]) ? node10022 : node9941;
										assign node9941 = (inp[2]) ? node9977 : node9942;
											assign node9942 = (inp[1]) ? node9962 : node9943;
												assign node9943 = (inp[15]) ? node9951 : node9944;
													assign node9944 = (inp[14]) ? node9948 : node9945;
														assign node9945 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node9948 = (inp[5]) ? 4'b1100 : 4'b1000;
													assign node9951 = (inp[5]) ? node9957 : node9952;
														assign node9952 = (inp[11]) ? node9954 : 4'b1001;
															assign node9954 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node9957 = (inp[11]) ? 4'b1001 : node9958;
															assign node9958 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node9962 = (inp[15]) ? node9972 : node9963;
													assign node9963 = (inp[14]) ? node9967 : node9964;
														assign node9964 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node9967 = (inp[5]) ? node9969 : 4'b1100;
															assign node9969 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node9972 = (inp[5]) ? 4'b1100 : node9973;
														assign node9973 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node9977 = (inp[1]) ? node10007 : node9978;
												assign node9978 = (inp[15]) ? node9998 : node9979;
													assign node9979 = (inp[5]) ? node9993 : node9980;
														assign node9980 = (inp[9]) ? node9986 : node9981;
															assign node9981 = (inp[14]) ? node9983 : 4'b1101;
																assign node9983 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node9986 = (inp[11]) ? node9990 : node9987;
																assign node9987 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node9990 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node9993 = (inp[14]) ? 4'b1001 : node9994;
															assign node9994 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node9998 = (inp[11]) ? node10002 : node9999;
														assign node9999 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node10002 = (inp[5]) ? 4'b1100 : node10003;
															assign node10003 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node10007 = (inp[15]) ? node10013 : node10008;
													assign node10008 = (inp[5]) ? node10010 : 4'b1001;
														assign node10010 = (inp[14]) ? 4'b1101 : 4'b1001;
													assign node10013 = (inp[5]) ? node10017 : node10014;
														assign node10014 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node10017 = (inp[11]) ? 4'b1001 : node10018;
															assign node10018 = (inp[14]) ? 4'b1001 : 4'b1000;
										assign node10022 = (inp[2]) ? node10064 : node10023;
											assign node10023 = (inp[1]) ? node10051 : node10024;
												assign node10024 = (inp[5]) ? node10036 : node10025;
													assign node10025 = (inp[15]) ? node10031 : node10026;
														assign node10026 = (inp[14]) ? 4'b1010 : node10027;
															assign node10027 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node10031 = (inp[14]) ? 4'b1111 : node10032;
															assign node10032 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node10036 = (inp[15]) ? node10044 : node10037;
														assign node10037 = (inp[14]) ? node10041 : node10038;
															assign node10038 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node10041 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node10044 = (inp[9]) ? 4'b1010 : node10045;
															assign node10045 = (inp[11]) ? 4'b1010 : node10046;
																assign node10046 = (inp[14]) ? 4'b1010 : 4'b1011;
												assign node10051 = (inp[15]) ? node10059 : node10052;
													assign node10052 = (inp[14]) ? node10056 : node10053;
														assign node10053 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node10056 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node10059 = (inp[5]) ? 4'b1111 : node10060;
														assign node10060 = (inp[14]) ? 4'b1011 : 4'b1111;
											assign node10064 = (inp[1]) ? node10086 : node10065;
												assign node10065 = (inp[5]) ? node10077 : node10066;
													assign node10066 = (inp[14]) ? node10074 : node10067;
														assign node10067 = (inp[11]) ? node10071 : node10068;
															assign node10068 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node10071 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node10074 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node10077 = (inp[15]) ? node10081 : node10078;
														assign node10078 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node10081 = (inp[14]) ? 4'b1110 : node10082;
															assign node10082 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node10086 = (inp[15]) ? node10094 : node10087;
													assign node10087 = (inp[11]) ? 4'b1010 : node10088;
														assign node10088 = (inp[14]) ? node10090 : 4'b1010;
															assign node10090 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node10094 = (inp[14]) ? node10098 : node10095;
														assign node10095 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node10098 = (inp[5]) ? 4'b1010 : node10099;
															assign node10099 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node10103 = (inp[12]) ? node10199 : node10104;
										assign node10104 = (inp[2]) ? node10142 : node10105;
											assign node10105 = (inp[5]) ? node10123 : node10106;
												assign node10106 = (inp[1]) ? node10114 : node10107;
													assign node10107 = (inp[11]) ? 4'b1010 : node10108;
														assign node10108 = (inp[15]) ? node10110 : 4'b1010;
															assign node10110 = (inp[14]) ? 4'b1111 : 4'b1011;
													assign node10114 = (inp[15]) ? node10120 : node10115;
														assign node10115 = (inp[11]) ? node10117 : 4'b1110;
															assign node10117 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node10120 = (inp[14]) ? 4'b1010 : 4'b1110;
												assign node10123 = (inp[1]) ? node10131 : node10124;
													assign node10124 = (inp[14]) ? node10128 : node10125;
														assign node10125 = (inp[15]) ? 4'b1110 : 4'b1011;
														assign node10128 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node10131 = (inp[9]) ? 4'b1011 : node10132;
														assign node10132 = (inp[15]) ? node10136 : node10133;
															assign node10133 = (inp[14]) ? 4'b1011 : 4'b1111;
															assign node10136 = (inp[14]) ? node10138 : 4'b1011;
																assign node10138 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node10142 = (inp[1]) ? node10176 : node10143;
												assign node10143 = (inp[15]) ? node10163 : node10144;
													assign node10144 = (inp[5]) ? node10158 : node10145;
														assign node10145 = (inp[9]) ? node10151 : node10146;
															assign node10146 = (inp[11]) ? 4'b1111 : node10147;
																assign node10147 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node10151 = (inp[14]) ? node10155 : node10152;
																assign node10152 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node10155 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node10158 = (inp[14]) ? node10160 : 4'b1110;
															assign node10160 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node10163 = (inp[14]) ? node10171 : node10164;
														assign node10164 = (inp[5]) ? node10168 : node10165;
															assign node10165 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node10168 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node10171 = (inp[5]) ? node10173 : 4'b1011;
															assign node10173 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node10176 = (inp[15]) ? node10188 : node10177;
													assign node10177 = (inp[14]) ? node10183 : node10178;
														assign node10178 = (inp[11]) ? node10180 : 4'b1010;
															assign node10180 = (inp[5]) ? 4'b1011 : 4'b1010;
														assign node10183 = (inp[5]) ? node10185 : 4'b1010;
															assign node10185 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node10188 = (inp[5]) ? node10194 : node10189;
														assign node10189 = (inp[14]) ? node10191 : 4'b1011;
															assign node10191 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node10194 = (inp[14]) ? node10196 : 4'b1110;
															assign node10196 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node10199 = (inp[11]) ? node10267 : node10200;
											assign node10200 = (inp[2]) ? node10228 : node10201;
												assign node10201 = (inp[1]) ? node10215 : node10202;
													assign node10202 = (inp[14]) ? node10208 : node10203;
														assign node10203 = (inp[15]) ? 4'b1000 : node10204;
															assign node10204 = (inp[5]) ? 4'b1001 : 4'b1100;
														assign node10208 = (inp[15]) ? node10212 : node10209;
															assign node10209 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node10212 = (inp[5]) ? 4'b1001 : 4'b1100;
													assign node10215 = (inp[5]) ? node10223 : node10216;
														assign node10216 = (inp[15]) ? node10220 : node10217;
															assign node10217 = (inp[14]) ? 4'b1100 : 4'b1000;
															assign node10220 = (inp[14]) ? 4'b1000 : 4'b1101;
														assign node10223 = (inp[15]) ? 4'b1100 : node10224;
															assign node10224 = (inp[14]) ? 4'b1001 : 4'b1100;
												assign node10228 = (inp[15]) ? node10258 : node10229;
													assign node10229 = (inp[9]) ? node10243 : node10230;
														assign node10230 = (inp[5]) ? node10238 : node10231;
															assign node10231 = (inp[14]) ? node10235 : node10232;
																assign node10232 = (inp[1]) ? 4'b1101 : 4'b1000;
																assign node10235 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node10238 = (inp[14]) ? node10240 : 4'b1100;
																assign node10240 = (inp[1]) ? 4'b1100 : 4'b1001;
														assign node10243 = (inp[5]) ? node10251 : node10244;
															assign node10244 = (inp[1]) ? node10248 : node10245;
																assign node10245 = (inp[14]) ? 4'b1100 : 4'b1000;
																assign node10248 = (inp[14]) ? 4'b1000 : 4'b1101;
															assign node10251 = (inp[14]) ? node10255 : node10252;
																assign node10252 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node10255 = (inp[1]) ? 4'b1100 : 4'b1001;
													assign node10258 = (inp[1]) ? node10264 : node10259;
														assign node10259 = (inp[14]) ? node10261 : 4'b1101;
															assign node10261 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node10264 = (inp[14]) ? 4'b1101 : 4'b1001;
											assign node10267 = (inp[5]) ? node10303 : node10268;
												assign node10268 = (inp[14]) ? node10288 : node10269;
													assign node10269 = (inp[2]) ? node10277 : node10270;
														assign node10270 = (inp[1]) ? node10274 : node10271;
															assign node10271 = (inp[15]) ? 4'b1000 : 4'b1101;
															assign node10274 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node10277 = (inp[9]) ? node10283 : node10278;
															assign node10278 = (inp[1]) ? node10280 : 4'b1000;
																assign node10280 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node10283 = (inp[15]) ? node10285 : 4'b1101;
																assign node10285 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node10288 = (inp[1]) ? node10296 : node10289;
														assign node10289 = (inp[15]) ? node10293 : node10290;
															assign node10290 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node10293 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node10296 = (inp[15]) ? node10300 : node10297;
															assign node10297 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node10300 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node10303 = (inp[1]) ? node10315 : node10304;
													assign node10304 = (inp[15]) ? node10310 : node10305;
														assign node10305 = (inp[2]) ? node10307 : 4'b1101;
															assign node10307 = (inp[14]) ? 4'b1001 : 4'b1101;
														assign node10310 = (inp[14]) ? node10312 : 4'b1001;
															assign node10312 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node10315 = (inp[2]) ? node10323 : node10316;
														assign node10316 = (inp[14]) ? node10320 : node10317;
															assign node10317 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node10320 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node10323 = (inp[14]) ? node10325 : 4'b1000;
															assign node10325 = (inp[15]) ? 4'b1000 : 4'b1100;
							assign node10328 = (inp[13]) ? node10640 : node10329;
								assign node10329 = (inp[1]) ? node10465 : node10330;
									assign node10330 = (inp[2]) ? node10406 : node10331;
										assign node10331 = (inp[14]) ? node10349 : node10332;
											assign node10332 = (inp[4]) ? node10336 : node10333;
												assign node10333 = (inp[12]) ? 4'b1011 : 4'b1001;
												assign node10336 = (inp[12]) ? node10342 : node10337;
													assign node10337 = (inp[5]) ? node10339 : 4'b1011;
														assign node10339 = (inp[11]) ? 4'b1010 : 4'b1111;
													assign node10342 = (inp[5]) ? 4'b1000 : node10343;
														assign node10343 = (inp[15]) ? node10345 : 4'b1101;
															assign node10345 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node10349 = (inp[11]) ? node10377 : node10350;
												assign node10350 = (inp[5]) ? node10366 : node10351;
													assign node10351 = (inp[15]) ? node10359 : node10352;
														assign node10352 = (inp[4]) ? node10356 : node10353;
															assign node10353 = (inp[12]) ? 4'b1011 : 4'b1001;
															assign node10356 = (inp[12]) ? 4'b1001 : 4'b1011;
														assign node10359 = (inp[4]) ? node10363 : node10360;
															assign node10360 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node10363 = (inp[12]) ? 4'b1101 : 4'b1111;
													assign node10366 = (inp[4]) ? node10372 : node10367;
														assign node10367 = (inp[12]) ? 4'b1011 : node10368;
															assign node10368 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node10372 = (inp[15]) ? node10374 : 4'b1100;
															assign node10374 = (inp[12]) ? 4'b1000 : 4'b1010;
												assign node10377 = (inp[5]) ? node10393 : node10378;
													assign node10378 = (inp[15]) ? node10386 : node10379;
														assign node10379 = (inp[12]) ? node10383 : node10380;
															assign node10380 = (inp[4]) ? 4'b1010 : 4'b1000;
															assign node10383 = (inp[4]) ? 4'b1001 : 4'b1010;
														assign node10386 = (inp[4]) ? node10390 : node10387;
															assign node10387 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node10390 = (inp[12]) ? 4'b1101 : 4'b1110;
													assign node10393 = (inp[15]) ? node10399 : node10394;
														assign node10394 = (inp[12]) ? 4'b1011 : node10395;
															assign node10395 = (inp[4]) ? 4'b1111 : 4'b1100;
														assign node10399 = (inp[12]) ? node10403 : node10400;
															assign node10400 = (inp[4]) ? 4'b1011 : 4'b1001;
															assign node10403 = (inp[4]) ? 4'b1000 : 4'b1011;
										assign node10406 = (inp[4]) ? node10430 : node10407;
											assign node10407 = (inp[12]) ? node10419 : node10408;
												assign node10408 = (inp[14]) ? node10410 : 4'b1101;
													assign node10410 = (inp[5]) ? node10412 : 4'b1101;
														assign node10412 = (inp[15]) ? node10416 : node10413;
															assign node10413 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10416 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node10419 = (inp[14]) ? node10421 : 4'b1111;
													assign node10421 = (inp[11]) ? node10427 : node10422;
														assign node10422 = (inp[5]) ? 4'b1110 : node10423;
															assign node10423 = (inp[9]) ? 4'b1010 : 4'b1111;
														assign node10427 = (inp[15]) ? 4'b1011 : 4'b1111;
											assign node10430 = (inp[12]) ? node10446 : node10431;
												assign node10431 = (inp[5]) ? node10439 : node10432;
													assign node10432 = (inp[14]) ? node10434 : 4'b1110;
														assign node10434 = (inp[15]) ? node10436 : 4'b1110;
															assign node10436 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node10439 = (inp[15]) ? node10443 : node10440;
														assign node10440 = (inp[14]) ? 4'b1011 : 4'b1110;
														assign node10443 = (inp[14]) ? 4'b1111 : 4'b1011;
												assign node10446 = (inp[14]) ? node10456 : node10447;
													assign node10447 = (inp[5]) ? 4'b1101 : node10448;
														assign node10448 = (inp[11]) ? node10452 : node10449;
															assign node10449 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node10452 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node10456 = (inp[5]) ? node10460 : node10457;
														assign node10457 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node10460 = (inp[11]) ? node10462 : 4'b1000;
															assign node10462 = (inp[15]) ? 4'b1101 : 4'b1001;
									assign node10465 = (inp[2]) ? node10551 : node10466;
										assign node10466 = (inp[4]) ? node10500 : node10467;
											assign node10467 = (inp[12]) ? node10487 : node10468;
												assign node10468 = (inp[15]) ? node10478 : node10469;
													assign node10469 = (inp[5]) ? node10475 : node10470;
														assign node10470 = (inp[14]) ? node10472 : 4'b1101;
															assign node10472 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node10475 = (inp[14]) ? 4'b1001 : 4'b1101;
													assign node10478 = (inp[14]) ? node10482 : node10479;
														assign node10479 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node10482 = (inp[9]) ? 4'b1101 : node10483;
															assign node10483 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node10487 = (inp[14]) ? node10489 : 4'b1110;
													assign node10489 = (inp[15]) ? node10493 : node10490;
														assign node10490 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node10493 = (inp[11]) ? node10497 : node10494;
															assign node10494 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node10497 = (inp[5]) ? 4'b1110 : 4'b1010;
											assign node10500 = (inp[12]) ? node10530 : node10501;
												assign node10501 = (inp[5]) ? node10509 : node10502;
													assign node10502 = (inp[11]) ? 4'b1110 : node10503;
														assign node10503 = (inp[14]) ? node10505 : 4'b1111;
															assign node10505 = (inp[15]) ? 4'b1010 : 4'b1111;
													assign node10509 = (inp[11]) ? node10517 : node10510;
														assign node10510 = (inp[14]) ? node10514 : node10511;
															assign node10511 = (inp[15]) ? 4'b1010 : 4'b1111;
															assign node10514 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node10517 = (inp[9]) ? node10525 : node10518;
															assign node10518 = (inp[14]) ? node10522 : node10519;
																assign node10519 = (inp[15]) ? 4'b1011 : 4'b1110;
																assign node10522 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node10525 = (inp[14]) ? node10527 : 4'b1011;
																assign node10527 = (inp[15]) ? 4'b1110 : 4'b1011;
												assign node10530 = (inp[14]) ? node10542 : node10531;
													assign node10531 = (inp[5]) ? node10537 : node10532;
														assign node10532 = (inp[15]) ? 4'b1101 : node10533;
															assign node10533 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node10537 = (inp[11]) ? node10539 : 4'b1101;
															assign node10539 = (inp[15]) ? 4'b1100 : 4'b1101;
													assign node10542 = (inp[15]) ? node10546 : node10543;
														assign node10543 = (inp[5]) ? 4'b1001 : 4'b1100;
														assign node10546 = (inp[5]) ? node10548 : 4'b1001;
															assign node10548 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node10551 = (inp[4]) ? node10593 : node10552;
											assign node10552 = (inp[12]) ? node10572 : node10553;
												assign node10553 = (inp[15]) ? node10565 : node10554;
													assign node10554 = (inp[14]) ? node10558 : node10555;
														assign node10555 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node10558 = (inp[11]) ? node10562 : node10559;
															assign node10559 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node10562 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node10565 = (inp[11]) ? 4'b1000 : node10566;
														assign node10566 = (inp[5]) ? node10568 : 4'b1000;
															assign node10568 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node10572 = (inp[15]) ? node10584 : node10573;
													assign node10573 = (inp[5]) ? node10579 : node10574;
														assign node10574 = (inp[11]) ? node10576 : 4'b1010;
															assign node10576 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node10579 = (inp[14]) ? 4'b1011 : node10580;
															assign node10580 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node10584 = (inp[5]) ? node10588 : node10585;
														assign node10585 = (inp[14]) ? 4'b1111 : 4'b1011;
														assign node10588 = (inp[11]) ? 4'b1011 : node10589;
															assign node10589 = (inp[14]) ? 4'b1010 : 4'b1011;
											assign node10593 = (inp[12]) ? node10613 : node10594;
												assign node10594 = (inp[5]) ? node10604 : node10595;
													assign node10595 = (inp[14]) ? node10601 : node10596;
														assign node10596 = (inp[15]) ? 4'b1011 : node10597;
															assign node10597 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node10601 = (inp[11]) ? 4'b1111 : 4'b1011;
													assign node10604 = (inp[15]) ? node10608 : node10605;
														assign node10605 = (inp[14]) ? 4'b1111 : 4'b1011;
														assign node10608 = (inp[14]) ? 4'b1010 : node10609;
															assign node10609 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node10613 = (inp[15]) ? node10627 : node10614;
													assign node10614 = (inp[14]) ? node10622 : node10615;
														assign node10615 = (inp[5]) ? node10619 : node10616;
															assign node10616 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node10619 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node10622 = (inp[5]) ? node10624 : 4'b1000;
															assign node10624 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node10627 = (inp[14]) ? node10633 : node10628;
														assign node10628 = (inp[5]) ? 4'b1001 : node10629;
															assign node10629 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node10633 = (inp[5]) ? node10637 : node10634;
															assign node10634 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node10637 = (inp[11]) ? 4'b1001 : 4'b1000;
								assign node10640 = (inp[14]) ? node10794 : node10641;
									assign node10641 = (inp[12]) ? node10711 : node10642;
										assign node10642 = (inp[4]) ? node10674 : node10643;
											assign node10643 = (inp[15]) ? node10659 : node10644;
												assign node10644 = (inp[11]) ? node10652 : node10645;
													assign node10645 = (inp[2]) ? node10649 : node10646;
														assign node10646 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node10649 = (inp[1]) ? 4'b1000 : 4'b1101;
													assign node10652 = (inp[2]) ? node10656 : node10653;
														assign node10653 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node10656 = (inp[1]) ? 4'b1000 : 4'b1100;
												assign node10659 = (inp[11]) ? node10667 : node10660;
													assign node10660 = (inp[1]) ? node10664 : node10661;
														assign node10661 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node10664 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node10667 = (inp[2]) ? node10671 : node10668;
														assign node10668 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node10671 = (inp[1]) ? 4'b1000 : 4'b1101;
											assign node10674 = (inp[2]) ? node10692 : node10675;
												assign node10675 = (inp[5]) ? node10685 : node10676;
													assign node10676 = (inp[1]) ? 4'b1111 : node10677;
														assign node10677 = (inp[11]) ? node10681 : node10678;
															assign node10678 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node10681 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node10685 = (inp[15]) ? node10689 : node10686;
														assign node10686 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node10689 = (inp[1]) ? 4'b1010 : 4'b1111;
												assign node10692 = (inp[1]) ? node10704 : node10693;
													assign node10693 = (inp[15]) ? node10699 : node10694;
														assign node10694 = (inp[11]) ? 4'b1111 : node10695;
															assign node10695 = (inp[5]) ? 4'b1111 : 4'b1110;
														assign node10699 = (inp[5]) ? node10701 : 4'b1111;
															assign node10701 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node10704 = (inp[15]) ? node10708 : node10705;
														assign node10705 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node10708 = (inp[9]) ? 4'b1111 : 4'b1011;
										assign node10711 = (inp[4]) ? node10749 : node10712;
											assign node10712 = (inp[11]) ? node10728 : node10713;
												assign node10713 = (inp[15]) ? node10721 : node10714;
													assign node10714 = (inp[2]) ? node10718 : node10715;
														assign node10715 = (inp[1]) ? 4'b1110 : 4'b1011;
														assign node10718 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node10721 = (inp[2]) ? node10725 : node10722;
														assign node10722 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node10725 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node10728 = (inp[15]) ? node10736 : node10729;
													assign node10729 = (inp[1]) ? node10733 : node10730;
														assign node10730 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node10733 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node10736 = (inp[9]) ? node10742 : node10737;
														assign node10737 = (inp[2]) ? node10739 : 4'b1011;
															assign node10739 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node10742 = (inp[5]) ? node10744 : 4'b1011;
															assign node10744 = (inp[1]) ? node10746 : 4'b1011;
																assign node10746 = (inp[2]) ? 4'b1011 : 4'b1110;
											assign node10749 = (inp[2]) ? node10773 : node10750;
												assign node10750 = (inp[1]) ? node10762 : node10751;
													assign node10751 = (inp[5]) ? node10755 : node10752;
														assign node10752 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node10755 = (inp[15]) ? node10759 : node10756;
															assign node10756 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node10759 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node10762 = (inp[5]) ? node10768 : node10763;
														assign node10763 = (inp[15]) ? node10765 : 4'b1001;
															assign node10765 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node10768 = (inp[15]) ? 4'b1101 : node10769;
															assign node10769 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node10773 = (inp[5]) ? node10781 : node10774;
													assign node10774 = (inp[15]) ? node10778 : node10775;
														assign node10775 = (inp[1]) ? 4'b1100 : 4'b1001;
														assign node10778 = (inp[1]) ? 4'b1000 : 4'b1100;
													assign node10781 = (inp[1]) ? node10789 : node10782;
														assign node10782 = (inp[15]) ? node10786 : node10783;
															assign node10783 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node10786 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node10789 = (inp[15]) ? node10791 : 4'b1001;
															assign node10791 = (inp[11]) ? 4'b1001 : 4'b1000;
									assign node10794 = (inp[12]) ? node10886 : node10795;
										assign node10795 = (inp[4]) ? node10839 : node10796;
											assign node10796 = (inp[2]) ? node10818 : node10797;
												assign node10797 = (inp[1]) ? node10807 : node10798;
													assign node10798 = (inp[15]) ? node10802 : node10799;
														assign node10799 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node10802 = (inp[5]) ? node10804 : 4'b1000;
															assign node10804 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node10807 = (inp[5]) ? node10813 : node10808;
														assign node10808 = (inp[15]) ? node10810 : 4'b1101;
															assign node10810 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node10813 = (inp[15]) ? 4'b1101 : node10814;
															assign node10814 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node10818 = (inp[1]) ? node10830 : node10819;
													assign node10819 = (inp[15]) ? node10825 : node10820;
														assign node10820 = (inp[5]) ? 4'b1000 : node10821;
															assign node10821 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node10825 = (inp[5]) ? 4'b1101 : node10826;
															assign node10826 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node10830 = (inp[15]) ? node10834 : node10831;
														assign node10831 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node10834 = (inp[11]) ? node10836 : 4'b1000;
															assign node10836 = (inp[5]) ? 4'b1000 : 4'b1001;
											assign node10839 = (inp[5]) ? node10859 : node10840;
												assign node10840 = (inp[1]) ? node10850 : node10841;
													assign node10841 = (inp[15]) ? node10847 : node10842;
														assign node10842 = (inp[2]) ? node10844 : 4'b1011;
															assign node10844 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node10847 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node10850 = (inp[2]) ? node10854 : node10851;
														assign node10851 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node10854 = (inp[15]) ? node10856 : 4'b1011;
															assign node10856 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node10859 = (inp[11]) ? node10875 : node10860;
													assign node10860 = (inp[15]) ? node10868 : node10861;
														assign node10861 = (inp[1]) ? node10865 : node10862;
															assign node10862 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node10865 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node10868 = (inp[1]) ? node10872 : node10869;
															assign node10869 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node10872 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node10875 = (inp[2]) ? node10883 : node10876;
														assign node10876 = (inp[1]) ? node10880 : node10877;
															assign node10877 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node10880 = (inp[15]) ? 4'b1111 : 4'b1010;
														assign node10883 = (inp[15]) ? 4'b1110 : 4'b1111;
										assign node10886 = (inp[4]) ? node10930 : node10887;
											assign node10887 = (inp[2]) ? node10909 : node10888;
												assign node10888 = (inp[1]) ? node10900 : node10889;
													assign node10889 = (inp[15]) ? node10895 : node10890;
														assign node10890 = (inp[11]) ? 4'b1011 : node10891;
															assign node10891 = (inp[5]) ? 4'b1010 : 4'b1011;
														assign node10895 = (inp[5]) ? node10897 : 4'b1110;
															assign node10897 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node10900 = (inp[15]) ? node10906 : node10901;
														assign node10901 = (inp[5]) ? node10903 : 4'b1110;
															assign node10903 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node10906 = (inp[5]) ? 4'b1110 : 4'b1010;
												assign node10909 = (inp[1]) ? node10919 : node10910;
													assign node10910 = (inp[15]) ? node10916 : node10911;
														assign node10911 = (inp[11]) ? node10913 : 4'b1110;
															assign node10913 = (inp[5]) ? 4'b1110 : 4'b1111;
														assign node10916 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node10919 = (inp[5]) ? node10925 : node10920;
														assign node10920 = (inp[15]) ? node10922 : 4'b1011;
															assign node10922 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node10925 = (inp[11]) ? 4'b1011 : node10926;
															assign node10926 = (inp[15]) ? 4'b1011 : 4'b1010;
											assign node10930 = (inp[11]) ? node10962 : node10931;
												assign node10931 = (inp[5]) ? node10947 : node10932;
													assign node10932 = (inp[2]) ? node10940 : node10933;
														assign node10933 = (inp[1]) ? node10937 : node10934;
															assign node10934 = (inp[15]) ? 4'b1101 : 4'b1000;
															assign node10937 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node10940 = (inp[15]) ? node10944 : node10941;
															assign node10941 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node10944 = (inp[1]) ? 4'b1100 : 4'b1001;
													assign node10947 = (inp[15]) ? node10955 : node10948;
														assign node10948 = (inp[2]) ? node10952 : node10949;
															assign node10949 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node10952 = (inp[1]) ? 4'b1101 : 4'b1000;
														assign node10955 = (inp[2]) ? node10959 : node10956;
															assign node10956 = (inp[1]) ? 4'b1101 : 4'b1000;
															assign node10959 = (inp[1]) ? 4'b1001 : 4'b1101;
												assign node10962 = (inp[5]) ? node10986 : node10963;
													assign node10963 = (inp[15]) ? node10971 : node10964;
														assign node10964 = (inp[1]) ? node10968 : node10965;
															assign node10965 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node10968 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node10971 = (inp[9]) ? node10979 : node10972;
															assign node10972 = (inp[2]) ? node10976 : node10973;
																assign node10973 = (inp[1]) ? 4'b1000 : 4'b1100;
																assign node10976 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node10979 = (inp[1]) ? node10983 : node10980;
																assign node10980 = (inp[2]) ? 4'b1000 : 4'b1100;
																assign node10983 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node10986 = (inp[15]) ? node10994 : node10987;
														assign node10987 = (inp[1]) ? node10991 : node10988;
															assign node10988 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node10991 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node10994 = (inp[1]) ? node10998 : node10995;
															assign node10995 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node10998 = (inp[2]) ? 4'b1001 : 4'b1101;
						assign node11001 = (inp[0]) ? node11731 : node11002;
							assign node11002 = (inp[13]) ? node11340 : node11003;
								assign node11003 = (inp[1]) ? node11159 : node11004;
									assign node11004 = (inp[2]) ? node11082 : node11005;
										assign node11005 = (inp[4]) ? node11029 : node11006;
											assign node11006 = (inp[12]) ? node11018 : node11007;
												assign node11007 = (inp[15]) ? 4'b1001 : node11008;
													assign node11008 = (inp[5]) ? node11014 : node11009;
														assign node11009 = (inp[9]) ? 4'b1001 : node11010;
															assign node11010 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node11014 = (inp[14]) ? 4'b1101 : 4'b1001;
												assign node11018 = (inp[14]) ? node11020 : 4'b1011;
													assign node11020 = (inp[5]) ? 4'b1011 : node11021;
														assign node11021 = (inp[15]) ? node11025 : node11022;
															assign node11022 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node11025 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node11029 = (inp[12]) ? node11059 : node11030;
												assign node11030 = (inp[11]) ? node11046 : node11031;
													assign node11031 = (inp[5]) ? node11037 : node11032;
														assign node11032 = (inp[15]) ? node11034 : 4'b1011;
															assign node11034 = (inp[14]) ? 4'b1111 : 4'b1011;
														assign node11037 = (inp[9]) ? 4'b1010 : node11038;
															assign node11038 = (inp[15]) ? node11042 : node11039;
																assign node11039 = (inp[14]) ? 4'b1111 : 4'b1011;
																assign node11042 = (inp[14]) ? 4'b1010 : 4'b1111;
													assign node11046 = (inp[5]) ? node11052 : node11047;
														assign node11047 = (inp[14]) ? node11049 : 4'b1011;
															assign node11049 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node11052 = (inp[14]) ? node11056 : node11053;
															assign node11053 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node11056 = (inp[15]) ? 4'b1011 : 4'b1111;
												assign node11059 = (inp[5]) ? node11075 : node11060;
													assign node11060 = (inp[9]) ? node11068 : node11061;
														assign node11061 = (inp[14]) ? node11065 : node11062;
															assign node11062 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node11065 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node11068 = (inp[15]) ? node11072 : node11069;
															assign node11069 = (inp[11]) ? 4'b1101 : 4'b1001;
															assign node11072 = (inp[11]) ? 4'b1000 : 4'b1101;
													assign node11075 = (inp[15]) ? 4'b1000 : node11076;
														assign node11076 = (inp[14]) ? node11078 : 4'b1000;
															assign node11078 = (inp[11]) ? 4'b1101 : 4'b1100;
										assign node11082 = (inp[4]) ? node11110 : node11083;
											assign node11083 = (inp[12]) ? node11095 : node11084;
												assign node11084 = (inp[5]) ? node11086 : 4'b1101;
													assign node11086 = (inp[14]) ? node11088 : 4'b1101;
														assign node11088 = (inp[11]) ? node11092 : node11089;
															assign node11089 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node11092 = (inp[15]) ? 4'b1101 : 4'b1001;
												assign node11095 = (inp[14]) ? node11097 : 4'b1111;
													assign node11097 = (inp[11]) ? node11105 : node11098;
														assign node11098 = (inp[15]) ? node11102 : node11099;
															assign node11099 = (inp[5]) ? 4'b1110 : 4'b1111;
															assign node11102 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node11105 = (inp[5]) ? 4'b1111 : node11106;
															assign node11106 = (inp[15]) ? 4'b1011 : 4'b1111;
											assign node11110 = (inp[12]) ? node11128 : node11111;
												assign node11111 = (inp[5]) ? node11119 : node11112;
													assign node11112 = (inp[15]) ? node11114 : 4'b1110;
														assign node11114 = (inp[14]) ? node11116 : 4'b1110;
															assign node11116 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node11119 = (inp[14]) ? node11125 : node11120;
														assign node11120 = (inp[15]) ? 4'b1011 : node11121;
															assign node11121 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node11125 = (inp[15]) ? 4'b1111 : 4'b1011;
												assign node11128 = (inp[11]) ? node11144 : node11129;
													assign node11129 = (inp[15]) ? node11137 : node11130;
														assign node11130 = (inp[14]) ? node11134 : node11131;
															assign node11131 = (inp[5]) ? 4'b1101 : 4'b1000;
															assign node11134 = (inp[5]) ? 4'b1000 : 4'b1101;
														assign node11137 = (inp[5]) ? node11141 : node11138;
															assign node11138 = (inp[14]) ? 4'b1001 : 4'b1100;
															assign node11141 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node11144 = (inp[5]) ? node11154 : node11145;
														assign node11145 = (inp[9]) ? node11147 : 4'b1100;
															assign node11147 = (inp[15]) ? node11151 : node11148;
																assign node11148 = (inp[14]) ? 4'b1100 : 4'b1001;
																assign node11151 = (inp[14]) ? 4'b1001 : 4'b1101;
														assign node11154 = (inp[14]) ? node11156 : 4'b1101;
															assign node11156 = (inp[15]) ? 4'b1101 : 4'b1001;
									assign node11159 = (inp[2]) ? node11257 : node11160;
										assign node11160 = (inp[4]) ? node11210 : node11161;
											assign node11161 = (inp[12]) ? node11179 : node11162;
												assign node11162 = (inp[15]) ? node11170 : node11163;
													assign node11163 = (inp[14]) ? node11165 : 4'b1101;
														assign node11165 = (inp[11]) ? 4'b1100 : node11166;
															assign node11166 = (inp[5]) ? 4'b1001 : 4'b1101;
													assign node11170 = (inp[11]) ? node11176 : node11171;
														assign node11171 = (inp[14]) ? node11173 : 4'b1101;
															assign node11173 = (inp[5]) ? 4'b1100 : 4'b1101;
														assign node11176 = (inp[14]) ? 4'b1101 : 4'b1100;
												assign node11179 = (inp[15]) ? node11187 : node11180;
													assign node11180 = (inp[11]) ? node11182 : 4'b1110;
														assign node11182 = (inp[5]) ? 4'b1110 : node11183;
															assign node11183 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node11187 = (inp[5]) ? node11195 : node11188;
														assign node11188 = (inp[14]) ? node11192 : node11189;
															assign node11189 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node11192 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node11195 = (inp[9]) ? node11203 : node11196;
															assign node11196 = (inp[14]) ? node11200 : node11197;
																assign node11197 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node11200 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node11203 = (inp[14]) ? node11207 : node11204;
																assign node11204 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node11207 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node11210 = (inp[12]) ? node11234 : node11211;
												assign node11211 = (inp[14]) ? node11221 : node11212;
													assign node11212 = (inp[5]) ? node11214 : 4'b1111;
														assign node11214 = (inp[15]) ? node11218 : node11215;
															assign node11215 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node11218 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node11221 = (inp[15]) ? node11229 : node11222;
														assign node11222 = (inp[5]) ? node11226 : node11223;
															assign node11223 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node11226 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11229 = (inp[5]) ? 4'b1110 : node11230;
															assign node11230 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node11234 = (inp[5]) ? node11244 : node11235;
													assign node11235 = (inp[15]) ? node11241 : node11236;
														assign node11236 = (inp[14]) ? 4'b1100 : node11237;
															assign node11237 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node11241 = (inp[14]) ? 4'b1001 : 4'b1101;
													assign node11244 = (inp[15]) ? node11248 : node11245;
														assign node11245 = (inp[14]) ? 4'b1001 : 4'b1101;
														assign node11248 = (inp[9]) ? 4'b1101 : node11249;
															assign node11249 = (inp[11]) ? node11253 : node11250;
																assign node11250 = (inp[14]) ? 4'b1100 : 4'b1101;
																assign node11253 = (inp[14]) ? 4'b1101 : 4'b1100;
										assign node11257 = (inp[14]) ? node11295 : node11258;
											assign node11258 = (inp[4]) ? node11270 : node11259;
												assign node11259 = (inp[12]) ? node11265 : node11260;
													assign node11260 = (inp[15]) ? 4'b1000 : node11261;
														assign node11261 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node11265 = (inp[11]) ? 4'b1011 : node11266;
														assign node11266 = (inp[15]) ? 4'b1011 : 4'b1010;
												assign node11270 = (inp[12]) ? node11280 : node11271;
													assign node11271 = (inp[5]) ? node11277 : node11272;
														assign node11272 = (inp[15]) ? 4'b1011 : node11273;
															assign node11273 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11277 = (inp[15]) ? 4'b1110 : 4'b1011;
													assign node11280 = (inp[5]) ? node11288 : node11281;
														assign node11281 = (inp[15]) ? node11285 : node11282;
															assign node11282 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node11285 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node11288 = (inp[9]) ? 4'b1001 : node11289;
															assign node11289 = (inp[11]) ? 4'b1001 : node11290;
																assign node11290 = (inp[15]) ? 4'b1001 : 4'b1000;
											assign node11295 = (inp[4]) ? node11319 : node11296;
												assign node11296 = (inp[12]) ? node11310 : node11297;
													assign node11297 = (inp[15]) ? node11305 : node11298;
														assign node11298 = (inp[11]) ? node11302 : node11299;
															assign node11299 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node11302 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node11305 = (inp[11]) ? 4'b1000 : node11306;
															assign node11306 = (inp[5]) ? 4'b1001 : 4'b1000;
													assign node11310 = (inp[11]) ? node11314 : node11311;
														assign node11311 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node11314 = (inp[5]) ? 4'b1011 : node11315;
															assign node11315 = (inp[15]) ? 4'b1111 : 4'b1010;
												assign node11319 = (inp[12]) ? node11327 : node11320;
													assign node11320 = (inp[15]) ? node11324 : node11321;
														assign node11321 = (inp[5]) ? 4'b1111 : 4'b1010;
														assign node11324 = (inp[5]) ? 4'b1010 : 4'b1111;
													assign node11327 = (inp[15]) ? node11333 : node11328;
														assign node11328 = (inp[5]) ? node11330 : 4'b1000;
															assign node11330 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node11333 = (inp[5]) ? node11337 : node11334;
															assign node11334 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node11337 = (inp[11]) ? 4'b1001 : 4'b1000;
								assign node11340 = (inp[4]) ? node11512 : node11341;
									assign node11341 = (inp[12]) ? node11431 : node11342;
										assign node11342 = (inp[2]) ? node11384 : node11343;
											assign node11343 = (inp[1]) ? node11367 : node11344;
												assign node11344 = (inp[15]) ? node11352 : node11345;
													assign node11345 = (inp[14]) ? node11349 : node11346;
														assign node11346 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node11349 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node11352 = (inp[5]) ? node11358 : node11353;
														assign node11353 = (inp[14]) ? 4'b1000 : node11354;
															assign node11354 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node11358 = (inp[9]) ? node11360 : 4'b1001;
															assign node11360 = (inp[11]) ? node11364 : node11361;
																assign node11361 = (inp[14]) ? 4'b1001 : 4'b1000;
																assign node11364 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node11367 = (inp[15]) ? node11377 : node11368;
													assign node11368 = (inp[11]) ? node11374 : node11369;
														assign node11369 = (inp[14]) ? node11371 : 4'b1101;
															assign node11371 = (inp[5]) ? 4'b1000 : 4'b1101;
														assign node11374 = (inp[14]) ? 4'b1001 : 4'b1100;
													assign node11377 = (inp[14]) ? node11379 : 4'b1101;
														assign node11379 = (inp[11]) ? node11381 : 4'b1101;
															assign node11381 = (inp[5]) ? 4'b1101 : 4'b1100;
											assign node11384 = (inp[1]) ? node11408 : node11385;
												assign node11385 = (inp[15]) ? node11399 : node11386;
													assign node11386 = (inp[5]) ? node11394 : node11387;
														assign node11387 = (inp[11]) ? node11391 : node11388;
															assign node11388 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node11391 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node11394 = (inp[14]) ? 4'b1000 : node11395;
															assign node11395 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node11399 = (inp[11]) ? node11403 : node11400;
														assign node11400 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node11403 = (inp[5]) ? 4'b1101 : node11404;
															assign node11404 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node11408 = (inp[15]) ? node11414 : node11409;
													assign node11409 = (inp[5]) ? node11411 : 4'b1000;
														assign node11411 = (inp[14]) ? 4'b1100 : 4'b1000;
													assign node11414 = (inp[5]) ? 4'b1000 : node11415;
														assign node11415 = (inp[9]) ? node11423 : node11416;
															assign node11416 = (inp[14]) ? node11420 : node11417;
																assign node11417 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node11420 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node11423 = (inp[14]) ? node11427 : node11424;
																assign node11424 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node11427 = (inp[11]) ? 4'b1001 : 4'b1000;
										assign node11431 = (inp[2]) ? node11475 : node11432;
											assign node11432 = (inp[1]) ? node11452 : node11433;
												assign node11433 = (inp[15]) ? node11443 : node11434;
													assign node11434 = (inp[14]) ? node11438 : node11435;
														assign node11435 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node11438 = (inp[5]) ? node11440 : 4'b1011;
															assign node11440 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node11443 = (inp[14]) ? node11447 : node11444;
														assign node11444 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11447 = (inp[5]) ? node11449 : 4'b1110;
															assign node11449 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node11452 = (inp[15]) ? node11470 : node11453;
													assign node11453 = (inp[9]) ? node11463 : node11454;
														assign node11454 = (inp[11]) ? node11460 : node11455;
															assign node11455 = (inp[5]) ? node11457 : 4'b1110;
																assign node11457 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node11460 = (inp[5]) ? 4'b1110 : 4'b1111;
														assign node11463 = (inp[14]) ? node11467 : node11464;
															assign node11464 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node11467 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node11470 = (inp[14]) ? node11472 : 4'b1110;
														assign node11472 = (inp[5]) ? 4'b1110 : 4'b1010;
											assign node11475 = (inp[1]) ? node11493 : node11476;
												assign node11476 = (inp[15]) ? node11486 : node11477;
													assign node11477 = (inp[9]) ? node11479 : 4'b1110;
														assign node11479 = (inp[14]) ? node11483 : node11480;
															assign node11480 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node11483 = (inp[5]) ? 4'b1110 : 4'b1111;
													assign node11486 = (inp[14]) ? node11490 : node11487;
														assign node11487 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node11490 = (inp[5]) ? 4'b1111 : 4'b1011;
												assign node11493 = (inp[15]) ? node11503 : node11494;
													assign node11494 = (inp[5]) ? node11496 : 4'b1011;
														assign node11496 = (inp[9]) ? node11498 : 4'b1011;
															assign node11498 = (inp[14]) ? node11500 : 4'b1011;
																assign node11500 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node11503 = (inp[14]) ? node11507 : node11504;
														assign node11504 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11507 = (inp[5]) ? 4'b1011 : node11508;
															assign node11508 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node11512 = (inp[12]) ? node11632 : node11513;
										assign node11513 = (inp[5]) ? node11559 : node11514;
											assign node11514 = (inp[1]) ? node11540 : node11515;
												assign node11515 = (inp[2]) ? node11527 : node11516;
													assign node11516 = (inp[15]) ? node11522 : node11517;
														assign node11517 = (inp[11]) ? node11519 : 4'b1011;
															assign node11519 = (inp[14]) ? 4'b1011 : 4'b1010;
														assign node11522 = (inp[14]) ? 4'b1110 : node11523;
															assign node11523 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node11527 = (inp[15]) ? node11535 : node11528;
														assign node11528 = (inp[11]) ? node11532 : node11529;
															assign node11529 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node11532 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node11535 = (inp[14]) ? 4'b1010 : node11536;
															assign node11536 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node11540 = (inp[2]) ? node11550 : node11541;
													assign node11541 = (inp[14]) ? node11547 : node11542;
														assign node11542 = (inp[11]) ? node11544 : 4'b1111;
															assign node11544 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node11547 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node11550 = (inp[15]) ? node11552 : 4'b1011;
														assign node11552 = (inp[14]) ? node11556 : node11553;
															assign node11553 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node11556 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node11559 = (inp[11]) ? node11587 : node11560;
												assign node11560 = (inp[14]) ? node11574 : node11561;
													assign node11561 = (inp[2]) ? node11569 : node11562;
														assign node11562 = (inp[1]) ? node11566 : node11563;
															assign node11563 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node11566 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node11569 = (inp[1]) ? 4'b1111 : node11570;
															assign node11570 = (inp[15]) ? 4'b1010 : 4'b1111;
													assign node11574 = (inp[2]) ? node11580 : node11575;
														assign node11575 = (inp[15]) ? 4'b1110 : node11576;
															assign node11576 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node11580 = (inp[15]) ? node11584 : node11581;
															assign node11581 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node11584 = (inp[1]) ? 4'b1010 : 4'b1111;
												assign node11587 = (inp[14]) ? node11605 : node11588;
													assign node11588 = (inp[1]) ? node11596 : node11589;
														assign node11589 = (inp[2]) ? node11593 : node11590;
															assign node11590 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node11593 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node11596 = (inp[9]) ? 4'b1010 : node11597;
															assign node11597 = (inp[2]) ? node11601 : node11598;
																assign node11598 = (inp[15]) ? 4'b1010 : 4'b1110;
																assign node11601 = (inp[15]) ? 4'b1111 : 4'b1010;
													assign node11605 = (inp[9]) ? node11619 : node11606;
														assign node11606 = (inp[15]) ? node11612 : node11607;
															assign node11607 = (inp[2]) ? node11609 : 4'b1010;
																assign node11609 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node11612 = (inp[1]) ? node11616 : node11613;
																assign node11613 = (inp[2]) ? 4'b1110 : 4'b1011;
																assign node11616 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node11619 = (inp[1]) ? node11627 : node11620;
															assign node11620 = (inp[2]) ? node11624 : node11621;
																assign node11621 = (inp[15]) ? 4'b1011 : 4'b1111;
																assign node11624 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node11627 = (inp[2]) ? 4'b1111 : node11628;
																assign node11628 = (inp[15]) ? 4'b1111 : 4'b1010;
										assign node11632 = (inp[2]) ? node11682 : node11633;
											assign node11633 = (inp[1]) ? node11661 : node11634;
												assign node11634 = (inp[14]) ? node11646 : node11635;
													assign node11635 = (inp[5]) ? node11639 : node11636;
														assign node11636 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node11639 = (inp[11]) ? node11643 : node11640;
															assign node11640 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node11643 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node11646 = (inp[11]) ? node11652 : node11647;
														assign node11647 = (inp[5]) ? node11649 : 4'b1000;
															assign node11649 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node11652 = (inp[9]) ? node11654 : 4'b1001;
															assign node11654 = (inp[15]) ? node11658 : node11655;
																assign node11655 = (inp[5]) ? 4'b1100 : 4'b1001;
																assign node11658 = (inp[5]) ? 4'b1001 : 4'b1100;
												assign node11661 = (inp[5]) ? node11673 : node11662;
													assign node11662 = (inp[15]) ? node11666 : node11663;
														assign node11663 = (inp[14]) ? 4'b1101 : 4'b1001;
														assign node11666 = (inp[14]) ? node11670 : node11667;
															assign node11667 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node11670 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node11673 = (inp[15]) ? 4'b1101 : node11674;
														assign node11674 = (inp[14]) ? node11678 : node11675;
															assign node11675 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node11678 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node11682 = (inp[1]) ? node11712 : node11683;
												assign node11683 = (inp[14]) ? node11693 : node11684;
													assign node11684 = (inp[15]) ? node11688 : node11685;
														assign node11685 = (inp[5]) ? 4'b1100 : 4'b1001;
														assign node11688 = (inp[11]) ? node11690 : 4'b1100;
															assign node11690 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node11693 = (inp[11]) ? node11705 : node11694;
														assign node11694 = (inp[9]) ? node11700 : node11695;
															assign node11695 = (inp[5]) ? 4'b1000 : node11696;
																assign node11696 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node11700 = (inp[15]) ? node11702 : 4'b1101;
																assign node11702 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node11705 = (inp[5]) ? node11709 : node11706;
															assign node11706 = (inp[15]) ? 4'b1000 : 4'b1101;
															assign node11709 = (inp[15]) ? 4'b1101 : 4'b1000;
												assign node11712 = (inp[5]) ? node11722 : node11713;
													assign node11713 = (inp[15]) ? node11719 : node11714;
														assign node11714 = (inp[14]) ? node11716 : 4'b1100;
															assign node11716 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node11719 = (inp[14]) ? 4'b1100 : 4'b1000;
													assign node11722 = (inp[14]) ? node11728 : node11723;
														assign node11723 = (inp[15]) ? node11725 : 4'b1001;
															assign node11725 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node11728 = (inp[15]) ? 4'b1001 : 4'b1101;
							assign node11731 = (inp[13]) ? node12093 : node11732;
								assign node11732 = (inp[1]) ? node11882 : node11733;
									assign node11733 = (inp[2]) ? node11811 : node11734;
										assign node11734 = (inp[4]) ? node11762 : node11735;
											assign node11735 = (inp[12]) ? node11749 : node11736;
												assign node11736 = (inp[14]) ? node11738 : 4'b1000;
													assign node11738 = (inp[11]) ? node11744 : node11739;
														assign node11739 = (inp[5]) ? node11741 : 4'b1000;
															assign node11741 = (inp[15]) ? 4'b1000 : 4'b1100;
														assign node11744 = (inp[5]) ? node11746 : 4'b1001;
															assign node11746 = (inp[15]) ? 4'b1000 : 4'b1101;
												assign node11749 = (inp[14]) ? node11751 : 4'b1010;
													assign node11751 = (inp[11]) ? node11757 : node11752;
														assign node11752 = (inp[15]) ? node11754 : 4'b1010;
															assign node11754 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node11757 = (inp[5]) ? 4'b1010 : node11758;
															assign node11758 = (inp[15]) ? 4'b1111 : 4'b1011;
											assign node11762 = (inp[12]) ? node11786 : node11763;
												assign node11763 = (inp[5]) ? node11773 : node11764;
													assign node11764 = (inp[14]) ? node11766 : 4'b1010;
														assign node11766 = (inp[11]) ? node11770 : node11767;
															assign node11767 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node11770 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node11773 = (inp[15]) ? node11779 : node11774;
														assign node11774 = (inp[14]) ? 4'b1110 : node11775;
															assign node11775 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11779 = (inp[14]) ? node11783 : node11780;
															assign node11780 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node11783 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node11786 = (inp[5]) ? node11804 : node11787;
													assign node11787 = (inp[9]) ? node11797 : node11788;
														assign node11788 = (inp[11]) ? 4'b1100 : node11789;
															assign node11789 = (inp[14]) ? node11793 : node11790;
																assign node11790 = (inp[15]) ? 4'b1000 : 4'b1100;
																assign node11793 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node11797 = (inp[14]) ? node11801 : node11798;
															assign node11798 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node11801 = (inp[15]) ? 4'b1100 : 4'b1000;
													assign node11804 = (inp[15]) ? 4'b1001 : node11805;
														assign node11805 = (inp[14]) ? node11807 : 4'b1001;
															assign node11807 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node11811 = (inp[4]) ? node11835 : node11812;
											assign node11812 = (inp[12]) ? node11824 : node11813;
												assign node11813 = (inp[5]) ? node11815 : 4'b1100;
													assign node11815 = (inp[14]) ? node11817 : 4'b1100;
														assign node11817 = (inp[15]) ? node11821 : node11818;
															assign node11818 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node11821 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node11824 = (inp[14]) ? node11826 : 4'b1110;
													assign node11826 = (inp[15]) ? node11828 : 4'b1110;
														assign node11828 = (inp[11]) ? node11832 : node11829;
															assign node11829 = (inp[5]) ? 4'b1111 : 4'b1011;
															assign node11832 = (inp[5]) ? 4'b1110 : 4'b1010;
											assign node11835 = (inp[12]) ? node11853 : node11836;
												assign node11836 = (inp[5]) ? node11844 : node11837;
													assign node11837 = (inp[15]) ? node11839 : 4'b1111;
														assign node11839 = (inp[14]) ? node11841 : 4'b1111;
															assign node11841 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node11844 = (inp[15]) ? node11850 : node11845;
														assign node11845 = (inp[14]) ? 4'b1010 : node11846;
															assign node11846 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node11850 = (inp[14]) ? 4'b1110 : 4'b1010;
												assign node11853 = (inp[11]) ? node11871 : node11854;
													assign node11854 = (inp[15]) ? node11864 : node11855;
														assign node11855 = (inp[9]) ? 4'b1001 : node11856;
															assign node11856 = (inp[14]) ? node11860 : node11857;
																assign node11857 = (inp[5]) ? 4'b1100 : 4'b1001;
																assign node11860 = (inp[5]) ? 4'b1001 : 4'b1100;
														assign node11864 = (inp[5]) ? node11868 : node11865;
															assign node11865 = (inp[14]) ? 4'b1000 : 4'b1101;
															assign node11868 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node11871 = (inp[5]) ? node11877 : node11872;
														assign node11872 = (inp[15]) ? 4'b1000 : node11873;
															assign node11873 = (inp[14]) ? 4'b1101 : 4'b1000;
														assign node11877 = (inp[14]) ? node11879 : 4'b1100;
															assign node11879 = (inp[15]) ? 4'b1100 : 4'b1000;
									assign node11882 = (inp[2]) ? node11974 : node11883;
										assign node11883 = (inp[4]) ? node11925 : node11884;
											assign node11884 = (inp[12]) ? node11904 : node11885;
												assign node11885 = (inp[15]) ? node11893 : node11886;
													assign node11886 = (inp[14]) ? node11888 : 4'b1100;
														assign node11888 = (inp[5]) ? 4'b1000 : node11889;
															assign node11889 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node11893 = (inp[5]) ? node11899 : node11894;
														assign node11894 = (inp[11]) ? node11896 : 4'b1100;
															assign node11896 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node11899 = (inp[14]) ? node11901 : 4'b1100;
															assign node11901 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node11904 = (inp[15]) ? node11912 : node11905;
													assign node11905 = (inp[14]) ? node11907 : 4'b1111;
														assign node11907 = (inp[11]) ? node11909 : 4'b1111;
															assign node11909 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node11912 = (inp[5]) ? node11918 : node11913;
														assign node11913 = (inp[14]) ? node11915 : 4'b1111;
															assign node11915 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node11918 = (inp[14]) ? node11922 : node11919;
															assign node11919 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node11922 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node11925 = (inp[12]) ? node11953 : node11926;
												assign node11926 = (inp[15]) ? node11940 : node11927;
													assign node11927 = (inp[5]) ? node11933 : node11928;
														assign node11928 = (inp[14]) ? node11930 : 4'b1110;
															assign node11930 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node11933 = (inp[14]) ? node11937 : node11934;
															assign node11934 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node11937 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node11940 = (inp[14]) ? node11948 : node11941;
														assign node11941 = (inp[5]) ? node11945 : node11942;
															assign node11942 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node11945 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node11948 = (inp[5]) ? 4'b1111 : node11949;
															assign node11949 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node11953 = (inp[5]) ? node11963 : node11954;
													assign node11954 = (inp[15]) ? node11960 : node11955;
														assign node11955 = (inp[14]) ? 4'b1101 : node11956;
															assign node11956 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node11960 = (inp[14]) ? 4'b1000 : 4'b1100;
													assign node11963 = (inp[15]) ? node11967 : node11964;
														assign node11964 = (inp[14]) ? 4'b1000 : 4'b1100;
														assign node11967 = (inp[14]) ? node11971 : node11968;
															assign node11968 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node11971 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node11974 = (inp[14]) ? node12012 : node11975;
											assign node11975 = (inp[4]) ? node11987 : node11976;
												assign node11976 = (inp[12]) ? node11982 : node11977;
													assign node11977 = (inp[11]) ? 4'b1001 : node11978;
														assign node11978 = (inp[15]) ? 4'b1001 : 4'b1000;
													assign node11982 = (inp[15]) ? 4'b1010 : node11983;
														assign node11983 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node11987 = (inp[12]) ? node11999 : node11988;
													assign node11988 = (inp[5]) ? node11994 : node11989;
														assign node11989 = (inp[15]) ? 4'b1010 : node11990;
															assign node11990 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node11994 = (inp[15]) ? node11996 : 4'b1010;
															assign node11996 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node11999 = (inp[15]) ? node12007 : node12000;
														assign node12000 = (inp[5]) ? node12004 : node12001;
															assign node12001 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node12004 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node12007 = (inp[11]) ? 4'b1000 : node12008;
															assign node12008 = (inp[5]) ? 4'b1000 : 4'b1001;
											assign node12012 = (inp[9]) ? node12048 : node12013;
												assign node12013 = (inp[5]) ? node12029 : node12014;
													assign node12014 = (inp[15]) ? node12026 : node12015;
														assign node12015 = (inp[4]) ? node12023 : node12016;
															assign node12016 = (inp[12]) ? node12020 : node12017;
																assign node12017 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node12020 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node12023 = (inp[12]) ? 4'b1001 : 4'b1011;
														assign node12026 = (inp[4]) ? 4'b1110 : 4'b1001;
													assign node12029 = (inp[15]) ? node12039 : node12030;
														assign node12030 = (inp[12]) ? node12036 : node12031;
															assign node12031 = (inp[11]) ? node12033 : 4'b1101;
																assign node12033 = (inp[4]) ? 4'b1110 : 4'b1100;
															assign node12036 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node12039 = (inp[12]) ? node12043 : node12040;
															assign node12040 = (inp[4]) ? 4'b1011 : 4'b1001;
															assign node12043 = (inp[11]) ? 4'b1000 : node12044;
																assign node12044 = (inp[4]) ? 4'b1001 : 4'b1011;
												assign node12048 = (inp[4]) ? node12072 : node12049;
													assign node12049 = (inp[12]) ? node12061 : node12050;
														assign node12050 = (inp[15]) ? node12056 : node12051;
															assign node12051 = (inp[5]) ? node12053 : 4'b1000;
																assign node12053 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node12056 = (inp[5]) ? node12058 : 4'b1001;
																assign node12058 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node12061 = (inp[15]) ? node12067 : node12062;
															assign node12062 = (inp[5]) ? 4'b1010 : node12063;
																assign node12063 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node12067 = (inp[5]) ? node12069 : 4'b1110;
																assign node12069 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node12072 = (inp[12]) ? node12082 : node12073;
														assign node12073 = (inp[5]) ? node12079 : node12074;
															assign node12074 = (inp[15]) ? 4'b1110 : node12075;
																assign node12075 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node12079 = (inp[15]) ? 4'b1011 : 4'b1110;
														assign node12082 = (inp[11]) ? node12088 : node12083;
															assign node12083 = (inp[5]) ? 4'b1100 : node12084;
																assign node12084 = (inp[15]) ? 4'b1100 : 4'b1001;
															assign node12088 = (inp[5]) ? 4'b1101 : node12089;
																assign node12089 = (inp[15]) ? 4'b1101 : 4'b1001;
								assign node12093 = (inp[4]) ? node12239 : node12094;
									assign node12094 = (inp[12]) ? node12168 : node12095;
										assign node12095 = (inp[2]) ? node12131 : node12096;
											assign node12096 = (inp[1]) ? node12114 : node12097;
												assign node12097 = (inp[15]) ? node12105 : node12098;
													assign node12098 = (inp[5]) ? node12100 : 4'b1000;
														assign node12100 = (inp[14]) ? 4'b1100 : node12101;
															assign node12101 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node12105 = (inp[14]) ? node12109 : node12106;
														assign node12106 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node12109 = (inp[11]) ? 4'b1001 : node12110;
															assign node12110 = (inp[5]) ? 4'b1000 : 4'b1001;
												assign node12114 = (inp[15]) ? node12124 : node12115;
													assign node12115 = (inp[14]) ? node12119 : node12116;
														assign node12116 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node12119 = (inp[5]) ? node12121 : 4'b1100;
															assign node12121 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node12124 = (inp[11]) ? node12126 : 4'b1100;
														assign node12126 = (inp[5]) ? 4'b1100 : node12127;
															assign node12127 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node12131 = (inp[1]) ? node12149 : node12132;
												assign node12132 = (inp[15]) ? node12140 : node12133;
													assign node12133 = (inp[14]) ? node12137 : node12134;
														assign node12134 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node12137 = (inp[5]) ? 4'b1001 : 4'b1100;
													assign node12140 = (inp[11]) ? node12144 : node12141;
														assign node12141 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node12144 = (inp[14]) ? node12146 : 4'b1100;
															assign node12146 = (inp[5]) ? 4'b1100 : 4'b1101;
												assign node12149 = (inp[15]) ? node12155 : node12150;
													assign node12150 = (inp[5]) ? node12152 : 4'b1001;
														assign node12152 = (inp[14]) ? 4'b1101 : 4'b1001;
													assign node12155 = (inp[5]) ? node12163 : node12156;
														assign node12156 = (inp[11]) ? node12160 : node12157;
															assign node12157 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node12160 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node12163 = (inp[11]) ? 4'b1001 : node12164;
															assign node12164 = (inp[14]) ? 4'b1001 : 4'b1000;
										assign node12168 = (inp[2]) ? node12204 : node12169;
											assign node12169 = (inp[1]) ? node12189 : node12170;
												assign node12170 = (inp[14]) ? node12178 : node12171;
													assign node12171 = (inp[11]) ? node12175 : node12172;
														assign node12172 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node12175 = (inp[15]) ? 4'b1010 : 4'b1011;
													assign node12178 = (inp[5]) ? node12182 : node12179;
														assign node12179 = (inp[15]) ? 4'b1111 : 4'b1010;
														assign node12182 = (inp[15]) ? node12186 : node12183;
															assign node12183 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node12186 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node12189 = (inp[15]) ? node12199 : node12190;
													assign node12190 = (inp[11]) ? node12196 : node12191;
														assign node12191 = (inp[14]) ? node12193 : 4'b1111;
															assign node12193 = (inp[5]) ? 4'b1110 : 4'b1111;
														assign node12196 = (inp[14]) ? 4'b1111 : 4'b1110;
													assign node12199 = (inp[5]) ? 4'b1111 : node12200;
														assign node12200 = (inp[14]) ? 4'b1011 : 4'b1111;
											assign node12204 = (inp[1]) ? node12222 : node12205;
												assign node12205 = (inp[15]) ? node12215 : node12206;
													assign node12206 = (inp[14]) ? node12210 : node12207;
														assign node12207 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12210 = (inp[11]) ? node12212 : 4'b1111;
															assign node12212 = (inp[5]) ? 4'b1111 : 4'b1110;
													assign node12215 = (inp[14]) ? node12219 : node12216;
														assign node12216 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12219 = (inp[5]) ? 4'b1110 : 4'b1010;
												assign node12222 = (inp[15]) ? node12230 : node12223;
													assign node12223 = (inp[14]) ? node12225 : 4'b1010;
														assign node12225 = (inp[11]) ? 4'b1010 : node12226;
															assign node12226 = (inp[5]) ? 4'b1011 : 4'b1010;
													assign node12230 = (inp[14]) ? node12234 : node12231;
														assign node12231 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node12234 = (inp[5]) ? 4'b1010 : node12235;
															assign node12235 = (inp[11]) ? 4'b1111 : 4'b1110;
									assign node12239 = (inp[12]) ? node12337 : node12240;
										assign node12240 = (inp[5]) ? node12292 : node12241;
											assign node12241 = (inp[1]) ? node12273 : node12242;
												assign node12242 = (inp[2]) ? node12252 : node12243;
													assign node12243 = (inp[15]) ? node12247 : node12244;
														assign node12244 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12247 = (inp[14]) ? 4'b1111 : node12248;
															assign node12248 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node12252 = (inp[14]) ? node12268 : node12253;
														assign node12253 = (inp[9]) ? node12261 : node12254;
															assign node12254 = (inp[15]) ? node12258 : node12255;
																assign node12255 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node12258 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node12261 = (inp[15]) ? node12265 : node12262;
																assign node12262 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node12265 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12268 = (inp[15]) ? 4'b1011 : node12269;
															assign node12269 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node12273 = (inp[2]) ? node12283 : node12274;
													assign node12274 = (inp[14]) ? node12280 : node12275;
														assign node12275 = (inp[15]) ? 4'b1110 : node12276;
															assign node12276 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node12280 = (inp[15]) ? 4'b1010 : 4'b1110;
													assign node12283 = (inp[15]) ? node12285 : 4'b1010;
														assign node12285 = (inp[14]) ? node12289 : node12286;
															assign node12286 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node12289 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node12292 = (inp[1]) ? node12316 : node12293;
												assign node12293 = (inp[15]) ? node12305 : node12294;
													assign node12294 = (inp[2]) ? node12300 : node12295;
														assign node12295 = (inp[14]) ? node12297 : 4'b1011;
															assign node12297 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12300 = (inp[14]) ? node12302 : 4'b1110;
															assign node12302 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node12305 = (inp[2]) ? node12309 : node12306;
														assign node12306 = (inp[14]) ? 4'b1010 : 4'b1110;
														assign node12309 = (inp[14]) ? node12313 : node12310;
															assign node12310 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node12313 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node12316 = (inp[2]) ? node12326 : node12317;
													assign node12317 = (inp[14]) ? node12321 : node12318;
														assign node12318 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node12321 = (inp[15]) ? node12323 : 4'b1011;
															assign node12323 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node12326 = (inp[14]) ? node12332 : node12327;
														assign node12327 = (inp[15]) ? 4'b1110 : node12328;
															assign node12328 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12332 = (inp[11]) ? 4'b1010 : node12333;
															assign node12333 = (inp[15]) ? 4'b1011 : 4'b1111;
										assign node12337 = (inp[5]) ? node12385 : node12338;
											assign node12338 = (inp[2]) ? node12366 : node12339;
												assign node12339 = (inp[11]) ? node12353 : node12340;
													assign node12340 = (inp[1]) ? node12346 : node12341;
														assign node12341 = (inp[15]) ? node12343 : 4'b1001;
															assign node12343 = (inp[14]) ? 4'b1100 : 4'b1000;
														assign node12346 = (inp[15]) ? node12350 : node12347;
															assign node12347 = (inp[14]) ? 4'b1100 : 4'b1000;
															assign node12350 = (inp[14]) ? 4'b1000 : 4'b1101;
													assign node12353 = (inp[14]) ? node12361 : node12354;
														assign node12354 = (inp[1]) ? node12358 : node12355;
															assign node12355 = (inp[15]) ? 4'b1000 : 4'b1101;
															assign node12358 = (inp[15]) ? 4'b1100 : 4'b1000;
														assign node12361 = (inp[1]) ? node12363 : 4'b1000;
															assign node12363 = (inp[15]) ? 4'b1001 : 4'b1101;
												assign node12366 = (inp[1]) ? node12376 : node12367;
													assign node12367 = (inp[15]) ? node12371 : node12368;
														assign node12368 = (inp[14]) ? 4'b1100 : 4'b1000;
														assign node12371 = (inp[14]) ? node12373 : 4'b1101;
															assign node12373 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node12376 = (inp[15]) ? node12382 : node12377;
														assign node12377 = (inp[14]) ? node12379 : 4'b1101;
															assign node12379 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node12382 = (inp[14]) ? 4'b1101 : 4'b1001;
											assign node12385 = (inp[11]) ? node12415 : node12386;
												assign node12386 = (inp[1]) ? node12402 : node12387;
													assign node12387 = (inp[2]) ? node12395 : node12388;
														assign node12388 = (inp[14]) ? node12392 : node12389;
															assign node12389 = (inp[15]) ? 4'b1000 : 4'b1001;
															assign node12392 = (inp[15]) ? 4'b1001 : 4'b1101;
														assign node12395 = (inp[14]) ? node12399 : node12396;
															assign node12396 = (inp[15]) ? 4'b1101 : 4'b1100;
															assign node12399 = (inp[15]) ? 4'b1100 : 4'b1001;
													assign node12402 = (inp[15]) ? node12410 : node12403;
														assign node12403 = (inp[2]) ? node12407 : node12404;
															assign node12404 = (inp[14]) ? 4'b1001 : 4'b1100;
															assign node12407 = (inp[14]) ? 4'b1100 : 4'b1000;
														assign node12410 = (inp[14]) ? node12412 : 4'b1001;
															assign node12412 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node12415 = (inp[2]) ? node12431 : node12416;
													assign node12416 = (inp[1]) ? node12424 : node12417;
														assign node12417 = (inp[14]) ? node12421 : node12418;
															assign node12418 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node12421 = (inp[15]) ? 4'b1000 : 4'b1101;
														assign node12424 = (inp[14]) ? node12428 : node12425;
															assign node12425 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node12428 = (inp[15]) ? 4'b1100 : 4'b1000;
													assign node12431 = (inp[1]) ? node12433 : 4'b1100;
														assign node12433 = (inp[15]) ? 4'b1000 : node12434;
															assign node12434 = (inp[14]) ? 4'b1100 : 4'b1000;
					assign node12438 = (inp[5]) ? node14686 : node12439;
						assign node12439 = (inp[13]) ? node13727 : node12440;
							assign node12440 = (inp[9]) ? node13080 : node12441;
								assign node12441 = (inp[2]) ? node12751 : node12442;
									assign node12442 = (inp[1]) ? node12608 : node12443;
										assign node12443 = (inp[15]) ? node12529 : node12444;
											assign node12444 = (inp[14]) ? node12490 : node12445;
												assign node12445 = (inp[12]) ? node12465 : node12446;
													assign node12446 = (inp[4]) ? node12454 : node12447;
														assign node12447 = (inp[0]) ? node12451 : node12448;
															assign node12448 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node12451 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node12454 = (inp[11]) ? node12460 : node12455;
															assign node12455 = (inp[10]) ? node12457 : 4'b1011;
																assign node12457 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node12460 = (inp[0]) ? node12462 : 4'b1010;
																assign node12462 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node12465 = (inp[4]) ? node12481 : node12466;
														assign node12466 = (inp[10]) ? node12474 : node12467;
															assign node12467 = (inp[0]) ? node12471 : node12468;
																assign node12468 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node12471 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node12474 = (inp[0]) ? node12478 : node12475;
																assign node12475 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node12478 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12481 = (inp[11]) ? node12485 : node12482;
															assign node12482 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node12485 = (inp[0]) ? 4'b1000 : node12486;
																assign node12486 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node12490 = (inp[4]) ? node12508 : node12491;
													assign node12491 = (inp[12]) ? node12501 : node12492;
														assign node12492 = (inp[0]) ? node12494 : 4'b1001;
															assign node12494 = (inp[10]) ? node12498 : node12495;
																assign node12495 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node12498 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node12501 = (inp[0]) ? node12505 : node12502;
															assign node12502 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node12505 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node12508 = (inp[12]) ? node12520 : node12509;
														assign node12509 = (inp[10]) ? node12515 : node12510;
															assign node12510 = (inp[11]) ? 4'b1010 : node12511;
																assign node12511 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node12515 = (inp[11]) ? 4'b1011 : node12516;
																assign node12516 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node12520 = (inp[0]) ? node12522 : 4'b1001;
															assign node12522 = (inp[10]) ? node12526 : node12523;
																assign node12523 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node12526 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node12529 = (inp[14]) ? node12561 : node12530;
												assign node12530 = (inp[4]) ? node12546 : node12531;
													assign node12531 = (inp[12]) ? node12539 : node12532;
														assign node12532 = (inp[0]) ? node12536 : node12533;
															assign node12533 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node12536 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node12539 = (inp[10]) ? 4'b1110 : node12540;
															assign node12540 = (inp[0]) ? node12542 : 4'b1111;
																assign node12542 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node12546 = (inp[12]) ? node12556 : node12547;
														assign node12547 = (inp[0]) ? 4'b1011 : node12548;
															assign node12548 = (inp[11]) ? node12552 : node12549;
																assign node12549 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node12552 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node12556 = (inp[10]) ? 4'b1101 : node12557;
															assign node12557 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node12561 = (inp[12]) ? node12585 : node12562;
													assign node12562 = (inp[4]) ? node12574 : node12563;
														assign node12563 = (inp[11]) ? node12569 : node12564;
															assign node12564 = (inp[10]) ? node12566 : 4'b1000;
																assign node12566 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node12569 = (inp[0]) ? node12571 : 4'b1000;
																assign node12571 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node12574 = (inp[11]) ? node12580 : node12575;
															assign node12575 = (inp[0]) ? 4'b1010 : node12576;
																assign node12576 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node12580 = (inp[0]) ? 4'b1011 : node12581;
																assign node12581 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node12585 = (inp[4]) ? node12595 : node12586;
														assign node12586 = (inp[0]) ? node12588 : 4'b1011;
															assign node12588 = (inp[11]) ? node12592 : node12589;
																assign node12589 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node12592 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node12595 = (inp[11]) ? node12603 : node12596;
															assign node12596 = (inp[10]) ? node12600 : node12597;
																assign node12597 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node12600 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node12603 = (inp[10]) ? node12605 : 4'b1001;
																assign node12605 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node12608 = (inp[15]) ? node12680 : node12609;
											assign node12609 = (inp[12]) ? node12645 : node12610;
												assign node12610 = (inp[4]) ? node12630 : node12611;
													assign node12611 = (inp[10]) ? node12621 : node12612;
														assign node12612 = (inp[0]) ? node12618 : node12613;
															assign node12613 = (inp[14]) ? node12615 : 4'b1100;
																assign node12615 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node12618 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node12621 = (inp[0]) ? node12625 : node12622;
															assign node12622 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node12625 = (inp[11]) ? node12627 : 4'b1100;
																assign node12627 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node12630 = (inp[0]) ? node12636 : node12631;
														assign node12631 = (inp[10]) ? node12633 : 4'b1110;
															assign node12633 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node12636 = (inp[10]) ? node12642 : node12637;
															assign node12637 = (inp[11]) ? node12639 : 4'b1111;
																assign node12639 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node12642 = (inp[14]) ? 4'b1111 : 4'b1110;
												assign node12645 = (inp[4]) ? node12665 : node12646;
													assign node12646 = (inp[14]) ? node12658 : node12647;
														assign node12647 = (inp[11]) ? node12653 : node12648;
															assign node12648 = (inp[10]) ? 4'b1110 : node12649;
																assign node12649 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node12653 = (inp[0]) ? 4'b1111 : node12654;
																assign node12654 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node12658 = (inp[11]) ? 4'b1010 : node12659;
															assign node12659 = (inp[10]) ? 4'b1011 : node12660;
																assign node12660 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node12665 = (inp[0]) ? node12673 : node12666;
														assign node12666 = (inp[10]) ? node12668 : 4'b1100;
															assign node12668 = (inp[11]) ? node12670 : 4'b1101;
																assign node12670 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node12673 = (inp[10]) ? node12675 : 4'b1101;
															assign node12675 = (inp[11]) ? node12677 : 4'b1100;
																assign node12677 = (inp[14]) ? 4'b1101 : 4'b1100;
											assign node12680 = (inp[14]) ? node12714 : node12681;
												assign node12681 = (inp[4]) ? node12701 : node12682;
													assign node12682 = (inp[12]) ? node12690 : node12683;
														assign node12683 = (inp[10]) ? node12687 : node12684;
															assign node12684 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node12687 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node12690 = (inp[11]) ? node12696 : node12691;
															assign node12691 = (inp[0]) ? node12693 : 4'b1010;
																assign node12693 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node12696 = (inp[0]) ? node12698 : 4'b1011;
																assign node12698 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node12701 = (inp[12]) ? node12707 : node12702;
														assign node12702 = (inp[0]) ? 4'b1111 : node12703;
															assign node12703 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node12707 = (inp[0]) ? node12711 : node12708;
															assign node12708 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node12711 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node12714 = (inp[4]) ? node12736 : node12715;
													assign node12715 = (inp[12]) ? node12731 : node12716;
														assign node12716 = (inp[0]) ? node12724 : node12717;
															assign node12717 = (inp[11]) ? node12721 : node12718;
																assign node12718 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node12721 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node12724 = (inp[11]) ? node12728 : node12725;
																assign node12725 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node12728 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node12731 = (inp[0]) ? 4'b1110 : node12732;
															assign node12732 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node12736 = (inp[12]) ? node12744 : node12737;
														assign node12737 = (inp[10]) ? 4'b1111 : node12738;
															assign node12738 = (inp[11]) ? 4'b1111 : node12739;
																assign node12739 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node12744 = (inp[0]) ? node12746 : 4'b1101;
															assign node12746 = (inp[10]) ? 4'b1100 : node12747;
																assign node12747 = (inp[11]) ? 4'b1101 : 4'b1100;
									assign node12751 = (inp[1]) ? node12921 : node12752;
										assign node12752 = (inp[12]) ? node12832 : node12753;
											assign node12753 = (inp[4]) ? node12791 : node12754;
												assign node12754 = (inp[14]) ? node12770 : node12755;
													assign node12755 = (inp[15]) ? node12763 : node12756;
														assign node12756 = (inp[0]) ? node12760 : node12757;
															assign node12757 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node12760 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node12763 = (inp[11]) ? node12765 : 4'b1000;
															assign node12765 = (inp[10]) ? node12767 : 4'b1001;
																assign node12767 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node12770 = (inp[10]) ? node12780 : node12771;
														assign node12771 = (inp[0]) ? node12775 : node12772;
															assign node12772 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node12775 = (inp[11]) ? 4'b1101 : node12776;
																assign node12776 = (inp[15]) ? 4'b1100 : 4'b1101;
														assign node12780 = (inp[0]) ? node12786 : node12781;
															assign node12781 = (inp[11]) ? 4'b1101 : node12782;
																assign node12782 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node12786 = (inp[15]) ? node12788 : 4'b1100;
																assign node12788 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node12791 = (inp[15]) ? node12807 : node12792;
													assign node12792 = (inp[14]) ? node12800 : node12793;
														assign node12793 = (inp[0]) ? node12797 : node12794;
															assign node12794 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node12797 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node12800 = (inp[10]) ? node12804 : node12801;
															assign node12801 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node12804 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node12807 = (inp[11]) ? node12817 : node12808;
														assign node12808 = (inp[10]) ? node12810 : 4'b1110;
															assign node12810 = (inp[0]) ? node12814 : node12811;
																assign node12811 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node12814 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node12817 = (inp[10]) ? node12825 : node12818;
															assign node12818 = (inp[14]) ? node12822 : node12819;
																assign node12819 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node12822 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node12825 = (inp[14]) ? node12829 : node12826;
																assign node12826 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node12829 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node12832 = (inp[4]) ? node12876 : node12833;
												assign node12833 = (inp[11]) ? node12851 : node12834;
													assign node12834 = (inp[0]) ? node12840 : node12835;
														assign node12835 = (inp[10]) ? 4'b1010 : node12836;
															assign node12836 = (inp[15]) ? 4'b1011 : 4'b1110;
														assign node12840 = (inp[10]) ? node12846 : node12841;
															assign node12841 = (inp[14]) ? node12843 : 4'b1010;
																assign node12843 = (inp[15]) ? 4'b1110 : 4'b1010;
															assign node12846 = (inp[14]) ? node12848 : 4'b1110;
																assign node12848 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node12851 = (inp[15]) ? node12865 : node12852;
														assign node12852 = (inp[14]) ? node12860 : node12853;
															assign node12853 = (inp[10]) ? node12857 : node12854;
																assign node12854 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node12857 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node12860 = (inp[0]) ? 4'b1010 : node12861;
																assign node12861 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node12865 = (inp[14]) ? node12871 : node12866;
															assign node12866 = (inp[0]) ? node12868 : 4'b1010;
																assign node12868 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node12871 = (inp[0]) ? 4'b1110 : node12872;
																assign node12872 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node12876 = (inp[14]) ? node12898 : node12877;
													assign node12877 = (inp[15]) ? node12885 : node12878;
														assign node12878 = (inp[11]) ? node12880 : 4'b1100;
															assign node12880 = (inp[10]) ? 4'b1101 : node12881;
																assign node12881 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node12885 = (inp[11]) ? node12891 : node12886;
															assign node12886 = (inp[0]) ? node12888 : 4'b1001;
																assign node12888 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node12891 = (inp[0]) ? node12895 : node12892;
																assign node12892 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node12895 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node12898 = (inp[15]) ? node12906 : node12899;
														assign node12899 = (inp[0]) ? node12903 : node12900;
															assign node12900 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node12903 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node12906 = (inp[10]) ? node12914 : node12907;
															assign node12907 = (inp[11]) ? node12911 : node12908;
																assign node12908 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node12911 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node12914 = (inp[0]) ? node12918 : node12915;
																assign node12915 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node12918 = (inp[11]) ? 4'b1100 : 4'b1101;
										assign node12921 = (inp[12]) ? node12999 : node12922;
											assign node12922 = (inp[4]) ? node12956 : node12923;
												assign node12923 = (inp[15]) ? node12937 : node12924;
													assign node12924 = (inp[11]) ? node12926 : 4'b1000;
														assign node12926 = (inp[10]) ? node12932 : node12927;
															assign node12927 = (inp[0]) ? node12929 : 4'b1001;
																assign node12929 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node12932 = (inp[0]) ? node12934 : 4'b1000;
																assign node12934 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node12937 = (inp[14]) ? node12941 : node12938;
														assign node12938 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node12941 = (inp[10]) ? node12949 : node12942;
															assign node12942 = (inp[11]) ? node12946 : node12943;
																assign node12943 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node12946 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node12949 = (inp[0]) ? node12953 : node12950;
																assign node12950 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node12953 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node12956 = (inp[14]) ? node12980 : node12957;
													assign node12957 = (inp[0]) ? node12965 : node12958;
														assign node12958 = (inp[10]) ? 4'b1010 : node12959;
															assign node12959 = (inp[15]) ? node12961 : 4'b1010;
																assign node12961 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node12965 = (inp[10]) ? node12973 : node12966;
															assign node12966 = (inp[15]) ? node12970 : node12967;
																assign node12967 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node12970 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node12973 = (inp[11]) ? node12977 : node12974;
																assign node12974 = (inp[15]) ? 4'b1010 : 4'b1011;
																assign node12977 = (inp[15]) ? 4'b1011 : 4'b1010;
													assign node12980 = (inp[11]) ? node12992 : node12981;
														assign node12981 = (inp[0]) ? node12987 : node12982;
															assign node12982 = (inp[15]) ? node12984 : 4'b1011;
																assign node12984 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node12987 = (inp[15]) ? node12989 : 4'b1010;
																assign node12989 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node12992 = (inp[15]) ? 4'b1011 : node12993;
															assign node12993 = (inp[10]) ? node12995 : 4'b1011;
																assign node12995 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node12999 = (inp[4]) ? node13035 : node13000;
												assign node13000 = (inp[10]) ? node13020 : node13001;
													assign node13001 = (inp[0]) ? node13011 : node13002;
														assign node13002 = (inp[15]) ? node13006 : node13003;
															assign node13003 = (inp[14]) ? 4'b1110 : 4'b1010;
															assign node13006 = (inp[14]) ? 4'b1011 : node13007;
																assign node13007 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node13011 = (inp[15]) ? node13015 : node13012;
															assign node13012 = (inp[14]) ? 4'b1111 : 4'b1011;
															assign node13015 = (inp[14]) ? 4'b1010 : node13016;
																assign node13016 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node13020 = (inp[0]) ? node13028 : node13021;
														assign node13021 = (inp[14]) ? node13025 : node13022;
															assign node13022 = (inp[15]) ? 4'b1111 : 4'b1011;
															assign node13025 = (inp[15]) ? 4'b1010 : 4'b1111;
														assign node13028 = (inp[15]) ? node13032 : node13029;
															assign node13029 = (inp[14]) ? 4'b1110 : 4'b1010;
															assign node13032 = (inp[14]) ? 4'b1011 : 4'b1110;
												assign node13035 = (inp[15]) ? node13059 : node13036;
													assign node13036 = (inp[10]) ? node13052 : node13037;
														assign node13037 = (inp[0]) ? node13045 : node13038;
															assign node13038 = (inp[11]) ? node13042 : node13039;
																assign node13039 = (inp[14]) ? 4'b1000 : 4'b1001;
																assign node13042 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node13045 = (inp[14]) ? node13049 : node13046;
																assign node13046 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node13049 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node13052 = (inp[14]) ? 4'b1000 : node13053;
															assign node13053 = (inp[0]) ? node13055 : 4'b1000;
																assign node13055 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node13059 = (inp[14]) ? node13071 : node13060;
														assign node13060 = (inp[11]) ? node13066 : node13061;
															assign node13061 = (inp[10]) ? node13063 : 4'b1100;
																assign node13063 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node13066 = (inp[0]) ? 4'b1101 : node13067;
																assign node13067 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node13071 = (inp[0]) ? node13073 : 4'b1000;
															assign node13073 = (inp[10]) ? node13077 : node13074;
																assign node13074 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node13077 = (inp[11]) ? 4'b1000 : 4'b1001;
								assign node13080 = (inp[2]) ? node13400 : node13081;
									assign node13081 = (inp[1]) ? node13231 : node13082;
										assign node13082 = (inp[4]) ? node13160 : node13083;
											assign node13083 = (inp[12]) ? node13115 : node13084;
												assign node13084 = (inp[14]) ? node13098 : node13085;
													assign node13085 = (inp[15]) ? node13093 : node13086;
														assign node13086 = (inp[11]) ? 4'b1001 : node13087;
															assign node13087 = (inp[0]) ? node13089 : 4'b1000;
																assign node13089 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node13093 = (inp[0]) ? node13095 : 4'b1101;
															assign node13095 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node13098 = (inp[15]) ? node13108 : node13099;
														assign node13099 = (inp[10]) ? 4'b1000 : node13100;
															assign node13100 = (inp[0]) ? node13104 : node13101;
																assign node13101 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node13104 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node13108 = (inp[10]) ? node13112 : node13109;
															assign node13109 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node13112 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node13115 = (inp[11]) ? node13141 : node13116;
													assign node13116 = (inp[14]) ? node13130 : node13117;
														assign node13117 = (inp[15]) ? node13125 : node13118;
															assign node13118 = (inp[0]) ? node13122 : node13119;
																assign node13119 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node13122 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node13125 = (inp[0]) ? 4'b1110 : node13126;
																assign node13126 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node13130 = (inp[15]) ? node13136 : node13131;
															assign node13131 = (inp[0]) ? 4'b1111 : node13132;
																assign node13132 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node13136 = (inp[10]) ? 4'b1011 : node13137;
																assign node13137 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node13141 = (inp[14]) ? node13151 : node13142;
														assign node13142 = (inp[15]) ? node13144 : 4'b1011;
															assign node13144 = (inp[10]) ? node13148 : node13145;
																assign node13145 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node13148 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node13151 = (inp[15]) ? 4'b1010 : node13152;
															assign node13152 = (inp[10]) ? node13156 : node13153;
																assign node13153 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node13156 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node13160 = (inp[12]) ? node13190 : node13161;
												assign node13161 = (inp[15]) ? node13177 : node13162;
													assign node13162 = (inp[0]) ? node13166 : node13163;
														assign node13163 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node13166 = (inp[10]) ? node13172 : node13167;
															assign node13167 = (inp[14]) ? node13169 : 4'b1011;
																assign node13169 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node13172 = (inp[14]) ? node13174 : 4'b1010;
																assign node13174 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node13177 = (inp[11]) ? node13185 : node13178;
														assign node13178 = (inp[10]) ? node13182 : node13179;
															assign node13179 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node13182 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node13185 = (inp[0]) ? 4'b1010 : node13186;
															assign node13186 = (inp[14]) ? 4'b1011 : 4'b1010;
												assign node13190 = (inp[14]) ? node13208 : node13191;
													assign node13191 = (inp[15]) ? node13199 : node13192;
														assign node13192 = (inp[11]) ? node13194 : 4'b1000;
															assign node13194 = (inp[0]) ? node13196 : 4'b1001;
																assign node13196 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node13199 = (inp[11]) ? node13203 : node13200;
															assign node13200 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node13203 = (inp[10]) ? node13205 : 4'b1100;
																assign node13205 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node13208 = (inp[10]) ? node13220 : node13209;
														assign node13209 = (inp[0]) ? node13215 : node13210;
															assign node13210 = (inp[11]) ? node13212 : 4'b1001;
																assign node13212 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node13215 = (inp[15]) ? 4'b1000 : node13216;
																assign node13216 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node13220 = (inp[0]) ? node13226 : node13221;
															assign node13221 = (inp[15]) ? 4'b1000 : node13222;
																assign node13222 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node13226 = (inp[15]) ? 4'b1001 : node13227;
																assign node13227 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node13231 = (inp[12]) ? node13313 : node13232;
											assign node13232 = (inp[4]) ? node13272 : node13233;
												assign node13233 = (inp[15]) ? node13249 : node13234;
													assign node13234 = (inp[11]) ? node13242 : node13235;
														assign node13235 = (inp[10]) ? node13239 : node13236;
															assign node13236 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node13239 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node13242 = (inp[0]) ? 4'b1100 : node13243;
															assign node13243 = (inp[10]) ? node13245 : 4'b1100;
																assign node13245 = (inp[14]) ? 4'b1100 : 4'b1101;
													assign node13249 = (inp[14]) ? node13259 : node13250;
														assign node13250 = (inp[11]) ? 4'b1000 : node13251;
															assign node13251 = (inp[0]) ? node13255 : node13252;
																assign node13252 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node13255 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node13259 = (inp[10]) ? node13265 : node13260;
															assign node13260 = (inp[11]) ? 4'b1101 : node13261;
																assign node13261 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node13265 = (inp[11]) ? node13269 : node13266;
																assign node13266 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node13269 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node13272 = (inp[11]) ? node13288 : node13273;
													assign node13273 = (inp[0]) ? node13281 : node13274;
														assign node13274 = (inp[15]) ? node13278 : node13275;
															assign node13275 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node13278 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node13281 = (inp[10]) ? node13285 : node13282;
															assign node13282 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node13285 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node13288 = (inp[15]) ? node13298 : node13289;
														assign node13289 = (inp[10]) ? 4'b1110 : node13290;
															assign node13290 = (inp[14]) ? node13294 : node13291;
																assign node13291 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node13294 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node13298 = (inp[0]) ? node13306 : node13299;
															assign node13299 = (inp[10]) ? node13303 : node13300;
																assign node13300 = (inp[14]) ? 4'b1110 : 4'b1111;
																assign node13303 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node13306 = (inp[10]) ? node13310 : node13307;
																assign node13307 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node13310 = (inp[14]) ? 4'b1110 : 4'b1111;
											assign node13313 = (inp[4]) ? node13361 : node13314;
												assign node13314 = (inp[0]) ? node13336 : node13315;
													assign node13315 = (inp[10]) ? node13325 : node13316;
														assign node13316 = (inp[15]) ? node13322 : node13317;
															assign node13317 = (inp[14]) ? node13319 : 4'b1110;
																assign node13319 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node13322 = (inp[14]) ? 4'b1110 : 4'b1010;
														assign node13325 = (inp[14]) ? node13331 : node13326;
															assign node13326 = (inp[15]) ? 4'b1010 : node13327;
																assign node13327 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node13331 = (inp[15]) ? 4'b1111 : node13332;
																assign node13332 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node13336 = (inp[10]) ? node13348 : node13337;
														assign node13337 = (inp[15]) ? node13345 : node13338;
															assign node13338 = (inp[14]) ? node13342 : node13339;
																assign node13339 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node13342 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node13345 = (inp[14]) ? 4'b1111 : 4'b1011;
														assign node13348 = (inp[15]) ? node13356 : node13349;
															assign node13349 = (inp[14]) ? node13353 : node13350;
																assign node13350 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node13353 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node13356 = (inp[14]) ? 4'b1110 : node13357;
																assign node13357 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node13361 = (inp[14]) ? node13375 : node13362;
													assign node13362 = (inp[15]) ? node13368 : node13363;
														assign node13363 = (inp[10]) ? 4'b1100 : node13364;
															assign node13364 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node13368 = (inp[0]) ? node13372 : node13369;
															assign node13369 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node13372 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node13375 = (inp[15]) ? node13391 : node13376;
														assign node13376 = (inp[10]) ? node13384 : node13377;
															assign node13377 = (inp[11]) ? node13381 : node13378;
																assign node13378 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node13381 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node13384 = (inp[11]) ? node13388 : node13385;
																assign node13385 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node13388 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node13391 = (inp[11]) ? 4'b1100 : node13392;
															assign node13392 = (inp[0]) ? node13396 : node13393;
																assign node13393 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node13396 = (inp[10]) ? 4'b1101 : 4'b1100;
									assign node13400 = (inp[1]) ? node13556 : node13401;
										assign node13401 = (inp[15]) ? node13461 : node13402;
											assign node13402 = (inp[12]) ? node13426 : node13403;
												assign node13403 = (inp[4]) ? node13419 : node13404;
													assign node13404 = (inp[11]) ? node13412 : node13405;
														assign node13405 = (inp[10]) ? node13409 : node13406;
															assign node13406 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node13409 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node13412 = (inp[10]) ? node13416 : node13413;
															assign node13413 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node13416 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node13419 = (inp[10]) ? node13423 : node13420;
														assign node13420 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node13423 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node13426 = (inp[4]) ? node13446 : node13427;
													assign node13427 = (inp[14]) ? node13441 : node13428;
														assign node13428 = (inp[11]) ? node13436 : node13429;
															assign node13429 = (inp[10]) ? node13433 : node13430;
																assign node13430 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node13433 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node13436 = (inp[0]) ? 4'b1111 : node13437;
																assign node13437 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node13441 = (inp[0]) ? 4'b1011 : node13442;
															assign node13442 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node13446 = (inp[14]) ? node13454 : node13447;
														assign node13447 = (inp[10]) ? node13451 : node13448;
															assign node13448 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node13451 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node13454 = (inp[0]) ? node13458 : node13455;
															assign node13455 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node13458 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node13461 = (inp[14]) ? node13509 : node13462;
												assign node13462 = (inp[4]) ? node13484 : node13463;
													assign node13463 = (inp[12]) ? node13477 : node13464;
														assign node13464 = (inp[10]) ? node13472 : node13465;
															assign node13465 = (inp[11]) ? node13469 : node13466;
																assign node13466 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node13469 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node13472 = (inp[0]) ? 4'b1001 : node13473;
																assign node13473 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node13477 = (inp[0]) ? node13481 : node13478;
															assign node13478 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node13481 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node13484 = (inp[12]) ? node13500 : node13485;
														assign node13485 = (inp[10]) ? node13493 : node13486;
															assign node13486 = (inp[0]) ? node13490 : node13487;
																assign node13487 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node13490 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node13493 = (inp[11]) ? node13497 : node13494;
																assign node13494 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node13497 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node13500 = (inp[0]) ? 4'b1000 : node13501;
															assign node13501 = (inp[10]) ? node13505 : node13502;
																assign node13502 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node13505 = (inp[11]) ? 4'b1000 : 4'b1001;
												assign node13509 = (inp[10]) ? node13537 : node13510;
													assign node13510 = (inp[0]) ? node13522 : node13511;
														assign node13511 = (inp[12]) ? node13517 : node13512;
															assign node13512 = (inp[4]) ? node13514 : 4'b1100;
																assign node13514 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node13517 = (inp[4]) ? node13519 : 4'b1111;
																assign node13519 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node13522 = (inp[11]) ? node13530 : node13523;
															assign node13523 = (inp[4]) ? node13527 : node13524;
																assign node13524 = (inp[12]) ? 4'b1110 : 4'b1100;
																assign node13527 = (inp[12]) ? 4'b1100 : 4'b1111;
															assign node13530 = (inp[12]) ? node13534 : node13531;
																assign node13531 = (inp[4]) ? 4'b1110 : 4'b1101;
																assign node13534 = (inp[4]) ? 4'b1101 : 4'b1110;
													assign node13537 = (inp[4]) ? node13547 : node13538;
														assign node13538 = (inp[12]) ? 4'b1110 : node13539;
															assign node13539 = (inp[11]) ? node13543 : node13540;
																assign node13540 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node13543 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node13547 = (inp[12]) ? node13549 : 4'b1111;
															assign node13549 = (inp[11]) ? node13553 : node13550;
																assign node13550 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node13553 = (inp[0]) ? 4'b1100 : 4'b1101;
										assign node13556 = (inp[15]) ? node13646 : node13557;
											assign node13557 = (inp[4]) ? node13595 : node13558;
												assign node13558 = (inp[12]) ? node13582 : node13559;
													assign node13559 = (inp[10]) ? node13573 : node13560;
														assign node13560 = (inp[14]) ? node13566 : node13561;
															assign node13561 = (inp[11]) ? node13563 : 4'b1000;
																assign node13563 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node13566 = (inp[0]) ? node13570 : node13567;
																assign node13567 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node13570 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node13573 = (inp[11]) ? 4'b1001 : node13574;
															assign node13574 = (inp[14]) ? node13578 : node13575;
																assign node13575 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node13578 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node13582 = (inp[14]) ? node13588 : node13583;
														assign node13583 = (inp[0]) ? node13585 : 4'b1010;
															assign node13585 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node13588 = (inp[10]) ? node13592 : node13589;
															assign node13589 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node13592 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node13595 = (inp[12]) ? node13619 : node13596;
													assign node13596 = (inp[14]) ? node13608 : node13597;
														assign node13597 = (inp[0]) ? node13603 : node13598;
															assign node13598 = (inp[11]) ? 4'b1011 : node13599;
																assign node13599 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node13603 = (inp[11]) ? 4'b1010 : node13604;
																assign node13604 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node13608 = (inp[0]) ? node13614 : node13609;
															assign node13609 = (inp[10]) ? 4'b1010 : node13610;
																assign node13610 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node13614 = (inp[10]) ? 4'b1011 : node13615;
																assign node13615 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node13619 = (inp[11]) ? node13633 : node13620;
														assign node13620 = (inp[10]) ? node13626 : node13621;
															assign node13621 = (inp[14]) ? node13623 : 4'b1001;
																assign node13623 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node13626 = (inp[14]) ? node13630 : node13627;
																assign node13627 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node13630 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node13633 = (inp[10]) ? node13641 : node13634;
															assign node13634 = (inp[14]) ? node13638 : node13635;
																assign node13635 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node13638 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node13641 = (inp[0]) ? 4'b1000 : node13642;
																assign node13642 = (inp[14]) ? 4'b1000 : 4'b1001;
											assign node13646 = (inp[14]) ? node13690 : node13647;
												assign node13647 = (inp[12]) ? node13669 : node13648;
													assign node13648 = (inp[4]) ? node13656 : node13649;
														assign node13649 = (inp[10]) ? node13653 : node13650;
															assign node13650 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node13653 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node13656 = (inp[0]) ? node13662 : node13657;
															assign node13657 = (inp[11]) ? 4'b1011 : node13658;
																assign node13658 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node13662 = (inp[11]) ? node13666 : node13663;
																assign node13663 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node13666 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node13669 = (inp[4]) ? node13683 : node13670;
														assign node13670 = (inp[0]) ? node13678 : node13671;
															assign node13671 = (inp[10]) ? node13675 : node13672;
																assign node13672 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node13675 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node13678 = (inp[11]) ? 4'b1110 : node13679;
																assign node13679 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node13683 = (inp[0]) ? node13687 : node13684;
															assign node13684 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node13687 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node13690 = (inp[11]) ? node13710 : node13691;
													assign node13691 = (inp[0]) ? node13699 : node13692;
														assign node13692 = (inp[12]) ? node13696 : node13693;
															assign node13693 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node13696 = (inp[4]) ? 4'b1000 : 4'b1010;
														assign node13699 = (inp[10]) ? node13705 : node13700;
															assign node13700 = (inp[4]) ? node13702 : 4'b1001;
																assign node13702 = (inp[12]) ? 4'b1000 : 4'b1010;
															assign node13705 = (inp[12]) ? node13707 : 4'b1000;
																assign node13707 = (inp[4]) ? 4'b1001 : 4'b1011;
													assign node13710 = (inp[12]) ? node13720 : node13711;
														assign node13711 = (inp[4]) ? node13713 : 4'b1000;
															assign node13713 = (inp[0]) ? node13717 : node13714;
																assign node13714 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node13717 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node13720 = (inp[4]) ? 4'b1000 : node13721;
															assign node13721 = (inp[10]) ? 4'b1011 : node13722;
																assign node13722 = (inp[0]) ? 4'b1010 : 4'b1011;
							assign node13727 = (inp[4]) ? node14247 : node13728;
								assign node13728 = (inp[12]) ? node13992 : node13729;
									assign node13729 = (inp[15]) ? node13851 : node13730;
										assign node13730 = (inp[10]) ? node13784 : node13731;
											assign node13731 = (inp[11]) ? node13755 : node13732;
												assign node13732 = (inp[0]) ? node13746 : node13733;
													assign node13733 = (inp[14]) ? node13741 : node13734;
														assign node13734 = (inp[9]) ? node13736 : 4'b1100;
															assign node13736 = (inp[2]) ? 4'b1100 : node13737;
																assign node13737 = (inp[1]) ? 4'b1100 : 4'b1000;
														assign node13741 = (inp[2]) ? node13743 : 4'b1100;
															assign node13743 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node13746 = (inp[2]) ? node13750 : node13747;
														assign node13747 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node13750 = (inp[1]) ? 4'b1000 : node13751;
															assign node13751 = (inp[14]) ? 4'b1100 : 4'b1101;
												assign node13755 = (inp[0]) ? node13771 : node13756;
													assign node13756 = (inp[14]) ? node13764 : node13757;
														assign node13757 = (inp[1]) ? node13761 : node13758;
															assign node13758 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node13761 = (inp[2]) ? 4'b1001 : 4'b1101;
														assign node13764 = (inp[1]) ? node13768 : node13765;
															assign node13765 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node13768 = (inp[2]) ? 4'b1001 : 4'b1100;
													assign node13771 = (inp[14]) ? node13777 : node13772;
														assign node13772 = (inp[1]) ? 4'b1000 : node13773;
															assign node13773 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node13777 = (inp[1]) ? node13781 : node13778;
															assign node13778 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node13781 = (inp[2]) ? 4'b1000 : 4'b1101;
											assign node13784 = (inp[9]) ? node13816 : node13785;
												assign node13785 = (inp[11]) ? node13805 : node13786;
													assign node13786 = (inp[0]) ? node13796 : node13787;
														assign node13787 = (inp[2]) ? node13791 : node13788;
															assign node13788 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node13791 = (inp[1]) ? 4'b1000 : node13792;
																assign node13792 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node13796 = (inp[2]) ? node13800 : node13797;
															assign node13797 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node13800 = (inp[14]) ? node13802 : 4'b1100;
																assign node13802 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node13805 = (inp[1]) ? node13813 : node13806;
														assign node13806 = (inp[2]) ? node13808 : 4'b1000;
															assign node13808 = (inp[14]) ? node13810 : 4'b1100;
																assign node13810 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node13813 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node13816 = (inp[11]) ? node13836 : node13817;
													assign node13817 = (inp[1]) ? node13829 : node13818;
														assign node13818 = (inp[2]) ? node13822 : node13819;
															assign node13819 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node13822 = (inp[14]) ? node13826 : node13823;
																assign node13823 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node13826 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node13829 = (inp[2]) ? node13833 : node13830;
															assign node13830 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node13833 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node13836 = (inp[1]) ? node13842 : node13837;
														assign node13837 = (inp[2]) ? node13839 : 4'b1001;
															assign node13839 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node13842 = (inp[2]) ? 4'b1001 : node13843;
															assign node13843 = (inp[0]) ? node13847 : node13844;
																assign node13844 = (inp[14]) ? 4'b1101 : 4'b1100;
																assign node13847 = (inp[14]) ? 4'b1100 : 4'b1101;
										assign node13851 = (inp[11]) ? node13913 : node13852;
											assign node13852 = (inp[10]) ? node13884 : node13853;
												assign node13853 = (inp[0]) ? node13869 : node13854;
													assign node13854 = (inp[14]) ? node13862 : node13855;
														assign node13855 = (inp[1]) ? node13859 : node13856;
															assign node13856 = (inp[2]) ? 4'b1000 : 4'b1101;
															assign node13859 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node13862 = (inp[2]) ? node13866 : node13863;
															assign node13863 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node13866 = (inp[1]) ? 4'b1001 : 4'b1100;
													assign node13869 = (inp[1]) ? node13877 : node13870;
														assign node13870 = (inp[14]) ? node13874 : node13871;
															assign node13871 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node13874 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node13877 = (inp[2]) ? node13881 : node13878;
															assign node13878 = (inp[14]) ? 4'b1101 : 4'b1001;
															assign node13881 = (inp[14]) ? 4'b1000 : 4'b1101;
												assign node13884 = (inp[0]) ? node13900 : node13885;
													assign node13885 = (inp[14]) ? node13893 : node13886;
														assign node13886 = (inp[2]) ? node13890 : node13887;
															assign node13887 = (inp[1]) ? 4'b1001 : 4'b1100;
															assign node13890 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node13893 = (inp[9]) ? node13895 : 4'b1101;
															assign node13895 = (inp[2]) ? 4'b1000 : node13896;
																assign node13896 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node13900 = (inp[2]) ? node13906 : node13901;
														assign node13901 = (inp[1]) ? 4'b1000 : node13902;
															assign node13902 = (inp[14]) ? 4'b1000 : 4'b1101;
														assign node13906 = (inp[14]) ? node13910 : node13907;
															assign node13907 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node13910 = (inp[1]) ? 4'b1001 : 4'b1100;
											assign node13913 = (inp[14]) ? node13955 : node13914;
												assign node13914 = (inp[0]) ? node13940 : node13915;
													assign node13915 = (inp[9]) ? node13927 : node13916;
														assign node13916 = (inp[10]) ? node13922 : node13917;
															assign node13917 = (inp[1]) ? 4'b1001 : node13918;
																assign node13918 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node13922 = (inp[1]) ? node13924 : 4'b1001;
																assign node13924 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node13927 = (inp[10]) ? node13935 : node13928;
															assign node13928 = (inp[1]) ? node13932 : node13929;
																assign node13929 = (inp[2]) ? 4'b1000 : 4'b1100;
																assign node13932 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node13935 = (inp[1]) ? node13937 : 4'b1001;
																assign node13937 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node13940 = (inp[1]) ? node13948 : node13941;
														assign node13941 = (inp[2]) ? node13945 : node13942;
															assign node13942 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node13945 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node13948 = (inp[10]) ? node13952 : node13949;
															assign node13949 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node13952 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node13955 = (inp[1]) ? node13971 : node13956;
													assign node13956 = (inp[2]) ? node13962 : node13957;
														assign node13957 = (inp[10]) ? node13959 : 4'b1000;
															assign node13959 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node13962 = (inp[9]) ? 4'b1100 : node13963;
															assign node13963 = (inp[10]) ? node13967 : node13964;
																assign node13964 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node13967 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node13971 = (inp[2]) ? node13985 : node13972;
														assign node13972 = (inp[9]) ? node13978 : node13973;
															assign node13973 = (inp[0]) ? 4'b1100 : node13974;
																assign node13974 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node13978 = (inp[0]) ? node13982 : node13979;
																assign node13979 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node13982 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node13985 = (inp[9]) ? node13989 : node13986;
															assign node13986 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node13989 = (inp[0]) ? 4'b1000 : 4'b1001;
									assign node13992 = (inp[11]) ? node14114 : node13993;
										assign node13993 = (inp[14]) ? node14055 : node13994;
											assign node13994 = (inp[2]) ? node14026 : node13995;
												assign node13995 = (inp[10]) ? node14011 : node13996;
													assign node13996 = (inp[0]) ? node14004 : node13997;
														assign node13997 = (inp[15]) ? node14001 : node13998;
															assign node13998 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node14001 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node14004 = (inp[1]) ? node14008 : node14005;
															assign node14005 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node14008 = (inp[15]) ? 4'b1011 : 4'b1111;
													assign node14011 = (inp[0]) ? node14019 : node14012;
														assign node14012 = (inp[1]) ? node14016 : node14013;
															assign node14013 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node14016 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node14019 = (inp[1]) ? node14023 : node14020;
															assign node14020 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node14023 = (inp[15]) ? 4'b1010 : 4'b1110;
												assign node14026 = (inp[0]) ? node14042 : node14027;
													assign node14027 = (inp[10]) ? node14035 : node14028;
														assign node14028 = (inp[1]) ? node14032 : node14029;
															assign node14029 = (inp[15]) ? 4'b1010 : 4'b1111;
															assign node14032 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node14035 = (inp[1]) ? node14039 : node14036;
															assign node14036 = (inp[15]) ? 4'b1011 : 4'b1110;
															assign node14039 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node14042 = (inp[10]) ? node14048 : node14043;
														assign node14043 = (inp[15]) ? node14045 : 4'b1110;
															assign node14045 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node14048 = (inp[1]) ? node14052 : node14049;
															assign node14049 = (inp[15]) ? 4'b1010 : 4'b1111;
															assign node14052 = (inp[15]) ? 4'b1110 : 4'b1010;
											assign node14055 = (inp[0]) ? node14085 : node14056;
												assign node14056 = (inp[2]) ? node14072 : node14057;
													assign node14057 = (inp[10]) ? node14065 : node14058;
														assign node14058 = (inp[1]) ? node14062 : node14059;
															assign node14059 = (inp[15]) ? 4'b1010 : 4'b1111;
															assign node14062 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node14065 = (inp[1]) ? node14069 : node14066;
															assign node14066 = (inp[15]) ? 4'b1011 : 4'b1110;
															assign node14069 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node14072 = (inp[10]) ? node14080 : node14073;
														assign node14073 = (inp[15]) ? node14077 : node14074;
															assign node14074 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node14077 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node14080 = (inp[1]) ? 4'b1110 : node14081;
															assign node14081 = (inp[15]) ? 4'b1110 : 4'b1011;
												assign node14085 = (inp[10]) ? node14101 : node14086;
													assign node14086 = (inp[2]) ? node14094 : node14087;
														assign node14087 = (inp[15]) ? node14091 : node14088;
															assign node14088 = (inp[1]) ? 4'b1011 : 4'b1110;
															assign node14091 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node14094 = (inp[15]) ? node14098 : node14095;
															assign node14095 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node14098 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node14101 = (inp[2]) ? node14107 : node14102;
														assign node14102 = (inp[15]) ? node14104 : 4'b1010;
															assign node14104 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node14107 = (inp[15]) ? node14111 : node14108;
															assign node14108 = (inp[9]) ? 4'b1010 : 4'b1111;
															assign node14111 = (inp[1]) ? 4'b1011 : 4'b1111;
										assign node14114 = (inp[15]) ? node14174 : node14115;
											assign node14115 = (inp[1]) ? node14145 : node14116;
												assign node14116 = (inp[2]) ? node14132 : node14117;
													assign node14117 = (inp[14]) ? node14125 : node14118;
														assign node14118 = (inp[9]) ? node14120 : 4'b1010;
															assign node14120 = (inp[0]) ? node14122 : 4'b1011;
																assign node14122 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node14125 = (inp[10]) ? node14129 : node14126;
															assign node14126 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node14129 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node14132 = (inp[9]) ? node14138 : node14133;
														assign node14133 = (inp[0]) ? node14135 : 4'b1110;
															assign node14135 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node14138 = (inp[0]) ? node14142 : node14139;
															assign node14139 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node14142 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node14145 = (inp[14]) ? node14159 : node14146;
													assign node14146 = (inp[2]) ? node14154 : node14147;
														assign node14147 = (inp[0]) ? node14151 : node14148;
															assign node14148 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node14151 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node14154 = (inp[0]) ? node14156 : 4'b1010;
															assign node14156 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node14159 = (inp[2]) ? node14169 : node14160;
														assign node14160 = (inp[9]) ? node14162 : 4'b1011;
															assign node14162 = (inp[0]) ? node14166 : node14163;
																assign node14163 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node14166 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node14169 = (inp[10]) ? node14171 : 4'b1111;
															assign node14171 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node14174 = (inp[10]) ? node14218 : node14175;
												assign node14175 = (inp[0]) ? node14191 : node14176;
													assign node14176 = (inp[14]) ? node14184 : node14177;
														assign node14177 = (inp[2]) ? node14181 : node14178;
															assign node14178 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node14181 = (inp[1]) ? 4'b1110 : 4'b1011;
														assign node14184 = (inp[1]) ? node14188 : node14185;
															assign node14185 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node14188 = (inp[2]) ? 4'b1010 : 4'b1111;
													assign node14191 = (inp[9]) ? node14205 : node14192;
														assign node14192 = (inp[1]) ? node14200 : node14193;
															assign node14193 = (inp[2]) ? node14197 : node14194;
																assign node14194 = (inp[14]) ? 4'b1011 : 4'b1111;
																assign node14197 = (inp[14]) ? 4'b1111 : 4'b1010;
															assign node14200 = (inp[2]) ? 4'b1011 : node14201;
																assign node14201 = (inp[14]) ? 4'b1110 : 4'b1011;
														assign node14205 = (inp[14]) ? node14211 : node14206;
															assign node14206 = (inp[1]) ? 4'b1111 : node14207;
																assign node14207 = (inp[2]) ? 4'b1010 : 4'b1111;
															assign node14211 = (inp[2]) ? node14215 : node14212;
																assign node14212 = (inp[1]) ? 4'b1110 : 4'b1011;
																assign node14215 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node14218 = (inp[0]) ? node14232 : node14219;
													assign node14219 = (inp[1]) ? node14225 : node14220;
														assign node14220 = (inp[14]) ? 4'b1111 : node14221;
															assign node14221 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node14225 = (inp[14]) ? node14229 : node14226;
															assign node14226 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node14229 = (inp[2]) ? 4'b1011 : 4'b1110;
													assign node14232 = (inp[1]) ? node14240 : node14233;
														assign node14233 = (inp[2]) ? node14237 : node14234;
															assign node14234 = (inp[14]) ? 4'b1010 : 4'b1110;
															assign node14237 = (inp[14]) ? 4'b1110 : 4'b1011;
														assign node14240 = (inp[2]) ? node14244 : node14241;
															assign node14241 = (inp[14]) ? 4'b1111 : 4'b1010;
															assign node14244 = (inp[14]) ? 4'b1010 : 4'b1110;
								assign node14247 = (inp[12]) ? node14461 : node14248;
									assign node14248 = (inp[2]) ? node14388 : node14249;
										assign node14249 = (inp[1]) ? node14327 : node14250;
											assign node14250 = (inp[14]) ? node14286 : node14251;
												assign node14251 = (inp[15]) ? node14271 : node14252;
													assign node14252 = (inp[0]) ? node14260 : node14253;
														assign node14253 = (inp[11]) ? node14257 : node14254;
															assign node14254 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node14257 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node14260 = (inp[9]) ? node14266 : node14261;
															assign node14261 = (inp[11]) ? 4'b1011 : node14262;
																assign node14262 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node14266 = (inp[10]) ? 4'b1011 : node14267;
																assign node14267 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node14271 = (inp[9]) ? node14279 : node14272;
														assign node14272 = (inp[0]) ? node14276 : node14273;
															assign node14273 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node14276 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node14279 = (inp[10]) ? node14283 : node14280;
															assign node14280 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node14283 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node14286 = (inp[11]) ? node14310 : node14287;
													assign node14287 = (inp[15]) ? node14303 : node14288;
														assign node14288 = (inp[9]) ? node14296 : node14289;
															assign node14289 = (inp[0]) ? node14293 : node14290;
																assign node14290 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node14293 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node14296 = (inp[10]) ? node14300 : node14297;
																assign node14297 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node14300 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node14303 = (inp[0]) ? node14307 : node14304;
															assign node14304 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node14307 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node14310 = (inp[0]) ? node14318 : node14311;
														assign node14311 = (inp[10]) ? node14315 : node14312;
															assign node14312 = (inp[15]) ? 4'b1011 : 4'b1010;
															assign node14315 = (inp[15]) ? 4'b1010 : 4'b1011;
														assign node14318 = (inp[9]) ? node14320 : 4'b1011;
															assign node14320 = (inp[15]) ? node14324 : node14321;
																assign node14321 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node14324 = (inp[10]) ? 4'b1011 : 4'b1010;
											assign node14327 = (inp[11]) ? node14361 : node14328;
												assign node14328 = (inp[15]) ? node14342 : node14329;
													assign node14329 = (inp[9]) ? node14335 : node14330;
														assign node14330 = (inp[0]) ? node14332 : 4'b1110;
															assign node14332 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node14335 = (inp[0]) ? node14339 : node14336;
															assign node14336 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node14339 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node14342 = (inp[14]) ? node14354 : node14343;
														assign node14343 = (inp[9]) ? node14349 : node14344;
															assign node14344 = (inp[0]) ? node14346 : 4'b1111;
																assign node14346 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node14349 = (inp[0]) ? 4'b1110 : node14350;
																assign node14350 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node14354 = (inp[0]) ? node14358 : node14355;
															assign node14355 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node14358 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node14361 = (inp[15]) ? node14367 : node14362;
													assign node14362 = (inp[9]) ? node14364 : 4'b1111;
														assign node14364 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node14367 = (inp[14]) ? node14381 : node14368;
														assign node14368 = (inp[9]) ? node14376 : node14369;
															assign node14369 = (inp[10]) ? node14373 : node14370;
																assign node14370 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node14373 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node14376 = (inp[10]) ? node14378 : 4'b1110;
																assign node14378 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node14381 = (inp[10]) ? node14385 : node14382;
															assign node14382 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node14385 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node14388 = (inp[1]) ? node14438 : node14389;
											assign node14389 = (inp[0]) ? node14411 : node14390;
												assign node14390 = (inp[10]) ? node14400 : node14391;
													assign node14391 = (inp[15]) ? 4'b1111 : node14392;
														assign node14392 = (inp[14]) ? node14396 : node14393;
															assign node14393 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node14396 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node14400 = (inp[15]) ? 4'b1110 : node14401;
														assign node14401 = (inp[9]) ? node14407 : node14402;
															assign node14402 = (inp[11]) ? 4'b1110 : node14403;
																assign node14403 = (inp[14]) ? 4'b1111 : 4'b1110;
															assign node14407 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node14411 = (inp[10]) ? node14429 : node14412;
													assign node14412 = (inp[15]) ? 4'b1110 : node14413;
														assign node14413 = (inp[9]) ? node14421 : node14414;
															assign node14414 = (inp[14]) ? node14418 : node14415;
																assign node14415 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node14418 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node14421 = (inp[11]) ? node14425 : node14422;
																assign node14422 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node14425 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node14429 = (inp[15]) ? 4'b1111 : node14430;
														assign node14430 = (inp[11]) ? node14434 : node14431;
															assign node14431 = (inp[14]) ? 4'b1110 : 4'b1111;
															assign node14434 = (inp[14]) ? 4'b1111 : 4'b1110;
											assign node14438 = (inp[14]) ? node14454 : node14439;
												assign node14439 = (inp[15]) ? node14447 : node14440;
													assign node14440 = (inp[0]) ? node14444 : node14441;
														assign node14441 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node14444 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node14447 = (inp[10]) ? node14451 : node14448;
														assign node14448 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node14451 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node14454 = (inp[10]) ? node14458 : node14455;
													assign node14455 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node14458 = (inp[0]) ? 4'b1010 : 4'b1011;
									assign node14461 = (inp[1]) ? node14583 : node14462;
										assign node14462 = (inp[2]) ? node14528 : node14463;
											assign node14463 = (inp[15]) ? node14487 : node14464;
												assign node14464 = (inp[11]) ? node14472 : node14465;
													assign node14465 = (inp[10]) ? node14469 : node14466;
														assign node14466 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node14469 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node14472 = (inp[10]) ? node14480 : node14473;
														assign node14473 = (inp[14]) ? node14477 : node14474;
															assign node14474 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node14477 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node14480 = (inp[0]) ? node14484 : node14481;
															assign node14481 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node14484 = (inp[14]) ? 4'b1001 : 4'b1000;
												assign node14487 = (inp[14]) ? node14509 : node14488;
													assign node14488 = (inp[0]) ? node14496 : node14489;
														assign node14489 = (inp[9]) ? 4'b1101 : node14490;
															assign node14490 = (inp[10]) ? 4'b1101 : node14491;
																assign node14491 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node14496 = (inp[9]) ? node14504 : node14497;
															assign node14497 = (inp[10]) ? node14501 : node14498;
																assign node14498 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node14501 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node14504 = (inp[10]) ? node14506 : 4'b1100;
																assign node14506 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node14509 = (inp[9]) ? node14519 : node14510;
														assign node14510 = (inp[11]) ? 4'b1001 : node14511;
															assign node14511 = (inp[0]) ? node14515 : node14512;
																assign node14512 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node14515 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node14519 = (inp[0]) ? 4'b1000 : node14520;
															assign node14520 = (inp[10]) ? node14524 : node14521;
																assign node14521 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node14524 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node14528 = (inp[15]) ? node14564 : node14529;
												assign node14529 = (inp[0]) ? node14551 : node14530;
													assign node14530 = (inp[9]) ? node14542 : node14531;
														assign node14531 = (inp[11]) ? node14537 : node14532;
															assign node14532 = (inp[14]) ? 4'b1100 : node14533;
																assign node14533 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node14537 = (inp[10]) ? 4'b1101 : node14538;
																assign node14538 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node14542 = (inp[14]) ? 4'b1101 : node14543;
															assign node14543 = (inp[10]) ? node14547 : node14544;
																assign node14544 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node14547 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node14551 = (inp[14]) ? node14559 : node14552;
														assign node14552 = (inp[11]) ? node14556 : node14553;
															assign node14553 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node14556 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node14559 = (inp[11]) ? 4'b1100 : node14560;
															assign node14560 = (inp[10]) ? 4'b1101 : 4'b1100;
												assign node14564 = (inp[14]) ? node14578 : node14565;
													assign node14565 = (inp[9]) ? node14573 : node14566;
														assign node14566 = (inp[10]) ? node14570 : node14567;
															assign node14567 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node14570 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node14573 = (inp[10]) ? 4'b1001 : node14574;
															assign node14574 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node14578 = (inp[0]) ? 4'b1101 : node14579;
														assign node14579 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node14583 = (inp[2]) ? node14647 : node14584;
											assign node14584 = (inp[15]) ? node14624 : node14585;
												assign node14585 = (inp[9]) ? node14609 : node14586;
													assign node14586 = (inp[0]) ? node14598 : node14587;
														assign node14587 = (inp[10]) ? node14593 : node14588;
															assign node14588 = (inp[14]) ? 4'b1100 : node14589;
																assign node14589 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node14593 = (inp[11]) ? node14595 : 4'b1101;
																assign node14595 = (inp[14]) ? 4'b1101 : 4'b1100;
														assign node14598 = (inp[10]) ? node14604 : node14599;
															assign node14599 = (inp[14]) ? 4'b1101 : node14600;
																assign node14600 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node14604 = (inp[14]) ? 4'b1100 : node14605;
																assign node14605 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node14609 = (inp[14]) ? node14617 : node14610;
														assign node14610 = (inp[0]) ? 4'b1100 : node14611;
															assign node14611 = (inp[10]) ? node14613 : 4'b1100;
																assign node14613 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node14617 = (inp[10]) ? node14621 : node14618;
															assign node14618 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node14621 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node14624 = (inp[14]) ? node14640 : node14625;
													assign node14625 = (inp[0]) ? node14633 : node14626;
														assign node14626 = (inp[11]) ? node14630 : node14627;
															assign node14627 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node14630 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node14633 = (inp[11]) ? node14637 : node14634;
															assign node14634 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node14637 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node14640 = (inp[0]) ? node14644 : node14641;
														assign node14641 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node14644 = (inp[10]) ? 4'b1100 : 4'b1101;
											assign node14647 = (inp[14]) ? node14669 : node14648;
												assign node14648 = (inp[15]) ? node14656 : node14649;
													assign node14649 = (inp[10]) ? node14653 : node14650;
														assign node14650 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node14653 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node14656 = (inp[10]) ? node14664 : node14657;
														assign node14657 = (inp[0]) ? node14661 : node14658;
															assign node14658 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node14661 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node14664 = (inp[11]) ? node14666 : 4'b1101;
															assign node14666 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node14669 = (inp[15]) ? node14677 : node14670;
													assign node14670 = (inp[0]) ? node14674 : node14671;
														assign node14671 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node14674 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node14677 = (inp[9]) ? node14679 : 4'b1000;
														assign node14679 = (inp[0]) ? node14683 : node14680;
															assign node14680 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node14683 = (inp[10]) ? 4'b1000 : 4'b1001;
						assign node14686 = (inp[15]) ? node15620 : node14687;
							assign node14687 = (inp[14]) ? node15211 : node14688;
								assign node14688 = (inp[4]) ? node14912 : node14689;
									assign node14689 = (inp[12]) ? node14805 : node14690;
										assign node14690 = (inp[10]) ? node14744 : node14691;
											assign node14691 = (inp[0]) ? node14717 : node14692;
												assign node14692 = (inp[13]) ? node14708 : node14693;
													assign node14693 = (inp[11]) ? node14701 : node14694;
														assign node14694 = (inp[1]) ? node14698 : node14695;
															assign node14695 = (inp[2]) ? 4'b1001 : 4'b1101;
															assign node14698 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node14701 = (inp[1]) ? node14705 : node14702;
															assign node14702 = (inp[2]) ? 4'b1000 : 4'b1101;
															assign node14705 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node14708 = (inp[1]) ? node14714 : node14709;
														assign node14709 = (inp[2]) ? 4'b1000 : node14710;
															assign node14710 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node14714 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node14717 = (inp[13]) ? node14735 : node14718;
													assign node14718 = (inp[11]) ? node14728 : node14719;
														assign node14719 = (inp[9]) ? node14725 : node14720;
															assign node14720 = (inp[2]) ? node14722 : 4'b1000;
																assign node14722 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node14725 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node14728 = (inp[1]) ? node14732 : node14729;
															assign node14729 = (inp[2]) ? 4'b1001 : 4'b1100;
															assign node14732 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node14735 = (inp[1]) ? node14741 : node14736;
														assign node14736 = (inp[2]) ? 4'b1001 : node14737;
															assign node14737 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node14741 = (inp[2]) ? 4'b1101 : 4'b1001;
											assign node14744 = (inp[0]) ? node14772 : node14745;
												assign node14745 = (inp[11]) ? node14757 : node14746;
													assign node14746 = (inp[13]) ? node14754 : node14747;
														assign node14747 = (inp[1]) ? node14751 : node14748;
															assign node14748 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node14751 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node14754 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node14757 = (inp[13]) ? node14765 : node14758;
														assign node14758 = (inp[2]) ? node14762 : node14759;
															assign node14759 = (inp[1]) ? 4'b1001 : 4'b1100;
															assign node14762 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node14765 = (inp[2]) ? node14769 : node14766;
															assign node14766 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node14769 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node14772 = (inp[11]) ? node14790 : node14773;
													assign node14773 = (inp[13]) ? node14783 : node14774;
														assign node14774 = (inp[9]) ? node14776 : 4'b1101;
															assign node14776 = (inp[1]) ? node14780 : node14777;
																assign node14777 = (inp[2]) ? 4'b1001 : 4'b1101;
																assign node14780 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node14783 = (inp[2]) ? node14787 : node14784;
															assign node14784 = (inp[1]) ? 4'b1000 : 4'b1101;
															assign node14787 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node14790 = (inp[9]) ? node14800 : node14791;
														assign node14791 = (inp[1]) ? node14797 : node14792;
															assign node14792 = (inp[2]) ? 4'b1000 : node14793;
																assign node14793 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node14797 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node14800 = (inp[13]) ? 4'b1100 : node14801;
															assign node14801 = (inp[2]) ? 4'b1100 : 4'b1000;
										assign node14805 = (inp[2]) ? node14857 : node14806;
											assign node14806 = (inp[1]) ? node14836 : node14807;
												assign node14807 = (inp[9]) ? node14821 : node14808;
													assign node14808 = (inp[13]) ? 4'b1110 : node14809;
														assign node14809 = (inp[11]) ? node14815 : node14810;
															assign node14810 = (inp[10]) ? 4'b1110 : node14811;
																assign node14811 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node14815 = (inp[10]) ? 4'b1111 : node14816;
																assign node14816 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node14821 = (inp[0]) ? node14833 : node14822;
														assign node14822 = (inp[10]) ? node14828 : node14823;
															assign node14823 = (inp[13]) ? 4'b1110 : node14824;
																assign node14824 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node14828 = (inp[13]) ? 4'b1111 : node14829;
																assign node14829 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node14833 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node14836 = (inp[11]) ? node14844 : node14837;
													assign node14837 = (inp[10]) ? node14841 : node14838;
														assign node14838 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node14841 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node14844 = (inp[10]) ? node14852 : node14845;
														assign node14845 = (inp[0]) ? node14849 : node14846;
															assign node14846 = (inp[13]) ? 4'b1010 : 4'b1011;
															assign node14849 = (inp[13]) ? 4'b1011 : 4'b1010;
														assign node14852 = (inp[0]) ? 4'b1011 : node14853;
															assign node14853 = (inp[13]) ? 4'b1011 : 4'b1010;
											assign node14857 = (inp[1]) ? node14881 : node14858;
												assign node14858 = (inp[9]) ? node14868 : node14859;
													assign node14859 = (inp[11]) ? 4'b1011 : node14860;
														assign node14860 = (inp[0]) ? node14864 : node14861;
															assign node14861 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node14864 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node14868 = (inp[0]) ? node14878 : node14869;
														assign node14869 = (inp[10]) ? node14875 : node14870;
															assign node14870 = (inp[13]) ? node14872 : 4'b1010;
																assign node14872 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node14875 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node14878 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node14881 = (inp[9]) ? node14897 : node14882;
													assign node14882 = (inp[11]) ? node14890 : node14883;
														assign node14883 = (inp[10]) ? node14887 : node14884;
															assign node14884 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node14887 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node14890 = (inp[13]) ? 4'b1110 : node14891;
															assign node14891 = (inp[0]) ? node14893 : 4'b1110;
																assign node14893 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node14897 = (inp[0]) ? node14903 : node14898;
														assign node14898 = (inp[10]) ? node14900 : 4'b1111;
															assign node14900 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node14903 = (inp[10]) ? node14907 : node14904;
															assign node14904 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node14907 = (inp[13]) ? node14909 : 4'b1111;
																assign node14909 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node14912 = (inp[12]) ? node15070 : node14913;
										assign node14913 = (inp[1]) ? node14989 : node14914;
											assign node14914 = (inp[2]) ? node14948 : node14915;
												assign node14915 = (inp[11]) ? node14941 : node14916;
													assign node14916 = (inp[9]) ? node14932 : node14917;
														assign node14917 = (inp[10]) ? node14925 : node14918;
															assign node14918 = (inp[0]) ? node14922 : node14919;
																assign node14919 = (inp[13]) ? 4'b1110 : 4'b1111;
																assign node14922 = (inp[13]) ? 4'b1111 : 4'b1110;
															assign node14925 = (inp[13]) ? node14929 : node14926;
																assign node14926 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node14929 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node14932 = (inp[13]) ? node14934 : 4'b1111;
															assign node14934 = (inp[0]) ? node14938 : node14935;
																assign node14935 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node14938 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node14941 = (inp[0]) ? node14945 : node14942;
														assign node14942 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node14945 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node14948 = (inp[13]) ? node14964 : node14949;
													assign node14949 = (inp[9]) ? node14957 : node14950;
														assign node14950 = (inp[10]) ? node14954 : node14951;
															assign node14951 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node14954 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node14957 = (inp[0]) ? node14961 : node14958;
															assign node14958 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node14961 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node14964 = (inp[10]) ? node14974 : node14965;
														assign node14965 = (inp[9]) ? 4'b1011 : node14966;
															assign node14966 = (inp[11]) ? node14970 : node14967;
																assign node14967 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node14970 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node14974 = (inp[9]) ? node14982 : node14975;
															assign node14975 = (inp[11]) ? node14979 : node14976;
																assign node14976 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node14979 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node14982 = (inp[0]) ? node14986 : node14983;
																assign node14983 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node14986 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node14989 = (inp[2]) ? node15033 : node14990;
												assign node14990 = (inp[13]) ? node15018 : node14991;
													assign node14991 = (inp[9]) ? node15003 : node14992;
														assign node14992 = (inp[11]) ? node14998 : node14993;
															assign node14993 = (inp[10]) ? 4'b1011 : node14994;
																assign node14994 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node14998 = (inp[10]) ? node15000 : 4'b1011;
																assign node15000 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node15003 = (inp[11]) ? node15011 : node15004;
															assign node15004 = (inp[0]) ? node15008 : node15005;
																assign node15005 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node15008 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node15011 = (inp[10]) ? node15015 : node15012;
																assign node15012 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node15015 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node15018 = (inp[10]) ? node15026 : node15019;
														assign node15019 = (inp[0]) ? node15023 : node15020;
															assign node15020 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node15023 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node15026 = (inp[0]) ? node15030 : node15027;
															assign node15027 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node15030 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node15033 = (inp[9]) ? node15055 : node15034;
													assign node15034 = (inp[0]) ? node15044 : node15035;
														assign node15035 = (inp[10]) ? node15041 : node15036;
															assign node15036 = (inp[11]) ? node15038 : 4'b1111;
																assign node15038 = (inp[13]) ? 4'b1110 : 4'b1111;
															assign node15041 = (inp[13]) ? 4'b1111 : 4'b1110;
														assign node15044 = (inp[10]) ? node15050 : node15045;
															assign node15045 = (inp[13]) ? node15047 : 4'b1110;
																assign node15047 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node15050 = (inp[13]) ? node15052 : 4'b1111;
																assign node15052 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node15055 = (inp[11]) ? node15063 : node15056;
														assign node15056 = (inp[10]) ? node15060 : node15057;
															assign node15057 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node15060 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node15063 = (inp[0]) ? 4'b1111 : node15064;
															assign node15064 = (inp[13]) ? 4'b1111 : node15065;
																assign node15065 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node15070 = (inp[2]) ? node15140 : node15071;
											assign node15071 = (inp[1]) ? node15105 : node15072;
												assign node15072 = (inp[9]) ? node15088 : node15073;
													assign node15073 = (inp[11]) ? node15083 : node15074;
														assign node15074 = (inp[13]) ? node15076 : 4'b1000;
															assign node15076 = (inp[0]) ? node15080 : node15077;
																assign node15077 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node15080 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node15083 = (inp[0]) ? node15085 : 4'b1001;
															assign node15085 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node15088 = (inp[11]) ? node15098 : node15089;
														assign node15089 = (inp[0]) ? 4'b1000 : node15090;
															assign node15090 = (inp[13]) ? node15094 : node15091;
																assign node15091 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node15094 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node15098 = (inp[13]) ? 4'b1000 : node15099;
															assign node15099 = (inp[0]) ? node15101 : 4'b1000;
																assign node15101 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node15105 = (inp[13]) ? node15127 : node15106;
													assign node15106 = (inp[9]) ? node15114 : node15107;
														assign node15107 = (inp[11]) ? 4'b1101 : node15108;
															assign node15108 = (inp[0]) ? node15110 : 4'b1101;
																assign node15110 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node15114 = (inp[11]) ? node15120 : node15115;
															assign node15115 = (inp[0]) ? 4'b1101 : node15116;
																assign node15116 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node15120 = (inp[10]) ? node15124 : node15121;
																assign node15121 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node15124 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node15127 = (inp[9]) ? node15135 : node15128;
														assign node15128 = (inp[10]) ? node15132 : node15129;
															assign node15129 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node15132 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node15135 = (inp[0]) ? 4'b1100 : node15136;
															assign node15136 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node15140 = (inp[1]) ? node15164 : node15141;
												assign node15141 = (inp[10]) ? node15153 : node15142;
													assign node15142 = (inp[0]) ? node15148 : node15143;
														assign node15143 = (inp[11]) ? 4'b1100 : node15144;
															assign node15144 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node15148 = (inp[13]) ? 4'b1101 : node15149;
															assign node15149 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node15153 = (inp[0]) ? node15159 : node15154;
														assign node15154 = (inp[11]) ? 4'b1101 : node15155;
															assign node15155 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node15159 = (inp[11]) ? 4'b1100 : node15160;
															assign node15160 = (inp[13]) ? 4'b1100 : 4'b1101;
												assign node15164 = (inp[13]) ? node15190 : node15165;
													assign node15165 = (inp[11]) ? node15179 : node15166;
														assign node15166 = (inp[9]) ? node15172 : node15167;
															assign node15167 = (inp[10]) ? 4'b1001 : node15168;
																assign node15168 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node15172 = (inp[0]) ? node15176 : node15173;
																assign node15173 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node15176 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node15179 = (inp[9]) ? node15185 : node15180;
															assign node15180 = (inp[0]) ? 4'b1000 : node15181;
																assign node15181 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node15185 = (inp[10]) ? node15187 : 4'b1000;
																assign node15187 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node15190 = (inp[0]) ? node15200 : node15191;
														assign node15191 = (inp[9]) ? 4'b1001 : node15192;
															assign node15192 = (inp[11]) ? node15196 : node15193;
																assign node15193 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node15196 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node15200 = (inp[9]) ? node15206 : node15201;
															assign node15201 = (inp[10]) ? node15203 : 4'b1001;
																assign node15203 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node15206 = (inp[10]) ? 4'b1000 : node15207;
																assign node15207 = (inp[11]) ? 4'b1001 : 4'b1000;
								assign node15211 = (inp[4]) ? node15419 : node15212;
									assign node15212 = (inp[12]) ? node15302 : node15213;
										assign node15213 = (inp[0]) ? node15255 : node15214;
											assign node15214 = (inp[11]) ? node15240 : node15215;
												assign node15215 = (inp[10]) ? node15227 : node15216;
													assign node15216 = (inp[2]) ? node15222 : node15217;
														assign node15217 = (inp[13]) ? 4'b1100 : node15218;
															assign node15218 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node15222 = (inp[1]) ? node15224 : 4'b1100;
															assign node15224 = (inp[13]) ? 4'b1001 : 4'b1000;
													assign node15227 = (inp[13]) ? node15235 : node15228;
														assign node15228 = (inp[2]) ? node15232 : node15229;
															assign node15229 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node15232 = (inp[1]) ? 4'b1001 : 4'b1101;
														assign node15235 = (inp[1]) ? 4'b1101 : node15236;
															assign node15236 = (inp[2]) ? 4'b1101 : 4'b1001;
												assign node15240 = (inp[10]) ? node15250 : node15241;
													assign node15241 = (inp[2]) ? node15245 : node15242;
														assign node15242 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node15245 = (inp[1]) ? 4'b1000 : node15246;
															assign node15246 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node15250 = (inp[2]) ? 4'b1001 : node15251;
														assign node15251 = (inp[1]) ? 4'b1100 : 4'b1000;
											assign node15255 = (inp[2]) ? node15277 : node15256;
												assign node15256 = (inp[1]) ? node15268 : node15257;
													assign node15257 = (inp[10]) ? node15263 : node15258;
														assign node15258 = (inp[11]) ? 4'b1000 : node15259;
															assign node15259 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node15263 = (inp[13]) ? node15265 : 4'b1001;
															assign node15265 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node15268 = (inp[10]) ? node15274 : node15269;
														assign node15269 = (inp[13]) ? node15271 : 4'b1100;
															assign node15271 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node15274 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node15277 = (inp[1]) ? node15289 : node15278;
													assign node15278 = (inp[10]) ? node15284 : node15279;
														assign node15279 = (inp[11]) ? node15281 : 4'b1101;
															assign node15281 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node15284 = (inp[13]) ? 4'b1100 : node15285;
															assign node15285 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node15289 = (inp[10]) ? node15297 : node15290;
														assign node15290 = (inp[9]) ? 4'b1001 : node15291;
															assign node15291 = (inp[13]) ? node15293 : 4'b1001;
																assign node15293 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15297 = (inp[13]) ? node15299 : 4'b1000;
															assign node15299 = (inp[11]) ? 4'b1000 : 4'b1001;
										assign node15302 = (inp[13]) ? node15364 : node15303;
											assign node15303 = (inp[0]) ? node15335 : node15304;
												assign node15304 = (inp[10]) ? node15320 : node15305;
													assign node15305 = (inp[11]) ? node15313 : node15306;
														assign node15306 = (inp[9]) ? node15308 : 4'b1010;
															assign node15308 = (inp[2]) ? node15310 : 4'b1111;
																assign node15310 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node15313 = (inp[2]) ? node15317 : node15314;
															assign node15314 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node15317 = (inp[1]) ? 4'b1011 : 4'b1110;
													assign node15320 = (inp[11]) ? node15328 : node15321;
														assign node15321 = (inp[1]) ? node15325 : node15322;
															assign node15322 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node15325 = (inp[2]) ? 4'b1011 : 4'b1110;
														assign node15328 = (inp[2]) ? node15332 : node15329;
															assign node15329 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node15332 = (inp[1]) ? 4'b1010 : 4'b1111;
												assign node15335 = (inp[10]) ? node15347 : node15336;
													assign node15336 = (inp[2]) ? node15342 : node15337;
														assign node15337 = (inp[1]) ? 4'b1110 : node15338;
															assign node15338 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node15342 = (inp[1]) ? node15344 : 4'b1111;
															assign node15344 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node15347 = (inp[11]) ? node15357 : node15348;
														assign node15348 = (inp[9]) ? 4'b1010 : node15349;
															assign node15349 = (inp[2]) ? node15353 : node15350;
																assign node15350 = (inp[1]) ? 4'b1111 : 4'b1010;
																assign node15353 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node15357 = (inp[2]) ? node15361 : node15358;
															assign node15358 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node15361 = (inp[1]) ? 4'b1011 : 4'b1110;
											assign node15364 = (inp[10]) ? node15384 : node15365;
												assign node15365 = (inp[1]) ? node15377 : node15366;
													assign node15366 = (inp[2]) ? node15370 : node15367;
														assign node15367 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node15370 = (inp[11]) ? node15374 : node15371;
															assign node15371 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node15374 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node15377 = (inp[2]) ? node15381 : node15378;
														assign node15378 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node15381 = (inp[0]) ? 4'b1011 : 4'b1010;
												assign node15384 = (inp[0]) ? node15404 : node15385;
													assign node15385 = (inp[11]) ? node15399 : node15386;
														assign node15386 = (inp[9]) ? node15392 : node15387;
															assign node15387 = (inp[2]) ? 4'b1110 : node15388;
																assign node15388 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node15392 = (inp[2]) ? node15396 : node15393;
																assign node15393 = (inp[1]) ? 4'b1110 : 4'b1011;
																assign node15396 = (inp[1]) ? 4'b1011 : 4'b1110;
														assign node15399 = (inp[9]) ? node15401 : 4'b1011;
															assign node15401 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node15404 = (inp[11]) ? node15412 : node15405;
														assign node15405 = (inp[1]) ? node15409 : node15406;
															assign node15406 = (inp[2]) ? 4'b1111 : 4'b1010;
															assign node15409 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node15412 = (inp[1]) ? node15416 : node15413;
															assign node15413 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node15416 = (inp[9]) ? 4'b1111 : 4'b1010;
									assign node15419 = (inp[12]) ? node15529 : node15420;
										assign node15420 = (inp[0]) ? node15476 : node15421;
											assign node15421 = (inp[10]) ? node15453 : node15422;
												assign node15422 = (inp[11]) ? node15438 : node15423;
													assign node15423 = (inp[13]) ? node15431 : node15424;
														assign node15424 = (inp[9]) ? 4'b1010 : node15425;
															assign node15425 = (inp[2]) ? node15427 : 4'b1010;
																assign node15427 = (inp[1]) ? 4'b1010 : 4'b1111;
														assign node15431 = (inp[1]) ? node15435 : node15432;
															assign node15432 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node15435 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node15438 = (inp[13]) ? node15446 : node15439;
														assign node15439 = (inp[1]) ? node15443 : node15440;
															assign node15440 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node15443 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node15446 = (inp[2]) ? node15450 : node15447;
															assign node15447 = (inp[1]) ? 4'b1110 : 4'b1010;
															assign node15450 = (inp[1]) ? 4'b1010 : 4'b1111;
												assign node15453 = (inp[13]) ? node15467 : node15454;
													assign node15454 = (inp[11]) ? node15460 : node15455;
														assign node15455 = (inp[1]) ? node15457 : 4'b1110;
															assign node15457 = (inp[2]) ? 4'b1011 : 4'b1111;
														assign node15460 = (inp[1]) ? node15464 : node15461;
															assign node15461 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node15464 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node15467 = (inp[2]) ? node15471 : node15468;
														assign node15468 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node15471 = (inp[1]) ? 4'b1011 : node15472;
															assign node15472 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node15476 = (inp[10]) ? node15498 : node15477;
												assign node15477 = (inp[13]) ? node15491 : node15478;
													assign node15478 = (inp[11]) ? node15484 : node15479;
														assign node15479 = (inp[1]) ? 4'b1011 : node15480;
															assign node15480 = (inp[2]) ? 4'b1110 : 4'b1011;
														assign node15484 = (inp[2]) ? node15488 : node15485;
															assign node15485 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node15488 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node15491 = (inp[2]) ? node15495 : node15492;
														assign node15492 = (inp[1]) ? 4'b1111 : 4'b1011;
														assign node15495 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node15498 = (inp[13]) ? node15520 : node15499;
													assign node15499 = (inp[11]) ? node15509 : node15500;
														assign node15500 = (inp[9]) ? node15504 : node15501;
															assign node15501 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node15504 = (inp[2]) ? node15506 : 4'b1010;
																assign node15506 = (inp[1]) ? 4'b1010 : 4'b1111;
														assign node15509 = (inp[9]) ? node15515 : node15510;
															assign node15510 = (inp[2]) ? 4'b1011 : node15511;
																assign node15511 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node15515 = (inp[2]) ? node15517 : 4'b1111;
																assign node15517 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node15520 = (inp[2]) ? node15524 : node15521;
														assign node15521 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node15524 = (inp[1]) ? 4'b1010 : node15525;
															assign node15525 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node15529 = (inp[0]) ? node15573 : node15530;
											assign node15530 = (inp[10]) ? node15550 : node15531;
												assign node15531 = (inp[2]) ? node15543 : node15532;
													assign node15532 = (inp[1]) ? node15538 : node15533;
														assign node15533 = (inp[13]) ? 4'b1001 : node15534;
															assign node15534 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node15538 = (inp[11]) ? node15540 : 4'b1100;
															assign node15540 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node15543 = (inp[1]) ? node15545 : 4'b1100;
														assign node15545 = (inp[13]) ? 4'b1000 : node15546;
															assign node15546 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node15550 = (inp[1]) ? node15562 : node15551;
													assign node15551 = (inp[2]) ? node15557 : node15552;
														assign node15552 = (inp[11]) ? node15554 : 4'b1000;
															assign node15554 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node15557 = (inp[11]) ? 4'b1101 : node15558;
															assign node15558 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node15562 = (inp[2]) ? node15568 : node15563;
														assign node15563 = (inp[11]) ? node15565 : 4'b1101;
															assign node15565 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node15568 = (inp[13]) ? 4'b1001 : node15569;
															assign node15569 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node15573 = (inp[10]) ? node15597 : node15574;
												assign node15574 = (inp[2]) ? node15586 : node15575;
													assign node15575 = (inp[1]) ? node15581 : node15576;
														assign node15576 = (inp[13]) ? 4'b1000 : node15577;
															assign node15577 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15581 = (inp[13]) ? 4'b1101 : node15582;
															assign node15582 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node15586 = (inp[1]) ? node15592 : node15587;
														assign node15587 = (inp[11]) ? 4'b1101 : node15588;
															assign node15588 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node15592 = (inp[11]) ? node15594 : 4'b1001;
															assign node15594 = (inp[13]) ? 4'b1001 : 4'b1000;
												assign node15597 = (inp[2]) ? node15609 : node15598;
													assign node15598 = (inp[1]) ? node15604 : node15599;
														assign node15599 = (inp[11]) ? node15601 : 4'b1001;
															assign node15601 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node15604 = (inp[11]) ? node15606 : 4'b1100;
															assign node15606 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node15609 = (inp[1]) ? node15615 : node15610;
														assign node15610 = (inp[13]) ? node15612 : 4'b1100;
															assign node15612 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node15615 = (inp[11]) ? node15617 : 4'b1000;
															assign node15617 = (inp[13]) ? 4'b1000 : 4'b1001;
							assign node15620 = (inp[12]) ? node16104 : node15621;
								assign node15621 = (inp[4]) ? node15891 : node15622;
									assign node15622 = (inp[1]) ? node15762 : node15623;
										assign node15623 = (inp[11]) ? node15663 : node15624;
											assign node15624 = (inp[10]) ? node15648 : node15625;
												assign node15625 = (inp[0]) ? node15633 : node15626;
													assign node15626 = (inp[14]) ? node15630 : node15627;
														assign node15627 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node15630 = (inp[2]) ? 4'b1000 : 4'b1101;
													assign node15633 = (inp[9]) ? node15643 : node15634;
														assign node15634 = (inp[13]) ? 4'b1001 : node15635;
															assign node15635 = (inp[14]) ? node15639 : node15636;
																assign node15636 = (inp[2]) ? 4'b1100 : 4'b1000;
																assign node15639 = (inp[2]) ? 4'b1001 : 4'b1100;
														assign node15643 = (inp[14]) ? 4'b1100 : node15644;
															assign node15644 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node15648 = (inp[0]) ? node15656 : node15649;
													assign node15649 = (inp[14]) ? node15653 : node15650;
														assign node15650 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node15653 = (inp[2]) ? 4'b1001 : 4'b1100;
													assign node15656 = (inp[14]) ? node15660 : node15657;
														assign node15657 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node15660 = (inp[2]) ? 4'b1000 : 4'b1101;
											assign node15663 = (inp[10]) ? node15715 : node15664;
												assign node15664 = (inp[2]) ? node15688 : node15665;
													assign node15665 = (inp[14]) ? node15673 : node15666;
														assign node15666 = (inp[0]) ? node15670 : node15667;
															assign node15667 = (inp[13]) ? 4'b1001 : 4'b1000;
															assign node15670 = (inp[13]) ? 4'b1000 : 4'b1001;
														assign node15673 = (inp[9]) ? node15681 : node15674;
															assign node15674 = (inp[0]) ? node15678 : node15675;
																assign node15675 = (inp[13]) ? 4'b1100 : 4'b1101;
																assign node15678 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node15681 = (inp[0]) ? node15685 : node15682;
																assign node15682 = (inp[13]) ? 4'b1100 : 4'b1101;
																assign node15685 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node15688 = (inp[14]) ? node15702 : node15689;
														assign node15689 = (inp[9]) ? node15697 : node15690;
															assign node15690 = (inp[13]) ? node15694 : node15691;
																assign node15691 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node15694 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node15697 = (inp[0]) ? 4'b1100 : node15698;
																assign node15698 = (inp[13]) ? 4'b1101 : 4'b1100;
														assign node15702 = (inp[9]) ? node15708 : node15703;
															assign node15703 = (inp[13]) ? node15705 : 4'b1000;
																assign node15705 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node15708 = (inp[0]) ? node15712 : node15709;
																assign node15709 = (inp[13]) ? 4'b1001 : 4'b1000;
																assign node15712 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node15715 = (inp[2]) ? node15739 : node15716;
													assign node15716 = (inp[14]) ? node15732 : node15717;
														assign node15717 = (inp[9]) ? node15725 : node15718;
															assign node15718 = (inp[13]) ? node15722 : node15719;
																assign node15719 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node15722 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node15725 = (inp[13]) ? node15729 : node15726;
																assign node15726 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node15729 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node15732 = (inp[0]) ? node15736 : node15733;
															assign node15733 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node15736 = (inp[13]) ? 4'b1100 : 4'b1101;
													assign node15739 = (inp[14]) ? node15755 : node15740;
														assign node15740 = (inp[9]) ? node15748 : node15741;
															assign node15741 = (inp[0]) ? node15745 : node15742;
																assign node15742 = (inp[13]) ? 4'b1100 : 4'b1101;
																assign node15745 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node15748 = (inp[13]) ? node15752 : node15749;
																assign node15749 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node15752 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node15755 = (inp[0]) ? node15759 : node15756;
															assign node15756 = (inp[13]) ? 4'b1000 : 4'b1001;
															assign node15759 = (inp[13]) ? 4'b1001 : 4'b1000;
										assign node15762 = (inp[14]) ? node15816 : node15763;
											assign node15763 = (inp[2]) ? node15795 : node15764;
												assign node15764 = (inp[9]) ? node15774 : node15765;
													assign node15765 = (inp[11]) ? node15767 : 4'b1101;
														assign node15767 = (inp[0]) ? node15771 : node15768;
															assign node15768 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node15771 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node15774 = (inp[0]) ? node15786 : node15775;
														assign node15775 = (inp[10]) ? node15781 : node15776;
															assign node15776 = (inp[11]) ? 4'b1100 : node15777;
																assign node15777 = (inp[13]) ? 4'b1101 : 4'b1100;
															assign node15781 = (inp[11]) ? 4'b1101 : node15782;
																assign node15782 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node15786 = (inp[10]) ? node15790 : node15787;
															assign node15787 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node15790 = (inp[13]) ? node15792 : 4'b1100;
																assign node15792 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node15795 = (inp[0]) ? node15807 : node15796;
													assign node15796 = (inp[10]) ? node15802 : node15797;
														assign node15797 = (inp[13]) ? 4'b1000 : node15798;
															assign node15798 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node15802 = (inp[13]) ? 4'b1001 : node15803;
															assign node15803 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node15807 = (inp[10]) ? node15813 : node15808;
														assign node15808 = (inp[11]) ? node15810 : 4'b1001;
															assign node15810 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node15813 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node15816 = (inp[2]) ? node15848 : node15817;
												assign node15817 = (inp[13]) ? node15825 : node15818;
													assign node15818 = (inp[0]) ? node15822 : node15819;
														assign node15819 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node15822 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node15825 = (inp[11]) ? node15841 : node15826;
														assign node15826 = (inp[9]) ? node15834 : node15827;
															assign node15827 = (inp[10]) ? node15831 : node15828;
																assign node15828 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node15831 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node15834 = (inp[10]) ? node15838 : node15835;
																assign node15835 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node15838 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node15841 = (inp[0]) ? node15845 : node15842;
															assign node15842 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node15845 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node15848 = (inp[11]) ? node15870 : node15849;
													assign node15849 = (inp[0]) ? node15855 : node15850;
														assign node15850 = (inp[10]) ? 4'b1100 : node15851;
															assign node15851 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node15855 = (inp[9]) ? node15863 : node15856;
															assign node15856 = (inp[10]) ? node15860 : node15857;
																assign node15857 = (inp[13]) ? 4'b1101 : 4'b1100;
																assign node15860 = (inp[13]) ? 4'b1100 : 4'b1101;
															assign node15863 = (inp[13]) ? node15867 : node15864;
																assign node15864 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node15867 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node15870 = (inp[9]) ? node15878 : node15871;
														assign node15871 = (inp[0]) ? node15875 : node15872;
															assign node15872 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node15875 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node15878 = (inp[13]) ? node15884 : node15879;
															assign node15879 = (inp[0]) ? 4'b1100 : node15880;
																assign node15880 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node15884 = (inp[0]) ? node15888 : node15885;
																assign node15885 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node15888 = (inp[10]) ? 4'b1100 : 4'b1101;
									assign node15891 = (inp[1]) ? node15981 : node15892;
										assign node15892 = (inp[2]) ? node15928 : node15893;
											assign node15893 = (inp[10]) ? node15911 : node15894;
												assign node15894 = (inp[0]) ? node15902 : node15895;
													assign node15895 = (inp[13]) ? node15897 : 4'b1010;
														assign node15897 = (inp[14]) ? node15899 : 4'b1010;
															assign node15899 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node15902 = (inp[13]) ? node15904 : 4'b1011;
														assign node15904 = (inp[14]) ? node15908 : node15905;
															assign node15905 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node15908 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node15911 = (inp[0]) ? node15921 : node15912;
													assign node15912 = (inp[13]) ? node15914 : 4'b1011;
														assign node15914 = (inp[11]) ? node15918 : node15915;
															assign node15915 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node15918 = (inp[14]) ? 4'b1010 : 4'b1011;
													assign node15921 = (inp[13]) ? node15923 : 4'b1010;
														assign node15923 = (inp[14]) ? 4'b1011 : node15924;
															assign node15924 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node15928 = (inp[11]) ? node15960 : node15929;
												assign node15929 = (inp[13]) ? node15945 : node15930;
													assign node15930 = (inp[9]) ? node15932 : 4'b1111;
														assign node15932 = (inp[0]) ? node15938 : node15933;
															assign node15933 = (inp[14]) ? 4'b1111 : node15934;
																assign node15934 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node15938 = (inp[10]) ? node15942 : node15939;
																assign node15939 = (inp[14]) ? 4'b1111 : 4'b1110;
																assign node15942 = (inp[14]) ? 4'b1110 : 4'b1111;
													assign node15945 = (inp[0]) ? node15953 : node15946;
														assign node15946 = (inp[14]) ? node15950 : node15947;
															assign node15947 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node15950 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node15953 = (inp[14]) ? node15957 : node15954;
															assign node15954 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node15957 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node15960 = (inp[14]) ? node15968 : node15961;
													assign node15961 = (inp[10]) ? node15965 : node15962;
														assign node15962 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node15965 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node15968 = (inp[9]) ? node15976 : node15969;
														assign node15969 = (inp[13]) ? 4'b1110 : node15970;
															assign node15970 = (inp[10]) ? node15972 : 4'b1111;
																assign node15972 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node15976 = (inp[0]) ? 4'b1110 : node15977;
															assign node15977 = (inp[10]) ? 4'b1110 : 4'b1111;
										assign node15981 = (inp[2]) ? node16043 : node15982;
											assign node15982 = (inp[14]) ? node16022 : node15983;
												assign node15983 = (inp[9]) ? node16005 : node15984;
													assign node15984 = (inp[10]) ? node15994 : node15985;
														assign node15985 = (inp[11]) ? node15987 : 4'b1110;
															assign node15987 = (inp[13]) ? node15991 : node15988;
																assign node15988 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node15991 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node15994 = (inp[0]) ? node16000 : node15995;
															assign node15995 = (inp[13]) ? 4'b1111 : node15996;
																assign node15996 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node16000 = (inp[11]) ? node16002 : 4'b1110;
																assign node16002 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node16005 = (inp[11]) ? node16013 : node16006;
														assign node16006 = (inp[0]) ? node16010 : node16007;
															assign node16007 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node16010 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node16013 = (inp[0]) ? 4'b1111 : node16014;
															assign node16014 = (inp[13]) ? node16018 : node16015;
																assign node16015 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node16018 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node16022 = (inp[10]) ? node16034 : node16023;
													assign node16023 = (inp[0]) ? node16029 : node16024;
														assign node16024 = (inp[11]) ? 4'b1110 : node16025;
															assign node16025 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node16029 = (inp[11]) ? 4'b1111 : node16030;
															assign node16030 = (inp[13]) ? 4'b1111 : 4'b1110;
													assign node16034 = (inp[11]) ? 4'b1110 : node16035;
														assign node16035 = (inp[13]) ? node16039 : node16036;
															assign node16036 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node16039 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node16043 = (inp[9]) ? node16073 : node16044;
												assign node16044 = (inp[11]) ? node16062 : node16045;
													assign node16045 = (inp[0]) ? node16051 : node16046;
														assign node16046 = (inp[13]) ? 4'b1010 : node16047;
															assign node16047 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node16051 = (inp[13]) ? node16057 : node16052;
															assign node16052 = (inp[14]) ? node16054 : 4'b1010;
																assign node16054 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node16057 = (inp[14]) ? node16059 : 4'b1011;
																assign node16059 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node16062 = (inp[13]) ? 4'b1010 : node16063;
														assign node16063 = (inp[14]) ? node16065 : 4'b1010;
															assign node16065 = (inp[10]) ? node16069 : node16066;
																assign node16066 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node16069 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node16073 = (inp[10]) ? node16089 : node16074;
													assign node16074 = (inp[0]) ? node16082 : node16075;
														assign node16075 = (inp[11]) ? 4'b1010 : node16076;
															assign node16076 = (inp[13]) ? node16078 : 4'b1010;
																assign node16078 = (inp[14]) ? 4'b1010 : 4'b1011;
														assign node16082 = (inp[11]) ? 4'b1011 : node16083;
															assign node16083 = (inp[14]) ? 4'b1010 : node16084;
																assign node16084 = (inp[13]) ? 4'b1010 : 4'b1011;
													assign node16089 = (inp[0]) ? node16095 : node16090;
														assign node16090 = (inp[14]) ? 4'b1011 : node16091;
															assign node16091 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node16095 = (inp[11]) ? 4'b1010 : node16096;
															assign node16096 = (inp[13]) ? node16100 : node16097;
																assign node16097 = (inp[14]) ? 4'b1011 : 4'b1010;
																assign node16100 = (inp[14]) ? 4'b1010 : 4'b1011;
								assign node16104 = (inp[4]) ? node16296 : node16105;
									assign node16105 = (inp[10]) ? node16211 : node16106;
										assign node16106 = (inp[0]) ? node16164 : node16107;
											assign node16107 = (inp[13]) ? node16143 : node16108;
												assign node16108 = (inp[14]) ? node16130 : node16109;
													assign node16109 = (inp[11]) ? node16117 : node16110;
														assign node16110 = (inp[1]) ? node16114 : node16111;
															assign node16111 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node16114 = (inp[2]) ? 4'b1010 : 4'b1111;
														assign node16117 = (inp[9]) ? node16123 : node16118;
															assign node16118 = (inp[2]) ? node16120 : 4'b1110;
																assign node16120 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node16123 = (inp[2]) ? node16127 : node16124;
																assign node16124 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node16127 = (inp[1]) ? 4'b1010 : 4'b1110;
													assign node16130 = (inp[2]) ? node16136 : node16131;
														assign node16131 = (inp[1]) ? node16133 : 4'b1010;
															assign node16133 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node16136 = (inp[11]) ? node16140 : node16137;
															assign node16137 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node16140 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node16143 = (inp[2]) ? node16153 : node16144;
													assign node16144 = (inp[1]) ? 4'b1111 : node16145;
														assign node16145 = (inp[9]) ? node16147 : 4'b1011;
															assign node16147 = (inp[14]) ? node16149 : 4'b1010;
																assign node16149 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node16153 = (inp[1]) ? node16159 : node16154;
														assign node16154 = (inp[14]) ? 4'b1110 : node16155;
															assign node16155 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node16159 = (inp[14]) ? 4'b1010 : node16160;
															assign node16160 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node16164 = (inp[11]) ? node16198 : node16165;
												assign node16165 = (inp[14]) ? node16185 : node16166;
													assign node16166 = (inp[13]) ? node16174 : node16167;
														assign node16167 = (inp[2]) ? node16171 : node16168;
															assign node16168 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node16171 = (inp[1]) ? 4'b1011 : 4'b1111;
														assign node16174 = (inp[9]) ? node16180 : node16175;
															assign node16175 = (inp[1]) ? 4'b1010 : node16176;
																assign node16176 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node16180 = (inp[1]) ? node16182 : 4'b1010;
																assign node16182 = (inp[2]) ? 4'b1010 : 4'b1110;
													assign node16185 = (inp[2]) ? node16191 : node16186;
														assign node16186 = (inp[1]) ? node16188 : 4'b1011;
															assign node16188 = (inp[13]) ? 4'b1110 : 4'b1111;
														assign node16191 = (inp[13]) ? node16195 : node16192;
															assign node16192 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node16195 = (inp[1]) ? 4'b1011 : 4'b1111;
												assign node16198 = (inp[2]) ? node16208 : node16199;
													assign node16199 = (inp[1]) ? node16205 : node16200;
														assign node16200 = (inp[13]) ? node16202 : 4'b1011;
															assign node16202 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node16205 = (inp[13]) ? 4'b1110 : 4'b1111;
													assign node16208 = (inp[1]) ? 4'b1011 : 4'b1111;
										assign node16211 = (inp[0]) ? node16253 : node16212;
											assign node16212 = (inp[13]) ? node16234 : node16213;
												assign node16213 = (inp[11]) ? node16225 : node16214;
													assign node16214 = (inp[2]) ? node16220 : node16215;
														assign node16215 = (inp[1]) ? node16217 : 4'b1011;
															assign node16217 = (inp[14]) ? 4'b1111 : 4'b1110;
														assign node16220 = (inp[14]) ? 4'b1110 : node16221;
															assign node16221 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node16225 = (inp[1]) ? node16229 : node16226;
														assign node16226 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node16229 = (inp[2]) ? 4'b1011 : node16230;
															assign node16230 = (inp[14]) ? 4'b1110 : 4'b1111;
												assign node16234 = (inp[2]) ? node16242 : node16235;
													assign node16235 = (inp[1]) ? 4'b1110 : node16236;
														assign node16236 = (inp[14]) ? 4'b1010 : node16237;
															assign node16237 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node16242 = (inp[1]) ? node16248 : node16243;
														assign node16243 = (inp[14]) ? 4'b1111 : node16244;
															assign node16244 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node16248 = (inp[11]) ? 4'b1011 : node16249;
															assign node16249 = (inp[14]) ? 4'b1011 : 4'b1010;
											assign node16253 = (inp[13]) ? node16269 : node16254;
												assign node16254 = (inp[2]) ? node16258 : node16255;
													assign node16255 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node16258 = (inp[1]) ? node16264 : node16259;
														assign node16259 = (inp[11]) ? 4'b1110 : node16260;
															assign node16260 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node16264 = (inp[9]) ? 4'b1010 : node16265;
															assign node16265 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node16269 = (inp[2]) ? node16285 : node16270;
													assign node16270 = (inp[1]) ? 4'b1111 : node16271;
														assign node16271 = (inp[9]) ? node16279 : node16272;
															assign node16272 = (inp[11]) ? node16276 : node16273;
																assign node16273 = (inp[14]) ? 4'b1010 : 4'b1011;
																assign node16276 = (inp[14]) ? 4'b1011 : 4'b1010;
															assign node16279 = (inp[14]) ? node16281 : 4'b1010;
																assign node16281 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node16285 = (inp[1]) ? node16291 : node16286;
														assign node16286 = (inp[11]) ? 4'b1110 : node16287;
															assign node16287 = (inp[14]) ? 4'b1110 : 4'b1111;
														assign node16291 = (inp[11]) ? 4'b1010 : node16292;
															assign node16292 = (inp[14]) ? 4'b1010 : 4'b1011;
									assign node16296 = (inp[9]) ? node16430 : node16297;
										assign node16297 = (inp[10]) ? node16369 : node16298;
											assign node16298 = (inp[0]) ? node16330 : node16299;
												assign node16299 = (inp[1]) ? node16317 : node16300;
													assign node16300 = (inp[2]) ? node16310 : node16301;
														assign node16301 = (inp[13]) ? node16303 : 4'b1001;
															assign node16303 = (inp[11]) ? node16307 : node16304;
																assign node16304 = (inp[14]) ? 4'b1001 : 4'b1000;
																assign node16307 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node16310 = (inp[11]) ? 4'b1100 : node16311;
															assign node16311 = (inp[13]) ? 4'b1101 : node16312;
																assign node16312 = (inp[14]) ? 4'b1101 : 4'b1100;
													assign node16317 = (inp[2]) ? node16325 : node16318;
														assign node16318 = (inp[11]) ? node16320 : 4'b1100;
															assign node16320 = (inp[14]) ? 4'b1100 : node16321;
																assign node16321 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node16325 = (inp[11]) ? 4'b1000 : node16326;
															assign node16326 = (inp[13]) ? 4'b1000 : 4'b1001;
												assign node16330 = (inp[13]) ? node16348 : node16331;
													assign node16331 = (inp[2]) ? node16339 : node16332;
														assign node16332 = (inp[1]) ? node16334 : 4'b1000;
															assign node16334 = (inp[11]) ? 4'b1100 : node16335;
																assign node16335 = (inp[14]) ? 4'b1100 : 4'b1101;
														assign node16339 = (inp[1]) ? node16343 : node16340;
															assign node16340 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node16343 = (inp[14]) ? node16345 : 4'b1001;
																assign node16345 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node16348 = (inp[11]) ? node16360 : node16349;
														assign node16349 = (inp[2]) ? node16355 : node16350;
															assign node16350 = (inp[14]) ? 4'b1000 : node16351;
																assign node16351 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node16355 = (inp[1]) ? node16357 : 4'b1101;
																assign node16357 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node16360 = (inp[1]) ? node16366 : node16361;
															assign node16361 = (inp[14]) ? node16363 : 4'b1000;
																assign node16363 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node16366 = (inp[2]) ? 4'b1001 : 4'b1101;
											assign node16369 = (inp[11]) ? node16403 : node16370;
												assign node16370 = (inp[0]) ? node16384 : node16371;
													assign node16371 = (inp[1]) ? node16375 : node16372;
														assign node16372 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node16375 = (inp[2]) ? node16379 : node16376;
															assign node16376 = (inp[14]) ? 4'b1100 : 4'b1101;
															assign node16379 = (inp[13]) ? 4'b1000 : node16380;
																assign node16380 = (inp[14]) ? 4'b1000 : 4'b1001;
													assign node16384 = (inp[13]) ? node16392 : node16385;
														assign node16385 = (inp[14]) ? 4'b1001 : node16386;
															assign node16386 = (inp[1]) ? node16388 : 4'b1001;
																assign node16388 = (inp[2]) ? 4'b1000 : 4'b1100;
														assign node16392 = (inp[1]) ? node16398 : node16393;
															assign node16393 = (inp[2]) ? 4'b1100 : node16394;
																assign node16394 = (inp[14]) ? 4'b1001 : 4'b1000;
															assign node16398 = (inp[2]) ? node16400 : 4'b1100;
																assign node16400 = (inp[14]) ? 4'b1000 : 4'b1001;
												assign node16403 = (inp[0]) ? node16415 : node16404;
													assign node16404 = (inp[2]) ? node16412 : node16405;
														assign node16405 = (inp[1]) ? 4'b1101 : node16406;
															assign node16406 = (inp[14]) ? node16408 : 4'b1000;
																assign node16408 = (inp[13]) ? 4'b1001 : 4'b1000;
														assign node16412 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node16415 = (inp[2]) ? node16427 : node16416;
														assign node16416 = (inp[1]) ? node16422 : node16417;
															assign node16417 = (inp[13]) ? node16419 : 4'b1001;
																assign node16419 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node16422 = (inp[14]) ? 4'b1100 : node16423;
																assign node16423 = (inp[13]) ? 4'b1100 : 4'b1101;
														assign node16427 = (inp[1]) ? 4'b1000 : 4'b1100;
										assign node16430 = (inp[13]) ? node16500 : node16431;
											assign node16431 = (inp[1]) ? node16457 : node16432;
												assign node16432 = (inp[2]) ? node16440 : node16433;
													assign node16433 = (inp[0]) ? node16437 : node16434;
														assign node16434 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node16437 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node16440 = (inp[14]) ? node16448 : node16441;
														assign node16441 = (inp[0]) ? node16445 : node16442;
															assign node16442 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node16445 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node16448 = (inp[10]) ? node16450 : 4'b1101;
															assign node16450 = (inp[0]) ? node16454 : node16451;
																assign node16451 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node16454 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node16457 = (inp[2]) ? node16477 : node16458;
													assign node16458 = (inp[0]) ? node16466 : node16459;
														assign node16459 = (inp[10]) ? node16461 : 4'b1101;
															assign node16461 = (inp[14]) ? 4'b1101 : node16462;
																assign node16462 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node16466 = (inp[11]) ? node16472 : node16467;
															assign node16467 = (inp[14]) ? node16469 : 4'b1100;
																assign node16469 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node16472 = (inp[14]) ? node16474 : 4'b1101;
																assign node16474 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node16477 = (inp[0]) ? node16489 : node16478;
														assign node16478 = (inp[10]) ? node16484 : node16479;
															assign node16479 = (inp[14]) ? node16481 : 4'b1000;
																assign node16481 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node16484 = (inp[11]) ? 4'b1001 : node16485;
																assign node16485 = (inp[14]) ? 4'b1000 : 4'b1001;
														assign node16489 = (inp[10]) ? node16495 : node16490;
															assign node16490 = (inp[11]) ? 4'b1001 : node16491;
																assign node16491 = (inp[14]) ? 4'b1000 : 4'b1001;
															assign node16495 = (inp[11]) ? 4'b1000 : node16496;
																assign node16496 = (inp[14]) ? 4'b1001 : 4'b1000;
											assign node16500 = (inp[2]) ? node16534 : node16501;
												assign node16501 = (inp[1]) ? node16513 : node16502;
													assign node16502 = (inp[0]) ? 4'b1000 : node16503;
														assign node16503 = (inp[14]) ? node16505 : 4'b1000;
															assign node16505 = (inp[10]) ? node16509 : node16506;
																assign node16506 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node16509 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node16513 = (inp[11]) ? node16527 : node16514;
														assign node16514 = (inp[14]) ? node16522 : node16515;
															assign node16515 = (inp[0]) ? node16519 : node16516;
																assign node16516 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node16519 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node16522 = (inp[0]) ? 4'b1101 : node16523;
																assign node16523 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node16527 = (inp[14]) ? node16529 : 4'b1100;
															assign node16529 = (inp[10]) ? 4'b1100 : node16530;
																assign node16530 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node16534 = (inp[1]) ? node16546 : node16535;
													assign node16535 = (inp[10]) ? node16541 : node16536;
														assign node16536 = (inp[14]) ? node16538 : 4'b1101;
															assign node16538 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node16541 = (inp[0]) ? 4'b1100 : node16542;
															assign node16542 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node16546 = (inp[11]) ? node16554 : node16547;
														assign node16547 = (inp[0]) ? node16549 : 4'b1001;
															assign node16549 = (inp[10]) ? 4'b1001 : node16550;
																assign node16550 = (inp[14]) ? 4'b1001 : 4'b1000;
														assign node16554 = (inp[0]) ? node16558 : node16555;
															assign node16555 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node16558 = (inp[10]) ? 4'b1000 : 4'b1001;
			assign node16561 = (inp[14]) ? node23099 : node16562;
				assign node16562 = (inp[8]) ? node19914 : node16563;
					assign node16563 = (inp[12]) ? node17945 : node16564;
						assign node16564 = (inp[4]) ? node17276 : node16565;
							assign node16565 = (inp[11]) ? node16931 : node16566;
								assign node16566 = (inp[9]) ? node16742 : node16567;
									assign node16567 = (inp[2]) ? node16647 : node16568;
										assign node16568 = (inp[5]) ? node16600 : node16569;
											assign node16569 = (inp[13]) ? node16583 : node16570;
												assign node16570 = (inp[15]) ? node16574 : node16571;
													assign node16571 = (inp[7]) ? 4'b1010 : 4'b1000;
													assign node16574 = (inp[7]) ? node16580 : node16575;
														assign node16575 = (inp[1]) ? node16577 : 4'b1010;
															assign node16577 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node16580 = (inp[1]) ? 4'b1001 : 4'b1100;
												assign node16583 = (inp[0]) ? node16591 : node16584;
													assign node16584 = (inp[15]) ? node16588 : node16585;
														assign node16585 = (inp[7]) ? 4'b1110 : 4'b1100;
														assign node16588 = (inp[7]) ? 4'b1100 : 4'b1111;
													assign node16591 = (inp[15]) ? node16595 : node16592;
														assign node16592 = (inp[7]) ? 4'b1110 : 4'b1100;
														assign node16595 = (inp[1]) ? node16597 : 4'b1000;
															assign node16597 = (inp[7]) ? 4'b1100 : 4'b1110;
											assign node16600 = (inp[13]) ? node16616 : node16601;
												assign node16601 = (inp[15]) ? node16605 : node16602;
													assign node16602 = (inp[7]) ? 4'b1111 : 4'b1100;
													assign node16605 = (inp[7]) ? node16611 : node16606;
														assign node16606 = (inp[1]) ? node16608 : 4'b1110;
															assign node16608 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node16611 = (inp[1]) ? 4'b1100 : node16612;
															assign node16612 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node16616 = (inp[1]) ? node16632 : node16617;
													assign node16617 = (inp[7]) ? node16625 : node16618;
														assign node16618 = (inp[15]) ? node16622 : node16619;
															assign node16619 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node16622 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node16625 = (inp[15]) ? node16629 : node16626;
															assign node16626 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node16629 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node16632 = (inp[0]) ? node16640 : node16633;
														assign node16633 = (inp[7]) ? node16637 : node16634;
															assign node16634 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node16637 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node16640 = (inp[15]) ? node16644 : node16641;
															assign node16641 = (inp[7]) ? 4'b1010 : 4'b1001;
															assign node16644 = (inp[7]) ? 4'b1000 : 4'b1010;
										assign node16647 = (inp[0]) ? node16695 : node16648;
											assign node16648 = (inp[13]) ? node16670 : node16649;
												assign node16649 = (inp[5]) ? node16659 : node16650;
													assign node16650 = (inp[15]) ? node16654 : node16651;
														assign node16651 = (inp[7]) ? 4'b1010 : 4'b1000;
														assign node16654 = (inp[1]) ? node16656 : 4'b1100;
															assign node16656 = (inp[7]) ? 4'b1001 : 4'b1011;
													assign node16659 = (inp[15]) ? node16663 : node16660;
														assign node16660 = (inp[7]) ? 4'b1111 : 4'b1100;
														assign node16663 = (inp[7]) ? node16667 : node16664;
															assign node16664 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node16667 = (inp[1]) ? 4'b1100 : 4'b1000;
												assign node16670 = (inp[5]) ? node16680 : node16671;
													assign node16671 = (inp[15]) ? node16675 : node16672;
														assign node16672 = (inp[7]) ? 4'b1110 : 4'b1100;
														assign node16675 = (inp[7]) ? 4'b1000 : node16676;
															assign node16676 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node16680 = (inp[1]) ? node16688 : node16681;
														assign node16681 = (inp[15]) ? node16685 : node16682;
															assign node16682 = (inp[7]) ? 4'b1010 : 4'b1001;
															assign node16685 = (inp[7]) ? 4'b1101 : 4'b1010;
														assign node16688 = (inp[7]) ? node16692 : node16689;
															assign node16689 = (inp[15]) ? 4'b1010 : 4'b1001;
															assign node16692 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node16695 = (inp[7]) ? node16719 : node16696;
												assign node16696 = (inp[15]) ? node16710 : node16697;
													assign node16697 = (inp[1]) ? 4'b1001 : node16698;
														assign node16698 = (inp[10]) ? node16704 : node16699;
															assign node16699 = (inp[13]) ? node16701 : 4'b1001;
																assign node16701 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node16704 = (inp[5]) ? node16706 : 4'b1001;
																assign node16706 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node16710 = (inp[13]) ? node16714 : node16711;
														assign node16711 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node16714 = (inp[5]) ? node16716 : 4'b1110;
															assign node16716 = (inp[1]) ? 4'b1011 : 4'b1010;
												assign node16719 = (inp[15]) ? node16727 : node16720;
													assign node16720 = (inp[5]) ? node16724 : node16721;
														assign node16721 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node16724 = (inp[13]) ? 4'b1010 : 4'b1110;
													assign node16727 = (inp[13]) ? node16735 : node16728;
														assign node16728 = (inp[1]) ? node16732 : node16729;
															assign node16729 = (inp[5]) ? 4'b1000 : 4'b1101;
															assign node16732 = (inp[5]) ? 4'b1101 : 4'b1000;
														assign node16735 = (inp[5]) ? node16739 : node16736;
															assign node16736 = (inp[1]) ? 4'b1101 : 4'b1000;
															assign node16739 = (inp[1]) ? 4'b1000 : 4'b1101;
									assign node16742 = (inp[0]) ? node16832 : node16743;
										assign node16743 = (inp[7]) ? node16775 : node16744;
											assign node16744 = (inp[15]) ? node16754 : node16745;
												assign node16745 = (inp[5]) ? node16749 : node16746;
													assign node16746 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node16749 = (inp[13]) ? node16751 : 4'b1101;
														assign node16751 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node16754 = (inp[5]) ? node16764 : node16755;
													assign node16755 = (inp[13]) ? node16759 : node16756;
														assign node16756 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node16759 = (inp[2]) ? node16761 : 4'b1110;
															assign node16761 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node16764 = (inp[13]) ? node16770 : node16765;
														assign node16765 = (inp[2]) ? node16767 : 4'b1111;
															assign node16767 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node16770 = (inp[2]) ? 4'b1011 : node16771;
															assign node16771 = (inp[1]) ? 4'b1011 : 4'b1010;
											assign node16775 = (inp[15]) ? node16785 : node16776;
												assign node16776 = (inp[5]) ? node16780 : node16777;
													assign node16777 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node16780 = (inp[13]) ? node16782 : 4'b1110;
														assign node16782 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node16785 = (inp[2]) ? node16807 : node16786;
													assign node16786 = (inp[1]) ? node16794 : node16787;
														assign node16787 = (inp[5]) ? node16791 : node16788;
															assign node16788 = (inp[13]) ? 4'b1000 : 4'b1101;
															assign node16791 = (inp[13]) ? 4'b1101 : 4'b1000;
														assign node16794 = (inp[10]) ? node16802 : node16795;
															assign node16795 = (inp[13]) ? node16799 : node16796;
																assign node16796 = (inp[5]) ? 4'b1101 : 4'b1000;
																assign node16799 = (inp[5]) ? 4'b1000 : 4'b1101;
															assign node16802 = (inp[5]) ? 4'b1101 : node16803;
																assign node16803 = (inp[13]) ? 4'b1101 : 4'b1000;
													assign node16807 = (inp[10]) ? node16817 : node16808;
														assign node16808 = (inp[1]) ? node16810 : 4'b1001;
															assign node16810 = (inp[5]) ? node16814 : node16811;
																assign node16811 = (inp[13]) ? 4'b1101 : 4'b1000;
																assign node16814 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node16817 = (inp[5]) ? node16825 : node16818;
															assign node16818 = (inp[1]) ? node16822 : node16819;
																assign node16819 = (inp[13]) ? 4'b1001 : 4'b1101;
																assign node16822 = (inp[13]) ? 4'b1101 : 4'b1000;
															assign node16825 = (inp[13]) ? node16829 : node16826;
																assign node16826 = (inp[1]) ? 4'b1101 : 4'b1001;
																assign node16829 = (inp[1]) ? 4'b1001 : 4'b1100;
										assign node16832 = (inp[2]) ? node16878 : node16833;
											assign node16833 = (inp[7]) ? node16855 : node16834;
												assign node16834 = (inp[15]) ? node16842 : node16835;
													assign node16835 = (inp[5]) ? node16839 : node16836;
														assign node16836 = (inp[13]) ? 4'b1101 : 4'b1001;
														assign node16839 = (inp[13]) ? 4'b1000 : 4'b1101;
													assign node16842 = (inp[5]) ? node16850 : node16843;
														assign node16843 = (inp[13]) ? node16847 : node16844;
															assign node16844 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node16847 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node16850 = (inp[13]) ? 4'b1011 : node16851;
															assign node16851 = (inp[1]) ? 4'b1110 : 4'b1111;
												assign node16855 = (inp[15]) ? node16863 : node16856;
													assign node16856 = (inp[13]) ? node16860 : node16857;
														assign node16857 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node16860 = (inp[5]) ? 4'b1011 : 4'b1111;
													assign node16863 = (inp[1]) ? node16871 : node16864;
														assign node16864 = (inp[13]) ? node16868 : node16865;
															assign node16865 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node16868 = (inp[5]) ? 4'b1100 : 4'b1001;
														assign node16871 = (inp[5]) ? node16875 : node16872;
															assign node16872 = (inp[13]) ? 4'b1101 : 4'b1000;
															assign node16875 = (inp[13]) ? 4'b1001 : 4'b1101;
											assign node16878 = (inp[7]) ? node16896 : node16879;
												assign node16879 = (inp[15]) ? node16887 : node16880;
													assign node16880 = (inp[13]) ? node16884 : node16881;
														assign node16881 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node16884 = (inp[5]) ? 4'b1000 : 4'b1100;
													assign node16887 = (inp[13]) ? node16891 : node16888;
														assign node16888 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node16891 = (inp[5]) ? node16893 : 4'b1111;
															assign node16893 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node16896 = (inp[15]) ? node16904 : node16897;
													assign node16897 = (inp[5]) ? node16901 : node16898;
														assign node16898 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node16901 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node16904 = (inp[10]) ? node16918 : node16905;
														assign node16905 = (inp[1]) ? node16913 : node16906;
															assign node16906 = (inp[5]) ? node16910 : node16907;
																assign node16907 = (inp[13]) ? 4'b1001 : 4'b1100;
																assign node16910 = (inp[13]) ? 4'b1100 : 4'b1001;
															assign node16913 = (inp[13]) ? node16915 : 4'b1001;
																assign node16915 = (inp[5]) ? 4'b1001 : 4'b1100;
														assign node16918 = (inp[13]) ? node16926 : node16919;
															assign node16919 = (inp[5]) ? node16923 : node16920;
																assign node16920 = (inp[1]) ? 4'b1001 : 4'b1100;
																assign node16923 = (inp[1]) ? 4'b1100 : 4'b1001;
															assign node16926 = (inp[1]) ? 4'b1100 : node16927;
																assign node16927 = (inp[5]) ? 4'b1100 : 4'b1001;
								assign node16931 = (inp[9]) ? node17093 : node16932;
									assign node16932 = (inp[2]) ? node16998 : node16933;
										assign node16933 = (inp[15]) ? node16953 : node16934;
											assign node16934 = (inp[7]) ? node16944 : node16935;
												assign node16935 = (inp[5]) ? node16939 : node16936;
													assign node16936 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node16939 = (inp[13]) ? node16941 : 4'b1101;
														assign node16941 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node16944 = (inp[5]) ? node16948 : node16945;
													assign node16945 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node16948 = (inp[13]) ? node16950 : 4'b1110;
														assign node16950 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node16953 = (inp[7]) ? node16975 : node16954;
												assign node16954 = (inp[5]) ? node16966 : node16955;
													assign node16955 = (inp[13]) ? node16961 : node16956;
														assign node16956 = (inp[1]) ? node16958 : 4'b1011;
															assign node16958 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node16961 = (inp[0]) ? node16963 : 4'b1110;
															assign node16963 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node16966 = (inp[13]) ? node16970 : node16967;
														assign node16967 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node16970 = (inp[0]) ? 4'b1011 : node16971;
															assign node16971 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node16975 = (inp[13]) ? node16985 : node16976;
													assign node16976 = (inp[1]) ? node16982 : node16977;
														assign node16977 = (inp[5]) ? node16979 : 4'b1101;
															assign node16979 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node16982 = (inp[5]) ? 4'b1101 : 4'b1000;
													assign node16985 = (inp[1]) ? node16993 : node16986;
														assign node16986 = (inp[5]) ? node16990 : node16987;
															assign node16987 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node16990 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node16993 = (inp[5]) ? node16995 : 4'b1101;
															assign node16995 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node16998 = (inp[0]) ? node17052 : node16999;
											assign node16999 = (inp[13]) ? node17025 : node17000;
												assign node17000 = (inp[5]) ? node17014 : node17001;
													assign node17001 = (inp[1]) ? node17009 : node17002;
														assign node17002 = (inp[15]) ? node17006 : node17003;
															assign node17003 = (inp[7]) ? 4'b1011 : 4'b1001;
															assign node17006 = (inp[7]) ? 4'b1101 : 4'b1011;
														assign node17009 = (inp[15]) ? node17011 : 4'b1011;
															assign node17011 = (inp[7]) ? 4'b1000 : 4'b1010;
													assign node17014 = (inp[7]) ? node17020 : node17015;
														assign node17015 = (inp[15]) ? node17017 : 4'b1101;
															assign node17017 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node17020 = (inp[15]) ? node17022 : 4'b1110;
															assign node17022 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node17025 = (inp[5]) ? node17037 : node17026;
													assign node17026 = (inp[15]) ? node17030 : node17027;
														assign node17027 = (inp[7]) ? 4'b1111 : 4'b1101;
														assign node17030 = (inp[7]) ? node17034 : node17031;
															assign node17031 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node17034 = (inp[1]) ? 4'b1101 : 4'b1001;
													assign node17037 = (inp[1]) ? node17045 : node17038;
														assign node17038 = (inp[15]) ? node17042 : node17039;
															assign node17039 = (inp[7]) ? 4'b1011 : 4'b1000;
															assign node17042 = (inp[7]) ? 4'b1100 : 4'b1011;
														assign node17045 = (inp[15]) ? node17049 : node17046;
															assign node17046 = (inp[10]) ? 4'b1011 : 4'b1000;
															assign node17049 = (inp[7]) ? 4'b1001 : 4'b1011;
											assign node17052 = (inp[7]) ? node17070 : node17053;
												assign node17053 = (inp[15]) ? node17061 : node17054;
													assign node17054 = (inp[13]) ? node17058 : node17055;
														assign node17055 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node17058 = (inp[5]) ? 4'b1000 : 4'b1100;
													assign node17061 = (inp[13]) ? node17065 : node17062;
														assign node17062 = (inp[5]) ? 4'b1110 : 4'b1010;
														assign node17065 = (inp[5]) ? node17067 : 4'b1111;
															assign node17067 = (inp[1]) ? 4'b1010 : 4'b1011;
												assign node17070 = (inp[15]) ? node17078 : node17071;
													assign node17071 = (inp[5]) ? node17075 : node17072;
														assign node17072 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node17075 = (inp[13]) ? 4'b1011 : 4'b1111;
													assign node17078 = (inp[1]) ? node17086 : node17079;
														assign node17079 = (inp[13]) ? node17083 : node17080;
															assign node17080 = (inp[5]) ? 4'b1001 : 4'b1100;
															assign node17083 = (inp[5]) ? 4'b1100 : 4'b1001;
														assign node17086 = (inp[13]) ? node17090 : node17087;
															assign node17087 = (inp[5]) ? 4'b1100 : 4'b1001;
															assign node17090 = (inp[5]) ? 4'b1001 : 4'b1100;
									assign node17093 = (inp[0]) ? node17169 : node17094;
										assign node17094 = (inp[5]) ? node17120 : node17095;
											assign node17095 = (inp[13]) ? node17105 : node17096;
												assign node17096 = (inp[7]) ? node17100 : node17097;
													assign node17097 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node17100 = (inp[15]) ? node17102 : 4'b1010;
														assign node17102 = (inp[1]) ? 4'b1001 : 4'b1100;
												assign node17105 = (inp[15]) ? node17109 : node17106;
													assign node17106 = (inp[7]) ? 4'b1110 : 4'b1100;
													assign node17109 = (inp[7]) ? node17115 : node17110;
														assign node17110 = (inp[2]) ? node17112 : 4'b1111;
															assign node17112 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node17115 = (inp[1]) ? 4'b1100 : node17116;
															assign node17116 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node17120 = (inp[13]) ? node17136 : node17121;
												assign node17121 = (inp[7]) ? node17129 : node17122;
													assign node17122 = (inp[15]) ? node17124 : 4'b1100;
														assign node17124 = (inp[2]) ? node17126 : 4'b1110;
															assign node17126 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node17129 = (inp[15]) ? node17131 : 4'b1111;
														assign node17131 = (inp[1]) ? 4'b1100 : node17132;
															assign node17132 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node17136 = (inp[1]) ? node17156 : node17137;
													assign node17137 = (inp[10]) ? node17149 : node17138;
														assign node17138 = (inp[2]) ? node17142 : node17139;
															assign node17139 = (inp[7]) ? 4'b1100 : 4'b1000;
															assign node17142 = (inp[7]) ? node17146 : node17143;
																assign node17143 = (inp[15]) ? 4'b1010 : 4'b1001;
																assign node17146 = (inp[15]) ? 4'b1101 : 4'b1010;
														assign node17149 = (inp[2]) ? node17151 : 4'b1011;
															assign node17151 = (inp[7]) ? node17153 : 4'b1010;
																assign node17153 = (inp[15]) ? 4'b1101 : 4'b1010;
													assign node17156 = (inp[15]) ? node17164 : node17157;
														assign node17157 = (inp[7]) ? node17161 : node17158;
															assign node17158 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node17161 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node17164 = (inp[7]) ? node17166 : 4'b1010;
															assign node17166 = (inp[2]) ? 4'b1000 : 4'b1001;
										assign node17169 = (inp[2]) ? node17223 : node17170;
											assign node17170 = (inp[5]) ? node17188 : node17171;
												assign node17171 = (inp[13]) ? node17179 : node17172;
													assign node17172 = (inp[15]) ? node17176 : node17173;
														assign node17173 = (inp[7]) ? 4'b1010 : 4'b1000;
														assign node17176 = (inp[7]) ? 4'b1001 : 4'b1011;
													assign node17179 = (inp[15]) ? node17183 : node17180;
														assign node17180 = (inp[7]) ? 4'b1110 : 4'b1100;
														assign node17183 = (inp[1]) ? node17185 : 4'b1111;
															assign node17185 = (inp[7]) ? 4'b1100 : 4'b1110;
												assign node17188 = (inp[13]) ? node17204 : node17189;
													assign node17189 = (inp[1]) ? node17197 : node17190;
														assign node17190 = (inp[15]) ? node17194 : node17191;
															assign node17191 = (inp[7]) ? 4'b1111 : 4'b1100;
															assign node17194 = (inp[7]) ? 4'b1000 : 4'b1110;
														assign node17197 = (inp[10]) ? node17199 : 4'b1111;
															assign node17199 = (inp[7]) ? node17201 : 4'b1100;
																assign node17201 = (inp[15]) ? 4'b1100 : 4'b1111;
													assign node17204 = (inp[1]) ? node17216 : node17205;
														assign node17205 = (inp[10]) ? node17209 : node17206;
															assign node17206 = (inp[7]) ? 4'b1101 : 4'b1001;
															assign node17209 = (inp[15]) ? node17213 : node17210;
																assign node17210 = (inp[7]) ? 4'b1010 : 4'b1001;
																assign node17213 = (inp[7]) ? 4'b1101 : 4'b1010;
														assign node17216 = (inp[15]) ? node17220 : node17217;
															assign node17217 = (inp[7]) ? 4'b1010 : 4'b1001;
															assign node17220 = (inp[7]) ? 4'b1000 : 4'b1010;
											assign node17223 = (inp[15]) ? node17245 : node17224;
												assign node17224 = (inp[7]) ? node17238 : node17225;
													assign node17225 = (inp[1]) ? node17233 : node17226;
														assign node17226 = (inp[5]) ? node17230 : node17227;
															assign node17227 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node17230 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node17233 = (inp[13]) ? 4'b1101 : node17234;
															assign node17234 = (inp[5]) ? 4'b1101 : 4'b1001;
													assign node17238 = (inp[5]) ? node17242 : node17239;
														assign node17239 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node17242 = (inp[13]) ? 4'b1010 : 4'b1110;
												assign node17245 = (inp[7]) ? node17255 : node17246;
													assign node17246 = (inp[13]) ? node17250 : node17247;
														assign node17247 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node17250 = (inp[5]) ? node17252 : 4'b1110;
															assign node17252 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node17255 = (inp[5]) ? node17267 : node17256;
														assign node17256 = (inp[10]) ? node17262 : node17257;
															assign node17257 = (inp[1]) ? node17259 : 4'b1101;
																assign node17259 = (inp[13]) ? 4'b1101 : 4'b1000;
															assign node17262 = (inp[1]) ? 4'b1000 : node17263;
																assign node17263 = (inp[13]) ? 4'b1000 : 4'b1101;
														assign node17267 = (inp[10]) ? node17273 : node17268;
															assign node17268 = (inp[13]) ? node17270 : 4'b1000;
																assign node17270 = (inp[1]) ? 4'b1000 : 4'b1101;
															assign node17273 = (inp[1]) ? 4'b1101 : 4'b1000;
							assign node17276 = (inp[9]) ? node17630 : node17277;
								assign node17277 = (inp[11]) ? node17445 : node17278;
									assign node17278 = (inp[0]) ? node17378 : node17279;
										assign node17279 = (inp[2]) ? node17339 : node17280;
											assign node17280 = (inp[7]) ? node17318 : node17281;
												assign node17281 = (inp[15]) ? node17289 : node17282;
													assign node17282 = (inp[13]) ? node17286 : node17283;
														assign node17283 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node17286 = (inp[5]) ? 4'b1001 : 4'b1100;
													assign node17289 = (inp[10]) ? node17303 : node17290;
														assign node17290 = (inp[13]) ? node17296 : node17291;
															assign node17291 = (inp[1]) ? node17293 : 4'b1110;
																assign node17293 = (inp[5]) ? 4'b1011 : 4'b1110;
															assign node17296 = (inp[5]) ? node17300 : node17297;
																assign node17297 = (inp[1]) ? 4'b1010 : 4'b1111;
																assign node17300 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node17303 = (inp[5]) ? node17311 : node17304;
															assign node17304 = (inp[13]) ? node17308 : node17305;
																assign node17305 = (inp[1]) ? 4'b1110 : 4'b1010;
																assign node17308 = (inp[1]) ? 4'b1010 : 4'b1111;
															assign node17311 = (inp[13]) ? node17315 : node17312;
																assign node17312 = (inp[1]) ? 4'b1011 : 4'b1110;
																assign node17315 = (inp[1]) ? 4'b1110 : 4'b1010;
												assign node17318 = (inp[15]) ? node17326 : node17319;
													assign node17319 = (inp[5]) ? node17323 : node17320;
														assign node17320 = (inp[13]) ? 4'b1110 : 4'b1010;
														assign node17323 = (inp[13]) ? 4'b1010 : 4'b1111;
													assign node17326 = (inp[5]) ? node17334 : node17327;
														assign node17327 = (inp[13]) ? node17331 : node17328;
															assign node17328 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node17331 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node17334 = (inp[13]) ? node17336 : 4'b1100;
															assign node17336 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node17339 = (inp[13]) ? node17361 : node17340;
												assign node17340 = (inp[5]) ? node17350 : node17341;
													assign node17341 = (inp[15]) ? node17345 : node17342;
														assign node17342 = (inp[7]) ? 4'b1011 : 4'b1001;
														assign node17345 = (inp[7]) ? 4'b1000 : node17346;
															assign node17346 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node17350 = (inp[7]) ? node17356 : node17351;
														assign node17351 = (inp[15]) ? node17353 : 4'b1100;
															assign node17353 = (inp[1]) ? 4'b1011 : 4'b1110;
														assign node17356 = (inp[15]) ? node17358 : 4'b1111;
															assign node17358 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node17361 = (inp[5]) ? node17371 : node17362;
													assign node17362 = (inp[7]) ? node17368 : node17363;
														assign node17363 = (inp[15]) ? node17365 : 4'b1101;
															assign node17365 = (inp[1]) ? 4'b1011 : 4'b1110;
														assign node17368 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node17371 = (inp[15]) ? node17375 : node17372;
														assign node17372 = (inp[7]) ? 4'b1011 : 4'b1000;
														assign node17375 = (inp[7]) ? 4'b1001 : 4'b1011;
										assign node17378 = (inp[5]) ? node17412 : node17379;
											assign node17379 = (inp[13]) ? node17395 : node17380;
												assign node17380 = (inp[15]) ? node17384 : node17381;
													assign node17381 = (inp[7]) ? 4'b1010 : 4'b1000;
													assign node17384 = (inp[7]) ? node17390 : node17385;
														assign node17385 = (inp[1]) ? node17387 : 4'b1010;
															assign node17387 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node17390 = (inp[2]) ? node17392 : 4'b1001;
															assign node17392 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node17395 = (inp[1]) ? node17405 : node17396;
													assign node17396 = (inp[15]) ? node17400 : node17397;
														assign node17397 = (inp[7]) ? 4'b1110 : 4'b1100;
														assign node17400 = (inp[7]) ? node17402 : 4'b1111;
															assign node17402 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node17405 = (inp[15]) ? node17409 : node17406;
														assign node17406 = (inp[7]) ? 4'b1110 : 4'b1100;
														assign node17409 = (inp[7]) ? 4'b1100 : 4'b1010;
											assign node17412 = (inp[13]) ? node17434 : node17413;
												assign node17413 = (inp[7]) ? node17425 : node17414;
													assign node17414 = (inp[15]) ? node17418 : node17415;
														assign node17415 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node17418 = (inp[1]) ? node17422 : node17419;
															assign node17419 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node17422 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node17425 = (inp[15]) ? node17429 : node17426;
														assign node17426 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node17429 = (inp[2]) ? 4'b1100 : node17430;
															assign node17430 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node17434 = (inp[7]) ? node17442 : node17435;
													assign node17435 = (inp[15]) ? node17437 : 4'b1001;
														assign node17437 = (inp[1]) ? node17439 : 4'b1010;
															assign node17439 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node17442 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node17445 = (inp[0]) ? node17547 : node17446;
										assign node17446 = (inp[7]) ? node17498 : node17447;
											assign node17447 = (inp[15]) ? node17461 : node17448;
												assign node17448 = (inp[13]) ? node17454 : node17449;
													assign node17449 = (inp[5]) ? 4'b1101 : node17450;
														assign node17450 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node17454 = (inp[5]) ? node17458 : node17455;
														assign node17455 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node17458 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node17461 = (inp[2]) ? node17485 : node17462;
													assign node17462 = (inp[10]) ? node17478 : node17463;
														assign node17463 = (inp[5]) ? node17471 : node17464;
															assign node17464 = (inp[1]) ? node17468 : node17465;
																assign node17465 = (inp[13]) ? 4'b1110 : 4'b1011;
																assign node17468 = (inp[13]) ? 4'b1011 : 4'b1111;
															assign node17471 = (inp[1]) ? node17475 : node17472;
																assign node17472 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node17475 = (inp[13]) ? 4'b1111 : 4'b1010;
														assign node17478 = (inp[5]) ? node17480 : 4'b1011;
															assign node17480 = (inp[13]) ? node17482 : 4'b1111;
																assign node17482 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node17485 = (inp[1]) ? node17493 : node17486;
														assign node17486 = (inp[5]) ? node17490 : node17487;
															assign node17487 = (inp[13]) ? 4'b1111 : 4'b1010;
															assign node17490 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node17493 = (inp[10]) ? 4'b1111 : node17494;
															assign node17494 = (inp[5]) ? 4'b1010 : 4'b1111;
											assign node17498 = (inp[15]) ? node17528 : node17499;
												assign node17499 = (inp[2]) ? node17507 : node17500;
													assign node17500 = (inp[5]) ? node17504 : node17501;
														assign node17501 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node17504 = (inp[13]) ? 4'b1011 : 4'b1110;
													assign node17507 = (inp[1]) ? node17515 : node17508;
														assign node17508 = (inp[5]) ? node17512 : node17509;
															assign node17509 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node17512 = (inp[13]) ? 4'b1010 : 4'b1110;
														assign node17515 = (inp[10]) ? node17521 : node17516;
															assign node17516 = (inp[13]) ? node17518 : 4'b1010;
																assign node17518 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node17521 = (inp[13]) ? node17525 : node17522;
																assign node17522 = (inp[5]) ? 4'b1110 : 4'b1010;
																assign node17525 = (inp[5]) ? 4'b1010 : 4'b1110;
												assign node17528 = (inp[13]) ? node17540 : node17529;
													assign node17529 = (inp[5]) ? node17535 : node17530;
														assign node17530 = (inp[2]) ? 4'b1001 : node17531;
															assign node17531 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node17535 = (inp[1]) ? 4'b1101 : node17536;
															assign node17536 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node17540 = (inp[5]) ? node17542 : 4'b1100;
														assign node17542 = (inp[2]) ? 4'b1000 : node17543;
															assign node17543 = (inp[1]) ? 4'b1001 : 4'b1000;
										assign node17547 = (inp[7]) ? node17595 : node17548;
											assign node17548 = (inp[15]) ? node17558 : node17549;
												assign node17549 = (inp[5]) ? node17553 : node17550;
													assign node17550 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node17553 = (inp[13]) ? 4'b1000 : node17554;
														assign node17554 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node17558 = (inp[2]) ? node17580 : node17559;
													assign node17559 = (inp[1]) ? node17573 : node17560;
														assign node17560 = (inp[10]) ? node17566 : node17561;
															assign node17561 = (inp[13]) ? node17563 : 4'b1110;
																assign node17563 = (inp[5]) ? 4'b1011 : 4'b1110;
															assign node17566 = (inp[13]) ? node17570 : node17567;
																assign node17567 = (inp[5]) ? 4'b1110 : 4'b1011;
																assign node17570 = (inp[5]) ? 4'b1011 : 4'b1110;
														assign node17573 = (inp[5]) ? node17577 : node17574;
															assign node17574 = (inp[13]) ? 4'b1011 : 4'b1110;
															assign node17577 = (inp[13]) ? 4'b1110 : 4'b1011;
													assign node17580 = (inp[13]) ? node17588 : node17581;
														assign node17581 = (inp[5]) ? node17585 : node17582;
															assign node17582 = (inp[1]) ? 4'b1111 : 4'b1011;
															assign node17585 = (inp[10]) ? 4'b1111 : 4'b1010;
														assign node17588 = (inp[1]) ? node17592 : node17589;
															assign node17589 = (inp[5]) ? 4'b1011 : 4'b1110;
															assign node17592 = (inp[5]) ? 4'b1111 : 4'b1011;
											assign node17595 = (inp[15]) ? node17613 : node17596;
												assign node17596 = (inp[1]) ? node17606 : node17597;
													assign node17597 = (inp[5]) ? node17601 : node17598;
														assign node17598 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node17601 = (inp[13]) ? 4'b1011 : node17602;
															assign node17602 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node17606 = (inp[13]) ? node17610 : node17607;
														assign node17607 = (inp[5]) ? 4'b1111 : 4'b1011;
														assign node17610 = (inp[5]) ? 4'b1011 : 4'b1111;
												assign node17613 = (inp[13]) ? node17625 : node17614;
													assign node17614 = (inp[5]) ? node17620 : node17615;
														assign node17615 = (inp[2]) ? node17617 : 4'b1000;
															assign node17617 = (inp[1]) ? 4'b1000 : 4'b1001;
														assign node17620 = (inp[2]) ? 4'b1101 : node17621;
															assign node17621 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node17625 = (inp[5]) ? node17627 : 4'b1101;
														assign node17627 = (inp[2]) ? 4'b1000 : 4'b1001;
								assign node17630 = (inp[11]) ? node17780 : node17631;
									assign node17631 = (inp[2]) ? node17697 : node17632;
										assign node17632 = (inp[5]) ? node17666 : node17633;
											assign node17633 = (inp[13]) ? node17649 : node17634;
												assign node17634 = (inp[15]) ? node17638 : node17635;
													assign node17635 = (inp[7]) ? 4'b1011 : 4'b1001;
													assign node17638 = (inp[7]) ? node17644 : node17639;
														assign node17639 = (inp[1]) ? node17641 : 4'b1011;
															assign node17641 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node17644 = (inp[1]) ? 4'b1000 : node17645;
															assign node17645 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node17649 = (inp[1]) ? node17659 : node17650;
													assign node17650 = (inp[15]) ? node17654 : node17651;
														assign node17651 = (inp[7]) ? 4'b1111 : 4'b1101;
														assign node17654 = (inp[7]) ? node17656 : 4'b1110;
															assign node17656 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node17659 = (inp[7]) ? node17663 : node17660;
														assign node17660 = (inp[15]) ? 4'b1011 : 4'b1101;
														assign node17663 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node17666 = (inp[13]) ? node17684 : node17667;
												assign node17667 = (inp[15]) ? node17675 : node17668;
													assign node17668 = (inp[7]) ? node17672 : node17669;
														assign node17669 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node17672 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node17675 = (inp[7]) ? node17679 : node17676;
														assign node17676 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node17679 = (inp[1]) ? node17681 : 4'b1101;
															assign node17681 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node17684 = (inp[7]) ? node17690 : node17685;
													assign node17685 = (inp[15]) ? node17687 : 4'b1000;
														assign node17687 = (inp[1]) ? 4'b1110 : 4'b1011;
													assign node17690 = (inp[15]) ? node17692 : 4'b1011;
														assign node17692 = (inp[1]) ? 4'b1001 : node17693;
															assign node17693 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node17697 = (inp[7]) ? node17737 : node17698;
											assign node17698 = (inp[15]) ? node17720 : node17699;
												assign node17699 = (inp[0]) ? node17707 : node17700;
													assign node17700 = (inp[5]) ? node17704 : node17701;
														assign node17701 = (inp[13]) ? 4'b1100 : 4'b1000;
														assign node17704 = (inp[13]) ? 4'b1001 : 4'b1101;
													assign node17707 = (inp[1]) ? node17713 : node17708;
														assign node17708 = (inp[13]) ? 4'b1101 : node17709;
															assign node17709 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node17713 = (inp[13]) ? node17717 : node17714;
															assign node17714 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node17717 = (inp[5]) ? 4'b1000 : 4'b1101;
												assign node17720 = (inp[13]) ? node17730 : node17721;
													assign node17721 = (inp[1]) ? node17727 : node17722;
														assign node17722 = (inp[5]) ? 4'b1111 : node17723;
															assign node17723 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node17727 = (inp[5]) ? 4'b1010 : 4'b1111;
													assign node17730 = (inp[5]) ? 4'b1111 : node17731;
														assign node17731 = (inp[1]) ? 4'b1010 : node17732;
															assign node17732 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node17737 = (inp[15]) ? node17761 : node17738;
												assign node17738 = (inp[0]) ? node17754 : node17739;
													assign node17739 = (inp[10]) ? node17747 : node17740;
														assign node17740 = (inp[13]) ? node17744 : node17741;
															assign node17741 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node17744 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node17747 = (inp[13]) ? node17751 : node17748;
															assign node17748 = (inp[5]) ? 4'b1110 : 4'b1010;
															assign node17751 = (inp[5]) ? 4'b1010 : 4'b1110;
													assign node17754 = (inp[13]) ? node17758 : node17755;
														assign node17755 = (inp[5]) ? 4'b1110 : 4'b1011;
														assign node17758 = (inp[5]) ? 4'b1011 : 4'b1111;
												assign node17761 = (inp[13]) ? node17769 : node17762;
													assign node17762 = (inp[5]) ? node17766 : node17763;
														assign node17763 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node17766 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node17769 = (inp[5]) ? node17775 : node17770;
														assign node17770 = (inp[0]) ? node17772 : 4'b1100;
															assign node17772 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node17775 = (inp[1]) ? node17777 : 4'b1000;
															assign node17777 = (inp[0]) ? 4'b1001 : 4'b1000;
									assign node17780 = (inp[5]) ? node17848 : node17781;
										assign node17781 = (inp[13]) ? node17817 : node17782;
											assign node17782 = (inp[15]) ? node17794 : node17783;
												assign node17783 = (inp[7]) ? node17789 : node17784;
													assign node17784 = (inp[0]) ? 4'b1000 : node17785;
														assign node17785 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node17789 = (inp[0]) ? 4'b1010 : node17790;
														assign node17790 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node17794 = (inp[7]) ? node17804 : node17795;
													assign node17795 = (inp[1]) ? node17801 : node17796;
														assign node17796 = (inp[0]) ? 4'b1010 : node17797;
															assign node17797 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node17801 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node17804 = (inp[0]) ? node17812 : node17805;
														assign node17805 = (inp[10]) ? 4'b1000 : node17806;
															assign node17806 = (inp[2]) ? 4'b1000 : node17807;
																assign node17807 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node17812 = (inp[1]) ? 4'b1001 : node17813;
															assign node17813 = (inp[10]) ? 4'b1001 : 4'b1000;
											assign node17817 = (inp[15]) ? node17829 : node17818;
												assign node17818 = (inp[7]) ? node17824 : node17819;
													assign node17819 = (inp[0]) ? 4'b1100 : node17820;
														assign node17820 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node17824 = (inp[2]) ? node17826 : 4'b1110;
														assign node17826 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node17829 = (inp[7]) ? node17841 : node17830;
													assign node17830 = (inp[1]) ? node17836 : node17831;
														assign node17831 = (inp[0]) ? 4'b1111 : node17832;
															assign node17832 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node17836 = (inp[2]) ? node17838 : 4'b1010;
															assign node17838 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node17841 = (inp[1]) ? 4'b1100 : node17842;
														assign node17842 = (inp[2]) ? 4'b1101 : node17843;
															assign node17843 = (inp[0]) ? 4'b1100 : 4'b1101;
										assign node17848 = (inp[13]) ? node17882 : node17849;
											assign node17849 = (inp[7]) ? node17865 : node17850;
												assign node17850 = (inp[15]) ? node17856 : node17851;
													assign node17851 = (inp[2]) ? 4'b1100 : node17852;
														assign node17852 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node17856 = (inp[1]) ? node17862 : node17857;
														assign node17857 = (inp[2]) ? 4'b1110 : node17858;
															assign node17858 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node17862 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node17865 = (inp[15]) ? node17871 : node17866;
													assign node17866 = (inp[0]) ? node17868 : 4'b1111;
														assign node17868 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node17871 = (inp[0]) ? node17877 : node17872;
														assign node17872 = (inp[2]) ? node17874 : 4'b1100;
															assign node17874 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node17877 = (inp[2]) ? 4'b1100 : node17878;
															assign node17878 = (inp[1]) ? 4'b1101 : 4'b1100;
											assign node17882 = (inp[1]) ? node17924 : node17883;
												assign node17883 = (inp[10]) ? node17905 : node17884;
													assign node17884 = (inp[2]) ? node17892 : node17885;
														assign node17885 = (inp[7]) ? node17889 : node17886;
															assign node17886 = (inp[15]) ? 4'b1010 : 4'b1001;
															assign node17889 = (inp[15]) ? 4'b1001 : 4'b1010;
														assign node17892 = (inp[15]) ? node17900 : node17893;
															assign node17893 = (inp[7]) ? node17897 : node17894;
																assign node17894 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node17897 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node17900 = (inp[7]) ? 4'b1001 : node17901;
																assign node17901 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node17905 = (inp[7]) ? node17913 : node17906;
														assign node17906 = (inp[15]) ? 4'b1011 : node17907;
															assign node17907 = (inp[0]) ? 4'b1001 : node17908;
																assign node17908 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node17913 = (inp[15]) ? node17919 : node17914;
															assign node17914 = (inp[0]) ? 4'b1010 : node17915;
																assign node17915 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node17919 = (inp[2]) ? 4'b1001 : node17920;
																assign node17920 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node17924 = (inp[7]) ? node17934 : node17925;
													assign node17925 = (inp[15]) ? node17929 : node17926;
														assign node17926 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node17929 = (inp[0]) ? node17931 : 4'b1110;
															assign node17931 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node17934 = (inp[15]) ? node17940 : node17935;
														assign node17935 = (inp[0]) ? 4'b1010 : node17936;
															assign node17936 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node17940 = (inp[2]) ? node17942 : 4'b1000;
															assign node17942 = (inp[10]) ? 4'b1001 : 4'b1000;
						assign node17945 = (inp[7]) ? node18923 : node17946;
							assign node17946 = (inp[15]) ? node18492 : node17947;
								assign node17947 = (inp[1]) ? node18273 : node17948;
									assign node17948 = (inp[10]) ? node18120 : node17949;
										assign node17949 = (inp[13]) ? node18037 : node17950;
											assign node17950 = (inp[0]) ? node17990 : node17951;
												assign node17951 = (inp[2]) ? node17967 : node17952;
													assign node17952 = (inp[4]) ? node17960 : node17953;
														assign node17953 = (inp[11]) ? node17957 : node17954;
															assign node17954 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node17957 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node17960 = (inp[5]) ? node17964 : node17961;
															assign node17961 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node17964 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node17967 = (inp[9]) ? node17975 : node17968;
														assign node17968 = (inp[11]) ? node17972 : node17969;
															assign node17969 = (inp[4]) ? 4'b1101 : 4'b1000;
															assign node17972 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node17975 = (inp[11]) ? node17983 : node17976;
															assign node17976 = (inp[4]) ? node17980 : node17977;
																assign node17977 = (inp[5]) ? 4'b1101 : 4'b1001;
																assign node17980 = (inp[5]) ? 4'b1001 : 4'b1100;
															assign node17983 = (inp[5]) ? node17987 : node17984;
																assign node17984 = (inp[4]) ? 4'b1101 : 4'b1000;
																assign node17987 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node17990 = (inp[2]) ? node18018 : node17991;
													assign node17991 = (inp[4]) ? node18007 : node17992;
														assign node17992 = (inp[5]) ? node18000 : node17993;
															assign node17993 = (inp[11]) ? node17997 : node17994;
																assign node17994 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node17997 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node18000 = (inp[11]) ? node18004 : node18001;
																assign node18001 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node18004 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node18007 = (inp[5]) ? node18013 : node18008;
															assign node18008 = (inp[11]) ? 4'b1100 : node18009;
																assign node18009 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node18013 = (inp[9]) ? 4'b1000 : node18014;
																assign node18014 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node18018 = (inp[4]) ? node18028 : node18019;
														assign node18019 = (inp[5]) ? 4'b1100 : node18020;
															assign node18020 = (inp[9]) ? node18024 : node18021;
																assign node18021 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node18024 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node18028 = (inp[5]) ? node18030 : 4'b1101;
															assign node18030 = (inp[9]) ? node18034 : node18031;
																assign node18031 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node18034 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node18037 = (inp[11]) ? node18083 : node18038;
												assign node18038 = (inp[2]) ? node18060 : node18039;
													assign node18039 = (inp[4]) ? node18051 : node18040;
														assign node18040 = (inp[5]) ? node18044 : node18041;
															assign node18041 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node18044 = (inp[0]) ? node18048 : node18045;
																assign node18045 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node18048 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node18051 = (inp[5]) ? node18057 : node18052;
															assign node18052 = (inp[9]) ? 4'b1000 : node18053;
																assign node18053 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node18057 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node18060 = (inp[0]) ? node18068 : node18061;
														assign node18061 = (inp[4]) ? node18063 : 4'b1000;
															assign node18063 = (inp[5]) ? 4'b1101 : node18064;
																assign node18064 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node18068 = (inp[9]) ? node18076 : node18069;
															assign node18069 = (inp[5]) ? node18073 : node18070;
																assign node18070 = (inp[4]) ? 4'b1000 : 4'b1101;
																assign node18073 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node18076 = (inp[4]) ? node18080 : node18077;
																assign node18077 = (inp[5]) ? 4'b1000 : 4'b1100;
																assign node18080 = (inp[5]) ? 4'b1100 : 4'b1001;
												assign node18083 = (inp[0]) ? node18101 : node18084;
													assign node18084 = (inp[9]) ? node18094 : node18085;
														assign node18085 = (inp[5]) ? node18089 : node18086;
															assign node18086 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node18089 = (inp[4]) ? node18091 : 4'b1000;
																assign node18091 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node18094 = (inp[5]) ? node18098 : node18095;
															assign node18095 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node18098 = (inp[4]) ? 4'b1101 : 4'b1000;
													assign node18101 = (inp[9]) ? node18113 : node18102;
														assign node18102 = (inp[2]) ? node18108 : node18103;
															assign node18103 = (inp[4]) ? node18105 : 4'b1000;
																assign node18105 = (inp[5]) ? 4'b1100 : 4'b1000;
															assign node18108 = (inp[4]) ? 4'b1100 : node18109;
																assign node18109 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node18113 = (inp[2]) ? node18115 : 4'b1101;
															assign node18115 = (inp[4]) ? 4'b1000 : node18116;
																assign node18116 = (inp[5]) ? 4'b1001 : 4'b1101;
										assign node18120 = (inp[9]) ? node18194 : node18121;
											assign node18121 = (inp[11]) ? node18165 : node18122;
												assign node18122 = (inp[5]) ? node18142 : node18123;
													assign node18123 = (inp[2]) ? node18131 : node18124;
														assign node18124 = (inp[13]) ? node18128 : node18125;
															assign node18125 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node18128 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node18131 = (inp[4]) ? node18137 : node18132;
															assign node18132 = (inp[13]) ? 4'b1101 : node18133;
																assign node18133 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node18137 = (inp[13]) ? 4'b1000 : node18138;
																assign node18138 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node18142 = (inp[0]) ? node18158 : node18143;
														assign node18143 = (inp[2]) ? node18151 : node18144;
															assign node18144 = (inp[4]) ? node18148 : node18145;
																assign node18145 = (inp[13]) ? 4'b1000 : 4'b1100;
																assign node18148 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node18151 = (inp[13]) ? node18155 : node18152;
																assign node18152 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node18155 = (inp[4]) ? 4'b1100 : 4'b1001;
														assign node18158 = (inp[4]) ? node18162 : node18159;
															assign node18159 = (inp[13]) ? 4'b1001 : 4'b1100;
															assign node18162 = (inp[13]) ? 4'b1101 : 4'b1001;
												assign node18165 = (inp[5]) ? node18183 : node18166;
													assign node18166 = (inp[13]) ? node18174 : node18167;
														assign node18167 = (inp[4]) ? node18169 : 4'b1001;
															assign node18169 = (inp[2]) ? node18171 : 4'b1101;
																assign node18171 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node18174 = (inp[4]) ? node18178 : node18175;
															assign node18175 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node18178 = (inp[0]) ? node18180 : 4'b1001;
																assign node18180 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node18183 = (inp[4]) ? node18189 : node18184;
														assign node18184 = (inp[13]) ? node18186 : 4'b1101;
															assign node18186 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node18189 = (inp[13]) ? node18191 : 4'b1000;
															assign node18191 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node18194 = (inp[0]) ? node18228 : node18195;
												assign node18195 = (inp[11]) ? node18215 : node18196;
													assign node18196 = (inp[5]) ? node18204 : node18197;
														assign node18197 = (inp[4]) ? node18201 : node18198;
															assign node18198 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node18201 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node18204 = (inp[13]) ? node18208 : node18205;
															assign node18205 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node18208 = (inp[4]) ? node18212 : node18209;
																assign node18209 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node18212 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node18215 = (inp[2]) ? node18221 : node18216;
														assign node18216 = (inp[5]) ? 4'b1101 : node18217;
															assign node18217 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node18221 = (inp[4]) ? node18223 : 4'b1000;
															assign node18223 = (inp[5]) ? 4'b1000 : node18224;
																assign node18224 = (inp[13]) ? 4'b1000 : 4'b1101;
												assign node18228 = (inp[11]) ? node18254 : node18229;
													assign node18229 = (inp[5]) ? node18241 : node18230;
														assign node18230 = (inp[2]) ? node18236 : node18231;
															assign node18231 = (inp[4]) ? 4'b1000 : node18232;
																assign node18232 = (inp[13]) ? 4'b1101 : 4'b1001;
															assign node18236 = (inp[4]) ? node18238 : 4'b1000;
																assign node18238 = (inp[13]) ? 4'b1001 : 4'b1101;
														assign node18241 = (inp[2]) ? node18247 : node18242;
															assign node18242 = (inp[4]) ? 4'b1000 : node18243;
																assign node18243 = (inp[13]) ? 4'b1000 : 4'b1101;
															assign node18247 = (inp[4]) ? node18251 : node18248;
																assign node18248 = (inp[13]) ? 4'b1000 : 4'b1100;
																assign node18251 = (inp[13]) ? 4'b1100 : 4'b1000;
													assign node18254 = (inp[5]) ? node18266 : node18255;
														assign node18255 = (inp[2]) ? node18259 : node18256;
															assign node18256 = (inp[13]) ? 4'b1100 : 4'b1000;
															assign node18259 = (inp[4]) ? node18263 : node18260;
																assign node18260 = (inp[13]) ? 4'b1101 : 4'b1001;
																assign node18263 = (inp[13]) ? 4'b1000 : 4'b1100;
														assign node18266 = (inp[13]) ? node18270 : node18267;
															assign node18267 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node18270 = (inp[4]) ? 4'b1101 : 4'b1001;
									assign node18273 = (inp[13]) ? node18401 : node18274;
										assign node18274 = (inp[2]) ? node18328 : node18275;
											assign node18275 = (inp[5]) ? node18297 : node18276;
												assign node18276 = (inp[4]) ? node18284 : node18277;
													assign node18277 = (inp[9]) ? node18281 : node18278;
														assign node18278 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node18281 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node18284 = (inp[0]) ? node18290 : node18285;
														assign node18285 = (inp[11]) ? 4'b1001 : node18286;
															assign node18286 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node18290 = (inp[11]) ? node18294 : node18291;
															assign node18291 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node18294 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node18297 = (inp[4]) ? node18321 : node18298;
													assign node18298 = (inp[10]) ? node18312 : node18299;
														assign node18299 = (inp[0]) ? node18307 : node18300;
															assign node18300 = (inp[11]) ? node18304 : node18301;
																assign node18301 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node18304 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node18307 = (inp[11]) ? node18309 : 4'b1000;
																assign node18309 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node18312 = (inp[11]) ? node18314 : 4'b1001;
															assign node18314 = (inp[9]) ? node18318 : node18315;
																assign node18315 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node18318 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node18321 = (inp[11]) ? node18325 : node18322;
														assign node18322 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node18325 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node18328 = (inp[11]) ? node18358 : node18329;
												assign node18329 = (inp[4]) ? node18341 : node18330;
													assign node18330 = (inp[5]) ? node18338 : node18331;
														assign node18331 = (inp[0]) ? node18335 : node18332;
															assign node18332 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node18335 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node18338 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node18341 = (inp[5]) ? node18345 : node18342;
														assign node18342 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node18345 = (inp[10]) ? node18353 : node18346;
															assign node18346 = (inp[9]) ? node18350 : node18347;
																assign node18347 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node18350 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node18353 = (inp[0]) ? node18355 : 4'b1101;
																assign node18355 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node18358 = (inp[10]) ? node18378 : node18359;
													assign node18359 = (inp[9]) ? node18367 : node18360;
														assign node18360 = (inp[4]) ? node18364 : node18361;
															assign node18361 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node18364 = (inp[5]) ? 4'b1101 : 4'b1000;
														assign node18367 = (inp[5]) ? node18373 : node18368;
															assign node18368 = (inp[4]) ? 4'b1001 : node18369;
																assign node18369 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node18373 = (inp[4]) ? node18375 : 4'b1000;
																assign node18375 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node18378 = (inp[0]) ? node18392 : node18379;
														assign node18379 = (inp[9]) ? node18385 : node18380;
															assign node18380 = (inp[5]) ? 4'b1100 : node18381;
																assign node18381 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node18385 = (inp[4]) ? node18389 : node18386;
																assign node18386 = (inp[5]) ? 4'b1000 : 4'b1101;
																assign node18389 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node18392 = (inp[9]) ? 4'b1100 : node18393;
															assign node18393 = (inp[5]) ? node18397 : node18394;
																assign node18394 = (inp[4]) ? 4'b1000 : 4'b1101;
																assign node18397 = (inp[4]) ? 4'b1101 : 4'b1001;
										assign node18401 = (inp[9]) ? node18445 : node18402;
											assign node18402 = (inp[11]) ? node18422 : node18403;
												assign node18403 = (inp[0]) ? node18415 : node18404;
													assign node18404 = (inp[5]) ? node18410 : node18405;
														assign node18405 = (inp[4]) ? 4'b1101 : node18406;
															assign node18406 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node18410 = (inp[4]) ? 4'b1000 : node18411;
															assign node18411 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node18415 = (inp[4]) ? node18419 : node18416;
														assign node18416 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node18419 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node18422 = (inp[0]) ? node18434 : node18423;
													assign node18423 = (inp[5]) ? node18429 : node18424;
														assign node18424 = (inp[4]) ? 4'b1100 : node18425;
															assign node18425 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node18429 = (inp[4]) ? 4'b1001 : node18430;
															assign node18430 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node18434 = (inp[4]) ? node18438 : node18435;
														assign node18435 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node18438 = (inp[5]) ? node18442 : node18439;
															assign node18439 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node18442 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node18445 = (inp[11]) ? node18469 : node18446;
												assign node18446 = (inp[4]) ? node18458 : node18447;
													assign node18447 = (inp[5]) ? node18453 : node18448;
														assign node18448 = (inp[0]) ? 4'b1001 : node18449;
															assign node18449 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node18453 = (inp[0]) ? 4'b1101 : node18454;
															assign node18454 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node18458 = (inp[5]) ? node18464 : node18459;
														assign node18459 = (inp[2]) ? 4'b1100 : node18460;
															assign node18460 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node18464 = (inp[2]) ? 4'b1001 : node18465;
															assign node18465 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node18469 = (inp[0]) ? node18481 : node18470;
													assign node18470 = (inp[5]) ? node18476 : node18471;
														assign node18471 = (inp[4]) ? 4'b1101 : node18472;
															assign node18472 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node18476 = (inp[4]) ? 4'b1000 : node18477;
															assign node18477 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node18481 = (inp[4]) ? node18485 : node18482;
														assign node18482 = (inp[5]) ? 4'b1100 : 4'b1000;
														assign node18485 = (inp[5]) ? node18489 : node18486;
															assign node18486 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node18489 = (inp[2]) ? 4'b1000 : 4'b1001;
								assign node18492 = (inp[5]) ? node18698 : node18493;
									assign node18493 = (inp[13]) ? node18589 : node18494;
										assign node18494 = (inp[1]) ? node18542 : node18495;
											assign node18495 = (inp[9]) ? node18517 : node18496;
												assign node18496 = (inp[11]) ? node18508 : node18497;
													assign node18497 = (inp[0]) ? node18499 : 4'b1010;
														assign node18499 = (inp[10]) ? node18505 : node18500;
															assign node18500 = (inp[2]) ? node18502 : 4'b1010;
																assign node18502 = (inp[4]) ? 4'b1010 : 4'b1011;
															assign node18505 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node18508 = (inp[0]) ? node18510 : 4'b1011;
														assign node18510 = (inp[10]) ? 4'b1010 : node18511;
															assign node18511 = (inp[2]) ? node18513 : 4'b1010;
																assign node18513 = (inp[4]) ? 4'b1011 : 4'b1010;
												assign node18517 = (inp[11]) ? node18533 : node18518;
													assign node18518 = (inp[0]) ? node18520 : 4'b1011;
														assign node18520 = (inp[10]) ? node18528 : node18521;
															assign node18521 = (inp[2]) ? node18525 : node18522;
																assign node18522 = (inp[4]) ? 4'b1010 : 4'b1011;
																assign node18525 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node18528 = (inp[2]) ? node18530 : 4'b1011;
																assign node18530 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node18533 = (inp[0]) ? node18535 : 4'b1010;
														assign node18535 = (inp[2]) ? node18539 : node18536;
															assign node18536 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node18539 = (inp[4]) ? 4'b1010 : 4'b1011;
											assign node18542 = (inp[4]) ? node18566 : node18543;
												assign node18543 = (inp[11]) ? node18555 : node18544;
													assign node18544 = (inp[9]) ? node18550 : node18545;
														assign node18545 = (inp[0]) ? 4'b1110 : node18546;
															assign node18546 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node18550 = (inp[2]) ? 4'b1111 : node18551;
															assign node18551 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node18555 = (inp[9]) ? node18561 : node18556;
														assign node18556 = (inp[2]) ? 4'b1111 : node18557;
															assign node18557 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node18561 = (inp[2]) ? 4'b1110 : node18562;
															assign node18562 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node18566 = (inp[11]) ? node18578 : node18567;
													assign node18567 = (inp[9]) ? node18573 : node18568;
														assign node18568 = (inp[2]) ? node18570 : 4'b1010;
															assign node18570 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node18573 = (inp[0]) ? 4'b1011 : node18574;
															assign node18574 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node18578 = (inp[9]) ? node18584 : node18579;
														assign node18579 = (inp[2]) ? node18581 : 4'b1011;
															assign node18581 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node18584 = (inp[2]) ? node18586 : 4'b1010;
															assign node18586 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node18589 = (inp[1]) ? node18651 : node18590;
											assign node18590 = (inp[10]) ? node18622 : node18591;
												assign node18591 = (inp[0]) ? node18599 : node18592;
													assign node18592 = (inp[9]) ? node18596 : node18593;
														assign node18593 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node18596 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node18599 = (inp[2]) ? node18607 : node18600;
														assign node18600 = (inp[11]) ? node18602 : 4'b1111;
															assign node18602 = (inp[4]) ? 4'b1111 : node18603;
																assign node18603 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node18607 = (inp[4]) ? node18615 : node18608;
															assign node18608 = (inp[11]) ? node18612 : node18609;
																assign node18609 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node18612 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node18615 = (inp[11]) ? node18619 : node18616;
																assign node18616 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node18619 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node18622 = (inp[9]) ? node18640 : node18623;
													assign node18623 = (inp[11]) ? node18633 : node18624;
														assign node18624 = (inp[0]) ? node18626 : 4'b1111;
															assign node18626 = (inp[2]) ? node18630 : node18627;
																assign node18627 = (inp[4]) ? 4'b1110 : 4'b1111;
																assign node18630 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node18633 = (inp[4]) ? 4'b1110 : node18634;
															assign node18634 = (inp[0]) ? node18636 : 4'b1110;
																assign node18636 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node18640 = (inp[11]) ? node18646 : node18641;
														assign node18641 = (inp[0]) ? node18643 : 4'b1110;
															assign node18643 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node18646 = (inp[0]) ? node18648 : 4'b1111;
															assign node18648 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node18651 = (inp[4]) ? node18677 : node18652;
												assign node18652 = (inp[0]) ? node18660 : node18653;
													assign node18653 = (inp[9]) ? node18657 : node18654;
														assign node18654 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node18657 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node18660 = (inp[11]) ? node18672 : node18661;
														assign node18661 = (inp[10]) ? node18667 : node18662;
															assign node18662 = (inp[2]) ? 4'b1010 : node18663;
																assign node18663 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node18667 = (inp[2]) ? node18669 : 4'b1011;
																assign node18669 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node18672 = (inp[2]) ? node18674 : 4'b1011;
															assign node18674 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node18677 = (inp[2]) ? node18685 : node18678;
													assign node18678 = (inp[9]) ? node18682 : node18679;
														assign node18679 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node18682 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node18685 = (inp[11]) ? 4'b1111 : node18686;
														assign node18686 = (inp[10]) ? node18692 : node18687;
															assign node18687 = (inp[9]) ? 4'b1111 : node18688;
																assign node18688 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node18692 = (inp[0]) ? node18694 : 4'b1110;
																assign node18694 = (inp[9]) ? 4'b1110 : 4'b1111;
									assign node18698 = (inp[13]) ? node18798 : node18699;
										assign node18699 = (inp[4]) ? node18743 : node18700;
											assign node18700 = (inp[1]) ? node18724 : node18701;
												assign node18701 = (inp[9]) ? node18713 : node18702;
													assign node18702 = (inp[11]) ? node18708 : node18703;
														assign node18703 = (inp[0]) ? node18705 : 4'b1110;
															assign node18705 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node18708 = (inp[2]) ? node18710 : 4'b1111;
															assign node18710 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node18713 = (inp[11]) ? node18719 : node18714;
														assign node18714 = (inp[2]) ? node18716 : 4'b1111;
															assign node18716 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node18719 = (inp[2]) ? node18721 : 4'b1110;
															assign node18721 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node18724 = (inp[9]) ? node18736 : node18725;
													assign node18725 = (inp[11]) ? node18731 : node18726;
														assign node18726 = (inp[0]) ? node18728 : 4'b1010;
															assign node18728 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node18731 = (inp[2]) ? node18733 : 4'b1011;
															assign node18733 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node18736 = (inp[11]) ? 4'b1010 : node18737;
														assign node18737 = (inp[0]) ? node18739 : 4'b1011;
															assign node18739 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node18743 = (inp[11]) ? node18767 : node18744;
												assign node18744 = (inp[0]) ? node18756 : node18745;
													assign node18745 = (inp[9]) ? node18751 : node18746;
														assign node18746 = (inp[2]) ? 4'b1110 : node18747;
															assign node18747 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node18751 = (inp[1]) ? 4'b1111 : node18752;
															assign node18752 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node18756 = (inp[9]) ? node18762 : node18757;
														assign node18757 = (inp[1]) ? node18759 : 4'b1111;
															assign node18759 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node18762 = (inp[2]) ? node18764 : 4'b1110;
															assign node18764 = (inp[1]) ? 4'b1111 : 4'b1110;
												assign node18767 = (inp[10]) ? node18779 : node18768;
													assign node18768 = (inp[9]) ? node18772 : node18769;
														assign node18769 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node18772 = (inp[2]) ? node18774 : 4'b1111;
															assign node18774 = (inp[0]) ? node18776 : 4'b1110;
																assign node18776 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node18779 = (inp[9]) ? node18791 : node18780;
														assign node18780 = (inp[2]) ? node18786 : node18781;
															assign node18781 = (inp[0]) ? 4'b1110 : node18782;
																assign node18782 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node18786 = (inp[1]) ? 4'b1111 : node18787;
																assign node18787 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node18791 = (inp[0]) ? 4'b1111 : node18792;
															assign node18792 = (inp[1]) ? 4'b1110 : node18793;
																assign node18793 = (inp[2]) ? 4'b1110 : 4'b1111;
										assign node18798 = (inp[4]) ? node18864 : node18799;
											assign node18799 = (inp[1]) ? node18835 : node18800;
												assign node18800 = (inp[2]) ? node18822 : node18801;
													assign node18801 = (inp[10]) ? node18809 : node18802;
														assign node18802 = (inp[0]) ? node18804 : 4'b1011;
															assign node18804 = (inp[11]) ? 4'b1010 : node18805;
																assign node18805 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node18809 = (inp[9]) ? node18815 : node18810;
															assign node18810 = (inp[0]) ? node18812 : 4'b1010;
																assign node18812 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node18815 = (inp[11]) ? node18819 : node18816;
																assign node18816 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node18819 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node18822 = (inp[0]) ? node18828 : node18823;
														assign node18823 = (inp[9]) ? node18825 : 4'b1011;
															assign node18825 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node18828 = (inp[10]) ? 4'b1011 : node18829;
															assign node18829 = (inp[9]) ? 4'b1011 : node18830;
																assign node18830 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node18835 = (inp[0]) ? node18841 : node18836;
													assign node18836 = (inp[9]) ? 4'b1111 : node18837;
														assign node18837 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node18841 = (inp[9]) ? node18849 : node18842;
														assign node18842 = (inp[11]) ? node18846 : node18843;
															assign node18843 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node18846 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node18849 = (inp[10]) ? node18857 : node18850;
															assign node18850 = (inp[11]) ? node18854 : node18851;
																assign node18851 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node18854 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node18857 = (inp[11]) ? node18861 : node18858;
																assign node18858 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node18861 = (inp[2]) ? 4'b1110 : 4'b1111;
											assign node18864 = (inp[2]) ? node18902 : node18865;
												assign node18865 = (inp[10]) ? node18887 : node18866;
													assign node18866 = (inp[0]) ? node18874 : node18867;
														assign node18867 = (inp[9]) ? node18871 : node18868;
															assign node18868 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node18871 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node18874 = (inp[1]) ? node18882 : node18875;
															assign node18875 = (inp[9]) ? node18879 : node18876;
																assign node18876 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node18879 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node18882 = (inp[11]) ? 4'b1011 : node18883;
																assign node18883 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node18887 = (inp[1]) ? node18895 : node18888;
														assign node18888 = (inp[0]) ? node18890 : 4'b1011;
															assign node18890 = (inp[11]) ? 4'b1011 : node18891;
																assign node18891 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node18895 = (inp[9]) ? node18899 : node18896;
															assign node18896 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node18899 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node18902 = (inp[9]) ? node18912 : node18903;
													assign node18903 = (inp[11]) ? node18909 : node18904;
														assign node18904 = (inp[0]) ? 4'b1010 : node18905;
															assign node18905 = (inp[1]) ? 4'b1011 : 4'b1010;
														assign node18909 = (inp[1]) ? 4'b1010 : 4'b1011;
													assign node18912 = (inp[11]) ? node18918 : node18913;
														assign node18913 = (inp[0]) ? 4'b1011 : node18914;
															assign node18914 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node18918 = (inp[1]) ? node18920 : 4'b1010;
															assign node18920 = (inp[0]) ? 4'b1010 : 4'b1011;
							assign node18923 = (inp[15]) ? node19433 : node18924;
								assign node18924 = (inp[4]) ? node19218 : node18925;
									assign node18925 = (inp[2]) ? node19071 : node18926;
										assign node18926 = (inp[11]) ? node19002 : node18927;
											assign node18927 = (inp[0]) ? node18949 : node18928;
												assign node18928 = (inp[5]) ? node18942 : node18929;
													assign node18929 = (inp[9]) ? node18937 : node18930;
														assign node18930 = (inp[1]) ? node18934 : node18931;
															assign node18931 = (inp[13]) ? 4'b1110 : 4'b1010;
															assign node18934 = (inp[13]) ? 4'b1010 : 4'b1111;
														assign node18937 = (inp[1]) ? 4'b1110 : node18938;
															assign node18938 = (inp[13]) ? 4'b1111 : 4'b1011;
													assign node18942 = (inp[9]) ? node18944 : 4'b1111;
														assign node18944 = (inp[1]) ? node18946 : 4'b1011;
															assign node18946 = (inp[13]) ? 4'b1110 : 4'b1010;
												assign node18949 = (inp[10]) ? node18975 : node18950;
													assign node18950 = (inp[1]) ? node18964 : node18951;
														assign node18951 = (inp[13]) ? node18959 : node18952;
															assign node18952 = (inp[5]) ? node18956 : node18953;
																assign node18953 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node18956 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node18959 = (inp[5]) ? node18961 : 4'b1111;
																assign node18961 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node18964 = (inp[13]) ? node18970 : node18965;
															assign node18965 = (inp[5]) ? node18967 : 4'b1111;
																assign node18967 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node18970 = (inp[5]) ? 4'b1111 : node18971;
																assign node18971 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node18975 = (inp[5]) ? node18987 : node18976;
														assign node18976 = (inp[9]) ? node18982 : node18977;
															assign node18977 = (inp[1]) ? 4'b1110 : node18978;
																assign node18978 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node18982 = (inp[1]) ? node18984 : 4'b1110;
																assign node18984 = (inp[13]) ? 4'b1011 : 4'b1111;
														assign node18987 = (inp[9]) ? node18995 : node18988;
															assign node18988 = (inp[1]) ? node18992 : node18989;
																assign node18989 = (inp[13]) ? 4'b1010 : 4'b1110;
																assign node18992 = (inp[13]) ? 4'b1111 : 4'b1011;
															assign node18995 = (inp[1]) ? node18999 : node18996;
																assign node18996 = (inp[13]) ? 4'b1011 : 4'b1111;
																assign node18999 = (inp[13]) ? 4'b1110 : 4'b1010;
											assign node19002 = (inp[0]) ? node19024 : node19003;
												assign node19003 = (inp[9]) ? node19015 : node19004;
													assign node19004 = (inp[1]) ? node19010 : node19005;
														assign node19005 = (inp[5]) ? 4'b1011 : node19006;
															assign node19006 = (inp[13]) ? 4'b1111 : 4'b1011;
														assign node19010 = (inp[13]) ? node19012 : 4'b1110;
															assign node19012 = (inp[5]) ? 4'b1110 : 4'b1011;
													assign node19015 = (inp[5]) ? node19017 : 4'b1010;
														assign node19017 = (inp[13]) ? node19021 : node19018;
															assign node19018 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node19021 = (inp[1]) ? 4'b1111 : 4'b1010;
												assign node19024 = (inp[10]) ? node19046 : node19025;
													assign node19025 = (inp[13]) ? node19039 : node19026;
														assign node19026 = (inp[1]) ? node19032 : node19027;
															assign node19027 = (inp[5]) ? node19029 : 4'b1011;
																assign node19029 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node19032 = (inp[5]) ? node19036 : node19033;
																assign node19033 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node19036 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node19039 = (inp[9]) ? 4'b1111 : node19040;
															assign node19040 = (inp[1]) ? 4'b1011 : node19041;
																assign node19041 = (inp[5]) ? 4'b1011 : 4'b1110;
													assign node19046 = (inp[13]) ? node19056 : node19047;
														assign node19047 = (inp[9]) ? 4'b1011 : node19048;
															assign node19048 = (inp[5]) ? node19052 : node19049;
																assign node19049 = (inp[1]) ? 4'b1111 : 4'b1010;
																assign node19052 = (inp[1]) ? 4'b1010 : 4'b1111;
														assign node19056 = (inp[1]) ? node19064 : node19057;
															assign node19057 = (inp[5]) ? node19061 : node19058;
																assign node19058 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node19061 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node19064 = (inp[5]) ? node19068 : node19065;
																assign node19065 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node19068 = (inp[9]) ? 4'b1111 : 4'b1110;
										assign node19071 = (inp[13]) ? node19137 : node19072;
											assign node19072 = (inp[0]) ? node19106 : node19073;
												assign node19073 = (inp[10]) ? node19089 : node19074;
													assign node19074 = (inp[5]) ? node19082 : node19075;
														assign node19075 = (inp[9]) ? node19079 : node19076;
															assign node19076 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node19079 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node19082 = (inp[1]) ? 4'b1011 : node19083;
															assign node19083 = (inp[9]) ? node19085 : 4'b1111;
																assign node19085 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node19089 = (inp[5]) ? node19103 : node19090;
														assign node19090 = (inp[1]) ? node19096 : node19091;
															assign node19091 = (inp[9]) ? 4'b1010 : node19092;
																assign node19092 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node19096 = (inp[9]) ? node19100 : node19097;
																assign node19097 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node19100 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node19103 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node19106 = (inp[9]) ? node19122 : node19107;
													assign node19107 = (inp[11]) ? node19115 : node19108;
														assign node19108 = (inp[5]) ? node19112 : node19109;
															assign node19109 = (inp[1]) ? 4'b1110 : 4'b1011;
															assign node19112 = (inp[1]) ? 4'b1010 : 4'b1110;
														assign node19115 = (inp[5]) ? node19119 : node19116;
															assign node19116 = (inp[1]) ? 4'b1111 : 4'b1010;
															assign node19119 = (inp[1]) ? 4'b1011 : 4'b1111;
													assign node19122 = (inp[11]) ? node19130 : node19123;
														assign node19123 = (inp[1]) ? node19127 : node19124;
															assign node19124 = (inp[5]) ? 4'b1111 : 4'b1010;
															assign node19127 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node19130 = (inp[1]) ? node19134 : node19131;
															assign node19131 = (inp[5]) ? 4'b1110 : 4'b1011;
															assign node19134 = (inp[5]) ? 4'b1010 : 4'b1110;
											assign node19137 = (inp[1]) ? node19183 : node19138;
												assign node19138 = (inp[5]) ? node19160 : node19139;
													assign node19139 = (inp[10]) ? node19147 : node19140;
														assign node19140 = (inp[9]) ? node19144 : node19141;
															assign node19141 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node19144 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node19147 = (inp[0]) ? node19153 : node19148;
															assign node19148 = (inp[9]) ? 4'b1110 : node19149;
																assign node19149 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node19153 = (inp[11]) ? node19157 : node19154;
																assign node19154 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node19157 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node19160 = (inp[10]) ? node19170 : node19161;
														assign node19161 = (inp[0]) ? 4'b1010 : node19162;
															assign node19162 = (inp[9]) ? node19166 : node19163;
																assign node19163 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node19166 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node19170 = (inp[11]) ? node19178 : node19171;
															assign node19171 = (inp[9]) ? node19175 : node19172;
																assign node19172 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node19175 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node19178 = (inp[9]) ? 4'b1011 : node19179;
																assign node19179 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node19183 = (inp[5]) ? node19197 : node19184;
													assign node19184 = (inp[11]) ? node19190 : node19185;
														assign node19185 = (inp[0]) ? 4'b1011 : node19186;
															assign node19186 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node19190 = (inp[9]) ? node19194 : node19191;
															assign node19191 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node19194 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node19197 = (inp[10]) ? node19209 : node19198;
														assign node19198 = (inp[9]) ? node19204 : node19199;
															assign node19199 = (inp[0]) ? 4'b1111 : node19200;
																assign node19200 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node19204 = (inp[11]) ? node19206 : 4'b1110;
																assign node19206 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node19209 = (inp[9]) ? 4'b1111 : node19210;
															assign node19210 = (inp[11]) ? node19214 : node19211;
																assign node19211 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node19214 = (inp[0]) ? 4'b1111 : 4'b1110;
									assign node19218 = (inp[13]) ? node19320 : node19219;
										assign node19219 = (inp[0]) ? node19267 : node19220;
											assign node19220 = (inp[1]) ? node19242 : node19221;
												assign node19221 = (inp[5]) ? node19229 : node19222;
													assign node19222 = (inp[11]) ? node19226 : node19223;
														assign node19223 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node19226 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node19229 = (inp[10]) ? node19237 : node19230;
														assign node19230 = (inp[11]) ? node19234 : node19231;
															assign node19231 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node19234 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node19237 = (inp[11]) ? 4'b1010 : node19238;
															assign node19238 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node19242 = (inp[5]) ? node19260 : node19243;
													assign node19243 = (inp[10]) ? node19251 : node19244;
														assign node19244 = (inp[9]) ? 4'b1010 : node19245;
															assign node19245 = (inp[2]) ? 4'b1011 : node19246;
																assign node19246 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node19251 = (inp[11]) ? node19253 : 4'b1011;
															assign node19253 = (inp[9]) ? node19257 : node19254;
																assign node19254 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node19257 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node19260 = (inp[9]) ? node19264 : node19261;
														assign node19261 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node19264 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node19267 = (inp[9]) ? node19295 : node19268;
												assign node19268 = (inp[11]) ? node19282 : node19269;
													assign node19269 = (inp[5]) ? node19275 : node19270;
														assign node19270 = (inp[1]) ? 4'b1010 : node19271;
															assign node19271 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node19275 = (inp[1]) ? node19279 : node19276;
															assign node19276 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node19279 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node19282 = (inp[1]) ? node19290 : node19283;
														assign node19283 = (inp[2]) ? node19287 : node19284;
															assign node19284 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node19287 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node19290 = (inp[5]) ? node19292 : 4'b1011;
															assign node19292 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node19295 = (inp[11]) ? node19309 : node19296;
													assign node19296 = (inp[1]) ? node19304 : node19297;
														assign node19297 = (inp[2]) ? node19301 : node19298;
															assign node19298 = (inp[5]) ? 4'b1010 : 4'b1110;
															assign node19301 = (inp[5]) ? 4'b1011 : 4'b1111;
														assign node19304 = (inp[5]) ? node19306 : 4'b1011;
															assign node19306 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node19309 = (inp[1]) ? node19317 : node19310;
														assign node19310 = (inp[2]) ? node19314 : node19311;
															assign node19311 = (inp[5]) ? 4'b1011 : 4'b1111;
															assign node19314 = (inp[5]) ? 4'b1010 : 4'b1110;
														assign node19317 = (inp[5]) ? 4'b1110 : 4'b1010;
										assign node19320 = (inp[5]) ? node19382 : node19321;
											assign node19321 = (inp[1]) ? node19335 : node19322;
												assign node19322 = (inp[9]) ? node19330 : node19323;
													assign node19323 = (inp[11]) ? node19325 : 4'b1011;
														assign node19325 = (inp[2]) ? node19327 : 4'b1010;
															assign node19327 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node19330 = (inp[0]) ? node19332 : 4'b1010;
														assign node19332 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node19335 = (inp[10]) ? node19361 : node19336;
													assign node19336 = (inp[0]) ? node19350 : node19337;
														assign node19337 = (inp[11]) ? node19343 : node19338;
															assign node19338 = (inp[2]) ? 4'b1110 : node19339;
																assign node19339 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node19343 = (inp[2]) ? node19347 : node19344;
																assign node19344 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node19347 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node19350 = (inp[2]) ? node19356 : node19351;
															assign node19351 = (inp[9]) ? 4'b1111 : node19352;
																assign node19352 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node19356 = (inp[11]) ? node19358 : 4'b1111;
																assign node19358 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node19361 = (inp[0]) ? node19375 : node19362;
														assign node19362 = (inp[9]) ? node19368 : node19363;
															assign node19363 = (inp[2]) ? 4'b1111 : node19364;
																assign node19364 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node19368 = (inp[11]) ? node19372 : node19369;
																assign node19369 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node19372 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node19375 = (inp[9]) ? node19379 : node19376;
															assign node19376 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node19379 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node19382 = (inp[1]) ? node19404 : node19383;
												assign node19383 = (inp[9]) ? node19393 : node19384;
													assign node19384 = (inp[11]) ? node19388 : node19385;
														assign node19385 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node19388 = (inp[2]) ? 4'b1111 : node19389;
															assign node19389 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node19393 = (inp[11]) ? node19399 : node19394;
														assign node19394 = (inp[0]) ? node19396 : 4'b1111;
															assign node19396 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node19399 = (inp[0]) ? node19401 : 4'b1110;
															assign node19401 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node19404 = (inp[0]) ? node19420 : node19405;
													assign node19405 = (inp[9]) ? node19413 : node19406;
														assign node19406 = (inp[10]) ? 4'b1011 : node19407;
															assign node19407 = (inp[11]) ? 4'b1011 : node19408;
																assign node19408 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node19413 = (inp[2]) ? node19417 : node19414;
															assign node19414 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node19417 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node19420 = (inp[2]) ? node19426 : node19421;
														assign node19421 = (inp[11]) ? 4'b1011 : node19422;
															assign node19422 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node19426 = (inp[9]) ? node19430 : node19427;
															assign node19427 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node19430 = (inp[11]) ? 4'b1010 : 4'b1011;
								assign node19433 = (inp[1]) ? node19733 : node19434;
									assign node19434 = (inp[0]) ? node19588 : node19435;
										assign node19435 = (inp[4]) ? node19515 : node19436;
											assign node19436 = (inp[5]) ? node19486 : node19437;
												assign node19437 = (inp[13]) ? node19457 : node19438;
													assign node19438 = (inp[10]) ? node19452 : node19439;
														assign node19439 = (inp[2]) ? node19447 : node19440;
															assign node19440 = (inp[9]) ? node19444 : node19441;
																assign node19441 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node19444 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node19447 = (inp[9]) ? node19449 : 4'b1001;
																assign node19449 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19452 = (inp[11]) ? node19454 : 4'b1000;
															assign node19454 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node19457 = (inp[2]) ? node19473 : node19458;
														assign node19458 = (inp[10]) ? node19466 : node19459;
															assign node19459 = (inp[9]) ? node19463 : node19460;
																assign node19460 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node19463 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node19466 = (inp[11]) ? node19470 : node19467;
																assign node19467 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node19470 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node19473 = (inp[10]) ? node19479 : node19474;
															assign node19474 = (inp[9]) ? node19476 : 4'b1101;
																assign node19476 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node19479 = (inp[9]) ? node19483 : node19480;
																assign node19480 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node19483 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node19486 = (inp[13]) ? node19494 : node19487;
													assign node19487 = (inp[9]) ? node19491 : node19488;
														assign node19488 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node19491 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node19494 = (inp[11]) ? node19508 : node19495;
														assign node19495 = (inp[10]) ? node19503 : node19496;
															assign node19496 = (inp[2]) ? node19500 : node19497;
																assign node19497 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node19500 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node19503 = (inp[9]) ? 4'b1001 : node19504;
																assign node19504 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node19508 = (inp[2]) ? node19512 : node19509;
															assign node19509 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node19512 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node19515 = (inp[11]) ? node19559 : node19516;
												assign node19516 = (inp[10]) ? node19540 : node19517;
													assign node19517 = (inp[2]) ? node19531 : node19518;
														assign node19518 = (inp[9]) ? node19524 : node19519;
															assign node19519 = (inp[13]) ? 4'b1000 : node19520;
																assign node19520 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node19524 = (inp[13]) ? node19528 : node19525;
																assign node19525 = (inp[5]) ? 4'b1000 : 4'b1100;
																assign node19528 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node19531 = (inp[9]) ? node19535 : node19532;
															assign node19532 = (inp[13]) ? 4'b1101 : 4'b1000;
															assign node19535 = (inp[13]) ? 4'b1001 : node19536;
																assign node19536 = (inp[5]) ? 4'b1001 : 4'b1101;
													assign node19540 = (inp[9]) ? node19552 : node19541;
														assign node19541 = (inp[13]) ? node19547 : node19542;
															assign node19542 = (inp[2]) ? 4'b1100 : node19543;
																assign node19543 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node19547 = (inp[5]) ? node19549 : 4'b1000;
																assign node19549 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node19552 = (inp[5]) ? node19556 : node19553;
															assign node19553 = (inp[13]) ? 4'b1001 : 4'b1100;
															assign node19556 = (inp[2]) ? 4'b1100 : 4'b1000;
												assign node19559 = (inp[5]) ? node19569 : node19560;
													assign node19560 = (inp[13]) ? node19566 : node19561;
														assign node19561 = (inp[9]) ? node19563 : 4'b1100;
															assign node19563 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node19566 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node19569 = (inp[13]) ? node19577 : node19570;
														assign node19570 = (inp[9]) ? node19574 : node19571;
															assign node19571 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node19574 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node19577 = (inp[10]) ? node19583 : node19578;
															assign node19578 = (inp[9]) ? 4'b1100 : node19579;
																assign node19579 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node19583 = (inp[9]) ? node19585 : 4'b1100;
																assign node19585 = (inp[2]) ? 4'b1101 : 4'b1100;
										assign node19588 = (inp[4]) ? node19656 : node19589;
											assign node19589 = (inp[13]) ? node19629 : node19590;
												assign node19590 = (inp[5]) ? node19610 : node19591;
													assign node19591 = (inp[2]) ? node19599 : node19592;
														assign node19592 = (inp[11]) ? node19596 : node19593;
															assign node19593 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node19596 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node19599 = (inp[10]) ? node19605 : node19600;
															assign node19600 = (inp[9]) ? node19602 : 4'b1000;
																assign node19602 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node19605 = (inp[11]) ? 4'b1001 : node19606;
																assign node19606 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node19610 = (inp[2]) ? node19624 : node19611;
														assign node19611 = (inp[10]) ? node19619 : node19612;
															assign node19612 = (inp[11]) ? node19616 : node19613;
																assign node19613 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node19616 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node19619 = (inp[11]) ? 4'b1101 : node19620;
																assign node19620 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node19624 = (inp[11]) ? 4'b1100 : node19625;
															assign node19625 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node19629 = (inp[5]) ? node19645 : node19630;
													assign node19630 = (inp[9]) ? node19638 : node19631;
														assign node19631 = (inp[2]) ? node19635 : node19632;
															assign node19632 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node19635 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node19638 = (inp[2]) ? node19642 : node19639;
															assign node19639 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node19642 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node19645 = (inp[2]) ? node19651 : node19646;
														assign node19646 = (inp[11]) ? node19648 : 4'b1000;
															assign node19648 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node19651 = (inp[11]) ? node19653 : 4'b1001;
															assign node19653 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node19656 = (inp[2]) ? node19682 : node19657;
												assign node19657 = (inp[9]) ? node19669 : node19658;
													assign node19658 = (inp[11]) ? node19666 : node19659;
														assign node19659 = (inp[5]) ? node19663 : node19660;
															assign node19660 = (inp[13]) ? 4'b1001 : 4'b1101;
															assign node19663 = (inp[13]) ? 4'b1100 : 4'b1001;
														assign node19666 = (inp[13]) ? 4'b1101 : 4'b1100;
													assign node19669 = (inp[11]) ? node19675 : node19670;
														assign node19670 = (inp[13]) ? 4'b1101 : node19671;
															assign node19671 = (inp[5]) ? 4'b1000 : 4'b1100;
														assign node19675 = (inp[13]) ? node19679 : node19676;
															assign node19676 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node19679 = (inp[5]) ? 4'b1100 : 4'b1001;
												assign node19682 = (inp[10]) ? node19710 : node19683;
													assign node19683 = (inp[13]) ? node19697 : node19684;
														assign node19684 = (inp[5]) ? node19690 : node19685;
															assign node19685 = (inp[11]) ? 4'b1101 : node19686;
																assign node19686 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node19690 = (inp[9]) ? node19694 : node19691;
																assign node19691 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node19694 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node19697 = (inp[5]) ? node19703 : node19698;
															assign node19698 = (inp[11]) ? 4'b1000 : node19699;
																assign node19699 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node19703 = (inp[11]) ? node19707 : node19704;
																assign node19704 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node19707 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node19710 = (inp[9]) ? node19722 : node19711;
														assign node19711 = (inp[11]) ? node19717 : node19712;
															assign node19712 = (inp[13]) ? 4'b1000 : node19713;
																assign node19713 = (inp[5]) ? 4'b1001 : 4'b1101;
															assign node19717 = (inp[13]) ? node19719 : 4'b1000;
																assign node19719 = (inp[5]) ? 4'b1101 : 4'b1001;
														assign node19722 = (inp[11]) ? node19728 : node19723;
															assign node19723 = (inp[13]) ? node19725 : 4'b1100;
																assign node19725 = (inp[5]) ? 4'b1101 : 4'b1001;
															assign node19728 = (inp[13]) ? 4'b1100 : node19729;
																assign node19729 = (inp[5]) ? 4'b1001 : 4'b1101;
									assign node19733 = (inp[9]) ? node19823 : node19734;
										assign node19734 = (inp[11]) ? node19782 : node19735;
											assign node19735 = (inp[4]) ? node19763 : node19736;
												assign node19736 = (inp[0]) ? node19748 : node19737;
													assign node19737 = (inp[13]) ? node19745 : node19738;
														assign node19738 = (inp[5]) ? node19742 : node19739;
															assign node19739 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node19742 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node19745 = (inp[5]) ? 4'b1001 : 4'b1101;
													assign node19748 = (inp[2]) ? node19756 : node19749;
														assign node19749 = (inp[5]) ? node19753 : node19750;
															assign node19750 = (inp[13]) ? 4'b1100 : 4'b1001;
															assign node19753 = (inp[13]) ? 4'b1001 : 4'b1100;
														assign node19756 = (inp[5]) ? node19760 : node19757;
															assign node19757 = (inp[13]) ? 4'b1100 : 4'b1001;
															assign node19760 = (inp[13]) ? 4'b1000 : 4'b1100;
												assign node19763 = (inp[5]) ? node19775 : node19764;
													assign node19764 = (inp[13]) ? node19770 : node19765;
														assign node19765 = (inp[2]) ? node19767 : 4'b1001;
															assign node19767 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node19770 = (inp[2]) ? node19772 : 4'b1100;
															assign node19772 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node19775 = (inp[13]) ? node19777 : 4'b1100;
														assign node19777 = (inp[0]) ? 4'b1000 : node19778;
															assign node19778 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node19782 = (inp[2]) ? node19806 : node19783;
												assign node19783 = (inp[13]) ? node19797 : node19784;
													assign node19784 = (inp[5]) ? node19790 : node19785;
														assign node19785 = (inp[4]) ? 4'b1000 : node19786;
															assign node19786 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node19790 = (inp[4]) ? node19794 : node19791;
															assign node19791 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node19794 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node19797 = (inp[5]) ? node19803 : node19798;
														assign node19798 = (inp[0]) ? 4'b1101 : node19799;
															assign node19799 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node19803 = (inp[4]) ? 4'b1001 : 4'b1000;
												assign node19806 = (inp[5]) ? node19818 : node19807;
													assign node19807 = (inp[13]) ? node19813 : node19808;
														assign node19808 = (inp[0]) ? 4'b1000 : node19809;
															assign node19809 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node19813 = (inp[4]) ? node19815 : 4'b1101;
															assign node19815 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node19818 = (inp[13]) ? node19820 : 4'b1101;
														assign node19820 = (inp[0]) ? 4'b1001 : 4'b1000;
										assign node19823 = (inp[11]) ? node19865 : node19824;
											assign node19824 = (inp[2]) ? node19850 : node19825;
												assign node19825 = (inp[13]) ? node19841 : node19826;
													assign node19826 = (inp[5]) ? node19828 : 4'b1000;
														assign node19828 = (inp[10]) ? node19836 : node19829;
															assign node19829 = (inp[4]) ? node19833 : node19830;
																assign node19830 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node19833 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node19836 = (inp[4]) ? node19838 : 4'b1100;
																assign node19838 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node19841 = (inp[5]) ? node19847 : node19842;
														assign node19842 = (inp[0]) ? 4'b1101 : node19843;
															assign node19843 = (inp[4]) ? 4'b1101 : 4'b1100;
														assign node19847 = (inp[4]) ? 4'b1001 : 4'b1000;
												assign node19850 = (inp[13]) ? node19856 : node19851;
													assign node19851 = (inp[5]) ? 4'b1101 : node19852;
														assign node19852 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node19856 = (inp[5]) ? node19862 : node19857;
														assign node19857 = (inp[0]) ? 4'b1101 : node19858;
															assign node19858 = (inp[4]) ? 4'b1100 : 4'b1101;
														assign node19862 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node19865 = (inp[13]) ? node19891 : node19866;
												assign node19866 = (inp[5]) ? node19876 : node19867;
													assign node19867 = (inp[0]) ? 4'b1001 : node19868;
														assign node19868 = (inp[4]) ? node19872 : node19869;
															assign node19869 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node19872 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node19876 = (inp[2]) ? 4'b1100 : node19877;
														assign node19877 = (inp[10]) ? node19885 : node19878;
															assign node19878 = (inp[4]) ? node19882 : node19879;
																assign node19879 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node19882 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node19885 = (inp[4]) ? 4'b1101 : node19886;
																assign node19886 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node19891 = (inp[5]) ? node19903 : node19892;
													assign node19892 = (inp[0]) ? 4'b1100 : node19893;
														assign node19893 = (inp[10]) ? node19897 : node19894;
															assign node19894 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node19897 = (inp[4]) ? 4'b1100 : node19898;
																assign node19898 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node19903 = (inp[0]) ? node19909 : node19904;
														assign node19904 = (inp[2]) ? 4'b1001 : node19905;
															assign node19905 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node19909 = (inp[4]) ? 4'b1000 : node19910;
															assign node19910 = (inp[2]) ? 4'b1000 : 4'b1001;
					assign node19914 = (inp[13]) ? node21458 : node19915;
						assign node19915 = (inp[5]) ? node20861 : node19916;
							assign node19916 = (inp[1]) ? node20398 : node19917;
								assign node19917 = (inp[10]) ? node20173 : node19918;
									assign node19918 = (inp[2]) ? node20018 : node19919;
										assign node19919 = (inp[15]) ? node19961 : node19920;
											assign node19920 = (inp[4]) ? node19944 : node19921;
												assign node19921 = (inp[12]) ? node19929 : node19922;
													assign node19922 = (inp[11]) ? node19926 : node19923;
														assign node19923 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node19926 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node19929 = (inp[7]) ? node19937 : node19930;
														assign node19930 = (inp[11]) ? node19934 : node19931;
															assign node19931 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node19934 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node19937 = (inp[11]) ? node19941 : node19938;
															assign node19938 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node19941 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node19944 = (inp[12]) ? node19952 : node19945;
													assign node19945 = (inp[11]) ? node19949 : node19946;
														assign node19946 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node19949 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node19952 = (inp[7]) ? 4'b0010 : node19953;
														assign node19953 = (inp[0]) ? node19957 : node19954;
															assign node19954 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node19957 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node19961 = (inp[4]) ? node19999 : node19962;
												assign node19962 = (inp[12]) ? node19982 : node19963;
													assign node19963 = (inp[7]) ? node19969 : node19964;
														assign node19964 = (inp[11]) ? 4'b0010 : node19965;
															assign node19965 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node19969 = (inp[9]) ? node19977 : node19970;
															assign node19970 = (inp[0]) ? node19974 : node19971;
																assign node19971 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node19974 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node19977 = (inp[0]) ? 4'b0111 : node19978;
																assign node19978 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node19982 = (inp[0]) ? node19992 : node19983;
														assign node19983 = (inp[9]) ? 4'b0010 : node19984;
															assign node19984 = (inp[11]) ? node19988 : node19985;
																assign node19985 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node19988 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node19992 = (inp[11]) ? node19996 : node19993;
															assign node19993 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node19996 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node19999 = (inp[7]) ? node20009 : node20000;
													assign node20000 = (inp[12]) ? 4'b0000 : node20001;
														assign node20001 = (inp[11]) ? node20005 : node20002;
															assign node20002 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node20005 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node20009 = (inp[0]) ? 4'b0000 : node20010;
														assign node20010 = (inp[12]) ? node20014 : node20011;
															assign node20011 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20014 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node20018 = (inp[12]) ? node20090 : node20019;
											assign node20019 = (inp[15]) ? node20051 : node20020;
												assign node20020 = (inp[4]) ? node20036 : node20021;
													assign node20021 = (inp[7]) ? node20029 : node20022;
														assign node20022 = (inp[0]) ? node20026 : node20023;
															assign node20023 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20026 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node20029 = (inp[11]) ? node20033 : node20030;
															assign node20030 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node20033 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node20036 = (inp[7]) ? node20042 : node20037;
														assign node20037 = (inp[11]) ? 4'b0010 : node20038;
															assign node20038 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node20042 = (inp[9]) ? node20044 : 4'b0010;
															assign node20044 = (inp[11]) ? node20048 : node20045;
																assign node20045 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node20048 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node20051 = (inp[4]) ? node20071 : node20052;
													assign node20052 = (inp[7]) ? node20064 : node20053;
														assign node20053 = (inp[9]) ? node20059 : node20054;
															assign node20054 = (inp[11]) ? 4'b0010 : node20055;
																assign node20055 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node20059 = (inp[11]) ? node20061 : 4'b0010;
																assign node20061 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node20064 = (inp[0]) ? node20068 : node20065;
															assign node20065 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node20068 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node20071 = (inp[7]) ? node20081 : node20072;
														assign node20072 = (inp[9]) ? 4'b0100 : node20073;
															assign node20073 = (inp[11]) ? node20077 : node20074;
																assign node20074 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node20077 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node20081 = (inp[9]) ? node20087 : node20082;
															assign node20082 = (inp[11]) ? 4'b0000 : node20083;
																assign node20083 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node20087 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node20090 = (inp[15]) ? node20134 : node20091;
												assign node20091 = (inp[4]) ? node20111 : node20092;
													assign node20092 = (inp[7]) ? node20100 : node20093;
														assign node20093 = (inp[11]) ? node20097 : node20094;
															assign node20094 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node20097 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node20100 = (inp[9]) ? node20106 : node20101;
															assign node20101 = (inp[11]) ? 4'b0100 : node20102;
																assign node20102 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node20106 = (inp[0]) ? 4'b0101 : node20107;
																assign node20107 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node20111 = (inp[7]) ? node20119 : node20112;
														assign node20112 = (inp[11]) ? node20116 : node20113;
															assign node20113 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node20116 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node20119 = (inp[9]) ? node20127 : node20120;
															assign node20120 = (inp[0]) ? node20124 : node20121;
																assign node20121 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node20124 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node20127 = (inp[11]) ? node20131 : node20128;
																assign node20128 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node20131 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node20134 = (inp[4]) ? node20156 : node20135;
													assign node20135 = (inp[9]) ? node20149 : node20136;
														assign node20136 = (inp[0]) ? node20142 : node20137;
															assign node20137 = (inp[7]) ? 4'b0011 : node20138;
																assign node20138 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node20142 = (inp[11]) ? node20146 : node20143;
																assign node20143 = (inp[7]) ? 4'b0010 : 4'b0011;
																assign node20146 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node20149 = (inp[7]) ? node20151 : 4'b0011;
															assign node20151 = (inp[0]) ? 4'b0011 : node20152;
																assign node20152 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node20156 = (inp[0]) ? node20166 : node20157;
														assign node20157 = (inp[9]) ? node20159 : 4'b0000;
															assign node20159 = (inp[7]) ? node20163 : node20160;
																assign node20160 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node20163 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node20166 = (inp[11]) ? node20170 : node20167;
															assign node20167 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node20170 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node20173 = (inp[2]) ? node20299 : node20174;
										assign node20174 = (inp[7]) ? node20222 : node20175;
											assign node20175 = (inp[4]) ? node20191 : node20176;
												assign node20176 = (inp[15]) ? node20184 : node20177;
													assign node20177 = (inp[0]) ? node20181 : node20178;
														assign node20178 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node20181 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node20184 = (inp[11]) ? node20188 : node20185;
														assign node20185 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node20188 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node20191 = (inp[15]) ? node20207 : node20192;
													assign node20192 = (inp[12]) ? node20200 : node20193;
														assign node20193 = (inp[11]) ? node20197 : node20194;
															assign node20194 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node20197 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node20200 = (inp[11]) ? node20204 : node20201;
															assign node20201 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node20204 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node20207 = (inp[12]) ? node20215 : node20208;
														assign node20208 = (inp[0]) ? node20212 : node20209;
															assign node20209 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node20212 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node20215 = (inp[11]) ? node20219 : node20216;
															assign node20216 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node20219 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node20222 = (inp[4]) ? node20260 : node20223;
												assign node20223 = (inp[15]) ? node20239 : node20224;
													assign node20224 = (inp[12]) ? node20232 : node20225;
														assign node20225 = (inp[11]) ? node20229 : node20226;
															assign node20226 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node20229 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node20232 = (inp[0]) ? node20236 : node20233;
															assign node20233 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node20236 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node20239 = (inp[12]) ? node20253 : node20240;
														assign node20240 = (inp[9]) ? node20246 : node20241;
															assign node20241 = (inp[0]) ? node20243 : 4'b0110;
																assign node20243 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node20246 = (inp[11]) ? node20250 : node20247;
																assign node20247 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node20250 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node20253 = (inp[11]) ? node20257 : node20254;
															assign node20254 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node20257 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node20260 = (inp[15]) ? node20282 : node20261;
													assign node20261 = (inp[12]) ? node20269 : node20262;
														assign node20262 = (inp[0]) ? node20266 : node20263;
															assign node20263 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node20266 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node20269 = (inp[9]) ? node20275 : node20270;
															assign node20270 = (inp[0]) ? node20272 : 4'b0010;
																assign node20272 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node20275 = (inp[11]) ? node20279 : node20276;
																assign node20276 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node20279 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node20282 = (inp[9]) ? node20288 : node20283;
														assign node20283 = (inp[11]) ? 4'b0000 : node20284;
															assign node20284 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node20288 = (inp[0]) ? node20294 : node20289;
															assign node20289 = (inp[11]) ? node20291 : 4'b0001;
																assign node20291 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node20294 = (inp[11]) ? node20296 : 4'b0000;
																assign node20296 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node20299 = (inp[11]) ? node20347 : node20300;
											assign node20300 = (inp[4]) ? node20322 : node20301;
												assign node20301 = (inp[15]) ? node20311 : node20302;
													assign node20302 = (inp[7]) ? node20306 : node20303;
														assign node20303 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node20306 = (inp[12]) ? node20308 : 4'b0000;
															assign node20308 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node20311 = (inp[0]) ? node20315 : node20312;
														assign node20312 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node20315 = (inp[12]) ? node20319 : node20316;
															assign node20316 = (inp[7]) ? 4'b0111 : 4'b0011;
															assign node20319 = (inp[7]) ? 4'b0010 : 4'b0011;
												assign node20322 = (inp[15]) ? node20332 : node20323;
													assign node20323 = (inp[7]) ? 4'b0010 : node20324;
														assign node20324 = (inp[0]) ? node20328 : node20325;
															assign node20325 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node20328 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node20332 = (inp[7]) ? node20340 : node20333;
														assign node20333 = (inp[12]) ? node20337 : node20334;
															assign node20334 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node20337 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node20340 = (inp[0]) ? node20344 : node20341;
															assign node20341 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node20344 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node20347 = (inp[15]) ? node20373 : node20348;
												assign node20348 = (inp[4]) ? node20360 : node20349;
													assign node20349 = (inp[7]) ? node20353 : node20350;
														assign node20350 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node20353 = (inp[12]) ? node20357 : node20354;
															assign node20354 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node20357 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node20360 = (inp[7]) ? node20366 : node20361;
														assign node20361 = (inp[12]) ? node20363 : 4'b0011;
															assign node20363 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node20366 = (inp[12]) ? node20370 : node20367;
															assign node20367 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node20370 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node20373 = (inp[4]) ? node20383 : node20374;
													assign node20374 = (inp[7]) ? node20378 : node20375;
														assign node20375 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node20378 = (inp[12]) ? node20380 : 4'b0111;
															assign node20380 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node20383 = (inp[7]) ? node20391 : node20384;
														assign node20384 = (inp[12]) ? node20388 : node20385;
															assign node20385 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node20388 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node20391 = (inp[12]) ? node20395 : node20392;
															assign node20392 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node20395 = (inp[0]) ? 4'b0001 : 4'b0000;
								assign node20398 = (inp[10]) ? node20632 : node20399;
									assign node20399 = (inp[0]) ? node20523 : node20400;
										assign node20400 = (inp[7]) ? node20466 : node20401;
											assign node20401 = (inp[4]) ? node20435 : node20402;
												assign node20402 = (inp[15]) ? node20416 : node20403;
													assign node20403 = (inp[2]) ? node20409 : node20404;
														assign node20404 = (inp[12]) ? 4'b0100 : node20405;
															assign node20405 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node20409 = (inp[11]) ? node20413 : node20410;
															assign node20410 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node20413 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node20416 = (inp[12]) ? node20428 : node20417;
														assign node20417 = (inp[9]) ? node20423 : node20418;
															assign node20418 = (inp[2]) ? 4'b0110 : node20419;
																assign node20419 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node20423 = (inp[2]) ? node20425 : 4'b0110;
																assign node20425 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node20428 = (inp[2]) ? node20432 : node20429;
															assign node20429 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node20432 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node20435 = (inp[15]) ? node20445 : node20436;
													assign node20436 = (inp[12]) ? node20442 : node20437;
														assign node20437 = (inp[2]) ? 4'b0110 : node20438;
															assign node20438 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node20442 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node20445 = (inp[12]) ? node20459 : node20446;
														assign node20446 = (inp[9]) ? node20452 : node20447;
															assign node20447 = (inp[11]) ? 4'b0000 : node20448;
																assign node20448 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node20452 = (inp[2]) ? node20456 : node20453;
																assign node20453 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node20456 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node20459 = (inp[11]) ? node20463 : node20460;
															assign node20460 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node20463 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node20466 = (inp[4]) ? node20486 : node20467;
												assign node20467 = (inp[15]) ? node20475 : node20468;
													assign node20468 = (inp[12]) ? node20472 : node20469;
														assign node20469 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node20472 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node20475 = (inp[12]) ? node20479 : node20476;
														assign node20476 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node20479 = (inp[2]) ? node20483 : node20480;
															assign node20480 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node20483 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node20486 = (inp[15]) ? node20500 : node20487;
													assign node20487 = (inp[12]) ? node20495 : node20488;
														assign node20488 = (inp[11]) ? node20492 : node20489;
															assign node20489 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node20492 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node20495 = (inp[11]) ? node20497 : 4'b0110;
															assign node20497 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node20500 = (inp[12]) ? node20514 : node20501;
														assign node20501 = (inp[9]) ? node20509 : node20502;
															assign node20502 = (inp[11]) ? node20506 : node20503;
																assign node20503 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node20506 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node20509 = (inp[2]) ? 4'b0101 : node20510;
																assign node20510 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node20514 = (inp[9]) ? node20516 : 4'b0100;
															assign node20516 = (inp[2]) ? node20520 : node20517;
																assign node20517 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node20520 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node20523 = (inp[12]) ? node20573 : node20524;
											assign node20524 = (inp[15]) ? node20548 : node20525;
												assign node20525 = (inp[4]) ? node20529 : node20526;
													assign node20526 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node20529 = (inp[9]) ? node20539 : node20530;
														assign node20530 = (inp[7]) ? 4'b0110 : node20531;
															assign node20531 = (inp[11]) ? node20535 : node20532;
																assign node20532 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node20535 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node20539 = (inp[7]) ? 4'b0111 : node20540;
															assign node20540 = (inp[2]) ? node20544 : node20541;
																assign node20541 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node20544 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node20548 = (inp[4]) ? node20560 : node20549;
													assign node20549 = (inp[7]) ? node20557 : node20550;
														assign node20550 = (inp[9]) ? node20552 : 4'b0110;
															assign node20552 = (inp[11]) ? 4'b0111 : node20553;
																assign node20553 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node20557 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node20560 = (inp[7]) ? node20568 : node20561;
														assign node20561 = (inp[11]) ? node20565 : node20562;
															assign node20562 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node20565 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node20568 = (inp[11]) ? node20570 : 4'b0101;
															assign node20570 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node20573 = (inp[15]) ? node20593 : node20574;
												assign node20574 = (inp[4]) ? node20582 : node20575;
													assign node20575 = (inp[7]) ? node20579 : node20576;
														assign node20576 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node20579 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node20582 = (inp[7]) ? node20586 : node20583;
														assign node20583 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node20586 = (inp[11]) ? node20590 : node20587;
															assign node20587 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node20590 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node20593 = (inp[4]) ? node20609 : node20594;
													assign node20594 = (inp[2]) ? node20602 : node20595;
														assign node20595 = (inp[7]) ? node20599 : node20596;
															assign node20596 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node20599 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node20602 = (inp[7]) ? node20606 : node20603;
															assign node20603 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node20606 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node20609 = (inp[2]) ? node20623 : node20610;
														assign node20610 = (inp[9]) ? node20618 : node20611;
															assign node20611 = (inp[11]) ? node20615 : node20612;
																assign node20612 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node20615 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node20618 = (inp[11]) ? node20620 : 4'b0101;
																assign node20620 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node20623 = (inp[9]) ? 4'b0100 : node20624;
															assign node20624 = (inp[11]) ? node20628 : node20625;
																assign node20625 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node20628 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node20632 = (inp[2]) ? node20736 : node20633;
										assign node20633 = (inp[0]) ? node20685 : node20634;
											assign node20634 = (inp[11]) ? node20660 : node20635;
												assign node20635 = (inp[15]) ? node20649 : node20636;
													assign node20636 = (inp[4]) ? node20644 : node20637;
														assign node20637 = (inp[7]) ? node20641 : node20638;
															assign node20638 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node20641 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node20644 = (inp[7]) ? 4'b0110 : node20645;
															assign node20645 = (inp[12]) ? 4'b0011 : 4'b0110;
													assign node20649 = (inp[4]) ? node20655 : node20650;
														assign node20650 = (inp[7]) ? 4'b0110 : node20651;
															assign node20651 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node20655 = (inp[7]) ? 4'b0101 : node20656;
															assign node20656 = (inp[12]) ? 4'b0100 : 4'b0001;
												assign node20660 = (inp[15]) ? node20670 : node20661;
													assign node20661 = (inp[4]) ? node20667 : node20662;
														assign node20662 = (inp[12]) ? node20664 : 4'b0101;
															assign node20664 = (inp[7]) ? 4'b0001 : 4'b0100;
														assign node20667 = (inp[9]) ? 4'b0111 : 4'b0010;
													assign node20670 = (inp[4]) ? node20678 : node20671;
														assign node20671 = (inp[7]) ? node20675 : node20672;
															assign node20672 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node20675 = (inp[12]) ? 4'b0111 : 4'b0010;
														assign node20678 = (inp[12]) ? node20682 : node20679;
															assign node20679 = (inp[7]) ? 4'b0100 : 4'b0000;
															assign node20682 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node20685 = (inp[11]) ? node20711 : node20686;
												assign node20686 = (inp[15]) ? node20698 : node20687;
													assign node20687 = (inp[4]) ? node20693 : node20688;
														assign node20688 = (inp[12]) ? node20690 : 4'b0101;
															assign node20690 = (inp[7]) ? 4'b0001 : 4'b0100;
														assign node20693 = (inp[7]) ? 4'b0111 : node20694;
															assign node20694 = (inp[12]) ? 4'b0010 : 4'b0111;
													assign node20698 = (inp[4]) ? node20706 : node20699;
														assign node20699 = (inp[7]) ? node20703 : node20700;
															assign node20700 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node20703 = (inp[12]) ? 4'b0111 : 4'b0010;
														assign node20706 = (inp[12]) ? node20708 : 4'b0000;
															assign node20708 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node20711 = (inp[15]) ? node20723 : node20712;
													assign node20712 = (inp[4]) ? node20718 : node20713;
														assign node20713 = (inp[12]) ? node20715 : 4'b0100;
															assign node20715 = (inp[7]) ? 4'b0000 : 4'b0101;
														assign node20718 = (inp[12]) ? node20720 : 4'b0110;
															assign node20720 = (inp[7]) ? 4'b0110 : 4'b0011;
													assign node20723 = (inp[4]) ? node20731 : node20724;
														assign node20724 = (inp[7]) ? node20728 : node20725;
															assign node20725 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node20728 = (inp[12]) ? 4'b0110 : 4'b0011;
														assign node20731 = (inp[7]) ? 4'b0101 : node20732;
															assign node20732 = (inp[12]) ? 4'b0100 : 4'b0001;
										assign node20736 = (inp[7]) ? node20798 : node20737;
											assign node20737 = (inp[4]) ? node20765 : node20738;
												assign node20738 = (inp[15]) ? node20750 : node20739;
													assign node20739 = (inp[9]) ? node20741 : 4'b0101;
														assign node20741 = (inp[0]) ? node20743 : 4'b0101;
															assign node20743 = (inp[12]) ? node20747 : node20744;
																assign node20744 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node20747 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node20750 = (inp[0]) ? node20758 : node20751;
														assign node20751 = (inp[11]) ? node20755 : node20752;
															assign node20752 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node20755 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node20758 = (inp[11]) ? node20762 : node20759;
															assign node20759 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node20762 = (inp[12]) ? 4'b0110 : 4'b0111;
												assign node20765 = (inp[15]) ? node20781 : node20766;
													assign node20766 = (inp[12]) ? node20774 : node20767;
														assign node20767 = (inp[0]) ? node20771 : node20768;
															assign node20768 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node20771 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node20774 = (inp[11]) ? node20778 : node20775;
															assign node20775 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node20778 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node20781 = (inp[12]) ? node20791 : node20782;
														assign node20782 = (inp[9]) ? node20788 : node20783;
															assign node20783 = (inp[0]) ? node20785 : 4'b0000;
																assign node20785 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node20788 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node20791 = (inp[11]) ? node20795 : node20792;
															assign node20792 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node20795 = (inp[0]) ? 4'b0101 : 4'b0100;
											assign node20798 = (inp[4]) ? node20830 : node20799;
												assign node20799 = (inp[15]) ? node20815 : node20800;
													assign node20800 = (inp[12]) ? node20808 : node20801;
														assign node20801 = (inp[0]) ? node20805 : node20802;
															assign node20802 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node20805 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node20808 = (inp[0]) ? node20812 : node20809;
															assign node20809 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node20812 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node20815 = (inp[12]) ? node20823 : node20816;
														assign node20816 = (inp[0]) ? node20820 : node20817;
															assign node20817 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node20820 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node20823 = (inp[0]) ? node20827 : node20824;
															assign node20824 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node20827 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node20830 = (inp[15]) ? node20842 : node20831;
													assign node20831 = (inp[12]) ? node20837 : node20832;
														assign node20832 = (inp[0]) ? node20834 : 4'b0110;
															assign node20834 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node20837 = (inp[11]) ? 4'b0111 : node20838;
															assign node20838 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node20842 = (inp[12]) ? node20852 : node20843;
														assign node20843 = (inp[9]) ? node20845 : 4'b0100;
															assign node20845 = (inp[0]) ? node20849 : node20846;
																assign node20846 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node20849 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node20852 = (inp[9]) ? 4'b0101 : node20853;
															assign node20853 = (inp[11]) ? node20857 : node20854;
																assign node20854 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node20857 = (inp[0]) ? 4'b0100 : 4'b0101;
							assign node20861 = (inp[1]) ? node21033 : node20862;
								assign node20862 = (inp[11]) ? node20956 : node20863;
									assign node20863 = (inp[0]) ? node20919 : node20864;
										assign node20864 = (inp[2]) ? node20892 : node20865;
											assign node20865 = (inp[4]) ? node20879 : node20866;
												assign node20866 = (inp[15]) ? node20874 : node20867;
													assign node20867 = (inp[12]) ? node20871 : node20868;
														assign node20868 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node20871 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node20874 = (inp[12]) ? 4'b0110 : node20875;
														assign node20875 = (inp[7]) ? 4'b0011 : 4'b0110;
												assign node20879 = (inp[15]) ? node20887 : node20880;
													assign node20880 = (inp[12]) ? node20884 : node20881;
														assign node20881 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node20884 = (inp[7]) ? 4'b0110 : 4'b0011;
													assign node20887 = (inp[12]) ? 4'b0101 : node20888;
														assign node20888 = (inp[7]) ? 4'b0100 : 4'b0001;
											assign node20892 = (inp[12]) ? node20908 : node20893;
												assign node20893 = (inp[7]) ? node20901 : node20894;
													assign node20894 = (inp[15]) ? node20898 : node20895;
														assign node20895 = (inp[4]) ? 4'b0110 : 4'b0100;
														assign node20898 = (inp[4]) ? 4'b0000 : 4'b0110;
													assign node20901 = (inp[15]) ? node20905 : node20902;
														assign node20902 = (inp[4]) ? 4'b0111 : 4'b0101;
														assign node20905 = (inp[4]) ? 4'b0101 : 4'b0010;
												assign node20908 = (inp[15]) ? node20916 : node20909;
													assign node20909 = (inp[4]) ? node20913 : node20910;
														assign node20910 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node20913 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node20916 = (inp[4]) ? 4'b0100 : 4'b0110;
										assign node20919 = (inp[12]) ? node20941 : node20920;
											assign node20920 = (inp[7]) ? node20930 : node20921;
												assign node20921 = (inp[15]) ? node20925 : node20922;
													assign node20922 = (inp[4]) ? 4'b0111 : 4'b0101;
													assign node20925 = (inp[4]) ? node20927 : 4'b0111;
														assign node20927 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node20930 = (inp[15]) ? node20934 : node20931;
													assign node20931 = (inp[4]) ? 4'b0110 : 4'b0100;
													assign node20934 = (inp[4]) ? node20938 : node20935;
														assign node20935 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node20938 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node20941 = (inp[15]) ? node20951 : node20942;
												assign node20942 = (inp[4]) ? node20946 : node20943;
													assign node20943 = (inp[7]) ? 4'b0001 : 4'b0101;
													assign node20946 = (inp[7]) ? 4'b0111 : node20947;
														assign node20947 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node20951 = (inp[4]) ? node20953 : 4'b0111;
													assign node20953 = (inp[2]) ? 4'b0101 : 4'b0100;
									assign node20956 = (inp[0]) ? node20994 : node20957;
										assign node20957 = (inp[7]) ? node20973 : node20958;
											assign node20958 = (inp[4]) ? node20962 : node20959;
												assign node20959 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node20962 = (inp[15]) ? node20968 : node20963;
													assign node20963 = (inp[12]) ? node20965 : 4'b0111;
														assign node20965 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node20968 = (inp[12]) ? node20970 : 4'b0001;
														assign node20970 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node20973 = (inp[12]) ? node20985 : node20974;
												assign node20974 = (inp[15]) ? node20978 : node20975;
													assign node20975 = (inp[4]) ? 4'b0110 : 4'b0100;
													assign node20978 = (inp[4]) ? node20982 : node20979;
														assign node20979 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node20982 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node20985 = (inp[4]) ? node20989 : node20986;
													assign node20986 = (inp[15]) ? 4'b0111 : 4'b0001;
													assign node20989 = (inp[15]) ? node20991 : 4'b0111;
														assign node20991 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node20994 = (inp[7]) ? node21012 : node20995;
											assign node20995 = (inp[4]) ? node20999 : node20996;
												assign node20996 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node20999 = (inp[15]) ? node21005 : node21000;
													assign node21000 = (inp[12]) ? node21002 : 4'b0110;
														assign node21002 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node21005 = (inp[12]) ? node21009 : node21006;
														assign node21006 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node21009 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node21012 = (inp[12]) ? node21024 : node21013;
												assign node21013 = (inp[15]) ? node21017 : node21014;
													assign node21014 = (inp[4]) ? 4'b0111 : 4'b0101;
													assign node21017 = (inp[4]) ? node21021 : node21018;
														assign node21018 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node21021 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node21024 = (inp[4]) ? node21028 : node21025;
													assign node21025 = (inp[15]) ? 4'b0110 : 4'b0000;
													assign node21028 = (inp[15]) ? node21030 : 4'b0110;
														assign node21030 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node21033 = (inp[0]) ? node21275 : node21034;
									assign node21034 = (inp[10]) ? node21196 : node21035;
										assign node21035 = (inp[9]) ? node21105 : node21036;
											assign node21036 = (inp[12]) ? node21070 : node21037;
												assign node21037 = (inp[11]) ? node21051 : node21038;
													assign node21038 = (inp[4]) ? node21044 : node21039;
														assign node21039 = (inp[15]) ? node21041 : 4'b0001;
															assign node21041 = (inp[7]) ? 4'b0110 : 4'b0011;
														assign node21044 = (inp[2]) ? node21048 : node21045;
															assign node21045 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node21048 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node21051 = (inp[15]) ? node21061 : node21052;
														assign node21052 = (inp[4]) ? node21054 : 4'b0000;
															assign node21054 = (inp[2]) ? node21058 : node21055;
																assign node21055 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node21058 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node21061 = (inp[4]) ? node21065 : node21062;
															assign node21062 = (inp[7]) ? 4'b0111 : 4'b0010;
															assign node21065 = (inp[7]) ? node21067 : 4'b0100;
																assign node21067 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node21070 = (inp[15]) ? node21096 : node21071;
													assign node21071 = (inp[4]) ? node21081 : node21072;
														assign node21072 = (inp[7]) ? node21078 : node21073;
															assign node21073 = (inp[2]) ? 4'b0000 : node21074;
																assign node21074 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node21078 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node21081 = (inp[7]) ? node21089 : node21082;
															assign node21082 = (inp[11]) ? node21086 : node21083;
																assign node21083 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node21086 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node21089 = (inp[11]) ? node21093 : node21090;
																assign node21090 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node21093 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node21096 = (inp[4]) ? node21100 : node21097;
														assign node21097 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node21100 = (inp[11]) ? 4'b0001 : node21101;
															assign node21101 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node21105 = (inp[2]) ? node21153 : node21106;
												assign node21106 = (inp[4]) ? node21132 : node21107;
													assign node21107 = (inp[15]) ? node21119 : node21108;
														assign node21108 = (inp[11]) ? node21114 : node21109;
															assign node21109 = (inp[7]) ? 4'b0001 : node21110;
																assign node21110 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node21114 = (inp[12]) ? 4'b0000 : node21115;
																assign node21115 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node21119 = (inp[7]) ? node21125 : node21120;
															assign node21120 = (inp[12]) ? 4'b0011 : node21121;
																assign node21121 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node21125 = (inp[11]) ? node21129 : node21126;
																assign node21126 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node21129 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node21132 = (inp[15]) ? node21142 : node21133;
														assign node21133 = (inp[11]) ? node21139 : node21134;
															assign node21134 = (inp[12]) ? 4'b0110 : node21135;
																assign node21135 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node21139 = (inp[7]) ? 4'b0011 : 4'b0111;
														assign node21142 = (inp[11]) ? node21148 : node21143;
															assign node21143 = (inp[7]) ? 4'b0001 : node21144;
																assign node21144 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node21148 = (inp[7]) ? 4'b0000 : node21149;
																assign node21149 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node21153 = (inp[11]) ? node21173 : node21154;
													assign node21154 = (inp[15]) ? node21164 : node21155;
														assign node21155 = (inp[4]) ? 4'b0010 : node21156;
															assign node21156 = (inp[7]) ? node21160 : node21157;
																assign node21157 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node21160 = (inp[12]) ? 4'b0101 : 4'b0000;
														assign node21164 = (inp[4]) ? 4'b0000 : node21165;
															assign node21165 = (inp[7]) ? node21169 : node21166;
																assign node21166 = (inp[12]) ? 4'b0010 : 4'b0011;
																assign node21169 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node21173 = (inp[15]) ? node21185 : node21174;
														assign node21174 = (inp[4]) ? node21182 : node21175;
															assign node21175 = (inp[7]) ? node21179 : node21176;
																assign node21176 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node21179 = (inp[12]) ? 4'b0100 : 4'b0001;
															assign node21182 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node21185 = (inp[4]) ? node21191 : node21186;
															assign node21186 = (inp[7]) ? 4'b0111 : node21187;
																assign node21187 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node21191 = (inp[7]) ? 4'b0001 : node21192;
																assign node21192 = (inp[12]) ? 4'b0001 : 4'b0100;
										assign node21196 = (inp[12]) ? node21238 : node21197;
											assign node21197 = (inp[15]) ? node21221 : node21198;
												assign node21198 = (inp[4]) ? node21208 : node21199;
													assign node21199 = (inp[9]) ? 4'b0000 : node21200;
														assign node21200 = (inp[2]) ? 4'b0001 : node21201;
															assign node21201 = (inp[7]) ? node21203 : 4'b0001;
																assign node21203 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node21208 = (inp[11]) ? node21216 : node21209;
														assign node21209 = (inp[7]) ? node21213 : node21210;
															assign node21210 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node21213 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node21216 = (inp[7]) ? node21218 : 4'b0011;
															assign node21218 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node21221 = (inp[4]) ? node21229 : node21222;
													assign node21222 = (inp[7]) ? node21226 : node21223;
														assign node21223 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node21226 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node21229 = (inp[7]) ? node21233 : node21230;
														assign node21230 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node21233 = (inp[2]) ? 4'b0000 : node21234;
															assign node21234 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node21238 = (inp[15]) ? node21264 : node21239;
												assign node21239 = (inp[4]) ? node21249 : node21240;
													assign node21240 = (inp[7]) ? node21246 : node21241;
														assign node21241 = (inp[11]) ? node21243 : 4'b0000;
															assign node21243 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node21246 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node21249 = (inp[7]) ? node21257 : node21250;
														assign node21250 = (inp[11]) ? node21254 : node21251;
															assign node21251 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node21254 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node21257 = (inp[2]) ? node21261 : node21258;
															assign node21258 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node21261 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node21264 = (inp[4]) ? node21268 : node21265;
													assign node21265 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node21268 = (inp[2]) ? node21272 : node21269;
														assign node21269 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node21272 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node21275 = (inp[7]) ? node21395 : node21276;
										assign node21276 = (inp[4]) ? node21332 : node21277;
											assign node21277 = (inp[15]) ? node21301 : node21278;
												assign node21278 = (inp[11]) ? node21294 : node21279;
													assign node21279 = (inp[9]) ? node21287 : node21280;
														assign node21280 = (inp[12]) ? node21284 : node21281;
															assign node21281 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node21284 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node21287 = (inp[12]) ? node21291 : node21288;
															assign node21288 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node21291 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node21294 = (inp[2]) ? node21298 : node21295;
														assign node21295 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node21298 = (inp[12]) ? 4'b0000 : 4'b0001;
												assign node21301 = (inp[10]) ? node21317 : node21302;
													assign node21302 = (inp[9]) ? node21310 : node21303;
														assign node21303 = (inp[11]) ? node21307 : node21304;
															assign node21304 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node21307 = (inp[12]) ? 4'b0010 : 4'b0011;
														assign node21310 = (inp[2]) ? 4'b0011 : node21311;
															assign node21311 = (inp[12]) ? 4'b0010 : node21312;
																assign node21312 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node21317 = (inp[2]) ? node21325 : node21318;
														assign node21318 = (inp[12]) ? node21322 : node21319;
															assign node21319 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node21322 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node21325 = (inp[11]) ? node21329 : node21326;
															assign node21326 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node21329 = (inp[12]) ? 4'b0010 : 4'b0011;
											assign node21332 = (inp[15]) ? node21376 : node21333;
												assign node21333 = (inp[12]) ? node21357 : node21334;
													assign node21334 = (inp[9]) ? node21344 : node21335;
														assign node21335 = (inp[10]) ? node21337 : 4'b0011;
															assign node21337 = (inp[2]) ? node21341 : node21338;
																assign node21338 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node21341 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node21344 = (inp[10]) ? node21350 : node21345;
															assign node21345 = (inp[2]) ? node21347 : 4'b0010;
																assign node21347 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node21350 = (inp[2]) ? node21354 : node21351;
																assign node21351 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node21354 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node21357 = (inp[9]) ? node21371 : node21358;
														assign node21358 = (inp[10]) ? node21366 : node21359;
															assign node21359 = (inp[11]) ? node21363 : node21360;
																assign node21360 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node21363 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node21366 = (inp[11]) ? 4'b0110 : node21367;
																assign node21367 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node21371 = (inp[11]) ? node21373 : 4'b0110;
															assign node21373 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node21376 = (inp[12]) ? node21380 : node21377;
													assign node21377 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node21380 = (inp[9]) ? node21388 : node21381;
														assign node21381 = (inp[2]) ? node21385 : node21382;
															assign node21382 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node21385 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node21388 = (inp[2]) ? node21392 : node21389;
															assign node21389 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node21392 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node21395 = (inp[4]) ? node21423 : node21396;
											assign node21396 = (inp[15]) ? node21416 : node21397;
												assign node21397 = (inp[12]) ? node21413 : node21398;
													assign node21398 = (inp[10]) ? node21406 : node21399;
														assign node21399 = (inp[9]) ? 4'b0001 : node21400;
															assign node21400 = (inp[2]) ? node21402 : 4'b0001;
																assign node21402 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node21406 = (inp[2]) ? node21410 : node21407;
															assign node21407 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node21410 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node21413 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node21416 = (inp[12]) ? node21420 : node21417;
													assign node21417 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node21420 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node21423 = (inp[15]) ? node21451 : node21424;
												assign node21424 = (inp[10]) ? node21432 : node21425;
													assign node21425 = (inp[11]) ? node21429 : node21426;
														assign node21426 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node21429 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node21432 = (inp[12]) ? node21444 : node21433;
														assign node21433 = (inp[9]) ? node21439 : node21434;
															assign node21434 = (inp[11]) ? 4'b0010 : node21435;
																assign node21435 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node21439 = (inp[11]) ? node21441 : 4'b0010;
																assign node21441 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node21444 = (inp[2]) ? node21448 : node21445;
															assign node21445 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node21448 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node21451 = (inp[11]) ? node21455 : node21452;
													assign node21452 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node21455 = (inp[2]) ? 4'b0000 : 4'b0001;
						assign node21458 = (inp[5]) ? node22194 : node21459;
							assign node21459 = (inp[1]) ? node21741 : node21460;
								assign node21460 = (inp[0]) ? node21574 : node21461;
									assign node21461 = (inp[2]) ? node21519 : node21462;
										assign node21462 = (inp[11]) ? node21492 : node21463;
											assign node21463 = (inp[15]) ? node21477 : node21464;
												assign node21464 = (inp[4]) ? node21470 : node21465;
													assign node21465 = (inp[12]) ? node21467 : 4'b0000;
														assign node21467 = (inp[7]) ? 4'b0101 : 4'b0000;
													assign node21470 = (inp[7]) ? node21474 : node21471;
														assign node21471 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node21474 = (inp[12]) ? 4'b0011 : 4'b0010;
												assign node21477 = (inp[4]) ? node21485 : node21478;
													assign node21478 = (inp[12]) ? node21482 : node21479;
														assign node21479 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node21482 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node21485 = (inp[12]) ? node21489 : node21486;
														assign node21486 = (inp[7]) ? 4'b0000 : 4'b0101;
														assign node21489 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node21492 = (inp[15]) ? node21506 : node21493;
												assign node21493 = (inp[4]) ? node21499 : node21494;
													assign node21494 = (inp[12]) ? node21496 : 4'b0001;
														assign node21496 = (inp[7]) ? 4'b0100 : 4'b0001;
													assign node21499 = (inp[7]) ? node21503 : node21500;
														assign node21500 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node21503 = (inp[12]) ? 4'b0010 : 4'b0011;
												assign node21506 = (inp[4]) ? node21512 : node21507;
													assign node21507 = (inp[7]) ? node21509 : 4'b0010;
														assign node21509 = (inp[12]) ? 4'b0011 : 4'b0110;
													assign node21512 = (inp[12]) ? node21516 : node21513;
														assign node21513 = (inp[7]) ? 4'b0001 : 4'b0100;
														assign node21516 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node21519 = (inp[11]) ? node21547 : node21520;
											assign node21520 = (inp[12]) ? node21532 : node21521;
												assign node21521 = (inp[15]) ? node21525 : node21522;
													assign node21522 = (inp[4]) ? 4'b0010 : 4'b0001;
													assign node21525 = (inp[4]) ? node21529 : node21526;
														assign node21526 = (inp[7]) ? 4'b0110 : 4'b0010;
														assign node21529 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node21532 = (inp[15]) ? node21540 : node21533;
													assign node21533 = (inp[4]) ? node21537 : node21534;
														assign node21534 = (inp[7]) ? 4'b0101 : 4'b0001;
														assign node21537 = (inp[7]) ? 4'b0011 : 4'b0110;
													assign node21540 = (inp[4]) ? node21544 : node21541;
														assign node21541 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node21544 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node21547 = (inp[15]) ? node21559 : node21548;
												assign node21548 = (inp[4]) ? node21554 : node21549;
													assign node21549 = (inp[12]) ? node21551 : 4'b0000;
														assign node21551 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node21554 = (inp[12]) ? node21556 : 4'b0011;
														assign node21556 = (inp[7]) ? 4'b0010 : 4'b0111;
												assign node21559 = (inp[4]) ? node21567 : node21560;
													assign node21560 = (inp[12]) ? node21564 : node21561;
														assign node21561 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node21564 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node21567 = (inp[12]) ? node21571 : node21568;
														assign node21568 = (inp[7]) ? 4'b0000 : 4'b0100;
														assign node21571 = (inp[7]) ? 4'b0001 : 4'b0000;
									assign node21574 = (inp[15]) ? node21628 : node21575;
										assign node21575 = (inp[4]) ? node21617 : node21576;
											assign node21576 = (inp[7]) ? node21592 : node21577;
												assign node21577 = (inp[10]) ? node21585 : node21578;
													assign node21578 = (inp[2]) ? node21582 : node21579;
														assign node21579 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node21582 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node21585 = (inp[2]) ? node21589 : node21586;
														assign node21586 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node21589 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node21592 = (inp[12]) ? node21614 : node21593;
													assign node21593 = (inp[10]) ? node21599 : node21594;
														assign node21594 = (inp[11]) ? 4'b0001 : node21595;
															assign node21595 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node21599 = (inp[9]) ? node21607 : node21600;
															assign node21600 = (inp[11]) ? node21604 : node21601;
																assign node21601 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node21604 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node21607 = (inp[11]) ? node21611 : node21608;
																assign node21608 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node21611 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node21614 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node21617 = (inp[11]) ? node21623 : node21618;
												assign node21618 = (inp[12]) ? node21620 : 4'b0011;
													assign node21620 = (inp[7]) ? 4'b0010 : 4'b0111;
												assign node21623 = (inp[12]) ? node21625 : 4'b0010;
													assign node21625 = (inp[7]) ? 4'b0011 : 4'b0110;
										assign node21628 = (inp[4]) ? node21672 : node21629;
											assign node21629 = (inp[7]) ? node21651 : node21630;
												assign node21630 = (inp[12]) ? node21638 : node21631;
													assign node21631 = (inp[11]) ? node21635 : node21632;
														assign node21632 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node21635 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node21638 = (inp[9]) ? node21646 : node21639;
														assign node21639 = (inp[2]) ? node21643 : node21640;
															assign node21640 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node21643 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node21646 = (inp[10]) ? 4'b0011 : node21647;
															assign node21647 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node21651 = (inp[12]) ? node21665 : node21652;
													assign node21652 = (inp[9]) ? node21660 : node21653;
														assign node21653 = (inp[2]) ? node21657 : node21654;
															assign node21654 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node21657 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node21660 = (inp[11]) ? node21662 : 4'b0111;
															assign node21662 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node21665 = (inp[2]) ? node21669 : node21666;
														assign node21666 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node21669 = (inp[11]) ? 4'b0011 : 4'b0010;
											assign node21672 = (inp[7]) ? node21692 : node21673;
												assign node21673 = (inp[12]) ? node21677 : node21674;
													assign node21674 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node21677 = (inp[9]) ? node21685 : node21678;
														assign node21678 = (inp[11]) ? node21682 : node21679;
															assign node21679 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node21682 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node21685 = (inp[2]) ? node21689 : node21686;
															assign node21686 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node21689 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node21692 = (inp[10]) ? node21722 : node21693;
													assign node21693 = (inp[11]) ? node21709 : node21694;
														assign node21694 = (inp[9]) ? node21702 : node21695;
															assign node21695 = (inp[2]) ? node21699 : node21696;
																assign node21696 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node21699 = (inp[12]) ? 4'b0001 : 4'b0000;
															assign node21702 = (inp[2]) ? node21706 : node21703;
																assign node21703 = (inp[12]) ? 4'b0000 : 4'b0001;
																assign node21706 = (inp[12]) ? 4'b0001 : 4'b0000;
														assign node21709 = (inp[9]) ? node21717 : node21710;
															assign node21710 = (inp[2]) ? node21714 : node21711;
																assign node21711 = (inp[12]) ? 4'b0001 : 4'b0000;
																assign node21714 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node21717 = (inp[2]) ? 4'b0001 : node21718;
																assign node21718 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node21722 = (inp[9]) ? node21734 : node21723;
														assign node21723 = (inp[2]) ? node21729 : node21724;
															assign node21724 = (inp[12]) ? 4'b0001 : node21725;
																assign node21725 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node21729 = (inp[11]) ? node21731 : 4'b0000;
																assign node21731 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node21734 = (inp[12]) ? 4'b0000 : node21735;
															assign node21735 = (inp[11]) ? node21737 : 4'b0000;
																assign node21737 = (inp[2]) ? 4'b0001 : 4'b0000;
								assign node21741 = (inp[10]) ? node21931 : node21742;
									assign node21742 = (inp[0]) ? node21836 : node21743;
										assign node21743 = (inp[11]) ? node21781 : node21744;
											assign node21744 = (inp[7]) ? node21766 : node21745;
												assign node21745 = (inp[12]) ? node21757 : node21746;
													assign node21746 = (inp[2]) ? node21752 : node21747;
														assign node21747 = (inp[15]) ? 4'b0000 : node21748;
															assign node21748 = (inp[4]) ? 4'b0110 : 4'b0100;
														assign node21752 = (inp[4]) ? 4'b0110 : node21753;
															assign node21753 = (inp[15]) ? 4'b0110 : 4'b0101;
													assign node21757 = (inp[15]) ? node21763 : node21758;
														assign node21758 = (inp[4]) ? node21760 : 4'b0101;
															assign node21760 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node21763 = (inp[4]) ? 4'b0101 : 4'b0111;
												assign node21766 = (inp[4]) ? node21778 : node21767;
													assign node21767 = (inp[15]) ? node21773 : node21768;
														assign node21768 = (inp[2]) ? node21770 : 4'b0100;
															assign node21770 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node21773 = (inp[12]) ? 4'b0110 : node21774;
															assign node21774 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node21778 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node21781 = (inp[2]) ? node21809 : node21782;
												assign node21782 = (inp[12]) ? node21794 : node21783;
													assign node21783 = (inp[15]) ? node21787 : node21784;
														assign node21784 = (inp[4]) ? 4'b0111 : 4'b0101;
														assign node21787 = (inp[4]) ? node21791 : node21788;
															assign node21788 = (inp[7]) ? 4'b0011 : 4'b0111;
															assign node21791 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node21794 = (inp[7]) ? node21802 : node21795;
														assign node21795 = (inp[15]) ? node21799 : node21796;
															assign node21796 = (inp[9]) ? 4'b0011 : 4'b0100;
															assign node21799 = (inp[4]) ? 4'b0100 : 4'b0110;
														assign node21802 = (inp[15]) ? node21806 : node21803;
															assign node21803 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node21806 = (inp[4]) ? 4'b0101 : 4'b0111;
												assign node21809 = (inp[4]) ? node21823 : node21810;
													assign node21810 = (inp[15]) ? node21816 : node21811;
														assign node21811 = (inp[12]) ? node21813 : 4'b0100;
															assign node21813 = (inp[7]) ? 4'b0000 : 4'b0101;
														assign node21816 = (inp[12]) ? node21820 : node21817;
															assign node21817 = (inp[7]) ? 4'b0010 : 4'b0111;
															assign node21820 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node21823 = (inp[15]) ? node21829 : node21824;
														assign node21824 = (inp[12]) ? node21826 : 4'b0111;
															assign node21826 = (inp[7]) ? 4'b0111 : 4'b0010;
														assign node21829 = (inp[12]) ? node21833 : node21830;
															assign node21830 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node21833 = (inp[7]) ? 4'b0101 : 4'b0100;
										assign node21836 = (inp[11]) ? node21892 : node21837;
											assign node21837 = (inp[2]) ? node21863 : node21838;
												assign node21838 = (inp[7]) ? node21852 : node21839;
													assign node21839 = (inp[4]) ? node21845 : node21840;
														assign node21840 = (inp[15]) ? 4'b0110 : node21841;
															assign node21841 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node21845 = (inp[15]) ? node21849 : node21846;
															assign node21846 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node21849 = (inp[12]) ? 4'b0100 : 4'b0001;
													assign node21852 = (inp[4]) ? node21860 : node21853;
														assign node21853 = (inp[15]) ? node21857 : node21854;
															assign node21854 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node21857 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node21860 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node21863 = (inp[4]) ? node21879 : node21864;
													assign node21864 = (inp[15]) ? node21872 : node21865;
														assign node21865 = (inp[7]) ? node21869 : node21866;
															assign node21866 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node21869 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node21872 = (inp[12]) ? node21876 : node21873;
															assign node21873 = (inp[7]) ? 4'b0010 : 4'b0111;
															assign node21876 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node21879 = (inp[15]) ? node21885 : node21880;
														assign node21880 = (inp[12]) ? node21882 : 4'b0111;
															assign node21882 = (inp[7]) ? 4'b0111 : 4'b0010;
														assign node21885 = (inp[12]) ? node21889 : node21886;
															assign node21886 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node21889 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node21892 = (inp[4]) ? node21916 : node21893;
												assign node21893 = (inp[15]) ? node21907 : node21894;
													assign node21894 = (inp[2]) ? node21902 : node21895;
														assign node21895 = (inp[7]) ? node21899 : node21896;
															assign node21896 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node21899 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node21902 = (inp[12]) ? node21904 : 4'b0101;
															assign node21904 = (inp[9]) ? 4'b0100 : 4'b0001;
													assign node21907 = (inp[12]) ? node21913 : node21908;
														assign node21908 = (inp[7]) ? node21910 : 4'b0110;
															assign node21910 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node21913 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node21916 = (inp[15]) ? node21924 : node21917;
													assign node21917 = (inp[12]) ? node21919 : 4'b0110;
														assign node21919 = (inp[7]) ? 4'b0110 : node21920;
															assign node21920 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node21924 = (inp[12]) ? node21928 : node21925;
														assign node21925 = (inp[7]) ? 4'b0100 : 4'b0000;
														assign node21928 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node21931 = (inp[2]) ? node22091 : node21932;
										assign node21932 = (inp[4]) ? node22012 : node21933;
											assign node21933 = (inp[15]) ? node21983 : node21934;
												assign node21934 = (inp[7]) ? node21956 : node21935;
													assign node21935 = (inp[0]) ? node21943 : node21936;
														assign node21936 = (inp[12]) ? node21940 : node21937;
															assign node21937 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node21940 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node21943 = (inp[9]) ? node21949 : node21944;
															assign node21944 = (inp[12]) ? node21946 : 4'b0100;
																assign node21946 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node21949 = (inp[12]) ? node21953 : node21950;
																assign node21950 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node21953 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node21956 = (inp[12]) ? node21968 : node21957;
														assign node21957 = (inp[9]) ? node21963 : node21958;
															assign node21958 = (inp[0]) ? node21960 : 4'b0101;
																assign node21960 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node21963 = (inp[11]) ? node21965 : 4'b0100;
																assign node21965 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node21968 = (inp[9]) ? node21976 : node21969;
															assign node21969 = (inp[0]) ? node21973 : node21970;
																assign node21970 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node21973 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node21976 = (inp[11]) ? node21980 : node21977;
																assign node21977 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node21980 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node21983 = (inp[12]) ? node21997 : node21984;
													assign node21984 = (inp[7]) ? node21990 : node21985;
														assign node21985 = (inp[11]) ? 4'b0110 : node21986;
															assign node21986 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node21990 = (inp[0]) ? node21994 : node21991;
															assign node21991 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node21994 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node21997 = (inp[11]) ? node22005 : node21998;
														assign node21998 = (inp[7]) ? node22002 : node21999;
															assign node21999 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node22002 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node22005 = (inp[7]) ? node22009 : node22006;
															assign node22006 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node22009 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node22012 = (inp[15]) ? node22040 : node22013;
												assign node22013 = (inp[12]) ? node22021 : node22014;
													assign node22014 = (inp[11]) ? node22018 : node22015;
														assign node22015 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node22018 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node22021 = (inp[7]) ? node22035 : node22022;
														assign node22022 = (inp[9]) ? node22028 : node22023;
															assign node22023 = (inp[11]) ? node22025 : 4'b0011;
																assign node22025 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node22028 = (inp[11]) ? node22032 : node22029;
																assign node22029 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node22032 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node22035 = (inp[0]) ? 4'b0110 : node22036;
															assign node22036 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node22040 = (inp[12]) ? node22070 : node22041;
													assign node22041 = (inp[7]) ? node22057 : node22042;
														assign node22042 = (inp[9]) ? node22050 : node22043;
															assign node22043 = (inp[0]) ? node22047 : node22044;
																assign node22044 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node22047 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node22050 = (inp[0]) ? node22054 : node22051;
																assign node22051 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node22054 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node22057 = (inp[9]) ? node22063 : node22058;
															assign node22058 = (inp[11]) ? 4'b0100 : node22059;
																assign node22059 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node22063 = (inp[11]) ? node22067 : node22064;
																assign node22064 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node22067 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node22070 = (inp[11]) ? node22076 : node22071;
														assign node22071 = (inp[7]) ? 4'b0101 : node22072;
															assign node22072 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node22076 = (inp[9]) ? node22084 : node22077;
															assign node22077 = (inp[7]) ? node22081 : node22078;
																assign node22078 = (inp[0]) ? 4'b0101 : 4'b0100;
																assign node22081 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node22084 = (inp[0]) ? node22088 : node22085;
																assign node22085 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node22088 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node22091 = (inp[0]) ? node22143 : node22092;
											assign node22092 = (inp[11]) ? node22116 : node22093;
												assign node22093 = (inp[4]) ? node22105 : node22094;
													assign node22094 = (inp[7]) ? node22102 : node22095;
														assign node22095 = (inp[15]) ? node22099 : node22096;
															assign node22096 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node22099 = (inp[12]) ? 4'b0111 : 4'b0110;
														assign node22102 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node22105 = (inp[15]) ? node22111 : node22106;
														assign node22106 = (inp[7]) ? 4'b0110 : node22107;
															assign node22107 = (inp[12]) ? 4'b0011 : 4'b0110;
														assign node22111 = (inp[7]) ? 4'b0100 : node22112;
															assign node22112 = (inp[12]) ? 4'b0101 : 4'b0000;
												assign node22116 = (inp[4]) ? node22130 : node22117;
													assign node22117 = (inp[15]) ? node22123 : node22118;
														assign node22118 = (inp[12]) ? node22120 : 4'b0100;
															assign node22120 = (inp[7]) ? 4'b0000 : 4'b0101;
														assign node22123 = (inp[7]) ? node22127 : node22124;
															assign node22124 = (inp[12]) ? 4'b0110 : 4'b0111;
															assign node22127 = (inp[12]) ? 4'b0111 : 4'b0010;
													assign node22130 = (inp[15]) ? node22136 : node22131;
														assign node22131 = (inp[12]) ? node22133 : 4'b0111;
															assign node22133 = (inp[7]) ? 4'b0111 : 4'b0010;
														assign node22136 = (inp[12]) ? node22140 : node22137;
															assign node22137 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node22140 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node22143 = (inp[11]) ? node22171 : node22144;
												assign node22144 = (inp[4]) ? node22158 : node22145;
													assign node22145 = (inp[15]) ? node22153 : node22146;
														assign node22146 = (inp[7]) ? node22150 : node22147;
															assign node22147 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node22150 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node22153 = (inp[12]) ? 4'b0111 : node22154;
															assign node22154 = (inp[7]) ? 4'b0010 : 4'b0111;
													assign node22158 = (inp[15]) ? node22164 : node22159;
														assign node22159 = (inp[7]) ? 4'b0111 : node22160;
															assign node22160 = (inp[12]) ? 4'b0010 : 4'b0111;
														assign node22164 = (inp[12]) ? node22168 : node22165;
															assign node22165 = (inp[7]) ? 4'b0101 : 4'b0001;
															assign node22168 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node22171 = (inp[4]) ? node22185 : node22172;
													assign node22172 = (inp[15]) ? node22178 : node22173;
														assign node22173 = (inp[12]) ? node22175 : 4'b0101;
															assign node22175 = (inp[7]) ? 4'b0001 : 4'b0100;
														assign node22178 = (inp[7]) ? node22182 : node22179;
															assign node22179 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node22182 = (inp[12]) ? 4'b0110 : 4'b0011;
													assign node22185 = (inp[15]) ? node22191 : node22186;
														assign node22186 = (inp[7]) ? 4'b0110 : node22187;
															assign node22187 = (inp[12]) ? 4'b0011 : 4'b0110;
														assign node22191 = (inp[7]) ? 4'b0100 : 4'b0101;
							assign node22194 = (inp[1]) ? node22650 : node22195;
								assign node22195 = (inp[10]) ? node22391 : node22196;
									assign node22196 = (inp[11]) ? node22282 : node22197;
										assign node22197 = (inp[0]) ? node22243 : node22198;
											assign node22198 = (inp[7]) ? node22216 : node22199;
												assign node22199 = (inp[4]) ? node22207 : node22200;
													assign node22200 = (inp[15]) ? node22204 : node22201;
														assign node22201 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node22204 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node22207 = (inp[15]) ? node22213 : node22208;
														assign node22208 = (inp[12]) ? 4'b0011 : node22209;
															assign node22209 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node22213 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node22216 = (inp[12]) ? node22228 : node22217;
													assign node22217 = (inp[15]) ? node22225 : node22218;
														assign node22218 = (inp[4]) ? node22222 : node22219;
															assign node22219 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node22222 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node22225 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node22228 = (inp[2]) ? node22236 : node22229;
														assign node22229 = (inp[15]) ? node22233 : node22230;
															assign node22230 = (inp[4]) ? 4'b0111 : 4'b0000;
															assign node22233 = (inp[4]) ? 4'b0100 : 4'b0111;
														assign node22236 = (inp[4]) ? node22240 : node22237;
															assign node22237 = (inp[15]) ? 4'b0110 : 4'b0001;
															assign node22240 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node22243 = (inp[7]) ? node22261 : node22244;
												assign node22244 = (inp[4]) ? node22252 : node22245;
													assign node22245 = (inp[15]) ? node22249 : node22246;
														assign node22246 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node22249 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node22252 = (inp[15]) ? node22258 : node22253;
														assign node22253 = (inp[12]) ? 4'b0010 : node22254;
															assign node22254 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node22258 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node22261 = (inp[4]) ? node22273 : node22262;
													assign node22262 = (inp[15]) ? node22270 : node22263;
														assign node22263 = (inp[12]) ? node22267 : node22264;
															assign node22264 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node22267 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node22270 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node22273 = (inp[15]) ? node22279 : node22274;
														assign node22274 = (inp[9]) ? 4'b0110 : node22275;
															assign node22275 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node22279 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node22282 = (inp[4]) ? node22330 : node22283;
											assign node22283 = (inp[15]) ? node22313 : node22284;
												assign node22284 = (inp[7]) ? node22300 : node22285;
													assign node22285 = (inp[12]) ? node22293 : node22286;
														assign node22286 = (inp[2]) ? node22290 : node22287;
															assign node22287 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node22290 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node22293 = (inp[0]) ? node22297 : node22294;
															assign node22294 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node22297 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node22300 = (inp[12]) ? node22306 : node22301;
														assign node22301 = (inp[0]) ? 4'b0100 : node22302;
															assign node22302 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node22306 = (inp[0]) ? node22310 : node22307;
															assign node22307 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node22310 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node22313 = (inp[12]) ? node22323 : node22314;
													assign node22314 = (inp[7]) ? node22320 : node22315;
														assign node22315 = (inp[0]) ? node22317 : 4'b0110;
															assign node22317 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node22320 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node22323 = (inp[2]) ? node22327 : node22324;
														assign node22324 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node22327 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node22330 = (inp[15]) ? node22368 : node22331;
												assign node22331 = (inp[12]) ? node22357 : node22332;
													assign node22332 = (inp[0]) ? node22348 : node22333;
														assign node22333 = (inp[9]) ? node22341 : node22334;
															assign node22334 = (inp[2]) ? node22338 : node22335;
																assign node22335 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node22338 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node22341 = (inp[7]) ? node22345 : node22342;
																assign node22342 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node22345 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node22348 = (inp[9]) ? 4'b0111 : node22349;
															assign node22349 = (inp[7]) ? node22353 : node22350;
																assign node22350 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node22353 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node22357 = (inp[7]) ? node22359 : 4'b0011;
														assign node22359 = (inp[9]) ? 4'b0111 : node22360;
															assign node22360 = (inp[2]) ? node22364 : node22361;
																assign node22361 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node22364 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node22368 = (inp[7]) ? node22376 : node22369;
													assign node22369 = (inp[12]) ? node22373 : node22370;
														assign node22370 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node22373 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node22376 = (inp[2]) ? node22384 : node22377;
														assign node22377 = (inp[0]) ? node22381 : node22378;
															assign node22378 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node22381 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node22384 = (inp[0]) ? node22388 : node22385;
															assign node22385 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node22388 = (inp[12]) ? 4'b0100 : 4'b0101;
									assign node22391 = (inp[0]) ? node22557 : node22392;
										assign node22392 = (inp[9]) ? node22470 : node22393;
											assign node22393 = (inp[4]) ? node22443 : node22394;
												assign node22394 = (inp[15]) ? node22420 : node22395;
													assign node22395 = (inp[12]) ? node22411 : node22396;
														assign node22396 = (inp[7]) ? node22404 : node22397;
															assign node22397 = (inp[2]) ? node22401 : node22398;
																assign node22398 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node22401 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node22404 = (inp[11]) ? node22408 : node22405;
																assign node22405 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node22408 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node22411 = (inp[7]) ? node22413 : 4'b0100;
															assign node22413 = (inp[2]) ? node22417 : node22414;
																assign node22414 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node22417 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node22420 = (inp[7]) ? node22434 : node22421;
														assign node22421 = (inp[12]) ? node22429 : node22422;
															assign node22422 = (inp[11]) ? node22426 : node22423;
																assign node22423 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node22426 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node22429 = (inp[2]) ? 4'b0111 : node22430;
																assign node22430 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node22434 = (inp[12]) ? node22438 : node22435;
															assign node22435 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node22438 = (inp[2]) ? 4'b0111 : node22439;
																assign node22439 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node22443 = (inp[15]) ? node22459 : node22444;
													assign node22444 = (inp[7]) ? node22450 : node22445;
														assign node22445 = (inp[12]) ? node22447 : 4'b0111;
															assign node22447 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node22450 = (inp[11]) ? 4'b0111 : node22451;
															assign node22451 = (inp[12]) ? node22455 : node22452;
																assign node22452 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node22455 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node22459 = (inp[11]) ? node22465 : node22460;
														assign node22460 = (inp[12]) ? 4'b0100 : node22461;
															assign node22461 = (inp[7]) ? 4'b0101 : 4'b0000;
														assign node22465 = (inp[12]) ? 4'b0101 : node22466;
															assign node22466 = (inp[7]) ? 4'b0100 : 4'b0001;
											assign node22470 = (inp[2]) ? node22510 : node22471;
												assign node22471 = (inp[11]) ? node22489 : node22472;
													assign node22472 = (inp[15]) ? node22482 : node22473;
														assign node22473 = (inp[4]) ? node22479 : node22474;
															assign node22474 = (inp[12]) ? node22476 : 4'b0101;
																assign node22476 = (inp[7]) ? 4'b0000 : 4'b0100;
															assign node22479 = (inp[7]) ? 4'b0110 : 4'b0011;
														assign node22482 = (inp[4]) ? 4'b0000 : node22483;
															assign node22483 = (inp[12]) ? 4'b0111 : node22484;
																assign node22484 = (inp[7]) ? 4'b0011 : 4'b0111;
													assign node22489 = (inp[15]) ? node22499 : node22490;
														assign node22490 = (inp[4]) ? node22494 : node22491;
															assign node22491 = (inp[7]) ? 4'b0001 : 4'b0101;
															assign node22494 = (inp[7]) ? node22496 : 4'b0110;
																assign node22496 = (inp[12]) ? 4'b0110 : 4'b0111;
														assign node22499 = (inp[4]) ? node22505 : node22500;
															assign node22500 = (inp[12]) ? 4'b0110 : node22501;
																assign node22501 = (inp[7]) ? 4'b0010 : 4'b0110;
															assign node22505 = (inp[7]) ? node22507 : 4'b0001;
																assign node22507 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node22510 = (inp[7]) ? node22530 : node22511;
													assign node22511 = (inp[4]) ? node22519 : node22512;
														assign node22512 = (inp[15]) ? node22516 : node22513;
															assign node22513 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node22516 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node22519 = (inp[15]) ? node22525 : node22520;
															assign node22520 = (inp[12]) ? node22522 : 4'b0110;
																assign node22522 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node22525 = (inp[11]) ? 4'b0001 : node22526;
																assign node22526 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node22530 = (inp[4]) ? node22542 : node22531;
														assign node22531 = (inp[15]) ? node22539 : node22532;
															assign node22532 = (inp[12]) ? node22536 : node22533;
																assign node22533 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node22536 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node22539 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node22542 = (inp[15]) ? node22550 : node22543;
															assign node22543 = (inp[11]) ? node22547 : node22544;
																assign node22544 = (inp[12]) ? 4'b0110 : 4'b0111;
																assign node22547 = (inp[12]) ? 4'b0111 : 4'b0110;
															assign node22550 = (inp[11]) ? node22554 : node22551;
																assign node22551 = (inp[12]) ? 4'b0100 : 4'b0101;
																assign node22554 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node22557 = (inp[11]) ? node22605 : node22558;
											assign node22558 = (inp[12]) ? node22586 : node22559;
												assign node22559 = (inp[15]) ? node22577 : node22560;
													assign node22560 = (inp[4]) ? node22568 : node22561;
														assign node22561 = (inp[7]) ? node22565 : node22562;
															assign node22562 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node22565 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node22568 = (inp[9]) ? 4'b0111 : node22569;
															assign node22569 = (inp[2]) ? node22573 : node22570;
																assign node22570 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node22573 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node22577 = (inp[4]) ? node22583 : node22578;
														assign node22578 = (inp[7]) ? 4'b0010 : node22579;
															assign node22579 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node22583 = (inp[7]) ? 4'b0100 : 4'b0001;
												assign node22586 = (inp[15]) ? node22600 : node22587;
													assign node22587 = (inp[4]) ? node22595 : node22588;
														assign node22588 = (inp[7]) ? node22592 : node22589;
															assign node22589 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node22592 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node22595 = (inp[7]) ? node22597 : 4'b0010;
															assign node22597 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node22600 = (inp[4]) ? 4'b0101 : node22601;
														assign node22601 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node22605 = (inp[2]) ? node22627 : node22606;
												assign node22606 = (inp[4]) ? node22616 : node22607;
													assign node22607 = (inp[15]) ? 4'b0111 : node22608;
														assign node22608 = (inp[12]) ? node22612 : node22609;
															assign node22609 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node22612 = (inp[7]) ? 4'b0000 : 4'b0100;
													assign node22616 = (inp[15]) ? node22624 : node22617;
														assign node22617 = (inp[12]) ? node22621 : node22618;
															assign node22618 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node22621 = (inp[7]) ? 4'b0111 : 4'b0011;
														assign node22624 = (inp[7]) ? 4'b0101 : 4'b0000;
												assign node22627 = (inp[15]) ? node22639 : node22628;
													assign node22628 = (inp[4]) ? node22632 : node22629;
														assign node22629 = (inp[7]) ? 4'b0001 : 4'b0101;
														assign node22632 = (inp[7]) ? node22636 : node22633;
															assign node22633 = (inp[12]) ? 4'b0011 : 4'b0110;
															assign node22636 = (inp[12]) ? 4'b0110 : 4'b0111;
													assign node22639 = (inp[4]) ? node22645 : node22640;
														assign node22640 = (inp[7]) ? node22642 : 4'b0110;
															assign node22642 = (inp[12]) ? 4'b0110 : 4'b0011;
														assign node22645 = (inp[12]) ? 4'b0100 : node22646;
															assign node22646 = (inp[7]) ? 4'b0101 : 4'b0000;
								assign node22650 = (inp[4]) ? node22914 : node22651;
									assign node22651 = (inp[15]) ? node22779 : node22652;
										assign node22652 = (inp[12]) ? node22726 : node22653;
											assign node22653 = (inp[2]) ? node22695 : node22654;
												assign node22654 = (inp[9]) ? node22674 : node22655;
													assign node22655 = (inp[10]) ? node22665 : node22656;
														assign node22656 = (inp[11]) ? 4'b0001 : node22657;
															assign node22657 = (inp[0]) ? node22661 : node22658;
																assign node22658 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node22661 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node22665 = (inp[0]) ? 4'b0000 : node22666;
															assign node22666 = (inp[7]) ? node22670 : node22667;
																assign node22667 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node22670 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node22674 = (inp[11]) ? node22682 : node22675;
														assign node22675 = (inp[0]) ? node22679 : node22676;
															assign node22676 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node22679 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node22682 = (inp[10]) ? node22690 : node22683;
															assign node22683 = (inp[7]) ? node22687 : node22684;
																assign node22684 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node22687 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node22690 = (inp[7]) ? 4'b0001 : node22691;
																assign node22691 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node22695 = (inp[0]) ? node22711 : node22696;
													assign node22696 = (inp[10]) ? node22704 : node22697;
														assign node22697 = (inp[9]) ? node22699 : 4'b0000;
															assign node22699 = (inp[11]) ? 4'b0000 : node22700;
																assign node22700 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node22704 = (inp[11]) ? node22708 : node22705;
															assign node22705 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node22708 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node22711 = (inp[10]) ? node22717 : node22712;
														assign node22712 = (inp[11]) ? node22714 : 4'b0001;
															assign node22714 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node22717 = (inp[9]) ? node22721 : node22718;
															assign node22718 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node22721 = (inp[11]) ? 4'b0000 : node22722;
																assign node22722 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node22726 = (inp[7]) ? node22740 : node22727;
												assign node22727 = (inp[2]) ? node22733 : node22728;
													assign node22728 = (inp[11]) ? 4'b0001 : node22729;
														assign node22729 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node22733 = (inp[0]) ? node22737 : node22734;
														assign node22734 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node22737 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node22740 = (inp[10]) ? node22766 : node22741;
													assign node22741 = (inp[9]) ? node22757 : node22742;
														assign node22742 = (inp[11]) ? node22750 : node22743;
															assign node22743 = (inp[0]) ? node22747 : node22744;
																assign node22744 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node22747 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node22750 = (inp[0]) ? node22754 : node22751;
																assign node22751 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node22754 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node22757 = (inp[2]) ? 4'b0100 : node22758;
															assign node22758 = (inp[11]) ? node22762 : node22759;
																assign node22759 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node22762 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node22766 = (inp[2]) ? node22774 : node22767;
														assign node22767 = (inp[0]) ? node22771 : node22768;
															assign node22768 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node22771 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node22774 = (inp[0]) ? node22776 : 4'b0101;
															assign node22776 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node22779 = (inp[12]) ? node22845 : node22780;
											assign node22780 = (inp[7]) ? node22818 : node22781;
												assign node22781 = (inp[9]) ? node22805 : node22782;
													assign node22782 = (inp[10]) ? node22796 : node22783;
														assign node22783 = (inp[11]) ? node22789 : node22784;
															assign node22784 = (inp[0]) ? node22786 : 4'b0010;
																assign node22786 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node22789 = (inp[0]) ? node22793 : node22790;
																assign node22790 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node22793 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node22796 = (inp[0]) ? node22798 : 4'b0011;
															assign node22798 = (inp[11]) ? node22802 : node22799;
																assign node22799 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node22802 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node22805 = (inp[11]) ? node22813 : node22806;
														assign node22806 = (inp[2]) ? node22810 : node22807;
															assign node22807 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node22810 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node22813 = (inp[0]) ? node22815 : 4'b0010;
															assign node22815 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node22818 = (inp[9]) ? node22832 : node22819;
													assign node22819 = (inp[0]) ? node22827 : node22820;
														assign node22820 = (inp[2]) ? node22824 : node22821;
															assign node22821 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node22824 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node22827 = (inp[2]) ? 4'b0110 : node22828;
															assign node22828 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node22832 = (inp[0]) ? node22840 : node22833;
														assign node22833 = (inp[2]) ? node22837 : node22834;
															assign node22834 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node22837 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node22840 = (inp[2]) ? 4'b0111 : node22841;
															assign node22841 = (inp[10]) ? 4'b0111 : 4'b0110;
											assign node22845 = (inp[10]) ? node22877 : node22846;
												assign node22846 = (inp[2]) ? node22864 : node22847;
													assign node22847 = (inp[7]) ? node22857 : node22848;
														assign node22848 = (inp[9]) ? node22850 : 4'b0010;
															assign node22850 = (inp[0]) ? node22854 : node22851;
																assign node22851 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node22854 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node22857 = (inp[0]) ? node22861 : node22858;
															assign node22858 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node22861 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node22864 = (inp[9]) ? node22870 : node22865;
														assign node22865 = (inp[7]) ? node22867 : 4'b0011;
															assign node22867 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node22870 = (inp[0]) ? node22874 : node22871;
															assign node22871 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node22874 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node22877 = (inp[2]) ? node22895 : node22878;
													assign node22878 = (inp[7]) ? node22888 : node22879;
														assign node22879 = (inp[9]) ? node22885 : node22880;
															assign node22880 = (inp[0]) ? node22882 : 4'b0011;
																assign node22882 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node22885 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node22888 = (inp[0]) ? node22892 : node22889;
															assign node22889 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node22892 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node22895 = (inp[7]) ? node22901 : node22896;
														assign node22896 = (inp[0]) ? node22898 : 4'b0010;
															assign node22898 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node22901 = (inp[9]) ? node22907 : node22902;
															assign node22902 = (inp[11]) ? node22904 : 4'b0010;
																assign node22904 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node22907 = (inp[0]) ? node22911 : node22908;
																assign node22908 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node22911 = (inp[11]) ? 4'b0010 : 4'b0011;
									assign node22914 = (inp[15]) ? node22986 : node22915;
										assign node22915 = (inp[7]) ? node22963 : node22916;
											assign node22916 = (inp[12]) ? node22948 : node22917;
												assign node22917 = (inp[10]) ? node22943 : node22918;
													assign node22918 = (inp[9]) ? node22928 : node22919;
														assign node22919 = (inp[2]) ? node22923 : node22920;
															assign node22920 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node22923 = (inp[0]) ? 4'b0010 : node22924;
																assign node22924 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node22928 = (inp[2]) ? node22936 : node22929;
															assign node22929 = (inp[0]) ? node22933 : node22930;
																assign node22930 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node22933 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node22936 = (inp[11]) ? node22940 : node22937;
																assign node22937 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node22940 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node22943 = (inp[2]) ? 4'b0011 : node22944;
														assign node22944 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node22948 = (inp[2]) ? node22956 : node22949;
													assign node22949 = (inp[0]) ? node22953 : node22950;
														assign node22950 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node22953 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node22956 = (inp[0]) ? node22960 : node22957;
														assign node22957 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node22960 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node22963 = (inp[10]) ? node22979 : node22964;
												assign node22964 = (inp[2]) ? node22972 : node22965;
													assign node22965 = (inp[0]) ? node22969 : node22966;
														assign node22966 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node22969 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node22972 = (inp[11]) ? node22976 : node22973;
														assign node22973 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node22976 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node22979 = (inp[0]) ? node22983 : node22980;
													assign node22980 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node22983 = (inp[11]) ? 4'b0010 : 4'b0011;
										assign node22986 = (inp[7]) ? node23050 : node22987;
											assign node22987 = (inp[12]) ? node23021 : node22988;
												assign node22988 = (inp[11]) ? node23006 : node22989;
													assign node22989 = (inp[9]) ? node22997 : node22990;
														assign node22990 = (inp[2]) ? node22994 : node22991;
															assign node22991 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node22994 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node22997 = (inp[10]) ? 4'b0100 : node22998;
															assign node22998 = (inp[2]) ? node23002 : node22999;
																assign node22999 = (inp[0]) ? 4'b0100 : 4'b0101;
																assign node23002 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node23006 = (inp[9]) ? node23014 : node23007;
														assign node23007 = (inp[0]) ? node23011 : node23008;
															assign node23008 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node23011 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node23014 = (inp[0]) ? node23018 : node23015;
															assign node23015 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node23018 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node23021 = (inp[10]) ? node23035 : node23022;
													assign node23022 = (inp[2]) ? node23028 : node23023;
														assign node23023 = (inp[0]) ? 4'b0000 : node23024;
															assign node23024 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node23028 = (inp[0]) ? node23032 : node23029;
															assign node23029 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node23032 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node23035 = (inp[2]) ? node23043 : node23036;
														assign node23036 = (inp[11]) ? node23040 : node23037;
															assign node23037 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node23040 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node23043 = (inp[11]) ? node23047 : node23044;
															assign node23044 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node23047 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node23050 = (inp[12]) ? node23086 : node23051;
												assign node23051 = (inp[9]) ? node23061 : node23052;
													assign node23052 = (inp[2]) ? node23054 : 4'b0001;
														assign node23054 = (inp[0]) ? node23058 : node23055;
															assign node23055 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node23058 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node23061 = (inp[2]) ? node23075 : node23062;
														assign node23062 = (inp[10]) ? node23068 : node23063;
															assign node23063 = (inp[0]) ? 4'b0000 : node23064;
																assign node23064 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node23068 = (inp[0]) ? node23072 : node23069;
																assign node23069 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node23072 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node23075 = (inp[10]) ? node23081 : node23076;
															assign node23076 = (inp[11]) ? node23078 : 4'b0001;
																assign node23078 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node23081 = (inp[0]) ? 4'b0001 : node23082;
																assign node23082 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node23086 = (inp[9]) ? node23094 : node23087;
													assign node23087 = (inp[11]) ? node23091 : node23088;
														assign node23088 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node23091 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node23094 = (inp[11]) ? node23096 : 4'b0000;
														assign node23096 = (inp[0]) ? 4'b0000 : 4'b0001;
				assign node23099 = (inp[4]) ? node25347 : node23100;
					assign node23100 = (inp[7]) ? node24236 : node23101;
						assign node23101 = (inp[8]) ? node23829 : node23102;
							assign node23102 = (inp[15]) ? node23408 : node23103;
								assign node23103 = (inp[12]) ? node23217 : node23104;
									assign node23104 = (inp[13]) ? node23128 : node23105;
										assign node23105 = (inp[9]) ? node23117 : node23106;
											assign node23106 = (inp[2]) ? node23112 : node23107;
												assign node23107 = (inp[0]) ? node23109 : 4'b0000;
													assign node23109 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node23112 = (inp[0]) ? node23114 : 4'b0001;
													assign node23114 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node23117 = (inp[2]) ? node23123 : node23118;
												assign node23118 = (inp[0]) ? node23120 : 4'b0001;
													assign node23120 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node23123 = (inp[0]) ? node23125 : 4'b0000;
													assign node23125 = (inp[5]) ? 4'b0001 : 4'b0000;
										assign node23128 = (inp[10]) ? node23176 : node23129;
											assign node23129 = (inp[11]) ? node23157 : node23130;
												assign node23130 = (inp[0]) ? node23136 : node23131;
													assign node23131 = (inp[9]) ? 4'b0100 : node23132;
														assign node23132 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node23136 = (inp[5]) ? node23152 : node23137;
														assign node23137 = (inp[1]) ? node23145 : node23138;
															assign node23138 = (inp[2]) ? node23142 : node23139;
																assign node23139 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node23142 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node23145 = (inp[9]) ? node23149 : node23146;
																assign node23146 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node23149 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node23152 = (inp[9]) ? node23154 : 4'b0100;
															assign node23154 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node23157 = (inp[9]) ? node23167 : node23158;
													assign node23158 = (inp[2]) ? node23164 : node23159;
														assign node23159 = (inp[0]) ? node23161 : 4'b0100;
															assign node23161 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node23164 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node23167 = (inp[2]) ? node23171 : node23168;
														assign node23168 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node23171 = (inp[0]) ? node23173 : 4'b0100;
															assign node23173 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node23176 = (inp[0]) ? node23192 : node23177;
												assign node23177 = (inp[1]) ? node23185 : node23178;
													assign node23178 = (inp[9]) ? node23182 : node23179;
														assign node23179 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node23182 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node23185 = (inp[2]) ? node23189 : node23186;
														assign node23186 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node23189 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node23192 = (inp[11]) ? node23208 : node23193;
													assign node23193 = (inp[5]) ? node23201 : node23194;
														assign node23194 = (inp[9]) ? node23198 : node23195;
															assign node23195 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node23198 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node23201 = (inp[2]) ? node23205 : node23202;
															assign node23202 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node23205 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node23208 = (inp[5]) ? node23210 : 4'b0100;
														assign node23210 = (inp[9]) ? node23214 : node23211;
															assign node23211 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node23214 = (inp[2]) ? 4'b0101 : 4'b0100;
									assign node23217 = (inp[13]) ? node23327 : node23218;
										assign node23218 = (inp[5]) ? node23262 : node23219;
											assign node23219 = (inp[9]) ? node23241 : node23220;
												assign node23220 = (inp[0]) ? node23228 : node23221;
													assign node23221 = (inp[2]) ? node23225 : node23222;
														assign node23222 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node23225 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node23228 = (inp[10]) ? node23234 : node23229;
														assign node23229 = (inp[1]) ? node23231 : 4'b0100;
															assign node23231 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node23234 = (inp[1]) ? node23238 : node23235;
															assign node23235 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node23238 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node23241 = (inp[0]) ? node23249 : node23242;
													assign node23242 = (inp[1]) ? node23246 : node23243;
														assign node23243 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node23246 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node23249 = (inp[10]) ? node23255 : node23250;
														assign node23250 = (inp[11]) ? 4'b0100 : node23251;
															assign node23251 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node23255 = (inp[2]) ? node23259 : node23256;
															assign node23256 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node23259 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node23262 = (inp[2]) ? node23296 : node23263;
												assign node23263 = (inp[0]) ? node23277 : node23264;
													assign node23264 = (inp[10]) ? node23272 : node23265;
														assign node23265 = (inp[1]) ? node23269 : node23266;
															assign node23266 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node23269 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node23272 = (inp[1]) ? node23274 : 4'b0100;
															assign node23274 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node23277 = (inp[11]) ? node23283 : node23278;
														assign node23278 = (inp[1]) ? node23280 : 4'b0101;
															assign node23280 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node23283 = (inp[10]) ? node23289 : node23284;
															assign node23284 = (inp[9]) ? node23286 : 4'b0101;
																assign node23286 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node23289 = (inp[9]) ? node23293 : node23290;
																assign node23290 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node23293 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node23296 = (inp[0]) ? node23310 : node23297;
													assign node23297 = (inp[11]) ? node23305 : node23298;
														assign node23298 = (inp[9]) ? node23302 : node23299;
															assign node23299 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node23302 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node23305 = (inp[9]) ? 4'b0101 : node23306;
															assign node23306 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node23310 = (inp[11]) ? node23318 : node23311;
														assign node23311 = (inp[9]) ? node23315 : node23312;
															assign node23312 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node23315 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node23318 = (inp[10]) ? node23320 : 4'b0100;
															assign node23320 = (inp[9]) ? node23324 : node23321;
																assign node23321 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node23324 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node23327 = (inp[2]) ? node23385 : node23328;
											assign node23328 = (inp[5]) ? node23358 : node23329;
												assign node23329 = (inp[9]) ? node23345 : node23330;
													assign node23330 = (inp[11]) ? node23338 : node23331;
														assign node23331 = (inp[0]) ? node23335 : node23332;
															assign node23332 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node23335 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node23338 = (inp[0]) ? node23342 : node23339;
															assign node23339 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node23342 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node23345 = (inp[10]) ? node23351 : node23346;
														assign node23346 = (inp[1]) ? node23348 : 4'b0001;
															assign node23348 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node23351 = (inp[11]) ? 4'b0001 : node23352;
															assign node23352 = (inp[1]) ? 4'b0001 : node23353;
																assign node23353 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node23358 = (inp[10]) ? node23374 : node23359;
													assign node23359 = (inp[0]) ? node23367 : node23360;
														assign node23360 = (inp[9]) ? node23364 : node23361;
															assign node23361 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node23364 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node23367 = (inp[9]) ? node23371 : node23368;
															assign node23368 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node23371 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node23374 = (inp[0]) ? node23380 : node23375;
														assign node23375 = (inp[1]) ? node23377 : 4'b0000;
															assign node23377 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node23380 = (inp[1]) ? 4'b0000 : node23381;
															assign node23381 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node23385 = (inp[1]) ? node23397 : node23386;
												assign node23386 = (inp[9]) ? node23392 : node23387;
													assign node23387 = (inp[0]) ? 4'b0000 : node23388;
														assign node23388 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node23392 = (inp[5]) ? 4'b0001 : node23393;
														assign node23393 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node23397 = (inp[9]) ? node23403 : node23398;
													assign node23398 = (inp[0]) ? 4'b0001 : node23399;
														assign node23399 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node23403 = (inp[5]) ? 4'b0000 : node23404;
														assign node23404 = (inp[0]) ? 4'b0000 : 4'b0001;
								assign node23408 = (inp[1]) ? node23642 : node23409;
									assign node23409 = (inp[5]) ? node23515 : node23410;
										assign node23410 = (inp[0]) ? node23484 : node23411;
											assign node23411 = (inp[13]) ? node23445 : node23412;
												assign node23412 = (inp[12]) ? node23432 : node23413;
													assign node23413 = (inp[10]) ? node23427 : node23414;
														assign node23414 = (inp[11]) ? node23420 : node23415;
															assign node23415 = (inp[2]) ? node23417 : 4'b0001;
																assign node23417 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node23420 = (inp[9]) ? node23424 : node23421;
																assign node23421 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node23424 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node23427 = (inp[2]) ? 4'b0000 : node23428;
															assign node23428 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node23432 = (inp[11]) ? node23438 : node23433;
														assign node23433 = (inp[2]) ? node23435 : 4'b0100;
															assign node23435 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node23438 = (inp[9]) ? node23442 : node23439;
															assign node23439 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node23442 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node23445 = (inp[12]) ? node23467 : node23446;
													assign node23446 = (inp[10]) ? node23454 : node23447;
														assign node23447 = (inp[2]) ? node23451 : node23448;
															assign node23448 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node23451 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node23454 = (inp[11]) ? node23460 : node23455;
															assign node23455 = (inp[2]) ? node23457 : 4'b0100;
																assign node23457 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node23460 = (inp[9]) ? node23464 : node23461;
																assign node23461 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node23464 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node23467 = (inp[11]) ? node23479 : node23468;
														assign node23468 = (inp[10]) ? node23474 : node23469;
															assign node23469 = (inp[9]) ? node23471 : 4'b0001;
																assign node23471 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node23474 = (inp[2]) ? node23476 : 4'b0001;
																assign node23476 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node23479 = (inp[2]) ? node23481 : 4'b0000;
															assign node23481 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node23484 = (inp[9]) ? node23500 : node23485;
												assign node23485 = (inp[2]) ? node23493 : node23486;
													assign node23486 = (inp[12]) ? node23490 : node23487;
														assign node23487 = (inp[13]) ? 4'b0101 : 4'b0000;
														assign node23490 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node23493 = (inp[13]) ? node23497 : node23494;
														assign node23494 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node23497 = (inp[12]) ? 4'b0001 : 4'b0100;
												assign node23500 = (inp[2]) ? node23508 : node23501;
													assign node23501 = (inp[13]) ? node23505 : node23502;
														assign node23502 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node23505 = (inp[12]) ? 4'b0001 : 4'b0100;
													assign node23508 = (inp[13]) ? node23512 : node23509;
														assign node23509 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node23512 = (inp[12]) ? 4'b0000 : 4'b0101;
										assign node23515 = (inp[12]) ? node23595 : node23516;
											assign node23516 = (inp[13]) ? node23552 : node23517;
												assign node23517 = (inp[0]) ? node23545 : node23518;
													assign node23518 = (inp[10]) ? node23530 : node23519;
														assign node23519 = (inp[11]) ? node23525 : node23520;
															assign node23520 = (inp[2]) ? node23522 : 4'b0001;
																assign node23522 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node23525 = (inp[9]) ? 4'b0001 : node23526;
																assign node23526 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node23530 = (inp[11]) ? node23538 : node23531;
															assign node23531 = (inp[2]) ? node23535 : node23532;
																assign node23532 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node23535 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node23538 = (inp[9]) ? node23542 : node23539;
																assign node23539 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node23542 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node23545 = (inp[9]) ? node23549 : node23546;
														assign node23546 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node23549 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node23552 = (inp[10]) ? node23570 : node23553;
													assign node23553 = (inp[2]) ? node23563 : node23554;
														assign node23554 = (inp[11]) ? node23556 : 4'b0100;
															assign node23556 = (inp[0]) ? node23560 : node23557;
																assign node23557 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node23560 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node23563 = (inp[9]) ? node23567 : node23564;
															assign node23564 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node23567 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node23570 = (inp[0]) ? node23580 : node23571;
														assign node23571 = (inp[11]) ? node23577 : node23572;
															assign node23572 = (inp[9]) ? node23574 : 4'b0100;
																assign node23574 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node23577 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node23580 = (inp[11]) ? node23588 : node23581;
															assign node23581 = (inp[2]) ? node23585 : node23582;
																assign node23582 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node23585 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node23588 = (inp[2]) ? node23592 : node23589;
																assign node23589 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node23592 = (inp[9]) ? 4'b0100 : 4'b0101;
											assign node23595 = (inp[13]) ? node23635 : node23596;
												assign node23596 = (inp[0]) ? node23620 : node23597;
													assign node23597 = (inp[10]) ? node23611 : node23598;
														assign node23598 = (inp[11]) ? node23606 : node23599;
															assign node23599 = (inp[9]) ? node23603 : node23600;
																assign node23600 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node23603 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node23606 = (inp[9]) ? 4'b0101 : node23607;
																assign node23607 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node23611 = (inp[11]) ? node23613 : 4'b0101;
															assign node23613 = (inp[2]) ? node23617 : node23614;
																assign node23614 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node23617 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node23620 = (inp[10]) ? node23628 : node23621;
														assign node23621 = (inp[9]) ? node23625 : node23622;
															assign node23622 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node23625 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node23628 = (inp[2]) ? node23632 : node23629;
															assign node23629 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node23632 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node23635 = (inp[2]) ? node23639 : node23636;
													assign node23636 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node23639 = (inp[9]) ? 4'b0000 : 4'b0001;
									assign node23642 = (inp[0]) ? node23716 : node23643;
										assign node23643 = (inp[12]) ? node23693 : node23644;
											assign node23644 = (inp[13]) ? node23680 : node23645;
												assign node23645 = (inp[9]) ? node23663 : node23646;
													assign node23646 = (inp[10]) ? node23658 : node23647;
														assign node23647 = (inp[11]) ? node23653 : node23648;
															assign node23648 = (inp[2]) ? node23650 : 4'b0100;
																assign node23650 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node23653 = (inp[5]) ? 4'b0101 : node23654;
																assign node23654 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node23658 = (inp[2]) ? node23660 : 4'b0101;
															assign node23660 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node23663 = (inp[11]) ? node23671 : node23664;
														assign node23664 = (inp[2]) ? node23668 : node23665;
															assign node23665 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node23668 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node23671 = (inp[10]) ? 4'b0100 : node23672;
															assign node23672 = (inp[2]) ? node23676 : node23673;
																assign node23673 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node23676 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node23680 = (inp[5]) ? node23686 : node23681;
													assign node23681 = (inp[9]) ? 4'b0001 : node23682;
														assign node23682 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node23686 = (inp[9]) ? node23690 : node23687;
														assign node23687 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node23690 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node23693 = (inp[13]) ? node23709 : node23694;
												assign node23694 = (inp[5]) ? node23702 : node23695;
													assign node23695 = (inp[2]) ? node23699 : node23696;
														assign node23696 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node23699 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node23702 = (inp[2]) ? node23706 : node23703;
														assign node23703 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node23706 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node23709 = (inp[2]) ? node23713 : node23710;
													assign node23710 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node23713 = (inp[9]) ? 4'b0101 : 4'b0100;
										assign node23716 = (inp[5]) ? node23798 : node23717;
											assign node23717 = (inp[11]) ? node23747 : node23718;
												assign node23718 = (inp[13]) ? node23730 : node23719;
													assign node23719 = (inp[12]) ? node23725 : node23720;
														assign node23720 = (inp[9]) ? node23722 : 4'b0100;
															assign node23722 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node23725 = (inp[2]) ? node23727 : 4'b0000;
															assign node23727 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node23730 = (inp[12]) ? node23742 : node23731;
														assign node23731 = (inp[10]) ? node23737 : node23732;
															assign node23732 = (inp[2]) ? node23734 : 4'b0001;
																assign node23734 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node23737 = (inp[9]) ? node23739 : 4'b0000;
																assign node23739 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node23742 = (inp[2]) ? node23744 : 4'b0100;
															assign node23744 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node23747 = (inp[10]) ? node23769 : node23748;
													assign node23748 = (inp[12]) ? node23758 : node23749;
														assign node23749 = (inp[13]) ? node23751 : 4'b0100;
															assign node23751 = (inp[9]) ? node23755 : node23752;
																assign node23752 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node23755 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node23758 = (inp[13]) ? node23764 : node23759;
															assign node23759 = (inp[9]) ? 4'b0000 : node23760;
																assign node23760 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node23764 = (inp[2]) ? 4'b0100 : node23765;
																assign node23765 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node23769 = (inp[12]) ? node23783 : node23770;
														assign node23770 = (inp[13]) ? node23776 : node23771;
															assign node23771 = (inp[9]) ? 4'b0101 : node23772;
																assign node23772 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node23776 = (inp[2]) ? node23780 : node23777;
																assign node23777 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node23780 = (inp[9]) ? 4'b0000 : 4'b0001;
														assign node23783 = (inp[13]) ? node23791 : node23784;
															assign node23784 = (inp[9]) ? node23788 : node23785;
																assign node23785 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node23788 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node23791 = (inp[2]) ? node23795 : node23792;
																assign node23792 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node23795 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node23798 = (inp[9]) ? node23814 : node23799;
												assign node23799 = (inp[2]) ? node23807 : node23800;
													assign node23800 = (inp[13]) ? node23804 : node23801;
														assign node23801 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node23804 = (inp[12]) ? 4'b0100 : 4'b0001;
													assign node23807 = (inp[12]) ? node23811 : node23808;
														assign node23808 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node23811 = (inp[13]) ? 4'b0101 : 4'b0000;
												assign node23814 = (inp[2]) ? node23822 : node23815;
													assign node23815 = (inp[13]) ? node23819 : node23816;
														assign node23816 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node23819 = (inp[12]) ? 4'b0101 : 4'b0000;
													assign node23822 = (inp[12]) ? node23826 : node23823;
														assign node23823 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node23826 = (inp[13]) ? 4'b0100 : 4'b0001;
							assign node23829 = (inp[10]) ? node24049 : node23830;
								assign node23830 = (inp[0]) ? node23940 : node23831;
									assign node23831 = (inp[2]) ? node23881 : node23832;
										assign node23832 = (inp[13]) ? node23848 : node23833;
											assign node23833 = (inp[1]) ? node23837 : node23834;
												assign node23834 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node23837 = (inp[12]) ? node23843 : node23838;
													assign node23838 = (inp[15]) ? node23840 : 4'b0110;
														assign node23840 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node23843 = (inp[15]) ? 4'b0010 : node23844;
														assign node23844 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node23848 = (inp[1]) ? node23870 : node23849;
												assign node23849 = (inp[12]) ? node23857 : node23850;
													assign node23850 = (inp[5]) ? node23854 : node23851;
														assign node23851 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node23854 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node23857 = (inp[11]) ? node23863 : node23858;
														assign node23858 = (inp[5]) ? 4'b0111 : node23859;
															assign node23859 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node23863 = (inp[5]) ? node23867 : node23864;
															assign node23864 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node23867 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node23870 = (inp[12]) ? node23876 : node23871;
													assign node23871 = (inp[15]) ? 4'b0110 : node23872;
														assign node23872 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node23876 = (inp[5]) ? 4'b0010 : node23877;
														assign node23877 = (inp[15]) ? 4'b0011 : 4'b0010;
										assign node23881 = (inp[13]) ? node23897 : node23882;
											assign node23882 = (inp[1]) ? node23886 : node23883;
												assign node23883 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node23886 = (inp[12]) ? node23892 : node23887;
													assign node23887 = (inp[5]) ? node23889 : 4'b0111;
														assign node23889 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node23892 = (inp[5]) ? 4'b0011 : node23893;
														assign node23893 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node23897 = (inp[1]) ? node23929 : node23898;
												assign node23898 = (inp[12]) ? node23922 : node23899;
													assign node23899 = (inp[9]) ? node23909 : node23900;
														assign node23900 = (inp[11]) ? node23902 : 4'b0011;
															assign node23902 = (inp[15]) ? node23906 : node23903;
																assign node23903 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node23906 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node23909 = (inp[11]) ? node23917 : node23910;
															assign node23910 = (inp[15]) ? node23914 : node23911;
																assign node23911 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node23914 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node23917 = (inp[5]) ? node23919 : 4'b0010;
																assign node23919 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node23922 = (inp[5]) ? node23926 : node23923;
														assign node23923 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node23926 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node23929 = (inp[12]) ? node23935 : node23930;
													assign node23930 = (inp[15]) ? 4'b0111 : node23931;
														assign node23931 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node23935 = (inp[5]) ? 4'b0011 : node23936;
														assign node23936 = (inp[15]) ? 4'b0010 : 4'b0011;
									assign node23940 = (inp[2]) ? node24002 : node23941;
										assign node23941 = (inp[13]) ? node23957 : node23942;
											assign node23942 = (inp[1]) ? node23946 : node23943;
												assign node23943 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node23946 = (inp[12]) ? node23952 : node23947;
													assign node23947 = (inp[5]) ? node23949 : 4'b0111;
														assign node23949 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node23952 = (inp[15]) ? 4'b0011 : node23953;
														assign node23953 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node23957 = (inp[1]) ? node23991 : node23958;
												assign node23958 = (inp[12]) ? node23974 : node23959;
													assign node23959 = (inp[11]) ? node23967 : node23960;
														assign node23960 = (inp[15]) ? node23964 : node23961;
															assign node23961 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node23964 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node23967 = (inp[15]) ? node23971 : node23968;
															assign node23968 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node23971 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node23974 = (inp[9]) ? node23980 : node23975;
														assign node23975 = (inp[5]) ? node23977 : 4'b0110;
															assign node23977 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node23980 = (inp[11]) ? node23986 : node23981;
															assign node23981 = (inp[5]) ? 4'b0111 : node23982;
																assign node23982 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node23986 = (inp[15]) ? 4'b0111 : node23987;
																assign node23987 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node23991 = (inp[12]) ? node23997 : node23992;
													assign node23992 = (inp[5]) ? node23994 : 4'b0111;
														assign node23994 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node23997 = (inp[15]) ? node23999 : 4'b0011;
														assign node23999 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node24002 = (inp[13]) ? node24016 : node24003;
											assign node24003 = (inp[1]) ? node24007 : node24004;
												assign node24004 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node24007 = (inp[12]) ? node24011 : node24008;
													assign node24008 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node24011 = (inp[15]) ? 4'b0010 : node24012;
														assign node24012 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node24016 = (inp[12]) ? node24036 : node24017;
												assign node24017 = (inp[1]) ? node24031 : node24018;
													assign node24018 = (inp[9]) ? node24026 : node24019;
														assign node24019 = (inp[15]) ? node24023 : node24020;
															assign node24020 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node24023 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node24026 = (inp[5]) ? 4'b0011 : node24027;
															assign node24027 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node24031 = (inp[15]) ? 4'b0110 : node24032;
														assign node24032 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node24036 = (inp[1]) ? node24044 : node24037;
													assign node24037 = (inp[5]) ? node24041 : node24038;
														assign node24038 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node24041 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node24044 = (inp[5]) ? 4'b0010 : node24045;
														assign node24045 = (inp[15]) ? 4'b0011 : 4'b0010;
								assign node24049 = (inp[2]) ? node24145 : node24050;
									assign node24050 = (inp[0]) ? node24104 : node24051;
										assign node24051 = (inp[13]) ? node24067 : node24052;
											assign node24052 = (inp[1]) ? node24056 : node24053;
												assign node24053 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node24056 = (inp[12]) ? node24062 : node24057;
													assign node24057 = (inp[15]) ? node24059 : 4'b0110;
														assign node24059 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node24062 = (inp[15]) ? 4'b0010 : node24063;
														assign node24063 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node24067 = (inp[1]) ? node24093 : node24068;
												assign node24068 = (inp[12]) ? node24076 : node24069;
													assign node24069 = (inp[15]) ? node24073 : node24070;
														assign node24070 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node24073 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node24076 = (inp[9]) ? node24084 : node24077;
														assign node24077 = (inp[5]) ? node24081 : node24078;
															assign node24078 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node24081 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node24084 = (inp[11]) ? 4'b0110 : node24085;
															assign node24085 = (inp[15]) ? node24089 : node24086;
																assign node24086 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node24089 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node24093 = (inp[12]) ? node24099 : node24094;
													assign node24094 = (inp[5]) ? node24096 : 4'b0110;
														assign node24096 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node24099 = (inp[5]) ? 4'b0010 : node24100;
														assign node24100 = (inp[15]) ? 4'b0011 : 4'b0010;
										assign node24104 = (inp[13]) ? node24120 : node24105;
											assign node24105 = (inp[1]) ? node24109 : node24106;
												assign node24106 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node24109 = (inp[12]) ? node24115 : node24110;
													assign node24110 = (inp[5]) ? node24112 : 4'b0111;
														assign node24112 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node24115 = (inp[15]) ? 4'b0011 : node24116;
														assign node24116 = (inp[5]) ? 4'b0011 : 4'b0010;
											assign node24120 = (inp[1]) ? node24136 : node24121;
												assign node24121 = (inp[12]) ? node24129 : node24122;
													assign node24122 = (inp[5]) ? node24126 : node24123;
														assign node24123 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node24126 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node24129 = (inp[5]) ? node24133 : node24130;
														assign node24130 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node24133 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node24136 = (inp[12]) ? node24140 : node24137;
													assign node24137 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node24140 = (inp[5]) ? 4'b0011 : node24141;
														assign node24141 = (inp[15]) ? 4'b0010 : 4'b0011;
									assign node24145 = (inp[0]) ? node24187 : node24146;
										assign node24146 = (inp[13]) ? node24162 : node24147;
											assign node24147 = (inp[1]) ? node24151 : node24148;
												assign node24148 = (inp[12]) ? 4'b0111 : 4'b0011;
												assign node24151 = (inp[12]) ? node24157 : node24152;
													assign node24152 = (inp[15]) ? node24154 : 4'b0111;
														assign node24154 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node24157 = (inp[5]) ? 4'b0011 : node24158;
														assign node24158 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node24162 = (inp[1]) ? node24176 : node24163;
												assign node24163 = (inp[12]) ? node24171 : node24164;
													assign node24164 = (inp[5]) ? node24168 : node24165;
														assign node24165 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node24168 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node24171 = (inp[5]) ? node24173 : 4'b0110;
														assign node24173 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node24176 = (inp[12]) ? node24182 : node24177;
													assign node24177 = (inp[5]) ? node24179 : 4'b0111;
														assign node24179 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node24182 = (inp[15]) ? node24184 : 4'b0011;
														assign node24184 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node24187 = (inp[13]) ? node24203 : node24188;
											assign node24188 = (inp[1]) ? node24192 : node24189;
												assign node24189 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node24192 = (inp[12]) ? node24198 : node24193;
													assign node24193 = (inp[15]) ? node24195 : 4'b0110;
														assign node24195 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node24198 = (inp[15]) ? 4'b0010 : node24199;
														assign node24199 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node24203 = (inp[1]) ? node24225 : node24204;
												assign node24204 = (inp[12]) ? node24218 : node24205;
													assign node24205 = (inp[9]) ? node24211 : node24206;
														assign node24206 = (inp[15]) ? 4'b0010 : node24207;
															assign node24207 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node24211 = (inp[5]) ? node24215 : node24212;
															assign node24212 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node24215 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node24218 = (inp[15]) ? node24222 : node24219;
														assign node24219 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node24222 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node24225 = (inp[12]) ? node24231 : node24226;
													assign node24226 = (inp[15]) ? 4'b0110 : node24227;
														assign node24227 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node24231 = (inp[15]) ? node24233 : 4'b0010;
														assign node24233 = (inp[5]) ? 4'b0010 : 4'b0011;
						assign node24236 = (inp[13]) ? node24838 : node24237;
							assign node24237 = (inp[12]) ? node24461 : node24238;
								assign node24238 = (inp[8]) ? node24334 : node24239;
									assign node24239 = (inp[15]) ? node24263 : node24240;
										assign node24240 = (inp[9]) ? node24252 : node24241;
											assign node24241 = (inp[2]) ? node24247 : node24242;
												assign node24242 = (inp[0]) ? 4'b0010 : node24243;
													assign node24243 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node24247 = (inp[5]) ? node24249 : 4'b0011;
													assign node24249 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node24252 = (inp[2]) ? node24258 : node24253;
												assign node24253 = (inp[5]) ? node24255 : 4'b0011;
													assign node24255 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node24258 = (inp[5]) ? node24260 : 4'b0010;
													assign node24260 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node24263 = (inp[1]) ? node24303 : node24264;
											assign node24264 = (inp[11]) ? node24286 : node24265;
												assign node24265 = (inp[2]) ? node24277 : node24266;
													assign node24266 = (inp[9]) ? node24272 : node24267;
														assign node24267 = (inp[5]) ? node24269 : 4'b0110;
															assign node24269 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node24272 = (inp[5]) ? node24274 : 4'b0111;
															assign node24274 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node24277 = (inp[9]) ? node24281 : node24278;
														assign node24278 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node24281 = (inp[0]) ? 4'b0110 : node24282;
															assign node24282 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node24286 = (inp[2]) ? node24298 : node24287;
													assign node24287 = (inp[9]) ? node24293 : node24288;
														assign node24288 = (inp[5]) ? node24290 : 4'b0110;
															assign node24290 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node24293 = (inp[0]) ? 4'b0111 : node24294;
															assign node24294 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node24298 = (inp[9]) ? node24300 : 4'b0111;
														assign node24300 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node24303 = (inp[5]) ? node24311 : node24304;
												assign node24304 = (inp[9]) ? node24308 : node24305;
													assign node24305 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node24308 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node24311 = (inp[2]) ? node24321 : node24312;
													assign node24312 = (inp[10]) ? node24314 : 4'b0011;
														assign node24314 = (inp[9]) ? node24318 : node24315;
															assign node24315 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node24318 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node24321 = (inp[10]) ? node24329 : node24322;
														assign node24322 = (inp[0]) ? node24326 : node24323;
															assign node24323 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node24326 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node24329 = (inp[0]) ? node24331 : 4'b0011;
															assign node24331 = (inp[9]) ? 4'b0011 : 4'b0010;
									assign node24334 = (inp[1]) ? node24378 : node24335;
										assign node24335 = (inp[15]) ? node24371 : node24336;
											assign node24336 = (inp[2]) ? node24352 : node24337;
												assign node24337 = (inp[10]) ? node24345 : node24338;
													assign node24338 = (inp[0]) ? node24342 : node24339;
														assign node24339 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node24342 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node24345 = (inp[5]) ? node24349 : node24346;
														assign node24346 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node24349 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node24352 = (inp[9]) ? node24366 : node24353;
													assign node24353 = (inp[11]) ? node24359 : node24354;
														assign node24354 = (inp[0]) ? 4'b0010 : node24355;
															assign node24355 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node24359 = (inp[10]) ? 4'b0011 : node24360;
															assign node24360 = (inp[0]) ? node24362 : 4'b0010;
																assign node24362 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node24366 = (inp[5]) ? node24368 : 4'b0010;
														assign node24368 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node24371 = (inp[2]) ? node24375 : node24372;
												assign node24372 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node24375 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node24378 = (inp[0]) ? node24406 : node24379;
											assign node24379 = (inp[5]) ? node24387 : node24380;
												assign node24380 = (inp[2]) ? node24384 : node24381;
													assign node24381 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node24384 = (inp[15]) ? 4'b0110 : 4'b0111;
												assign node24387 = (inp[11]) ? node24395 : node24388;
													assign node24388 = (inp[2]) ? node24392 : node24389;
														assign node24389 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node24392 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node24395 = (inp[10]) ? node24399 : node24396;
														assign node24396 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node24399 = (inp[2]) ? node24403 : node24400;
															assign node24400 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node24403 = (inp[15]) ? 4'b0111 : 4'b0110;
											assign node24406 = (inp[11]) ? node24426 : node24407;
												assign node24407 = (inp[15]) ? node24419 : node24408;
													assign node24408 = (inp[10]) ? node24414 : node24409;
														assign node24409 = (inp[5]) ? 4'b0111 : node24410;
															assign node24410 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node24414 = (inp[2]) ? node24416 : 4'b0110;
															assign node24416 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node24419 = (inp[5]) ? node24423 : node24420;
														assign node24420 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node24423 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node24426 = (inp[10]) ? node24442 : node24427;
													assign node24427 = (inp[15]) ? node24435 : node24428;
														assign node24428 = (inp[2]) ? node24432 : node24429;
															assign node24429 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node24432 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node24435 = (inp[5]) ? node24439 : node24436;
															assign node24436 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node24439 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node24442 = (inp[15]) ? node24452 : node24443;
														assign node24443 = (inp[9]) ? node24445 : 4'b0111;
															assign node24445 = (inp[5]) ? node24449 : node24446;
																assign node24446 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node24449 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node24452 = (inp[9]) ? node24454 : 4'b0110;
															assign node24454 = (inp[5]) ? node24458 : node24455;
																assign node24455 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node24458 = (inp[2]) ? 4'b0110 : 4'b0111;
								assign node24461 = (inp[1]) ? node24579 : node24462;
									assign node24462 = (inp[8]) ? node24556 : node24463;
										assign node24463 = (inp[15]) ? node24487 : node24464;
											assign node24464 = (inp[2]) ? node24476 : node24465;
												assign node24465 = (inp[9]) ? node24471 : node24466;
													assign node24466 = (inp[5]) ? 4'b0110 : node24467;
														assign node24467 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node24471 = (inp[5]) ? 4'b0111 : node24472;
														assign node24472 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node24476 = (inp[9]) ? node24482 : node24477;
													assign node24477 = (inp[0]) ? node24479 : 4'b0111;
														assign node24479 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node24482 = (inp[5]) ? 4'b0110 : node24483;
														assign node24483 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node24487 = (inp[5]) ? node24523 : node24488;
												assign node24488 = (inp[11]) ? node24502 : node24489;
													assign node24489 = (inp[10]) ? node24495 : node24490;
														assign node24490 = (inp[9]) ? node24492 : 4'b0011;
															assign node24492 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node24495 = (inp[2]) ? node24499 : node24496;
															assign node24496 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node24499 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node24502 = (inp[0]) ? node24510 : node24503;
														assign node24503 = (inp[9]) ? node24507 : node24504;
															assign node24504 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24507 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node24510 = (inp[10]) ? node24516 : node24511;
															assign node24511 = (inp[9]) ? 4'b0011 : node24512;
																assign node24512 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24516 = (inp[2]) ? node24520 : node24517;
																assign node24517 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node24520 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node24523 = (inp[11]) ? node24545 : node24524;
													assign node24524 = (inp[10]) ? node24532 : node24525;
														assign node24525 = (inp[9]) ? node24527 : 4'b0010;
															assign node24527 = (inp[2]) ? 4'b0010 : node24528;
																assign node24528 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node24532 = (inp[2]) ? node24540 : node24533;
															assign node24533 = (inp[9]) ? node24537 : node24534;
																assign node24534 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node24537 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node24540 = (inp[9]) ? node24542 : 4'b0011;
																assign node24542 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node24545 = (inp[2]) ? node24551 : node24546;
														assign node24546 = (inp[0]) ? 4'b0010 : node24547;
															assign node24547 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node24551 = (inp[0]) ? 4'b0011 : node24552;
															assign node24552 = (inp[9]) ? 4'b0010 : 4'b0011;
										assign node24556 = (inp[0]) ? node24568 : node24557;
											assign node24557 = (inp[2]) ? node24563 : node24558;
												assign node24558 = (inp[5]) ? 4'b0110 : node24559;
													assign node24559 = (inp[15]) ? 4'b0111 : 4'b0110;
												assign node24563 = (inp[15]) ? node24565 : 4'b0111;
													assign node24565 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node24568 = (inp[2]) ? node24574 : node24569;
												assign node24569 = (inp[15]) ? node24571 : 4'b0111;
													assign node24571 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node24574 = (inp[15]) ? node24576 : 4'b0110;
													assign node24576 = (inp[5]) ? 4'b0110 : 4'b0111;
									assign node24579 = (inp[8]) ? node24697 : node24580;
										assign node24580 = (inp[9]) ? node24640 : node24581;
											assign node24581 = (inp[10]) ? node24611 : node24582;
												assign node24582 = (inp[0]) ? node24596 : node24583;
													assign node24583 = (inp[11]) ? node24589 : node24584;
														assign node24584 = (inp[5]) ? 4'b0111 : node24585;
															assign node24585 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node24589 = (inp[2]) ? node24593 : node24590;
															assign node24590 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node24593 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node24596 = (inp[15]) ? node24602 : node24597;
														assign node24597 = (inp[2]) ? node24599 : 4'b0111;
															assign node24599 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node24602 = (inp[11]) ? node24604 : 4'b0111;
															assign node24604 = (inp[2]) ? node24608 : node24605;
																assign node24605 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node24608 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node24611 = (inp[0]) ? node24619 : node24612;
													assign node24612 = (inp[15]) ? node24616 : node24613;
														assign node24613 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node24616 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node24619 = (inp[2]) ? node24633 : node24620;
														assign node24620 = (inp[11]) ? node24626 : node24621;
															assign node24621 = (inp[15]) ? 4'b0111 : node24622;
																assign node24622 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node24626 = (inp[5]) ? node24630 : node24627;
																assign node24627 = (inp[15]) ? 4'b0111 : 4'b0110;
																assign node24630 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node24633 = (inp[15]) ? node24637 : node24634;
															assign node24634 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node24637 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node24640 = (inp[10]) ? node24674 : node24641;
												assign node24641 = (inp[11]) ? node24657 : node24642;
													assign node24642 = (inp[5]) ? node24650 : node24643;
														assign node24643 = (inp[15]) ? node24645 : 4'b0110;
															assign node24645 = (inp[0]) ? 4'b0110 : node24646;
																assign node24646 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node24650 = (inp[2]) ? node24654 : node24651;
															assign node24651 = (inp[15]) ? 4'b0111 : 4'b0110;
															assign node24654 = (inp[15]) ? 4'b0110 : 4'b0111;
													assign node24657 = (inp[2]) ? node24667 : node24658;
														assign node24658 = (inp[15]) ? node24664 : node24659;
															assign node24659 = (inp[5]) ? 4'b0110 : node24660;
																assign node24660 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node24664 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node24667 = (inp[15]) ? node24669 : 4'b0111;
															assign node24669 = (inp[5]) ? 4'b0110 : node24670;
																assign node24670 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node24674 = (inp[15]) ? node24686 : node24675;
													assign node24675 = (inp[2]) ? node24681 : node24676;
														assign node24676 = (inp[5]) ? 4'b0110 : node24677;
															assign node24677 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node24681 = (inp[0]) ? node24683 : 4'b0111;
															assign node24683 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node24686 = (inp[2]) ? node24692 : node24687;
														assign node24687 = (inp[0]) ? node24689 : 4'b0111;
															assign node24689 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node24692 = (inp[5]) ? 4'b0110 : node24693;
															assign node24693 = (inp[0]) ? 4'b0111 : 4'b0110;
										assign node24697 = (inp[0]) ? node24773 : node24698;
											assign node24698 = (inp[9]) ? node24732 : node24699;
												assign node24699 = (inp[11]) ? node24711 : node24700;
													assign node24700 = (inp[15]) ? node24702 : 4'b0011;
														assign node24702 = (inp[10]) ? 4'b0011 : node24703;
															assign node24703 = (inp[2]) ? node24707 : node24704;
																assign node24704 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node24707 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node24711 = (inp[2]) ? node24719 : node24712;
														assign node24712 = (inp[5]) ? node24716 : node24713;
															assign node24713 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node24716 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node24719 = (inp[10]) ? node24727 : node24720;
															assign node24720 = (inp[15]) ? node24724 : node24721;
																assign node24721 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node24724 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node24727 = (inp[15]) ? node24729 : 4'b0011;
																assign node24729 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node24732 = (inp[11]) ? node24756 : node24733;
													assign node24733 = (inp[10]) ? node24747 : node24734;
														assign node24734 = (inp[15]) ? node24740 : node24735;
															assign node24735 = (inp[5]) ? node24737 : 4'b0010;
																assign node24737 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24740 = (inp[5]) ? node24744 : node24741;
																assign node24741 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node24744 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node24747 = (inp[2]) ? node24749 : 4'b0010;
															assign node24749 = (inp[5]) ? node24753 : node24750;
																assign node24750 = (inp[15]) ? 4'b0010 : 4'b0011;
																assign node24753 = (inp[15]) ? 4'b0011 : 4'b0010;
													assign node24756 = (inp[10]) ? node24758 : 4'b0011;
														assign node24758 = (inp[5]) ? node24766 : node24759;
															assign node24759 = (inp[15]) ? node24763 : node24760;
																assign node24760 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node24763 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24766 = (inp[2]) ? node24770 : node24767;
																assign node24767 = (inp[15]) ? 4'b0010 : 4'b0011;
																assign node24770 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node24773 = (inp[9]) ? node24799 : node24774;
												assign node24774 = (inp[15]) ? node24782 : node24775;
													assign node24775 = (inp[2]) ? node24779 : node24776;
														assign node24776 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node24779 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node24782 = (inp[11]) ? node24792 : node24783;
														assign node24783 = (inp[10]) ? node24785 : 4'b0010;
															assign node24785 = (inp[5]) ? node24789 : node24786;
																assign node24786 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node24789 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node24792 = (inp[2]) ? node24796 : node24793;
															assign node24793 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node24796 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node24799 = (inp[11]) ? node24823 : node24800;
													assign node24800 = (inp[2]) ? node24808 : node24801;
														assign node24801 = (inp[5]) ? node24805 : node24802;
															assign node24802 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node24805 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node24808 = (inp[10]) ? node24816 : node24809;
															assign node24809 = (inp[5]) ? node24813 : node24810;
																assign node24810 = (inp[15]) ? 4'b0011 : 4'b0010;
																assign node24813 = (inp[15]) ? 4'b0010 : 4'b0011;
															assign node24816 = (inp[5]) ? node24820 : node24817;
																assign node24817 = (inp[15]) ? 4'b0011 : 4'b0010;
																assign node24820 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node24823 = (inp[15]) ? node24831 : node24824;
														assign node24824 = (inp[5]) ? node24828 : node24825;
															assign node24825 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24828 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node24831 = (inp[5]) ? node24835 : node24832;
															assign node24832 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node24835 = (inp[2]) ? 4'b0010 : 4'b0011;
							assign node24838 = (inp[12]) ? node25136 : node24839;
								assign node24839 = (inp[1]) ? node25025 : node24840;
									assign node24840 = (inp[8]) ? node24978 : node24841;
										assign node24841 = (inp[15]) ? node24911 : node24842;
											assign node24842 = (inp[10]) ? node24876 : node24843;
												assign node24843 = (inp[11]) ? node24865 : node24844;
													assign node24844 = (inp[9]) ? node24856 : node24845;
														assign node24845 = (inp[2]) ? node24851 : node24846;
															assign node24846 = (inp[0]) ? 4'b0110 : node24847;
																assign node24847 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node24851 = (inp[5]) ? node24853 : 4'b0111;
																assign node24853 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node24856 = (inp[2]) ? node24862 : node24857;
															assign node24857 = (inp[0]) ? 4'b0111 : node24858;
																assign node24858 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node24862 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node24865 = (inp[2]) ? node24867 : 4'b0111;
														assign node24867 = (inp[9]) ? node24873 : node24868;
															assign node24868 = (inp[5]) ? node24870 : 4'b0111;
																assign node24870 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node24873 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node24876 = (inp[5]) ? node24896 : node24877;
													assign node24877 = (inp[0]) ? node24889 : node24878;
														assign node24878 = (inp[11]) ? node24884 : node24879;
															assign node24879 = (inp[2]) ? node24881 : 4'b0110;
																assign node24881 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node24884 = (inp[9]) ? node24886 : 4'b0110;
																assign node24886 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node24889 = (inp[2]) ? node24893 : node24890;
															assign node24890 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node24893 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node24896 = (inp[9]) ? node24904 : node24897;
														assign node24897 = (inp[0]) ? node24901 : node24898;
															assign node24898 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node24901 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node24904 = (inp[0]) ? node24908 : node24905;
															assign node24905 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node24908 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node24911 = (inp[0]) ? node24949 : node24912;
												assign node24912 = (inp[11]) ? node24934 : node24913;
													assign node24913 = (inp[5]) ? node24927 : node24914;
														assign node24914 = (inp[10]) ? node24922 : node24915;
															assign node24915 = (inp[2]) ? node24919 : node24916;
																assign node24916 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node24919 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node24922 = (inp[2]) ? node24924 : 4'b0011;
																assign node24924 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node24927 = (inp[9]) ? node24931 : node24928;
															assign node24928 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node24931 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node24934 = (inp[5]) ? node24942 : node24935;
														assign node24935 = (inp[10]) ? 4'b0010 : node24936;
															assign node24936 = (inp[2]) ? 4'b0011 : node24937;
																assign node24937 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node24942 = (inp[2]) ? node24946 : node24943;
															assign node24943 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node24946 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node24949 = (inp[5]) ? node24969 : node24950;
													assign node24950 = (inp[10]) ? node24962 : node24951;
														assign node24951 = (inp[11]) ? node24957 : node24952;
															assign node24952 = (inp[9]) ? 4'b0010 : node24953;
																assign node24953 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node24957 = (inp[2]) ? 4'b0010 : node24958;
																assign node24958 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node24962 = (inp[9]) ? node24966 : node24963;
															assign node24963 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node24966 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node24969 = (inp[10]) ? 4'b0010 : node24970;
														assign node24970 = (inp[2]) ? node24974 : node24971;
															assign node24971 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node24974 = (inp[9]) ? 4'b0011 : 4'b0010;
										assign node24978 = (inp[9]) ? node25002 : node24979;
											assign node24979 = (inp[0]) ? node24991 : node24980;
												assign node24980 = (inp[2]) ? node24986 : node24981;
													assign node24981 = (inp[15]) ? node24983 : 4'b0010;
														assign node24983 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node24986 = (inp[5]) ? node24988 : 4'b0011;
														assign node24988 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node24991 = (inp[2]) ? node24997 : node24992;
													assign node24992 = (inp[5]) ? node24994 : 4'b0011;
														assign node24994 = (inp[15]) ? 4'b0010 : 4'b0011;
													assign node24997 = (inp[5]) ? node24999 : 4'b0010;
														assign node24999 = (inp[15]) ? 4'b0011 : 4'b0010;
											assign node25002 = (inp[2]) ? node25014 : node25003;
												assign node25003 = (inp[0]) ? node25009 : node25004;
													assign node25004 = (inp[15]) ? node25006 : 4'b0010;
														assign node25006 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node25009 = (inp[15]) ? node25011 : 4'b0011;
														assign node25011 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node25014 = (inp[0]) ? node25020 : node25015;
													assign node25015 = (inp[15]) ? node25017 : 4'b0011;
														assign node25017 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node25020 = (inp[5]) ? node25022 : 4'b0010;
														assign node25022 = (inp[15]) ? 4'b0011 : 4'b0010;
									assign node25025 = (inp[5]) ? node25113 : node25026;
										assign node25026 = (inp[15]) ? node25090 : node25027;
											assign node25027 = (inp[8]) ? node25061 : node25028;
												assign node25028 = (inp[10]) ? node25042 : node25029;
													assign node25029 = (inp[0]) ? node25035 : node25030;
														assign node25030 = (inp[2]) ? 4'b0111 : node25031;
															assign node25031 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node25035 = (inp[2]) ? node25039 : node25036;
															assign node25036 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node25039 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node25042 = (inp[11]) ? node25054 : node25043;
														assign node25043 = (inp[0]) ? node25049 : node25044;
															assign node25044 = (inp[9]) ? 4'b0111 : node25045;
																assign node25045 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node25049 = (inp[9]) ? node25051 : 4'b0111;
																assign node25051 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node25054 = (inp[9]) ? node25058 : node25055;
															assign node25055 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node25058 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node25061 = (inp[11]) ? node25069 : node25062;
													assign node25062 = (inp[2]) ? node25066 : node25063;
														assign node25063 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node25066 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node25069 = (inp[10]) ? node25083 : node25070;
														assign node25070 = (inp[9]) ? node25076 : node25071;
															assign node25071 = (inp[2]) ? 4'b0111 : node25072;
																assign node25072 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node25076 = (inp[2]) ? node25080 : node25077;
																assign node25077 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node25080 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node25083 = (inp[2]) ? node25087 : node25084;
															assign node25084 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node25087 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node25090 = (inp[2]) ? node25102 : node25091;
												assign node25091 = (inp[9]) ? node25097 : node25092;
													assign node25092 = (inp[0]) ? node25094 : 4'b0110;
														assign node25094 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node25097 = (inp[0]) ? 4'b0111 : node25098;
														assign node25098 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node25102 = (inp[9]) ? node25108 : node25103;
													assign node25103 = (inp[8]) ? node25105 : 4'b0111;
														assign node25105 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node25108 = (inp[8]) ? node25110 : 4'b0110;
														assign node25110 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node25113 = (inp[2]) ? node25125 : node25114;
											assign node25114 = (inp[0]) ? node25120 : node25115;
												assign node25115 = (inp[9]) ? 4'b0110 : node25116;
													assign node25116 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node25120 = (inp[9]) ? 4'b0111 : node25121;
													assign node25121 = (inp[8]) ? 4'b0111 : 4'b0110;
											assign node25125 = (inp[0]) ? node25131 : node25126;
												assign node25126 = (inp[9]) ? 4'b0111 : node25127;
													assign node25127 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node25131 = (inp[9]) ? 4'b0110 : node25132;
													assign node25132 = (inp[8]) ? 4'b0110 : 4'b0111;
								assign node25136 = (inp[1]) ? node25312 : node25137;
									assign node25137 = (inp[15]) ? node25265 : node25138;
										assign node25138 = (inp[8]) ? node25206 : node25139;
											assign node25139 = (inp[11]) ? node25173 : node25140;
												assign node25140 = (inp[5]) ? node25162 : node25141;
													assign node25141 = (inp[10]) ? node25155 : node25142;
														assign node25142 = (inp[0]) ? node25148 : node25143;
															assign node25143 = (inp[9]) ? node25145 : 4'b0011;
																assign node25145 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node25148 = (inp[2]) ? node25152 : node25149;
																assign node25149 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node25152 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node25155 = (inp[9]) ? node25159 : node25156;
															assign node25156 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node25159 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node25162 = (inp[9]) ? node25164 : 4'b0010;
														assign node25164 = (inp[10]) ? 4'b0010 : node25165;
															assign node25165 = (inp[2]) ? node25169 : node25166;
																assign node25166 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node25169 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node25173 = (inp[5]) ? node25181 : node25174;
													assign node25174 = (inp[9]) ? node25178 : node25175;
														assign node25175 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node25178 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node25181 = (inp[10]) ? node25197 : node25182;
														assign node25182 = (inp[0]) ? node25190 : node25183;
															assign node25183 = (inp[9]) ? node25187 : node25184;
																assign node25184 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node25187 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node25190 = (inp[2]) ? node25194 : node25191;
																assign node25191 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node25194 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node25197 = (inp[0]) ? node25199 : 4'b0011;
															assign node25199 = (inp[9]) ? node25203 : node25200;
																assign node25200 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node25203 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node25206 = (inp[10]) ? node25230 : node25207;
												assign node25207 = (inp[5]) ? node25215 : node25208;
													assign node25208 = (inp[2]) ? node25212 : node25209;
														assign node25209 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node25212 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node25215 = (inp[9]) ? node25223 : node25216;
														assign node25216 = (inp[2]) ? node25220 : node25217;
															assign node25217 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node25220 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node25223 = (inp[2]) ? node25227 : node25224;
															assign node25224 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node25227 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node25230 = (inp[9]) ? node25250 : node25231;
													assign node25231 = (inp[5]) ? node25245 : node25232;
														assign node25232 = (inp[11]) ? node25238 : node25233;
															assign node25233 = (inp[2]) ? 4'b0110 : node25234;
																assign node25234 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node25238 = (inp[2]) ? node25242 : node25239;
																assign node25239 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node25242 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node25245 = (inp[0]) ? 4'b0111 : node25246;
															assign node25246 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node25250 = (inp[11]) ? node25258 : node25251;
														assign node25251 = (inp[2]) ? 4'b0111 : node25252;
															assign node25252 = (inp[0]) ? 4'b0110 : node25253;
																assign node25253 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node25258 = (inp[2]) ? node25260 : 4'b0111;
															assign node25260 = (inp[0]) ? 4'b0111 : node25261;
																assign node25261 = (inp[5]) ? 4'b0111 : 4'b0110;
										assign node25265 = (inp[5]) ? node25289 : node25266;
											assign node25266 = (inp[9]) ? node25278 : node25267;
												assign node25267 = (inp[2]) ? node25273 : node25268;
													assign node25268 = (inp[0]) ? node25270 : 4'b0110;
														assign node25270 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node25273 = (inp[8]) ? node25275 : 4'b0111;
														assign node25275 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node25278 = (inp[2]) ? node25284 : node25279;
													assign node25279 = (inp[0]) ? 4'b0111 : node25280;
														assign node25280 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node25284 = (inp[8]) ? node25286 : 4'b0110;
														assign node25286 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node25289 = (inp[2]) ? node25301 : node25290;
												assign node25290 = (inp[0]) ? node25296 : node25291;
													assign node25291 = (inp[8]) ? 4'b0110 : node25292;
														assign node25292 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node25296 = (inp[9]) ? 4'b0111 : node25297;
														assign node25297 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node25301 = (inp[0]) ? node25307 : node25302;
													assign node25302 = (inp[9]) ? 4'b0111 : node25303;
														assign node25303 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node25307 = (inp[9]) ? 4'b0110 : node25308;
														assign node25308 = (inp[8]) ? 4'b0110 : 4'b0111;
									assign node25312 = (inp[9]) ? node25332 : node25313;
										assign node25313 = (inp[2]) ? node25323 : node25314;
											assign node25314 = (inp[0]) ? node25320 : node25315;
												assign node25315 = (inp[5]) ? node25317 : 4'b0010;
													assign node25317 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node25320 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node25323 = (inp[0]) ? node25329 : node25324;
												assign node25324 = (inp[8]) ? 4'b0011 : node25325;
													assign node25325 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node25329 = (inp[8]) ? 4'b0010 : 4'b0011;
										assign node25332 = (inp[2]) ? node25340 : node25333;
											assign node25333 = (inp[0]) ? 4'b0011 : node25334;
												assign node25334 = (inp[5]) ? 4'b0010 : node25335;
													assign node25335 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node25340 = (inp[0]) ? 4'b0010 : node25341;
												assign node25341 = (inp[5]) ? 4'b0011 : node25342;
													assign node25342 = (inp[8]) ? 4'b0011 : 4'b0010;
					assign node25347 = (inp[7]) ? node26175 : node25348;
						assign node25348 = (inp[8]) ? node25948 : node25349;
							assign node25349 = (inp[12]) ? node25555 : node25350;
								assign node25350 = (inp[13]) ? node25510 : node25351;
									assign node25351 = (inp[15]) ? node25433 : node25352;
										assign node25352 = (inp[10]) ? node25398 : node25353;
											assign node25353 = (inp[11]) ? node25385 : node25354;
												assign node25354 = (inp[2]) ? node25378 : node25355;
													assign node25355 = (inp[0]) ? node25365 : node25356;
														assign node25356 = (inp[1]) ? 4'b0011 : node25357;
															assign node25357 = (inp[9]) ? node25361 : node25358;
																assign node25358 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node25361 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node25365 = (inp[1]) ? node25371 : node25366;
															assign node25366 = (inp[9]) ? node25368 : 4'b0011;
																assign node25368 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node25371 = (inp[9]) ? node25375 : node25372;
																assign node25372 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node25375 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node25378 = (inp[9]) ? node25382 : node25379;
														assign node25379 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node25382 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node25385 = (inp[1]) ? node25391 : node25386;
													assign node25386 = (inp[9]) ? 4'b0010 : node25387;
														assign node25387 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node25391 = (inp[5]) ? node25395 : node25392;
														assign node25392 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node25395 = (inp[9]) ? 4'b0010 : 4'b0011;
											assign node25398 = (inp[11]) ? node25406 : node25399;
												assign node25399 = (inp[9]) ? node25403 : node25400;
													assign node25400 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node25403 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node25406 = (inp[2]) ? node25424 : node25407;
													assign node25407 = (inp[1]) ? node25415 : node25408;
														assign node25408 = (inp[5]) ? node25412 : node25409;
															assign node25409 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node25412 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node25415 = (inp[0]) ? node25417 : 4'b0011;
															assign node25417 = (inp[5]) ? node25421 : node25418;
																assign node25418 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node25421 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node25424 = (inp[1]) ? node25426 : 4'b0011;
														assign node25426 = (inp[9]) ? node25430 : node25427;
															assign node25427 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node25430 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node25433 = (inp[10]) ? node25473 : node25434;
											assign node25434 = (inp[1]) ? node25450 : node25435;
												assign node25435 = (inp[2]) ? node25443 : node25436;
													assign node25436 = (inp[5]) ? node25440 : node25437;
														assign node25437 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node25440 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node25443 = (inp[9]) ? node25447 : node25444;
														assign node25444 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node25447 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node25450 = (inp[5]) ? node25458 : node25451;
													assign node25451 = (inp[0]) ? node25455 : node25452;
														assign node25452 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node25455 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node25458 = (inp[11]) ? node25466 : node25459;
														assign node25459 = (inp[0]) ? node25463 : node25460;
															assign node25460 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node25463 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node25466 = (inp[9]) ? node25470 : node25467;
															assign node25467 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node25470 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node25473 = (inp[0]) ? node25481 : node25474;
												assign node25474 = (inp[5]) ? node25478 : node25475;
													assign node25475 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node25478 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node25481 = (inp[11]) ? node25501 : node25482;
													assign node25482 = (inp[5]) ? node25494 : node25483;
														assign node25483 = (inp[2]) ? node25489 : node25484;
															assign node25484 = (inp[9]) ? 4'b0110 : node25485;
																assign node25485 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node25489 = (inp[9]) ? node25491 : 4'b0110;
																assign node25491 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node25494 = (inp[9]) ? node25498 : node25495;
															assign node25495 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node25498 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node25501 = (inp[9]) ? node25505 : node25502;
														assign node25502 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node25505 = (inp[1]) ? 4'b0111 : node25506;
															assign node25506 = (inp[5]) ? 4'b0110 : 4'b0111;
									assign node25510 = (inp[15]) ? node25518 : node25511;
										assign node25511 = (inp[9]) ? node25515 : node25512;
											assign node25512 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node25515 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node25518 = (inp[1]) ? node25548 : node25519;
											assign node25519 = (inp[5]) ? node25527 : node25520;
												assign node25520 = (inp[0]) ? node25524 : node25521;
													assign node25521 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node25524 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node25527 = (inp[10]) ? node25535 : node25528;
													assign node25528 = (inp[9]) ? node25532 : node25529;
														assign node25529 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node25532 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node25535 = (inp[11]) ? node25541 : node25536;
														assign node25536 = (inp[9]) ? 4'b0011 : node25537;
															assign node25537 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node25541 = (inp[9]) ? node25545 : node25542;
															assign node25542 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node25545 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node25548 = (inp[5]) ? node25552 : node25549;
												assign node25549 = (inp[9]) ? 4'b0011 : 4'b0010;
												assign node25552 = (inp[9]) ? 4'b0010 : 4'b0011;
								assign node25555 = (inp[11]) ? node25687 : node25556;
									assign node25556 = (inp[9]) ? node25626 : node25557;
										assign node25557 = (inp[5]) ? node25599 : node25558;
											assign node25558 = (inp[15]) ? node25588 : node25559;
												assign node25559 = (inp[13]) ? node25581 : node25560;
													assign node25560 = (inp[2]) ? node25574 : node25561;
														assign node25561 = (inp[10]) ? node25569 : node25562;
															assign node25562 = (inp[1]) ? node25566 : node25563;
																assign node25563 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node25566 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node25569 = (inp[1]) ? node25571 : 4'b0010;
																assign node25571 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node25574 = (inp[1]) ? node25578 : node25575;
															assign node25575 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node25578 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node25581 = (inp[0]) ? node25585 : node25582;
														assign node25582 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node25585 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node25588 = (inp[13]) ? node25594 : node25589;
													assign node25589 = (inp[1]) ? 4'b0110 : node25590;
														assign node25590 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node25594 = (inp[1]) ? node25596 : 4'b0010;
														assign node25596 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node25599 = (inp[15]) ? node25615 : node25600;
												assign node25600 = (inp[13]) ? node25608 : node25601;
													assign node25601 = (inp[1]) ? node25605 : node25602;
														assign node25602 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node25605 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node25608 = (inp[0]) ? node25612 : node25609;
														assign node25609 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node25612 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node25615 = (inp[13]) ? node25621 : node25616;
													assign node25616 = (inp[1]) ? 4'b0111 : node25617;
														assign node25617 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node25621 = (inp[0]) ? 4'b0011 : node25622;
														assign node25622 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node25626 = (inp[5]) ? node25660 : node25627;
											assign node25627 = (inp[15]) ? node25649 : node25628;
												assign node25628 = (inp[13]) ? node25636 : node25629;
													assign node25629 = (inp[0]) ? node25633 : node25630;
														assign node25630 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node25633 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node25636 = (inp[2]) ? node25644 : node25637;
														assign node25637 = (inp[0]) ? node25641 : node25638;
															assign node25638 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node25641 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node25644 = (inp[10]) ? node25646 : 4'b0111;
															assign node25646 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node25649 = (inp[13]) ? node25655 : node25650;
													assign node25650 = (inp[0]) ? node25652 : 4'b0111;
														assign node25652 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node25655 = (inp[1]) ? node25657 : 4'b0011;
														assign node25657 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node25660 = (inp[15]) ? node25676 : node25661;
												assign node25661 = (inp[13]) ? node25669 : node25662;
													assign node25662 = (inp[0]) ? node25666 : node25663;
														assign node25663 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node25666 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node25669 = (inp[1]) ? node25673 : node25670;
														assign node25670 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node25673 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node25676 = (inp[13]) ? node25682 : node25677;
													assign node25677 = (inp[1]) ? 4'b0110 : node25678;
														assign node25678 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node25682 = (inp[1]) ? node25684 : 4'b0010;
														assign node25684 = (inp[0]) ? 4'b0010 : 4'b0011;
									assign node25687 = (inp[10]) ? node25803 : node25688;
										assign node25688 = (inp[15]) ? node25760 : node25689;
											assign node25689 = (inp[13]) ? node25727 : node25690;
												assign node25690 = (inp[1]) ? node25712 : node25691;
													assign node25691 = (inp[5]) ? node25697 : node25692;
														assign node25692 = (inp[9]) ? node25694 : 4'b0011;
															assign node25694 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node25697 = (inp[2]) ? node25705 : node25698;
															assign node25698 = (inp[9]) ? node25702 : node25699;
																assign node25699 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node25702 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node25705 = (inp[0]) ? node25709 : node25706;
																assign node25706 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node25709 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node25712 = (inp[9]) ? node25720 : node25713;
														assign node25713 = (inp[0]) ? node25717 : node25714;
															assign node25714 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node25717 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node25720 = (inp[0]) ? node25724 : node25721;
															assign node25721 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node25724 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node25727 = (inp[9]) ? node25745 : node25728;
													assign node25728 = (inp[0]) ? node25738 : node25729;
														assign node25729 = (inp[2]) ? node25735 : node25730;
															assign node25730 = (inp[1]) ? 4'b0111 : node25731;
																assign node25731 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node25735 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node25738 = (inp[1]) ? node25742 : node25739;
															assign node25739 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node25742 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node25745 = (inp[1]) ? node25755 : node25746;
														assign node25746 = (inp[2]) ? node25750 : node25747;
															assign node25747 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node25750 = (inp[0]) ? 4'b0111 : node25751;
																assign node25751 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node25755 = (inp[5]) ? node25757 : 4'b0111;
															assign node25757 = (inp[2]) ? 4'b0110 : 4'b0111;
											assign node25760 = (inp[13]) ? node25780 : node25761;
												assign node25761 = (inp[5]) ? node25773 : node25762;
													assign node25762 = (inp[9]) ? node25768 : node25763;
														assign node25763 = (inp[1]) ? 4'b0110 : node25764;
															assign node25764 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node25768 = (inp[0]) ? node25770 : 4'b0111;
															assign node25770 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node25773 = (inp[9]) ? node25775 : 4'b0111;
														assign node25775 = (inp[1]) ? 4'b0110 : node25776;
															assign node25776 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node25780 = (inp[9]) ? node25792 : node25781;
													assign node25781 = (inp[5]) ? node25787 : node25782;
														assign node25782 = (inp[0]) ? 4'b0010 : node25783;
															assign node25783 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node25787 = (inp[1]) ? node25789 : 4'b0011;
															assign node25789 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node25792 = (inp[5]) ? node25798 : node25793;
														assign node25793 = (inp[0]) ? 4'b0011 : node25794;
															assign node25794 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node25798 = (inp[1]) ? node25800 : 4'b0010;
															assign node25800 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node25803 = (inp[2]) ? node25873 : node25804;
											assign node25804 = (inp[15]) ? node25842 : node25805;
												assign node25805 = (inp[13]) ? node25825 : node25806;
													assign node25806 = (inp[0]) ? node25814 : node25807;
														assign node25807 = (inp[9]) ? node25809 : 4'b0010;
															assign node25809 = (inp[5]) ? node25811 : 4'b0010;
																assign node25811 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node25814 = (inp[1]) ? node25820 : node25815;
															assign node25815 = (inp[5]) ? 4'b0011 : node25816;
																assign node25816 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node25820 = (inp[9]) ? node25822 : 4'b0010;
																assign node25822 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node25825 = (inp[9]) ? node25837 : node25826;
														assign node25826 = (inp[0]) ? node25832 : node25827;
															assign node25827 = (inp[1]) ? 4'b0110 : node25828;
																assign node25828 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node25832 = (inp[5]) ? node25834 : 4'b0111;
																assign node25834 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node25837 = (inp[5]) ? 4'b0110 : node25838;
															assign node25838 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node25842 = (inp[13]) ? node25862 : node25843;
													assign node25843 = (inp[9]) ? node25851 : node25844;
														assign node25844 = (inp[5]) ? 4'b0111 : node25845;
															assign node25845 = (inp[1]) ? 4'b0110 : node25846;
																assign node25846 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node25851 = (inp[5]) ? node25857 : node25852;
															assign node25852 = (inp[0]) ? node25854 : 4'b0111;
																assign node25854 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node25857 = (inp[0]) ? node25859 : 4'b0110;
																assign node25859 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node25862 = (inp[5]) ? node25864 : 4'b0010;
														assign node25864 = (inp[9]) ? node25870 : node25865;
															assign node25865 = (inp[0]) ? 4'b0011 : node25866;
																assign node25866 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node25870 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node25873 = (inp[13]) ? node25909 : node25874;
												assign node25874 = (inp[15]) ? node25898 : node25875;
													assign node25875 = (inp[5]) ? node25889 : node25876;
														assign node25876 = (inp[0]) ? node25884 : node25877;
															assign node25877 = (inp[9]) ? node25881 : node25878;
																assign node25878 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node25881 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node25884 = (inp[1]) ? 4'b0011 : node25885;
																assign node25885 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node25889 = (inp[9]) ? node25891 : 4'b0010;
															assign node25891 = (inp[1]) ? node25895 : node25892;
																assign node25892 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node25895 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node25898 = (inp[5]) ? node25902 : node25899;
														assign node25899 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node25902 = (inp[9]) ? node25904 : 4'b0111;
															assign node25904 = (inp[0]) ? node25906 : 4'b0110;
																assign node25906 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node25909 = (inp[15]) ? node25929 : node25910;
													assign node25910 = (inp[9]) ? node25920 : node25911;
														assign node25911 = (inp[1]) ? 4'b0111 : node25912;
															assign node25912 = (inp[0]) ? node25916 : node25913;
																assign node25913 = (inp[5]) ? 4'b0111 : 4'b0110;
																assign node25916 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node25920 = (inp[1]) ? node25922 : 4'b0111;
															assign node25922 = (inp[5]) ? node25926 : node25923;
																assign node25923 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node25926 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node25929 = (inp[9]) ? node25939 : node25930;
														assign node25930 = (inp[5]) ? node25936 : node25931;
															assign node25931 = (inp[0]) ? 4'b0010 : node25932;
																assign node25932 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node25936 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node25939 = (inp[1]) ? node25941 : 4'b0011;
															assign node25941 = (inp[5]) ? node25945 : node25942;
																assign node25942 = (inp[0]) ? 4'b0011 : 4'b0010;
																assign node25945 = (inp[0]) ? 4'b0010 : 4'b0011;
							assign node25948 = (inp[5]) ? node25996 : node25949;
								assign node25949 = (inp[0]) ? node25973 : node25950;
									assign node25950 = (inp[12]) ? node25962 : node25951;
										assign node25951 = (inp[15]) ? node25955 : node25952;
											assign node25952 = (inp[1]) ? 4'b0100 : 4'b0000;
											assign node25955 = (inp[1]) ? node25959 : node25956;
												assign node25956 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node25959 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node25962 = (inp[15]) ? node25970 : node25963;
											assign node25963 = (inp[1]) ? node25967 : node25964;
												assign node25964 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node25967 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node25970 = (inp[1]) ? 4'b0000 : 4'b0100;
									assign node25973 = (inp[1]) ? node25985 : node25974;
										assign node25974 = (inp[15]) ? node25980 : node25975;
											assign node25975 = (inp[13]) ? node25977 : 4'b0001;
												assign node25977 = (inp[12]) ? 4'b0000 : 4'b0001;
											assign node25980 = (inp[13]) ? node25982 : 4'b0101;
												assign node25982 = (inp[12]) ? 4'b0101 : 4'b0100;
										assign node25985 = (inp[15]) ? node25991 : node25986;
											assign node25986 = (inp[12]) ? node25988 : 4'b0101;
												assign node25988 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node25991 = (inp[12]) ? 4'b0001 : node25992;
												assign node25992 = (inp[13]) ? 4'b0001 : 4'b0000;
								assign node25996 = (inp[0]) ? node26152 : node25997;
									assign node25997 = (inp[10]) ? node26071 : node25998;
										assign node25998 = (inp[9]) ? node26022 : node25999;
											assign node25999 = (inp[12]) ? node26011 : node26000;
												assign node26000 = (inp[15]) ? node26004 : node26001;
													assign node26001 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node26004 = (inp[1]) ? node26008 : node26005;
														assign node26005 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node26008 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node26011 = (inp[15]) ? node26019 : node26012;
													assign node26012 = (inp[1]) ? node26016 : node26013;
														assign node26013 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node26016 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node26019 = (inp[1]) ? 4'b0001 : 4'b0101;
											assign node26022 = (inp[11]) ? node26046 : node26023;
												assign node26023 = (inp[15]) ? node26035 : node26024;
													assign node26024 = (inp[1]) ? node26030 : node26025;
														assign node26025 = (inp[12]) ? node26027 : 4'b0001;
															assign node26027 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node26030 = (inp[12]) ? node26032 : 4'b0101;
															assign node26032 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node26035 = (inp[1]) ? node26041 : node26036;
														assign node26036 = (inp[12]) ? 4'b0101 : node26037;
															assign node26037 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node26041 = (inp[12]) ? 4'b0001 : node26042;
															assign node26042 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node26046 = (inp[1]) ? node26058 : node26047;
													assign node26047 = (inp[15]) ? node26053 : node26048;
														assign node26048 = (inp[13]) ? node26050 : 4'b0001;
															assign node26050 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node26053 = (inp[12]) ? 4'b0101 : node26054;
															assign node26054 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node26058 = (inp[15]) ? node26066 : node26059;
														assign node26059 = (inp[2]) ? 4'b0101 : node26060;
															assign node26060 = (inp[13]) ? 4'b0101 : node26061;
																assign node26061 = (inp[12]) ? 4'b0100 : 4'b0101;
														assign node26066 = (inp[13]) ? 4'b0001 : node26067;
															assign node26067 = (inp[12]) ? 4'b0001 : 4'b0000;
										assign node26071 = (inp[11]) ? node26129 : node26072;
											assign node26072 = (inp[2]) ? node26092 : node26073;
												assign node26073 = (inp[13]) ? node26085 : node26074;
													assign node26074 = (inp[1]) ? node26078 : node26075;
														assign node26075 = (inp[15]) ? 4'b0101 : 4'b0001;
														assign node26078 = (inp[15]) ? node26082 : node26079;
															assign node26079 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node26082 = (inp[12]) ? 4'b0001 : 4'b0000;
													assign node26085 = (inp[1]) ? node26089 : node26086;
														assign node26086 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node26089 = (inp[15]) ? 4'b0001 : 4'b0101;
												assign node26092 = (inp[9]) ? node26112 : node26093;
													assign node26093 = (inp[1]) ? node26103 : node26094;
														assign node26094 = (inp[15]) ? node26100 : node26095;
															assign node26095 = (inp[12]) ? node26097 : 4'b0001;
																assign node26097 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node26100 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node26103 = (inp[15]) ? node26107 : node26104;
															assign node26104 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node26107 = (inp[12]) ? 4'b0001 : node26108;
																assign node26108 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node26112 = (inp[1]) ? node26120 : node26113;
														assign node26113 = (inp[15]) ? node26117 : node26114;
															assign node26114 = (inp[12]) ? 4'b0000 : 4'b0001;
															assign node26117 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node26120 = (inp[15]) ? node26126 : node26121;
															assign node26121 = (inp[12]) ? node26123 : 4'b0101;
																assign node26123 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node26126 = (inp[12]) ? 4'b0001 : 4'b0000;
											assign node26129 = (inp[12]) ? node26141 : node26130;
												assign node26130 = (inp[15]) ? node26134 : node26131;
													assign node26131 = (inp[1]) ? 4'b0101 : 4'b0001;
													assign node26134 = (inp[1]) ? node26138 : node26135;
														assign node26135 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node26138 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node26141 = (inp[15]) ? node26149 : node26142;
													assign node26142 = (inp[1]) ? node26146 : node26143;
														assign node26143 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node26146 = (inp[13]) ? 4'b0101 : 4'b0100;
													assign node26149 = (inp[1]) ? 4'b0001 : 4'b0101;
									assign node26152 = (inp[12]) ? node26164 : node26153;
										assign node26153 = (inp[15]) ? node26157 : node26154;
											assign node26154 = (inp[1]) ? 4'b0100 : 4'b0000;
											assign node26157 = (inp[1]) ? node26161 : node26158;
												assign node26158 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node26161 = (inp[13]) ? 4'b0000 : 4'b0001;
										assign node26164 = (inp[15]) ? node26172 : node26165;
											assign node26165 = (inp[1]) ? node26169 : node26166;
												assign node26166 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node26169 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node26172 = (inp[1]) ? 4'b0000 : 4'b0100;
						assign node26175 = (inp[1]) ? node26361 : node26176;
							assign node26176 = (inp[8]) ? node26224 : node26177;
								assign node26177 = (inp[13]) ? node26201 : node26178;
									assign node26178 = (inp[9]) ? node26190 : node26179;
										assign node26179 = (inp[12]) ? node26185 : node26180;
											assign node26180 = (inp[0]) ? node26182 : 4'b0000;
												assign node26182 = (inp[15]) ? 4'b0001 : 4'b0000;
											assign node26185 = (inp[0]) ? node26187 : 4'b0001;
												assign node26187 = (inp[15]) ? 4'b0000 : 4'b0001;
										assign node26190 = (inp[12]) ? node26196 : node26191;
											assign node26191 = (inp[15]) ? node26193 : 4'b0001;
												assign node26193 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node26196 = (inp[0]) ? node26198 : 4'b0000;
												assign node26198 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node26201 = (inp[9]) ? node26213 : node26202;
										assign node26202 = (inp[12]) ? node26208 : node26203;
											assign node26203 = (inp[15]) ? node26205 : 4'b0100;
												assign node26205 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node26208 = (inp[15]) ? node26210 : 4'b0101;
												assign node26210 = (inp[0]) ? 4'b0101 : 4'b0100;
										assign node26213 = (inp[12]) ? node26219 : node26214;
											assign node26214 = (inp[0]) ? 4'b0101 : node26215;
												assign node26215 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node26219 = (inp[0]) ? 4'b0100 : node26220;
												assign node26220 = (inp[15]) ? 4'b0101 : 4'b0100;
								assign node26224 = (inp[13]) ? node26292 : node26225;
									assign node26225 = (inp[5]) ? node26233 : node26226;
										assign node26226 = (inp[0]) ? node26230 : node26227;
											assign node26227 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node26230 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node26233 = (inp[2]) ? node26263 : node26234;
											assign node26234 = (inp[15]) ? node26256 : node26235;
												assign node26235 = (inp[9]) ? node26243 : node26236;
													assign node26236 = (inp[0]) ? node26240 : node26237;
														assign node26237 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node26240 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node26243 = (inp[10]) ? node26249 : node26244;
														assign node26244 = (inp[12]) ? node26246 : 4'b0100;
															assign node26246 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node26249 = (inp[0]) ? node26253 : node26250;
															assign node26250 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node26253 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node26256 = (inp[0]) ? node26260 : node26257;
													assign node26257 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node26260 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node26263 = (inp[15]) ? node26271 : node26264;
												assign node26264 = (inp[12]) ? node26268 : node26265;
													assign node26265 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node26268 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node26271 = (inp[11]) ? node26281 : node26272;
													assign node26272 = (inp[9]) ? 4'b0100 : node26273;
														assign node26273 = (inp[0]) ? node26277 : node26274;
															assign node26274 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node26277 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node26281 = (inp[9]) ? node26285 : node26282;
														assign node26282 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node26285 = (inp[0]) ? node26289 : node26286;
															assign node26286 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node26289 = (inp[12]) ? 4'b0100 : 4'b0101;
									assign node26292 = (inp[11]) ? node26300 : node26293;
										assign node26293 = (inp[0]) ? node26297 : node26294;
											assign node26294 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node26297 = (inp[12]) ? 4'b0100 : 4'b0101;
										assign node26300 = (inp[5]) ? node26338 : node26301;
											assign node26301 = (inp[2]) ? node26331 : node26302;
												assign node26302 = (inp[10]) ? node26316 : node26303;
													assign node26303 = (inp[15]) ? node26309 : node26304;
														assign node26304 = (inp[12]) ? node26306 : 4'b0101;
															assign node26306 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node26309 = (inp[12]) ? node26313 : node26310;
															assign node26310 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node26313 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node26316 = (inp[9]) ? node26324 : node26317;
														assign node26317 = (inp[12]) ? node26321 : node26318;
															assign node26318 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node26321 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node26324 = (inp[0]) ? node26328 : node26325;
															assign node26325 = (inp[12]) ? 4'b0101 : 4'b0100;
															assign node26328 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node26331 = (inp[0]) ? node26335 : node26332;
													assign node26332 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node26335 = (inp[12]) ? 4'b0100 : 4'b0101;
											assign node26338 = (inp[15]) ? node26346 : node26339;
												assign node26339 = (inp[0]) ? node26343 : node26340;
													assign node26340 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node26343 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node26346 = (inp[9]) ? node26354 : node26347;
													assign node26347 = (inp[0]) ? node26351 : node26348;
														assign node26348 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node26351 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node26354 = (inp[12]) ? node26358 : node26355;
														assign node26355 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node26358 = (inp[0]) ? 4'b0100 : 4'b0101;
							assign node26361 = (inp[13]) ? node26493 : node26362;
								assign node26362 = (inp[8]) ? node26446 : node26363;
									assign node26363 = (inp[12]) ? node26371 : node26364;
										assign node26364 = (inp[15]) ? node26368 : node26365;
											assign node26365 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node26368 = (inp[9]) ? 4'b0100 : 4'b0101;
										assign node26371 = (inp[5]) ? node26417 : node26372;
											assign node26372 = (inp[11]) ? node26394 : node26373;
												assign node26373 = (inp[0]) ? node26387 : node26374;
													assign node26374 = (inp[2]) ? node26382 : node26375;
														assign node26375 = (inp[9]) ? node26379 : node26376;
															assign node26376 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node26379 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node26382 = (inp[9]) ? 4'b0100 : node26383;
															assign node26383 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node26387 = (inp[10]) ? 4'b0100 : node26388;
														assign node26388 = (inp[9]) ? node26390 : 4'b0100;
															assign node26390 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node26394 = (inp[10]) ? node26402 : node26395;
													assign node26395 = (inp[15]) ? node26399 : node26396;
														assign node26396 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node26399 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node26402 = (inp[2]) ? node26410 : node26403;
														assign node26403 = (inp[15]) ? node26407 : node26404;
															assign node26404 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node26407 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node26410 = (inp[9]) ? node26414 : node26411;
															assign node26411 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node26414 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node26417 = (inp[0]) ? node26425 : node26418;
												assign node26418 = (inp[9]) ? node26422 : node26419;
													assign node26419 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node26422 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node26425 = (inp[2]) ? node26431 : node26426;
													assign node26426 = (inp[15]) ? node26428 : 4'b0101;
														assign node26428 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node26431 = (inp[10]) ? node26437 : node26432;
														assign node26432 = (inp[15]) ? node26434 : 4'b0100;
															assign node26434 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node26437 = (inp[11]) ? 4'b0101 : node26438;
															assign node26438 = (inp[9]) ? node26442 : node26439;
																assign node26439 = (inp[15]) ? 4'b0101 : 4'b0100;
																assign node26442 = (inp[15]) ? 4'b0100 : 4'b0101;
									assign node26446 = (inp[12]) ? node26478 : node26447;
										assign node26447 = (inp[2]) ? node26455 : node26448;
											assign node26448 = (inp[0]) ? node26452 : node26449;
												assign node26449 = (inp[15]) ? 4'b0001 : 4'b0000;
												assign node26452 = (inp[15]) ? 4'b0000 : 4'b0001;
											assign node26455 = (inp[11]) ? node26463 : node26456;
												assign node26456 = (inp[15]) ? node26460 : node26457;
													assign node26457 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node26460 = (inp[0]) ? 4'b0000 : 4'b0001;
												assign node26463 = (inp[5]) ? node26471 : node26464;
													assign node26464 = (inp[15]) ? node26468 : node26465;
														assign node26465 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node26468 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node26471 = (inp[0]) ? node26475 : node26472;
														assign node26472 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node26475 = (inp[15]) ? 4'b0000 : 4'b0001;
										assign node26478 = (inp[2]) ? node26486 : node26479;
											assign node26479 = (inp[15]) ? node26483 : node26480;
												assign node26480 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node26483 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node26486 = (inp[15]) ? node26490 : node26487;
												assign node26487 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node26490 = (inp[0]) ? 4'b0000 : 4'b0001;
								assign node26493 = (inp[0]) ? node26499 : node26494;
									assign node26494 = (inp[9]) ? 4'b0001 : node26495;
										assign node26495 = (inp[8]) ? 4'b0001 : 4'b0000;
									assign node26499 = (inp[9]) ? 4'b0000 : node26500;
										assign node26500 = (inp[8]) ? 4'b0000 : 4'b0001;
		assign node26504 = (inp[8]) ? node40938 : node26505;
			assign node26505 = (inp[14]) ? node34509 : node26506;
				assign node26506 = (inp[5]) ? node30520 : node26507;
					assign node26507 = (inp[13]) ? node28431 : node26508;
						assign node26508 = (inp[6]) ? node27668 : node26509;
							assign node26509 = (inp[1]) ? node27087 : node26510;
								assign node26510 = (inp[2]) ? node26790 : node26511;
									assign node26511 = (inp[4]) ? node26659 : node26512;
										assign node26512 = (inp[7]) ? node26582 : node26513;
											assign node26513 = (inp[12]) ? node26545 : node26514;
												assign node26514 = (inp[15]) ? node26536 : node26515;
													assign node26515 = (inp[0]) ? node26521 : node26516;
														assign node26516 = (inp[10]) ? 4'b1000 : node26517;
															assign node26517 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node26521 = (inp[9]) ? node26529 : node26522;
															assign node26522 = (inp[10]) ? node26526 : node26523;
																assign node26523 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node26526 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node26529 = (inp[11]) ? node26533 : node26530;
																assign node26530 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node26533 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node26536 = (inp[0]) ? 4'b1001 : node26537;
														assign node26537 = (inp[9]) ? node26541 : node26538;
															assign node26538 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node26541 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node26545 = (inp[0]) ? node26567 : node26546;
													assign node26546 = (inp[15]) ? node26554 : node26547;
														assign node26547 = (inp[9]) ? node26551 : node26548;
															assign node26548 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node26551 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node26554 = (inp[11]) ? node26562 : node26555;
															assign node26555 = (inp[10]) ? node26559 : node26556;
																assign node26556 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node26559 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node26562 = (inp[10]) ? 4'b1011 : node26563;
																assign node26563 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node26567 = (inp[9]) ? node26575 : node26568;
														assign node26568 = (inp[11]) ? node26572 : node26569;
															assign node26569 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node26572 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node26575 = (inp[10]) ? node26579 : node26576;
															assign node26576 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node26579 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node26582 = (inp[12]) ? node26626 : node26583;
												assign node26583 = (inp[15]) ? node26607 : node26584;
													assign node26584 = (inp[11]) ? node26600 : node26585;
														assign node26585 = (inp[0]) ? node26593 : node26586;
															assign node26586 = (inp[9]) ? node26590 : node26587;
																assign node26587 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node26590 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node26593 = (inp[10]) ? node26597 : node26594;
																assign node26594 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node26597 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node26600 = (inp[9]) ? node26604 : node26601;
															assign node26601 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node26604 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node26607 = (inp[0]) ? node26613 : node26608;
														assign node26608 = (inp[10]) ? 4'b1111 : node26609;
															assign node26609 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node26613 = (inp[11]) ? node26619 : node26614;
															assign node26614 = (inp[9]) ? 4'b1110 : node26615;
																assign node26615 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node26619 = (inp[10]) ? node26623 : node26620;
																assign node26620 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node26623 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node26626 = (inp[15]) ? node26644 : node26627;
													assign node26627 = (inp[0]) ? node26637 : node26628;
														assign node26628 = (inp[11]) ? node26630 : 4'b1100;
															assign node26630 = (inp[10]) ? node26634 : node26631;
																assign node26631 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node26634 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node26637 = (inp[11]) ? 4'b1100 : node26638;
															assign node26638 = (inp[9]) ? node26640 : 4'b1101;
																assign node26640 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node26644 = (inp[9]) ? node26650 : node26645;
														assign node26645 = (inp[10]) ? 4'b1000 : node26646;
															assign node26646 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node26650 = (inp[10]) ? node26654 : node26651;
															assign node26651 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node26654 = (inp[11]) ? 4'b1001 : node26655;
																assign node26655 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node26659 = (inp[7]) ? node26723 : node26660;
											assign node26660 = (inp[0]) ? node26688 : node26661;
												assign node26661 = (inp[10]) ? node26679 : node26662;
													assign node26662 = (inp[9]) ? node26670 : node26663;
														assign node26663 = (inp[12]) ? node26667 : node26664;
															assign node26664 = (inp[15]) ? 4'b1100 : 4'b1010;
															assign node26667 = (inp[15]) ? 4'b1010 : 4'b1100;
														assign node26670 = (inp[12]) ? node26674 : node26671;
															assign node26671 = (inp[15]) ? 4'b1101 : 4'b1011;
															assign node26674 = (inp[15]) ? node26676 : 4'b1101;
																assign node26676 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node26679 = (inp[9]) ? 4'b1100 : node26680;
														assign node26680 = (inp[12]) ? node26682 : 4'b1101;
															assign node26682 = (inp[15]) ? node26684 : 4'b1101;
																assign node26684 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node26688 = (inp[12]) ? node26712 : node26689;
													assign node26689 = (inp[15]) ? node26703 : node26690;
														assign node26690 = (inp[10]) ? node26696 : node26691;
															assign node26691 = (inp[11]) ? 4'b1010 : node26692;
																assign node26692 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node26696 = (inp[9]) ? node26700 : node26697;
																assign node26697 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node26700 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node26703 = (inp[11]) ? node26705 : 4'b1100;
															assign node26705 = (inp[9]) ? node26709 : node26706;
																assign node26706 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node26709 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node26712 = (inp[15]) ? 4'b1011 : node26713;
														assign node26713 = (inp[11]) ? 4'b1101 : node26714;
															assign node26714 = (inp[10]) ? node26718 : node26715;
																assign node26715 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node26718 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node26723 = (inp[15]) ? node26759 : node26724;
												assign node26724 = (inp[12]) ? node26744 : node26725;
													assign node26725 = (inp[10]) ? node26733 : node26726;
														assign node26726 = (inp[9]) ? node26728 : 4'b1100;
															assign node26728 = (inp[11]) ? 4'b1101 : node26729;
																assign node26729 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node26733 = (inp[9]) ? node26739 : node26734;
															assign node26734 = (inp[11]) ? 4'b1101 : node26735;
																assign node26735 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node26739 = (inp[0]) ? node26741 : 4'b1100;
																assign node26741 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node26744 = (inp[10]) ? node26750 : node26745;
														assign node26745 = (inp[9]) ? 4'b1010 : node26746;
															assign node26746 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node26750 = (inp[11]) ? 4'b1010 : node26751;
															assign node26751 = (inp[0]) ? node26755 : node26752;
																assign node26752 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node26755 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node26759 = (inp[12]) ? node26775 : node26760;
													assign node26760 = (inp[0]) ? node26770 : node26761;
														assign node26761 = (inp[11]) ? 4'b1011 : node26762;
															assign node26762 = (inp[9]) ? node26766 : node26763;
																assign node26763 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node26766 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node26770 = (inp[9]) ? 4'b1010 : node26771;
															assign node26771 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node26775 = (inp[0]) ? node26783 : node26776;
														assign node26776 = (inp[11]) ? node26778 : 4'b1001;
															assign node26778 = (inp[10]) ? node26780 : 4'b1001;
																assign node26780 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node26783 = (inp[10]) ? node26787 : node26784;
															assign node26784 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node26787 = (inp[9]) ? 4'b1001 : 4'b1000;
									assign node26790 = (inp[15]) ? node26964 : node26791;
										assign node26791 = (inp[4]) ? node26865 : node26792;
											assign node26792 = (inp[7]) ? node26832 : node26793;
												assign node26793 = (inp[12]) ? node26811 : node26794;
													assign node26794 = (inp[0]) ? node26802 : node26795;
														assign node26795 = (inp[9]) ? node26799 : node26796;
															assign node26796 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node26799 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node26802 = (inp[9]) ? 4'b1101 : node26803;
															assign node26803 = (inp[11]) ? node26807 : node26804;
																assign node26804 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node26807 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node26811 = (inp[10]) ? node26821 : node26812;
														assign node26812 = (inp[0]) ? node26814 : 4'b1111;
															assign node26814 = (inp[11]) ? node26818 : node26815;
																assign node26815 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node26818 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node26821 = (inp[9]) ? node26827 : node26822;
															assign node26822 = (inp[0]) ? node26824 : 4'b1111;
																assign node26824 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node26827 = (inp[11]) ? 4'b1110 : node26828;
																assign node26828 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node26832 = (inp[12]) ? node26848 : node26833;
													assign node26833 = (inp[10]) ? node26843 : node26834;
														assign node26834 = (inp[9]) ? node26838 : node26835;
															assign node26835 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node26838 = (inp[0]) ? node26840 : 4'b1111;
																assign node26840 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node26843 = (inp[0]) ? 4'b1110 : node26844;
															assign node26844 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node26848 = (inp[10]) ? node26854 : node26849;
														assign node26849 = (inp[9]) ? node26851 : 4'b1001;
															assign node26851 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node26854 = (inp[9]) ? node26860 : node26855;
															assign node26855 = (inp[0]) ? node26857 : 4'b1000;
																assign node26857 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node26860 = (inp[11]) ? 4'b1001 : node26861;
																assign node26861 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node26865 = (inp[11]) ? node26919 : node26866;
												assign node26866 = (inp[0]) ? node26892 : node26867;
													assign node26867 = (inp[7]) ? node26883 : node26868;
														assign node26868 = (inp[12]) ? node26876 : node26869;
															assign node26869 = (inp[10]) ? node26873 : node26870;
																assign node26870 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node26873 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node26876 = (inp[9]) ? node26880 : node26877;
																assign node26877 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node26880 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node26883 = (inp[12]) ? node26885 : 4'b1000;
															assign node26885 = (inp[10]) ? node26889 : node26886;
																assign node26886 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node26889 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node26892 = (inp[10]) ? node26906 : node26893;
														assign node26893 = (inp[9]) ? node26899 : node26894;
															assign node26894 = (inp[12]) ? node26896 : 4'b1001;
																assign node26896 = (inp[7]) ? 4'b1111 : 4'b1001;
															assign node26899 = (inp[12]) ? node26903 : node26900;
																assign node26900 = (inp[7]) ? 4'b1000 : 4'b1111;
																assign node26903 = (inp[7]) ? 4'b1110 : 4'b1000;
														assign node26906 = (inp[9]) ? node26912 : node26907;
															assign node26907 = (inp[7]) ? node26909 : 4'b1111;
																assign node26909 = (inp[12]) ? 4'b1110 : 4'b1000;
															assign node26912 = (inp[12]) ? node26916 : node26913;
																assign node26913 = (inp[7]) ? 4'b1001 : 4'b1110;
																assign node26916 = (inp[7]) ? 4'b1111 : 4'b1001;
												assign node26919 = (inp[0]) ? node26941 : node26920;
													assign node26920 = (inp[10]) ? node26928 : node26921;
														assign node26921 = (inp[9]) ? 4'b1001 : node26922;
															assign node26922 = (inp[7]) ? 4'b1000 : node26923;
																assign node26923 = (inp[12]) ? 4'b1000 : 4'b1111;
														assign node26928 = (inp[9]) ? node26934 : node26929;
															assign node26929 = (inp[12]) ? node26931 : 4'b1001;
																assign node26931 = (inp[7]) ? 4'b1111 : 4'b1001;
															assign node26934 = (inp[12]) ? node26938 : node26935;
																assign node26935 = (inp[7]) ? 4'b1000 : 4'b1111;
																assign node26938 = (inp[7]) ? 4'b1110 : 4'b1000;
													assign node26941 = (inp[9]) ? node26955 : node26942;
														assign node26942 = (inp[10]) ? node26950 : node26943;
															assign node26943 = (inp[12]) ? node26947 : node26944;
																assign node26944 = (inp[7]) ? 4'b1001 : 4'b1111;
																assign node26947 = (inp[7]) ? 4'b1110 : 4'b1001;
															assign node26950 = (inp[7]) ? 4'b1111 : node26951;
																assign node26951 = (inp[12]) ? 4'b1000 : 4'b1110;
														assign node26955 = (inp[10]) ? node26959 : node26956;
															assign node26956 = (inp[7]) ? 4'b1111 : 4'b1000;
															assign node26959 = (inp[12]) ? 4'b1001 : node26960;
																assign node26960 = (inp[7]) ? 4'b1001 : 4'b1111;
										assign node26964 = (inp[12]) ? node27014 : node26965;
											assign node26965 = (inp[7]) ? node26989 : node26966;
												assign node26966 = (inp[4]) ? node26976 : node26967;
													assign node26967 = (inp[10]) ? node26969 : 4'b1101;
														assign node26969 = (inp[9]) ? 4'b1100 : node26970;
															assign node26970 = (inp[0]) ? node26972 : 4'b1101;
																assign node26972 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node26976 = (inp[11]) ? node26982 : node26977;
														assign node26977 = (inp[10]) ? 4'b1000 : node26978;
															assign node26978 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node26982 = (inp[9]) ? node26986 : node26983;
															assign node26983 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node26986 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node26989 = (inp[4]) ? node27001 : node26990;
													assign node26990 = (inp[11]) ? node26994 : node26991;
														assign node26991 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node26994 = (inp[10]) ? node26996 : 4'b1010;
															assign node26996 = (inp[9]) ? node26998 : 4'b1011;
																assign node26998 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node27001 = (inp[10]) ? node27007 : node27002;
														assign node27002 = (inp[9]) ? node27004 : 4'b1111;
															assign node27004 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node27007 = (inp[9]) ? 4'b1111 : node27008;
															assign node27008 = (inp[11]) ? node27010 : 4'b1110;
																assign node27010 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node27014 = (inp[7]) ? node27050 : node27015;
												assign node27015 = (inp[11]) ? node27031 : node27016;
													assign node27016 = (inp[0]) ? node27024 : node27017;
														assign node27017 = (inp[10]) ? node27019 : 4'b1111;
															assign node27019 = (inp[9]) ? node27021 : 4'b1111;
																assign node27021 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node27024 = (inp[9]) ? node27028 : node27025;
															assign node27025 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node27028 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node27031 = (inp[9]) ? node27043 : node27032;
														assign node27032 = (inp[10]) ? node27038 : node27033;
															assign node27033 = (inp[4]) ? node27035 : 4'b1110;
																assign node27035 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node27038 = (inp[4]) ? node27040 : 4'b1111;
																assign node27040 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node27043 = (inp[10]) ? node27045 : 4'b1111;
															assign node27045 = (inp[0]) ? node27047 : 4'b1110;
																assign node27047 = (inp[4]) ? 4'b1111 : 4'b1110;
												assign node27050 = (inp[9]) ? node27066 : node27051;
													assign node27051 = (inp[4]) ? node27057 : node27052;
														assign node27052 = (inp[10]) ? node27054 : 4'b1101;
															assign node27054 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node27057 = (inp[10]) ? node27061 : node27058;
															assign node27058 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node27061 = (inp[11]) ? node27063 : 4'b1101;
																assign node27063 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node27066 = (inp[4]) ? node27078 : node27067;
														assign node27067 = (inp[10]) ? node27073 : node27068;
															assign node27068 = (inp[11]) ? 4'b1100 : node27069;
																assign node27069 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node27073 = (inp[0]) ? node27075 : 4'b1101;
																assign node27075 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node27078 = (inp[10]) ? node27084 : node27079;
															assign node27079 = (inp[11]) ? node27081 : 4'b1101;
																assign node27081 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node27084 = (inp[0]) ? 4'b1100 : 4'b1101;
								assign node27087 = (inp[2]) ? node27373 : node27088;
									assign node27088 = (inp[7]) ? node27230 : node27089;
										assign node27089 = (inp[12]) ? node27151 : node27090;
											assign node27090 = (inp[4]) ? node27118 : node27091;
												assign node27091 = (inp[10]) ? node27111 : node27092;
													assign node27092 = (inp[9]) ? node27102 : node27093;
														assign node27093 = (inp[11]) ? node27099 : node27094;
															assign node27094 = (inp[0]) ? node27096 : 4'b1100;
																assign node27096 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node27099 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node27102 = (inp[0]) ? node27108 : node27103;
															assign node27103 = (inp[15]) ? node27105 : 4'b1101;
																assign node27105 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node27108 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node27111 = (inp[9]) ? 4'b1100 : node27112;
														assign node27112 = (inp[0]) ? node27114 : 4'b1101;
															assign node27114 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node27118 = (inp[15]) ? node27134 : node27119;
													assign node27119 = (inp[9]) ? node27125 : node27120;
														assign node27120 = (inp[10]) ? node27122 : 4'b1110;
															assign node27122 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node27125 = (inp[10]) ? node27131 : node27126;
															assign node27126 = (inp[11]) ? 4'b1111 : node27127;
																assign node27127 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node27131 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node27134 = (inp[10]) ? node27144 : node27135;
														assign node27135 = (inp[9]) ? node27141 : node27136;
															assign node27136 = (inp[11]) ? 4'b1001 : node27137;
																assign node27137 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node27141 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node27144 = (inp[0]) ? node27146 : 4'b1000;
															assign node27146 = (inp[9]) ? 4'b1000 : node27147;
																assign node27147 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node27151 = (inp[4]) ? node27185 : node27152;
												assign node27152 = (inp[0]) ? node27168 : node27153;
													assign node27153 = (inp[10]) ? node27163 : node27154;
														assign node27154 = (inp[9]) ? node27160 : node27155;
															assign node27155 = (inp[11]) ? node27157 : 4'b1111;
																assign node27157 = (inp[15]) ? 4'b1110 : 4'b1111;
															assign node27160 = (inp[15]) ? 4'b1111 : 4'b1110;
														assign node27163 = (inp[9]) ? 4'b1111 : node27164;
															assign node27164 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node27168 = (inp[11]) ? node27180 : node27169;
														assign node27169 = (inp[10]) ? node27175 : node27170;
															assign node27170 = (inp[9]) ? 4'b1111 : node27171;
																assign node27171 = (inp[15]) ? 4'b1111 : 4'b1110;
															assign node27175 = (inp[15]) ? 4'b1110 : node27176;
																assign node27176 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node27180 = (inp[9]) ? 4'b1110 : node27181;
															assign node27181 = (inp[10]) ? 4'b1110 : 4'b1111;
												assign node27185 = (inp[15]) ? node27215 : node27186;
													assign node27186 = (inp[0]) ? node27202 : node27187;
														assign node27187 = (inp[9]) ? node27195 : node27188;
															assign node27188 = (inp[10]) ? node27192 : node27189;
																assign node27189 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node27192 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node27195 = (inp[11]) ? node27199 : node27196;
																assign node27196 = (inp[10]) ? 4'b1101 : 4'b1100;
																assign node27199 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node27202 = (inp[11]) ? node27210 : node27203;
															assign node27203 = (inp[9]) ? node27207 : node27204;
																assign node27204 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node27207 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node27210 = (inp[9]) ? node27212 : 4'b1100;
																assign node27212 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node27215 = (inp[0]) ? node27221 : node27216;
														assign node27216 = (inp[9]) ? node27218 : 4'b1111;
															assign node27218 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node27221 = (inp[11]) ? 4'b1110 : node27222;
															assign node27222 = (inp[10]) ? node27226 : node27223;
																assign node27223 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node27226 = (inp[9]) ? 4'b1111 : 4'b1110;
										assign node27230 = (inp[12]) ? node27312 : node27231;
											assign node27231 = (inp[4]) ? node27275 : node27232;
												assign node27232 = (inp[15]) ? node27252 : node27233;
													assign node27233 = (inp[11]) ? node27245 : node27234;
														assign node27234 = (inp[0]) ? node27240 : node27235;
															assign node27235 = (inp[9]) ? 4'b1011 : node27236;
																assign node27236 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node27240 = (inp[10]) ? node27242 : 4'b1010;
																assign node27242 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node27245 = (inp[10]) ? 4'b1010 : node27246;
															assign node27246 = (inp[0]) ? 4'b1010 : node27247;
																assign node27247 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node27252 = (inp[0]) ? node27260 : node27253;
														assign node27253 = (inp[10]) ? node27257 : node27254;
															assign node27254 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node27257 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node27260 = (inp[10]) ? node27268 : node27261;
															assign node27261 = (inp[9]) ? node27265 : node27262;
																assign node27262 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node27265 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node27268 = (inp[9]) ? node27272 : node27269;
																assign node27269 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node27272 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node27275 = (inp[15]) ? node27293 : node27276;
													assign node27276 = (inp[9]) ? node27284 : node27277;
														assign node27277 = (inp[11]) ? node27281 : node27278;
															assign node27278 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node27281 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node27284 = (inp[10]) ? node27288 : node27285;
															assign node27285 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node27288 = (inp[0]) ? 4'b1000 : node27289;
																assign node27289 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node27293 = (inp[10]) ? node27303 : node27294;
														assign node27294 = (inp[9]) ? node27300 : node27295;
															assign node27295 = (inp[0]) ? 4'b1011 : node27296;
																assign node27296 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node27300 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node27303 = (inp[9]) ? node27309 : node27304;
															assign node27304 = (inp[11]) ? node27306 : 4'b1010;
																assign node27306 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node27309 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node27312 = (inp[4]) ? node27338 : node27313;
												assign node27313 = (inp[15]) ? node27329 : node27314;
													assign node27314 = (inp[0]) ? node27320 : node27315;
														assign node27315 = (inp[9]) ? node27317 : 4'b1000;
															assign node27317 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node27320 = (inp[9]) ? 4'b1001 : node27321;
															assign node27321 = (inp[10]) ? node27325 : node27322;
																assign node27322 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node27325 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node27329 = (inp[0]) ? 4'b1100 : node27330;
														assign node27330 = (inp[11]) ? 4'b1101 : node27331;
															assign node27331 = (inp[9]) ? node27333 : 4'b1100;
																assign node27333 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node27338 = (inp[15]) ? node27360 : node27339;
													assign node27339 = (inp[11]) ? node27355 : node27340;
														assign node27340 = (inp[0]) ? node27348 : node27341;
															assign node27341 = (inp[10]) ? node27345 : node27342;
																assign node27342 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node27345 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node27348 = (inp[9]) ? node27352 : node27349;
																assign node27349 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node27352 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node27355 = (inp[10]) ? node27357 : 4'b1111;
															assign node27357 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node27360 = (inp[9]) ? node27366 : node27361;
														assign node27361 = (inp[10]) ? node27363 : 4'b1101;
															assign node27363 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node27366 = (inp[10]) ? node27368 : 4'b1100;
															assign node27368 = (inp[0]) ? node27370 : 4'b1101;
																assign node27370 = (inp[11]) ? 4'b1101 : 4'b1100;
									assign node27373 = (inp[7]) ? node27509 : node27374;
										assign node27374 = (inp[12]) ? node27440 : node27375;
											assign node27375 = (inp[4]) ? node27409 : node27376;
												assign node27376 = (inp[15]) ? node27392 : node27377;
													assign node27377 = (inp[11]) ? node27385 : node27378;
														assign node27378 = (inp[10]) ? node27382 : node27379;
															assign node27379 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node27382 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node27385 = (inp[0]) ? node27387 : 4'b1001;
															assign node27387 = (inp[9]) ? node27389 : 4'b1001;
																assign node27389 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node27392 = (inp[10]) ? node27398 : node27393;
														assign node27393 = (inp[9]) ? 4'b1000 : node27394;
															assign node27394 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node27398 = (inp[9]) ? node27404 : node27399;
															assign node27399 = (inp[11]) ? 4'b1000 : node27400;
																assign node27400 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node27404 = (inp[11]) ? 4'b1001 : node27405;
																assign node27405 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node27409 = (inp[15]) ? node27423 : node27410;
													assign node27410 = (inp[10]) ? node27418 : node27411;
														assign node27411 = (inp[9]) ? node27415 : node27412;
															assign node27412 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node27415 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node27418 = (inp[9]) ? node27420 : 4'b1010;
															assign node27420 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node27423 = (inp[9]) ? node27429 : node27424;
														assign node27424 = (inp[10]) ? 4'b1101 : node27425;
															assign node27425 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node27429 = (inp[10]) ? node27435 : node27430;
															assign node27430 = (inp[11]) ? 4'b1101 : node27431;
																assign node27431 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node27435 = (inp[0]) ? node27437 : 4'b1100;
																assign node27437 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node27440 = (inp[4]) ? node27476 : node27441;
												assign node27441 = (inp[9]) ? node27461 : node27442;
													assign node27442 = (inp[0]) ? node27452 : node27443;
														assign node27443 = (inp[10]) ? node27449 : node27444;
															assign node27444 = (inp[11]) ? 4'b1010 : node27445;
																assign node27445 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node27449 = (inp[15]) ? 4'b1011 : 4'b1010;
														assign node27452 = (inp[15]) ? node27454 : 4'b1011;
															assign node27454 = (inp[10]) ? node27458 : node27455;
																assign node27455 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node27458 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node27461 = (inp[0]) ? node27467 : node27462;
														assign node27462 = (inp[11]) ? node27464 : 4'b1010;
															assign node27464 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node27467 = (inp[10]) ? node27473 : node27468;
															assign node27468 = (inp[15]) ? node27470 : 4'b1010;
																assign node27470 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node27473 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node27476 = (inp[15]) ? node27498 : node27477;
													assign node27477 = (inp[0]) ? node27485 : node27478;
														assign node27478 = (inp[10]) ? node27482 : node27479;
															assign node27479 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node27482 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node27485 = (inp[9]) ? node27493 : node27486;
															assign node27486 = (inp[11]) ? node27490 : node27487;
																assign node27487 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node27490 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node27493 = (inp[11]) ? 4'b1001 : node27494;
																assign node27494 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node27498 = (inp[11]) ? node27506 : node27499;
														assign node27499 = (inp[9]) ? node27503 : node27500;
															assign node27500 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node27503 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node27506 = (inp[0]) ? 4'b1011 : 4'b1010;
										assign node27509 = (inp[12]) ? node27599 : node27510;
											assign node27510 = (inp[4]) ? node27560 : node27511;
												assign node27511 = (inp[15]) ? node27533 : node27512;
													assign node27512 = (inp[10]) ? node27522 : node27513;
														assign node27513 = (inp[9]) ? node27519 : node27514;
															assign node27514 = (inp[0]) ? 4'b1110 : node27515;
																assign node27515 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node27519 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node27522 = (inp[9]) ? node27528 : node27523;
															assign node27523 = (inp[0]) ? 4'b1111 : node27524;
																assign node27524 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node27528 = (inp[11]) ? node27530 : 4'b1110;
																assign node27530 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node27533 = (inp[11]) ? node27547 : node27534;
														assign node27534 = (inp[0]) ? node27540 : node27535;
															assign node27535 = (inp[9]) ? node27537 : 4'b1010;
																assign node27537 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node27540 = (inp[10]) ? node27544 : node27541;
																assign node27541 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node27544 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node27547 = (inp[10]) ? node27553 : node27548;
															assign node27548 = (inp[0]) ? node27550 : 4'b1011;
																assign node27550 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node27553 = (inp[0]) ? node27557 : node27554;
																assign node27554 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node27557 = (inp[9]) ? 4'b1011 : 4'b1010;
												assign node27560 = (inp[15]) ? node27584 : node27561;
													assign node27561 = (inp[10]) ? node27573 : node27562;
														assign node27562 = (inp[9]) ? node27568 : node27563;
															assign node27563 = (inp[0]) ? 4'b1101 : node27564;
																assign node27564 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node27568 = (inp[0]) ? 4'b1100 : node27569;
																assign node27569 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node27573 = (inp[9]) ? node27579 : node27574;
															assign node27574 = (inp[0]) ? 4'b1100 : node27575;
																assign node27575 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node27579 = (inp[0]) ? 4'b1101 : node27580;
																assign node27580 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node27584 = (inp[9]) ? node27590 : node27585;
														assign node27585 = (inp[11]) ? node27587 : 4'b1110;
															assign node27587 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node27590 = (inp[0]) ? node27596 : node27591;
															assign node27591 = (inp[11]) ? node27593 : 4'b1111;
																assign node27593 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node27596 = (inp[10]) ? 4'b1110 : 4'b1111;
											assign node27599 = (inp[4]) ? node27629 : node27600;
												assign node27600 = (inp[15]) ? node27618 : node27601;
													assign node27601 = (inp[10]) ? node27613 : node27602;
														assign node27602 = (inp[9]) ? node27608 : node27603;
															assign node27603 = (inp[0]) ? node27605 : 4'b1100;
																assign node27605 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node27608 = (inp[11]) ? 4'b1101 : node27609;
																assign node27609 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node27613 = (inp[9]) ? 4'b1100 : node27614;
															assign node27614 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node27618 = (inp[9]) ? node27620 : 4'b1001;
														assign node27620 = (inp[0]) ? node27624 : node27621;
															assign node27621 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node27624 = (inp[11]) ? 4'b1001 : node27625;
																assign node27625 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node27629 = (inp[15]) ? node27651 : node27630;
													assign node27630 = (inp[10]) ? node27642 : node27631;
														assign node27631 = (inp[9]) ? node27637 : node27632;
															assign node27632 = (inp[0]) ? 4'b1011 : node27633;
																assign node27633 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node27637 = (inp[11]) ? node27639 : 4'b1010;
																assign node27639 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node27642 = (inp[9]) ? node27648 : node27643;
															assign node27643 = (inp[0]) ? 4'b1010 : node27644;
																assign node27644 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node27648 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node27651 = (inp[9]) ? node27657 : node27652;
														assign node27652 = (inp[10]) ? node27654 : 4'b1000;
															assign node27654 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node27657 = (inp[10]) ? node27663 : node27658;
															assign node27658 = (inp[11]) ? node27660 : 4'b1001;
																assign node27660 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node27663 = (inp[0]) ? 4'b1000 : node27664;
																assign node27664 = (inp[11]) ? 4'b1001 : 4'b1000;
							assign node27668 = (inp[12]) ? node28100 : node27669;
								assign node27669 = (inp[15]) ? node27911 : node27670;
									assign node27670 = (inp[7]) ? node27786 : node27671;
										assign node27671 = (inp[1]) ? node27725 : node27672;
											assign node27672 = (inp[10]) ? node27702 : node27673;
												assign node27673 = (inp[9]) ? node27685 : node27674;
													assign node27674 = (inp[4]) ? 4'b1000 : node27675;
														assign node27675 = (inp[11]) ? node27681 : node27676;
															assign node27676 = (inp[2]) ? 4'b1000 : node27677;
																assign node27677 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node27681 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node27685 = (inp[2]) ? node27693 : node27686;
														assign node27686 = (inp[11]) ? node27690 : node27687;
															assign node27687 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node27690 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node27693 = (inp[0]) ? node27697 : node27694;
															assign node27694 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node27697 = (inp[11]) ? node27699 : 4'b1000;
																assign node27699 = (inp[4]) ? 4'b1001 : 4'b1000;
												assign node27702 = (inp[2]) ? node27714 : node27703;
													assign node27703 = (inp[4]) ? 4'b1001 : node27704;
														assign node27704 = (inp[0]) ? node27706 : 4'b1001;
															assign node27706 = (inp[9]) ? node27710 : node27707;
																assign node27707 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node27710 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node27714 = (inp[9]) ? node27720 : node27715;
														assign node27715 = (inp[11]) ? node27717 : 4'b1001;
															assign node27717 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node27720 = (inp[11]) ? node27722 : 4'b1000;
															assign node27722 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node27725 = (inp[4]) ? node27749 : node27726;
												assign node27726 = (inp[9]) ? node27738 : node27727;
													assign node27727 = (inp[11]) ? node27733 : node27728;
														assign node27728 = (inp[2]) ? 4'b1100 : node27729;
															assign node27729 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node27733 = (inp[0]) ? node27735 : 4'b1101;
															assign node27735 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node27738 = (inp[11]) ? node27744 : node27739;
														assign node27739 = (inp[0]) ? node27741 : 4'b1101;
															assign node27741 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node27744 = (inp[0]) ? node27746 : 4'b1100;
															assign node27746 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node27749 = (inp[10]) ? node27767 : node27750;
													assign node27750 = (inp[11]) ? node27760 : node27751;
														assign node27751 = (inp[0]) ? node27755 : node27752;
															assign node27752 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node27755 = (inp[2]) ? node27757 : 4'b1000;
																assign node27757 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node27760 = (inp[2]) ? node27762 : 4'b1000;
															assign node27762 = (inp[0]) ? node27764 : 4'b1000;
																assign node27764 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node27767 = (inp[9]) ? node27779 : node27768;
														assign node27768 = (inp[11]) ? node27774 : node27769;
															assign node27769 = (inp[2]) ? node27771 : 4'b1000;
																assign node27771 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node27774 = (inp[2]) ? node27776 : 4'b1001;
																assign node27776 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node27779 = (inp[11]) ? node27781 : 4'b1001;
															assign node27781 = (inp[0]) ? node27783 : 4'b1000;
																assign node27783 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node27786 = (inp[1]) ? node27834 : node27787;
											assign node27787 = (inp[4]) ? node27815 : node27788;
												assign node27788 = (inp[0]) ? node27802 : node27789;
													assign node27789 = (inp[2]) ? node27795 : node27790;
														assign node27790 = (inp[11]) ? node27792 : 4'b1011;
															assign node27792 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node27795 = (inp[11]) ? node27799 : node27796;
															assign node27796 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node27799 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node27802 = (inp[2]) ? node27810 : node27803;
														assign node27803 = (inp[11]) ? node27807 : node27804;
															assign node27804 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node27807 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node27810 = (inp[9]) ? 4'b1011 : node27811;
															assign node27811 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node27815 = (inp[9]) ? node27827 : node27816;
													assign node27816 = (inp[11]) ? node27822 : node27817;
														assign node27817 = (inp[2]) ? 4'b1111 : node27818;
															assign node27818 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node27822 = (inp[2]) ? 4'b1110 : node27823;
															assign node27823 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node27827 = (inp[11]) ? node27829 : 4'b1110;
														assign node27829 = (inp[0]) ? 4'b1111 : node27830;
															assign node27830 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node27834 = (inp[10]) ? node27876 : node27835;
												assign node27835 = (inp[0]) ? node27855 : node27836;
													assign node27836 = (inp[9]) ? node27846 : node27837;
														assign node27837 = (inp[2]) ? node27841 : node27838;
															assign node27838 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node27841 = (inp[4]) ? 4'b1011 : node27842;
																assign node27842 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node27846 = (inp[11]) ? node27852 : node27847;
															assign node27847 = (inp[4]) ? 4'b1011 : node27848;
																assign node27848 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node27852 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node27855 = (inp[9]) ? node27867 : node27856;
														assign node27856 = (inp[11]) ? node27862 : node27857;
															assign node27857 = (inp[2]) ? node27859 : 4'b1010;
																assign node27859 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node27862 = (inp[2]) ? node27864 : 4'b1011;
																assign node27864 = (inp[4]) ? 4'b1010 : 4'b1011;
														assign node27867 = (inp[2]) ? node27869 : 4'b1010;
															assign node27869 = (inp[11]) ? node27873 : node27870;
																assign node27870 = (inp[4]) ? 4'b1010 : 4'b1011;
																assign node27873 = (inp[4]) ? 4'b1011 : 4'b1010;
												assign node27876 = (inp[0]) ? node27894 : node27877;
													assign node27877 = (inp[9]) ? node27883 : node27878;
														assign node27878 = (inp[11]) ? node27880 : 4'b1010;
															assign node27880 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node27883 = (inp[11]) ? node27889 : node27884;
															assign node27884 = (inp[2]) ? node27886 : 4'b1011;
																assign node27886 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node27889 = (inp[2]) ? node27891 : 4'b1010;
																assign node27891 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node27894 = (inp[9]) ? node27906 : node27895;
														assign node27895 = (inp[11]) ? node27901 : node27896;
															assign node27896 = (inp[2]) ? node27898 : 4'b1010;
																assign node27898 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node27901 = (inp[4]) ? node27903 : 4'b1011;
																assign node27903 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node27906 = (inp[11]) ? 4'b1010 : node27907;
															assign node27907 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node27911 = (inp[7]) ? node28001 : node27912;
										assign node27912 = (inp[11]) ? node27954 : node27913;
											assign node27913 = (inp[9]) ? node27931 : node27914;
												assign node27914 = (inp[1]) ? node27924 : node27915;
													assign node27915 = (inp[4]) ? node27921 : node27916;
														assign node27916 = (inp[2]) ? 4'b1010 : node27917;
															assign node27917 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node27921 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node27924 = (inp[4]) ? 4'b1010 : node27925;
														assign node27925 = (inp[0]) ? 4'b1110 : node27926;
															assign node27926 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node27931 = (inp[1]) ? node27943 : node27932;
													assign node27932 = (inp[4]) ? node27938 : node27933;
														assign node27933 = (inp[2]) ? 4'b1011 : node27934;
															assign node27934 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node27938 = (inp[0]) ? 4'b1110 : node27939;
															assign node27939 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node27943 = (inp[4]) ? node27949 : node27944;
														assign node27944 = (inp[2]) ? node27946 : 4'b1111;
															assign node27946 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node27949 = (inp[2]) ? 4'b1011 : node27950;
															assign node27950 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node27954 = (inp[9]) ? node27978 : node27955;
												assign node27955 = (inp[4]) ? node27967 : node27956;
													assign node27956 = (inp[1]) ? node27962 : node27957;
														assign node27957 = (inp[2]) ? 4'b1011 : node27958;
															assign node27958 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node27962 = (inp[0]) ? 4'b1111 : node27963;
															assign node27963 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node27967 = (inp[1]) ? node27973 : node27968;
														assign node27968 = (inp[2]) ? 4'b1110 : node27969;
															assign node27969 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node27973 = (inp[0]) ? 4'b1011 : node27974;
															assign node27974 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node27978 = (inp[4]) ? node27990 : node27979;
													assign node27979 = (inp[1]) ? node27985 : node27980;
														assign node27980 = (inp[2]) ? 4'b1010 : node27981;
															assign node27981 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node27985 = (inp[2]) ? node27987 : 4'b1110;
															assign node27987 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node27990 = (inp[1]) ? node27996 : node27991;
														assign node27991 = (inp[0]) ? 4'b1111 : node27992;
															assign node27992 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node27996 = (inp[10]) ? 4'b1010 : node27997;
															assign node27997 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node28001 = (inp[1]) ? node28057 : node28002;
											assign node28002 = (inp[4]) ? node28034 : node28003;
												assign node28003 = (inp[10]) ? node28021 : node28004;
													assign node28004 = (inp[9]) ? node28016 : node28005;
														assign node28005 = (inp[11]) ? node28011 : node28006;
															assign node28006 = (inp[2]) ? node28008 : 4'b1000;
																assign node28008 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node28011 = (inp[0]) ? 4'b1001 : node28012;
																assign node28012 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node28016 = (inp[11]) ? node28018 : 4'b1001;
															assign node28018 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node28021 = (inp[2]) ? node28029 : node28022;
														assign node28022 = (inp[11]) ? node28026 : node28023;
															assign node28023 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node28026 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node28029 = (inp[0]) ? node28031 : 4'b1000;
															assign node28031 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node28034 = (inp[9]) ? node28046 : node28035;
													assign node28035 = (inp[11]) ? node28041 : node28036;
														assign node28036 = (inp[2]) ? node28038 : 4'b1100;
															assign node28038 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node28041 = (inp[0]) ? node28043 : 4'b1101;
															assign node28043 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node28046 = (inp[11]) ? node28052 : node28047;
														assign node28047 = (inp[0]) ? node28049 : 4'b1101;
															assign node28049 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node28052 = (inp[0]) ? node28054 : 4'b1100;
															assign node28054 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node28057 = (inp[4]) ? node28077 : node28058;
												assign node28058 = (inp[9]) ? node28066 : node28059;
													assign node28059 = (inp[11]) ? 4'b1100 : node28060;
														assign node28060 = (inp[2]) ? 4'b1101 : node28061;
															assign node28061 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node28066 = (inp[11]) ? node28072 : node28067;
														assign node28067 = (inp[0]) ? node28069 : 4'b1100;
															assign node28069 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node28072 = (inp[0]) ? node28074 : 4'b1101;
															assign node28074 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node28077 = (inp[9]) ? node28089 : node28078;
													assign node28078 = (inp[11]) ? node28084 : node28079;
														assign node28079 = (inp[0]) ? node28081 : 4'b1001;
															assign node28081 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node28084 = (inp[0]) ? node28086 : 4'b1000;
															assign node28086 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node28089 = (inp[11]) ? node28095 : node28090;
														assign node28090 = (inp[2]) ? node28092 : 4'b1000;
															assign node28092 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node28095 = (inp[2]) ? node28097 : 4'b1001;
															assign node28097 = (inp[0]) ? 4'b1000 : 4'b1001;
								assign node28100 = (inp[15]) ? node28294 : node28101;
									assign node28101 = (inp[7]) ? node28203 : node28102;
										assign node28102 = (inp[4]) ? node28144 : node28103;
											assign node28103 = (inp[1]) ? node28123 : node28104;
												assign node28104 = (inp[9]) ? node28112 : node28105;
													assign node28105 = (inp[11]) ? node28107 : 4'b1000;
														assign node28107 = (inp[0]) ? node28109 : 4'b1001;
															assign node28109 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node28112 = (inp[11]) ? node28118 : node28113;
														assign node28113 = (inp[2]) ? 4'b1001 : node28114;
															assign node28114 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node28118 = (inp[0]) ? node28120 : 4'b1000;
															assign node28120 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node28123 = (inp[2]) ? node28131 : node28124;
													assign node28124 = (inp[9]) ? node28128 : node28125;
														assign node28125 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node28128 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node28131 = (inp[0]) ? node28137 : node28132;
														assign node28132 = (inp[9]) ? 4'b1000 : node28133;
															assign node28133 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node28137 = (inp[9]) ? node28141 : node28138;
															assign node28138 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node28141 = (inp[11]) ? 4'b1001 : 4'b1000;
											assign node28144 = (inp[1]) ? node28164 : node28145;
												assign node28145 = (inp[11]) ? node28155 : node28146;
													assign node28146 = (inp[9]) ? node28152 : node28147;
														assign node28147 = (inp[2]) ? node28149 : 4'b1000;
															assign node28149 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node28152 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node28155 = (inp[9]) ? node28161 : node28156;
														assign node28156 = (inp[0]) ? node28158 : 4'b1001;
															assign node28158 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node28161 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node28164 = (inp[2]) ? node28178 : node28165;
													assign node28165 = (inp[0]) ? node28171 : node28166;
														assign node28166 = (inp[9]) ? node28168 : 4'b1100;
															assign node28168 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node28171 = (inp[11]) ? node28175 : node28172;
															assign node28172 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node28175 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node28178 = (inp[10]) ? node28194 : node28179;
														assign node28179 = (inp[11]) ? node28187 : node28180;
															assign node28180 = (inp[9]) ? node28184 : node28181;
																assign node28181 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node28184 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node28187 = (inp[0]) ? node28191 : node28188;
																assign node28188 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node28191 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node28194 = (inp[0]) ? 4'b1100 : node28195;
															assign node28195 = (inp[11]) ? node28199 : node28196;
																assign node28196 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node28199 = (inp[9]) ? 4'b1101 : 4'b1100;
										assign node28203 = (inp[4]) ? node28247 : node28204;
											assign node28204 = (inp[1]) ? node28228 : node28205;
												assign node28205 = (inp[9]) ? node28217 : node28206;
													assign node28206 = (inp[11]) ? node28212 : node28207;
														assign node28207 = (inp[0]) ? 4'b1110 : node28208;
															assign node28208 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node28212 = (inp[2]) ? node28214 : 4'b1111;
															assign node28214 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node28217 = (inp[11]) ? node28223 : node28218;
														assign node28218 = (inp[0]) ? 4'b1111 : node28219;
															assign node28219 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node28223 = (inp[2]) ? node28225 : 4'b1110;
															assign node28225 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node28228 = (inp[11]) ? node28236 : node28229;
													assign node28229 = (inp[9]) ? node28233 : node28230;
														assign node28230 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node28233 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node28236 = (inp[9]) ? node28242 : node28237;
														assign node28237 = (inp[0]) ? node28239 : 4'b1011;
															assign node28239 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node28242 = (inp[0]) ? node28244 : 4'b1010;
															assign node28244 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node28247 = (inp[9]) ? node28271 : node28248;
												assign node28248 = (inp[11]) ? node28260 : node28249;
													assign node28249 = (inp[0]) ? node28255 : node28250;
														assign node28250 = (inp[2]) ? 4'b1010 : node28251;
															assign node28251 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node28255 = (inp[2]) ? node28257 : 4'b1010;
															assign node28257 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node28260 = (inp[1]) ? node28266 : node28261;
														assign node28261 = (inp[0]) ? 4'b1011 : node28262;
															assign node28262 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node28266 = (inp[2]) ? node28268 : 4'b1011;
															assign node28268 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node28271 = (inp[11]) ? node28283 : node28272;
													assign node28272 = (inp[10]) ? node28278 : node28273;
														assign node28273 = (inp[0]) ? node28275 : 4'b1011;
															assign node28275 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node28278 = (inp[0]) ? 4'b1011 : node28279;
															assign node28279 = (inp[1]) ? 4'b1011 : 4'b1010;
													assign node28283 = (inp[1]) ? node28289 : node28284;
														assign node28284 = (inp[0]) ? 4'b1010 : node28285;
															assign node28285 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node28289 = (inp[0]) ? node28291 : 4'b1010;
															assign node28291 = (inp[2]) ? 4'b1011 : 4'b1010;
									assign node28294 = (inp[7]) ? node28364 : node28295;
										assign node28295 = (inp[11]) ? node28323 : node28296;
											assign node28296 = (inp[9]) ? node28314 : node28297;
												assign node28297 = (inp[0]) ? node28299 : 4'b1010;
													assign node28299 = (inp[10]) ? node28307 : node28300;
														assign node28300 = (inp[2]) ? node28304 : node28301;
															assign node28301 = (inp[4]) ? 4'b1010 : 4'b1011;
															assign node28304 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node28307 = (inp[1]) ? 4'b1011 : node28308;
															assign node28308 = (inp[2]) ? 4'b1011 : node28309;
																assign node28309 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node28314 = (inp[0]) ? node28316 : 4'b1011;
													assign node28316 = (inp[2]) ? node28320 : node28317;
														assign node28317 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node28320 = (inp[4]) ? 4'b1010 : 4'b1011;
											assign node28323 = (inp[9]) ? node28339 : node28324;
												assign node28324 = (inp[0]) ? node28326 : 4'b1011;
													assign node28326 = (inp[1]) ? node28334 : node28327;
														assign node28327 = (inp[2]) ? node28331 : node28328;
															assign node28328 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node28331 = (inp[4]) ? 4'b1010 : 4'b1011;
														assign node28334 = (inp[4]) ? 4'b1010 : node28335;
															assign node28335 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node28339 = (inp[0]) ? node28341 : 4'b1010;
													assign node28341 = (inp[1]) ? node28357 : node28342;
														assign node28342 = (inp[10]) ? node28350 : node28343;
															assign node28343 = (inp[4]) ? node28347 : node28344;
																assign node28344 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node28347 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node28350 = (inp[4]) ? node28354 : node28351;
																assign node28351 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node28354 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node28357 = (inp[2]) ? node28361 : node28358;
															assign node28358 = (inp[4]) ? 4'b1010 : 4'b1011;
															assign node28361 = (inp[4]) ? 4'b1011 : 4'b1010;
										assign node28364 = (inp[9]) ? node28412 : node28365;
											assign node28365 = (inp[11]) ? node28391 : node28366;
												assign node28366 = (inp[0]) ? node28368 : 4'b1001;
													assign node28368 = (inp[10]) ? node28376 : node28369;
														assign node28369 = (inp[1]) ? node28371 : 4'b1000;
															assign node28371 = (inp[2]) ? 4'b1000 : node28372;
																assign node28372 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node28376 = (inp[1]) ? node28384 : node28377;
															assign node28377 = (inp[4]) ? node28381 : node28378;
																assign node28378 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node28381 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node28384 = (inp[2]) ? node28388 : node28385;
																assign node28385 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node28388 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node28391 = (inp[0]) ? node28393 : 4'b1000;
													assign node28393 = (inp[1]) ? node28401 : node28394;
														assign node28394 = (inp[2]) ? node28398 : node28395;
															assign node28395 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node28398 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node28401 = (inp[10]) ? node28407 : node28402;
															assign node28402 = (inp[4]) ? node28404 : 4'b1001;
																assign node28404 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node28407 = (inp[2]) ? node28409 : 4'b1001;
																assign node28409 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node28412 = (inp[11]) ? node28422 : node28413;
												assign node28413 = (inp[0]) ? node28415 : 4'b1000;
													assign node28415 = (inp[4]) ? node28419 : node28416;
														assign node28416 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node28419 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node28422 = (inp[0]) ? node28424 : 4'b1001;
													assign node28424 = (inp[2]) ? node28428 : node28425;
														assign node28425 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node28428 = (inp[4]) ? 4'b1000 : 4'b1001;
						assign node28431 = (inp[6]) ? node29607 : node28432;
							assign node28432 = (inp[9]) ? node29014 : node28433;
								assign node28433 = (inp[10]) ? node28729 : node28434;
									assign node28434 = (inp[11]) ? node28602 : node28435;
										assign node28435 = (inp[2]) ? node28517 : node28436;
											assign node28436 = (inp[1]) ? node28476 : node28437;
												assign node28437 = (inp[4]) ? node28451 : node28438;
													assign node28438 = (inp[15]) ? node28446 : node28439;
														assign node28439 = (inp[7]) ? node28443 : node28440;
															assign node28440 = (inp[12]) ? 4'b1110 : 4'b1100;
															assign node28443 = (inp[12]) ? 4'b1001 : 4'b1110;
														assign node28446 = (inp[7]) ? 4'b1100 : node28447;
															assign node28447 = (inp[12]) ? 4'b1111 : 4'b1101;
													assign node28451 = (inp[12]) ? node28465 : node28452;
														assign node28452 = (inp[7]) ? node28458 : node28453;
															assign node28453 = (inp[15]) ? node28455 : 4'b1110;
																assign node28455 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node28458 = (inp[15]) ? node28462 : node28459;
																assign node28459 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node28462 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node28465 = (inp[15]) ? node28471 : node28466;
															assign node28466 = (inp[7]) ? 4'b1111 : node28467;
																assign node28467 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node28471 = (inp[7]) ? 4'b1100 : node28472;
																assign node28472 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node28476 = (inp[7]) ? node28496 : node28477;
													assign node28477 = (inp[12]) ? node28489 : node28478;
														assign node28478 = (inp[15]) ? node28486 : node28479;
															assign node28479 = (inp[0]) ? node28483 : node28480;
																assign node28480 = (inp[4]) ? 4'b1011 : 4'b1001;
																assign node28483 = (inp[4]) ? 4'b1010 : 4'b1000;
															assign node28486 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node28489 = (inp[4]) ? node28493 : node28490;
															assign node28490 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node28493 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node28496 = (inp[12]) ? node28506 : node28497;
														assign node28497 = (inp[0]) ? node28503 : node28498;
															assign node28498 = (inp[15]) ? 4'b1111 : node28499;
																assign node28499 = (inp[4]) ? 4'b1101 : 4'b1111;
															assign node28503 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node28506 = (inp[4]) ? node28510 : node28507;
															assign node28507 = (inp[15]) ? 4'b1000 : 4'b1100;
															assign node28510 = (inp[15]) ? node28514 : node28511;
																assign node28511 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node28514 = (inp[0]) ? 4'b1000 : 4'b1001;
											assign node28517 = (inp[1]) ? node28567 : node28518;
												assign node28518 = (inp[7]) ? node28542 : node28519;
													assign node28519 = (inp[12]) ? node28531 : node28520;
														assign node28520 = (inp[4]) ? node28528 : node28521;
															assign node28521 = (inp[15]) ? node28525 : node28522;
																assign node28522 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node28525 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node28528 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node28531 = (inp[4]) ? node28539 : node28532;
															assign node28532 = (inp[15]) ? node28536 : node28533;
																assign node28533 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node28536 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node28539 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node28542 = (inp[12]) ? node28556 : node28543;
														assign node28543 = (inp[15]) ? node28551 : node28544;
															assign node28544 = (inp[4]) ? node28548 : node28545;
																assign node28545 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node28548 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node28551 = (inp[4]) ? 4'b1011 : node28552;
																assign node28552 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node28556 = (inp[15]) ? node28562 : node28557;
															assign node28557 = (inp[4]) ? node28559 : 4'b1101;
																assign node28559 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node28562 = (inp[4]) ? 4'b1000 : node28563;
																assign node28563 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node28567 = (inp[7]) ? node28589 : node28568;
													assign node28568 = (inp[12]) ? node28580 : node28569;
														assign node28569 = (inp[15]) ? node28575 : node28570;
															assign node28570 = (inp[4]) ? node28572 : 4'b1101;
																assign node28572 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node28575 = (inp[4]) ? node28577 : 4'b1100;
																assign node28577 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node28580 = (inp[15]) ? node28584 : node28581;
															assign node28581 = (inp[4]) ? 4'b1101 : 4'b1110;
															assign node28584 = (inp[0]) ? node28586 : 4'b1111;
																assign node28586 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node28589 = (inp[12]) ? node28595 : node28590;
														assign node28590 = (inp[4]) ? node28592 : 4'b1011;
															assign node28592 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28595 = (inp[15]) ? node28597 : 4'b1000;
															assign node28597 = (inp[4]) ? node28599 : 4'b1100;
																assign node28599 = (inp[0]) ? 4'b1101 : 4'b1100;
										assign node28602 = (inp[12]) ? node28666 : node28603;
											assign node28603 = (inp[7]) ? node28633 : node28604;
												assign node28604 = (inp[4]) ? node28620 : node28605;
													assign node28605 = (inp[15]) ? node28613 : node28606;
														assign node28606 = (inp[2]) ? node28610 : node28607;
															assign node28607 = (inp[1]) ? 4'b1001 : 4'b1101;
															assign node28610 = (inp[1]) ? 4'b1101 : 4'b1001;
														assign node28613 = (inp[2]) ? 4'b1000 : node28614;
															assign node28614 = (inp[1]) ? node28616 : 4'b1101;
																assign node28616 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node28620 = (inp[15]) ? node28626 : node28621;
														assign node28621 = (inp[2]) ? node28623 : 4'b1011;
															assign node28623 = (inp[1]) ? 4'b1110 : 4'b1010;
														assign node28626 = (inp[2]) ? node28630 : node28627;
															assign node28627 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node28630 = (inp[1]) ? 4'b1000 : 4'b1101;
												assign node28633 = (inp[15]) ? node28651 : node28634;
													assign node28634 = (inp[4]) ? node28642 : node28635;
														assign node28635 = (inp[2]) ? node28639 : node28636;
															assign node28636 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node28639 = (inp[1]) ? 4'b1010 : 4'b1011;
														assign node28642 = (inp[2]) ? node28646 : node28643;
															assign node28643 = (inp[1]) ? 4'b1101 : 4'b1001;
															assign node28646 = (inp[1]) ? node28648 : 4'b1100;
																assign node28648 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node28651 = (inp[1]) ? node28661 : node28652;
														assign node28652 = (inp[0]) ? node28658 : node28653;
															assign node28653 = (inp[2]) ? 4'b1010 : node28654;
																assign node28654 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node28658 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node28661 = (inp[4]) ? node28663 : 4'b1011;
															assign node28663 = (inp[0]) ? 4'b1111 : 4'b1011;
											assign node28666 = (inp[7]) ? node28700 : node28667;
												assign node28667 = (inp[4]) ? node28685 : node28668;
													assign node28668 = (inp[2]) ? node28678 : node28669;
														assign node28669 = (inp[1]) ? 4'b1010 : node28670;
															assign node28670 = (inp[15]) ? node28674 : node28671;
																assign node28671 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node28674 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node28678 = (inp[1]) ? node28682 : node28679;
															assign node28679 = (inp[15]) ? 4'b1010 : 4'b1011;
															assign node28682 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node28685 = (inp[15]) ? node28695 : node28686;
														assign node28686 = (inp[2]) ? node28690 : node28687;
															assign node28687 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node28690 = (inp[0]) ? node28692 : 4'b1100;
																assign node28692 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node28695 = (inp[2]) ? 4'b1111 : node28696;
															assign node28696 = (inp[1]) ? 4'b1010 : 4'b1110;
												assign node28700 = (inp[4]) ? node28720 : node28701;
													assign node28701 = (inp[2]) ? node28715 : node28702;
														assign node28702 = (inp[0]) ? node28708 : node28703;
															assign node28703 = (inp[1]) ? node28705 : 4'b1000;
																assign node28705 = (inp[15]) ? 4'b1001 : 4'b1101;
															assign node28708 = (inp[15]) ? node28712 : node28709;
																assign node28709 = (inp[1]) ? 4'b1100 : 4'b1001;
																assign node28712 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node28715 = (inp[1]) ? node28717 : 4'b1001;
															assign node28717 = (inp[15]) ? 4'b1101 : 4'b1001;
													assign node28720 = (inp[2]) ? node28726 : node28721;
														assign node28721 = (inp[1]) ? 4'b1011 : node28722;
															assign node28722 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node28726 = (inp[1]) ? 4'b1110 : 4'b1011;
									assign node28729 = (inp[11]) ? node28875 : node28730;
										assign node28730 = (inp[1]) ? node28804 : node28731;
											assign node28731 = (inp[2]) ? node28763 : node28732;
												assign node28732 = (inp[12]) ? node28746 : node28733;
													assign node28733 = (inp[15]) ? node28739 : node28734;
														assign node28734 = (inp[4]) ? 4'b1111 : node28735;
															assign node28735 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node28739 = (inp[4]) ? node28743 : node28740;
															assign node28740 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node28743 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node28746 = (inp[15]) ? node28756 : node28747;
														assign node28747 = (inp[7]) ? node28753 : node28748;
															assign node28748 = (inp[4]) ? node28750 : 4'b1111;
																assign node28750 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node28753 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node28756 = (inp[7]) ? 4'b1101 : node28757;
															assign node28757 = (inp[4]) ? node28759 : 4'b1110;
																assign node28759 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node28763 = (inp[12]) ? node28785 : node28764;
													assign node28764 = (inp[7]) ? node28774 : node28765;
														assign node28765 = (inp[4]) ? 4'b1010 : node28766;
															assign node28766 = (inp[0]) ? node28770 : node28767;
																assign node28767 = (inp[15]) ? 4'b1001 : 4'b1000;
																assign node28770 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node28774 = (inp[4]) ? node28782 : node28775;
															assign node28775 = (inp[15]) ? node28779 : node28776;
																assign node28776 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node28779 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node28782 = (inp[15]) ? 4'b1010 : 4'b1100;
													assign node28785 = (inp[7]) ? node28795 : node28786;
														assign node28786 = (inp[15]) ? node28792 : node28787;
															assign node28787 = (inp[4]) ? node28789 : 4'b1011;
																assign node28789 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node28792 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node28795 = (inp[15]) ? node28799 : node28796;
															assign node28796 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node28799 = (inp[4]) ? 4'b1001 : node28800;
																assign node28800 = (inp[0]) ? 4'b1001 : 4'b1000;
											assign node28804 = (inp[2]) ? node28832 : node28805;
												assign node28805 = (inp[7]) ? node28821 : node28806;
													assign node28806 = (inp[12]) ? node28816 : node28807;
														assign node28807 = (inp[15]) ? node28813 : node28808;
															assign node28808 = (inp[0]) ? 4'b1011 : node28809;
																assign node28809 = (inp[4]) ? 4'b1010 : 4'b1000;
															assign node28813 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node28816 = (inp[4]) ? node28818 : 4'b1010;
															assign node28818 = (inp[15]) ? 4'b1010 : 4'b1001;
													assign node28821 = (inp[12]) ? node28829 : node28822;
														assign node28822 = (inp[0]) ? 4'b1111 : node28823;
															assign node28823 = (inp[15]) ? 4'b1010 : node28824;
																assign node28824 = (inp[4]) ? 4'b1100 : 4'b1110;
														assign node28829 = (inp[15]) ? 4'b1001 : 4'b1101;
												assign node28832 = (inp[7]) ? node28854 : node28833;
													assign node28833 = (inp[12]) ? node28843 : node28834;
														assign node28834 = (inp[4]) ? node28840 : node28835;
															assign node28835 = (inp[15]) ? 4'b1101 : node28836;
																assign node28836 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node28840 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node28843 = (inp[15]) ? node28849 : node28844;
															assign node28844 = (inp[0]) ? node28846 : 4'b1111;
																assign node28846 = (inp[4]) ? 4'b1100 : 4'b1110;
															assign node28849 = (inp[0]) ? node28851 : 4'b1110;
																assign node28851 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node28854 = (inp[12]) ? node28864 : node28855;
														assign node28855 = (inp[4]) ? node28861 : node28856;
															assign node28856 = (inp[15]) ? node28858 : 4'b1010;
																assign node28858 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node28861 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node28864 = (inp[4]) ? node28868 : node28865;
															assign node28865 = (inp[15]) ? 4'b1101 : 4'b1001;
															assign node28868 = (inp[0]) ? node28872 : node28869;
																assign node28869 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node28872 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node28875 = (inp[7]) ? node28947 : node28876;
											assign node28876 = (inp[12]) ? node28906 : node28877;
												assign node28877 = (inp[15]) ? node28889 : node28878;
													assign node28878 = (inp[4]) ? node28884 : node28879;
														assign node28879 = (inp[1]) ? 4'b1100 : node28880;
															assign node28880 = (inp[0]) ? 4'b1000 : 4'b1100;
														assign node28884 = (inp[1]) ? 4'b1010 : node28885;
															assign node28885 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node28889 = (inp[0]) ? node28899 : node28890;
														assign node28890 = (inp[1]) ? node28894 : node28891;
															assign node28891 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node28894 = (inp[4]) ? 4'b1100 : node28895;
																assign node28895 = (inp[2]) ? 4'b1100 : 4'b1000;
														assign node28899 = (inp[2]) ? 4'b1001 : node28900;
															assign node28900 = (inp[4]) ? node28902 : 4'b1001;
																assign node28902 = (inp[1]) ? 4'b1101 : 4'b1001;
												assign node28906 = (inp[15]) ? node28920 : node28907;
													assign node28907 = (inp[4]) ? node28915 : node28908;
														assign node28908 = (inp[2]) ? 4'b1010 : node28909;
															assign node28909 = (inp[1]) ? 4'b1011 : node28910;
																assign node28910 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node28915 = (inp[2]) ? node28917 : 4'b1000;
															assign node28917 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node28920 = (inp[0]) ? node28934 : node28921;
														assign node28921 = (inp[4]) ? node28927 : node28922;
															assign node28922 = (inp[1]) ? node28924 : 4'b1011;
																assign node28924 = (inp[2]) ? 4'b1111 : 4'b1011;
															assign node28927 = (inp[2]) ? node28931 : node28928;
																assign node28928 = (inp[1]) ? 4'b1011 : 4'b1111;
																assign node28931 = (inp[1]) ? 4'b1110 : 4'b1011;
														assign node28934 = (inp[2]) ? node28942 : node28935;
															assign node28935 = (inp[1]) ? node28939 : node28936;
																assign node28936 = (inp[4]) ? 4'b1111 : 4'b1110;
																assign node28939 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node28942 = (inp[1]) ? 4'b1110 : node28943;
																assign node28943 = (inp[4]) ? 4'b1010 : 4'b1011;
											assign node28947 = (inp[12]) ? node28981 : node28948;
												assign node28948 = (inp[4]) ? node28962 : node28949;
													assign node28949 = (inp[15]) ? node28959 : node28950;
														assign node28950 = (inp[2]) ? node28954 : node28951;
															assign node28951 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node28954 = (inp[1]) ? node28956 : 4'b1010;
																assign node28956 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node28959 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node28962 = (inp[15]) ? node28970 : node28963;
														assign node28963 = (inp[2]) ? node28967 : node28964;
															assign node28964 = (inp[1]) ? 4'b1100 : 4'b1000;
															assign node28967 = (inp[1]) ? 4'b1000 : 4'b1101;
														assign node28970 = (inp[2]) ? node28974 : node28971;
															assign node28971 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node28974 = (inp[0]) ? node28978 : node28975;
																assign node28975 = (inp[1]) ? 4'b1010 : 4'b1011;
																assign node28978 = (inp[1]) ? 4'b1011 : 4'b1010;
												assign node28981 = (inp[15]) ? node28997 : node28982;
													assign node28982 = (inp[4]) ? node28990 : node28983;
														assign node28983 = (inp[0]) ? node28987 : node28984;
															assign node28984 = (inp[2]) ? 4'b1000 : 4'b1100;
															assign node28987 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node28990 = (inp[2]) ? node28994 : node28991;
															assign node28991 = (inp[1]) ? 4'b1010 : 4'b1111;
															assign node28994 = (inp[1]) ? 4'b1111 : 4'b1010;
													assign node28997 = (inp[0]) ? node29003 : node28998;
														assign node28998 = (inp[2]) ? 4'b1000 : node28999;
															assign node28999 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node29003 = (inp[2]) ? node29009 : node29004;
															assign node29004 = (inp[1]) ? 4'b1000 : node29005;
																assign node29005 = (inp[4]) ? 4'b1100 : 4'b1101;
															assign node29009 = (inp[1]) ? 4'b1101 : node29010;
																assign node29010 = (inp[4]) ? 4'b1001 : 4'b1000;
								assign node29014 = (inp[4]) ? node29320 : node29015;
									assign node29015 = (inp[7]) ? node29173 : node29016;
										assign node29016 = (inp[12]) ? node29086 : node29017;
											assign node29017 = (inp[2]) ? node29049 : node29018;
												assign node29018 = (inp[1]) ? node29030 : node29019;
													assign node29019 = (inp[10]) ? node29025 : node29020;
														assign node29020 = (inp[15]) ? 4'b1100 : node29021;
															assign node29021 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node29025 = (inp[0]) ? node29027 : 4'b1101;
															assign node29027 = (inp[15]) ? 4'b1101 : 4'b1100;
													assign node29030 = (inp[10]) ? node29038 : node29031;
														assign node29031 = (inp[11]) ? node29033 : 4'b1001;
															assign node29033 = (inp[0]) ? node29035 : 4'b1000;
																assign node29035 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node29038 = (inp[15]) ? node29044 : node29039;
															assign node29039 = (inp[0]) ? node29041 : 4'b1001;
																assign node29041 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node29044 = (inp[11]) ? node29046 : 4'b1000;
																assign node29046 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node29049 = (inp[1]) ? node29067 : node29050;
													assign node29050 = (inp[11]) ? node29060 : node29051;
														assign node29051 = (inp[0]) ? 4'b1000 : node29052;
															assign node29052 = (inp[10]) ? node29056 : node29053;
																assign node29053 = (inp[15]) ? 4'b1001 : 4'b1000;
																assign node29056 = (inp[15]) ? 4'b1000 : 4'b1001;
														assign node29060 = (inp[10]) ? node29064 : node29061;
															assign node29061 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node29064 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node29067 = (inp[11]) ? node29075 : node29068;
														assign node29068 = (inp[10]) ? 4'b1100 : node29069;
															assign node29069 = (inp[0]) ? 4'b1101 : node29070;
																assign node29070 = (inp[15]) ? 4'b1101 : 4'b1100;
														assign node29075 = (inp[10]) ? node29081 : node29076;
															assign node29076 = (inp[15]) ? node29078 : 4'b1100;
																assign node29078 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29081 = (inp[15]) ? node29083 : 4'b1101;
																assign node29083 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node29086 = (inp[10]) ? node29130 : node29087;
												assign node29087 = (inp[0]) ? node29107 : node29088;
													assign node29088 = (inp[15]) ? node29098 : node29089;
														assign node29089 = (inp[1]) ? node29095 : node29090;
															assign node29090 = (inp[2]) ? 4'b1010 : node29091;
																assign node29091 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29095 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node29098 = (inp[11]) ? node29102 : node29099;
															assign node29099 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node29102 = (inp[1]) ? 4'b1111 : node29103;
																assign node29103 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node29107 = (inp[15]) ? node29121 : node29108;
														assign node29108 = (inp[1]) ? node29114 : node29109;
															assign node29109 = (inp[2]) ? node29111 : 4'b1111;
																assign node29111 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node29114 = (inp[11]) ? node29118 : node29115;
																assign node29115 = (inp[2]) ? 4'b1110 : 4'b1010;
																assign node29118 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node29121 = (inp[2]) ? node29125 : node29122;
															assign node29122 = (inp[1]) ? 4'b1010 : 4'b1110;
															assign node29125 = (inp[11]) ? 4'b1011 : node29126;
																assign node29126 = (inp[1]) ? 4'b1110 : 4'b1010;
												assign node29130 = (inp[0]) ? node29156 : node29131;
													assign node29131 = (inp[11]) ? node29141 : node29132;
														assign node29132 = (inp[15]) ? node29134 : 4'b1110;
															assign node29134 = (inp[1]) ? node29138 : node29135;
																assign node29135 = (inp[2]) ? 4'b1010 : 4'b1111;
																assign node29138 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node29141 = (inp[15]) ? node29149 : node29142;
															assign node29142 = (inp[1]) ? node29146 : node29143;
																assign node29143 = (inp[2]) ? 4'b1011 : 4'b1111;
																assign node29146 = (inp[2]) ? 4'b1110 : 4'b1010;
															assign node29149 = (inp[2]) ? node29153 : node29150;
																assign node29150 = (inp[1]) ? 4'b1010 : 4'b1110;
																assign node29153 = (inp[1]) ? 4'b1110 : 4'b1010;
													assign node29156 = (inp[15]) ? node29166 : node29157;
														assign node29157 = (inp[1]) ? node29161 : node29158;
															assign node29158 = (inp[2]) ? 4'b1010 : 4'b1110;
															assign node29161 = (inp[2]) ? node29163 : 4'b1011;
																assign node29163 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node29166 = (inp[2]) ? node29170 : node29167;
															assign node29167 = (inp[1]) ? 4'b1011 : 4'b1111;
															assign node29170 = (inp[1]) ? 4'b1111 : 4'b1011;
										assign node29173 = (inp[12]) ? node29257 : node29174;
											assign node29174 = (inp[10]) ? node29214 : node29175;
												assign node29175 = (inp[1]) ? node29195 : node29176;
													assign node29176 = (inp[15]) ? node29186 : node29177;
														assign node29177 = (inp[2]) ? node29183 : node29178;
															assign node29178 = (inp[11]) ? node29180 : 4'b1111;
																assign node29180 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node29183 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node29186 = (inp[2]) ? node29190 : node29187;
															assign node29187 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node29190 = (inp[11]) ? 4'b1111 : node29191;
																assign node29191 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node29195 = (inp[0]) ? node29205 : node29196;
														assign node29196 = (inp[15]) ? node29202 : node29197;
															assign node29197 = (inp[2]) ? node29199 : 4'b1110;
																assign node29199 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node29202 = (inp[2]) ? 4'b1110 : 4'b1010;
														assign node29205 = (inp[15]) ? node29211 : node29206;
															assign node29206 = (inp[2]) ? 4'b1010 : node29207;
																assign node29207 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29211 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node29214 = (inp[1]) ? node29234 : node29215;
													assign node29215 = (inp[2]) ? node29225 : node29216;
														assign node29216 = (inp[15]) ? node29220 : node29217;
															assign node29217 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node29220 = (inp[0]) ? node29222 : 4'b1010;
																assign node29222 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node29225 = (inp[15]) ? node29231 : node29226;
															assign node29226 = (inp[11]) ? 4'b1011 : node29227;
																assign node29227 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node29231 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node29234 = (inp[0]) ? node29244 : node29235;
														assign node29235 = (inp[2]) ? node29239 : node29236;
															assign node29236 = (inp[15]) ? 4'b1011 : 4'b1111;
															assign node29239 = (inp[15]) ? 4'b1111 : node29240;
																assign node29240 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node29244 = (inp[11]) ? node29252 : node29245;
															assign node29245 = (inp[2]) ? node29249 : node29246;
																assign node29246 = (inp[15]) ? 4'b1010 : 4'b1110;
																assign node29249 = (inp[15]) ? 4'b1110 : 4'b1011;
															assign node29252 = (inp[15]) ? 4'b1111 : node29253;
																assign node29253 = (inp[2]) ? 4'b1011 : 4'b1111;
											assign node29257 = (inp[15]) ? node29291 : node29258;
												assign node29258 = (inp[0]) ? node29276 : node29259;
													assign node29259 = (inp[11]) ? node29267 : node29260;
														assign node29260 = (inp[2]) ? 4'b1001 : node29261;
															assign node29261 = (inp[1]) ? node29263 : 4'b1001;
																assign node29263 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node29267 = (inp[10]) ? node29271 : node29268;
															assign node29268 = (inp[1]) ? 4'b1000 : 4'b1101;
															assign node29271 = (inp[1]) ? 4'b1101 : node29272;
																assign node29272 = (inp[2]) ? 4'b1100 : 4'b1000;
													assign node29276 = (inp[10]) ? node29282 : node29277;
														assign node29277 = (inp[2]) ? node29279 : 4'b1000;
															assign node29279 = (inp[1]) ? 4'b1000 : 4'b1100;
														assign node29282 = (inp[1]) ? node29286 : node29283;
															assign node29283 = (inp[2]) ? 4'b1101 : 4'b1001;
															assign node29286 = (inp[2]) ? node29288 : 4'b1100;
																assign node29288 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node29291 = (inp[10]) ? node29305 : node29292;
													assign node29292 = (inp[0]) ? node29300 : node29293;
														assign node29293 = (inp[1]) ? node29295 : 4'b1000;
															assign node29295 = (inp[11]) ? 4'b1000 : node29296;
																assign node29296 = (inp[2]) ? 4'b1101 : 4'b1001;
														assign node29300 = (inp[2]) ? 4'b1101 : node29301;
															assign node29301 = (inp[1]) ? 4'b1001 : 4'b1101;
													assign node29305 = (inp[11]) ? node29313 : node29306;
														assign node29306 = (inp[2]) ? node29310 : node29307;
															assign node29307 = (inp[1]) ? 4'b1000 : 4'b1100;
															assign node29310 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node29313 = (inp[1]) ? node29315 : 4'b1001;
															assign node29315 = (inp[0]) ? 4'b1100 : node29316;
																assign node29316 = (inp[2]) ? 4'b1101 : 4'b1001;
									assign node29320 = (inp[12]) ? node29478 : node29321;
										assign node29321 = (inp[2]) ? node29401 : node29322;
											assign node29322 = (inp[7]) ? node29362 : node29323;
												assign node29323 = (inp[15]) ? node29341 : node29324;
													assign node29324 = (inp[1]) ? node29332 : node29325;
														assign node29325 = (inp[10]) ? node29329 : node29326;
															assign node29326 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29329 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node29332 = (inp[11]) ? node29338 : node29333;
															assign node29333 = (inp[10]) ? 4'b1010 : node29334;
																assign node29334 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node29338 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node29341 = (inp[1]) ? node29353 : node29342;
														assign node29342 = (inp[10]) ? node29348 : node29343;
															assign node29343 = (inp[0]) ? node29345 : 4'b1001;
																assign node29345 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node29348 = (inp[11]) ? 4'b1000 : node29349;
																assign node29349 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node29353 = (inp[10]) ? node29359 : node29354;
															assign node29354 = (inp[11]) ? node29356 : 4'b1101;
																assign node29356 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29359 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node29362 = (inp[15]) ? node29384 : node29363;
													assign node29363 = (inp[1]) ? node29373 : node29364;
														assign node29364 = (inp[10]) ? node29368 : node29365;
															assign node29365 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node29368 = (inp[0]) ? node29370 : 4'b1001;
																assign node29370 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node29373 = (inp[10]) ? node29379 : node29374;
															assign node29374 = (inp[11]) ? 4'b1100 : node29375;
																assign node29375 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node29379 = (inp[0]) ? node29381 : 4'b1101;
																assign node29381 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node29384 = (inp[1]) ? node29394 : node29385;
														assign node29385 = (inp[10]) ? node29391 : node29386;
															assign node29386 = (inp[11]) ? 4'b1111 : node29387;
																assign node29387 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node29391 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node29394 = (inp[10]) ? node29396 : 4'b1110;
															assign node29396 = (inp[11]) ? 4'b1111 : node29397;
																assign node29397 = (inp[0]) ? 4'b1110 : 4'b1111;
											assign node29401 = (inp[10]) ? node29441 : node29402;
												assign node29402 = (inp[15]) ? node29420 : node29403;
													assign node29403 = (inp[7]) ? node29415 : node29404;
														assign node29404 = (inp[1]) ? node29410 : node29405;
															assign node29405 = (inp[11]) ? 4'b1011 : node29406;
																assign node29406 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node29410 = (inp[11]) ? 4'b1111 : node29411;
																assign node29411 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node29415 = (inp[1]) ? 4'b1001 : node29416;
															assign node29416 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node29420 = (inp[7]) ? node29430 : node29421;
														assign node29421 = (inp[1]) ? node29427 : node29422;
															assign node29422 = (inp[0]) ? node29424 : 4'b1100;
																assign node29424 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node29427 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node29430 = (inp[1]) ? node29436 : node29431;
															assign node29431 = (inp[0]) ? 4'b1010 : node29432;
																assign node29432 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node29436 = (inp[0]) ? 4'b1011 : node29437;
																assign node29437 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node29441 = (inp[15]) ? node29457 : node29442;
													assign node29442 = (inp[7]) ? node29450 : node29443;
														assign node29443 = (inp[1]) ? 4'b1110 : node29444;
															assign node29444 = (inp[11]) ? 4'b1010 : node29445;
																assign node29445 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node29450 = (inp[1]) ? 4'b1000 : node29451;
															assign node29451 = (inp[0]) ? node29453 : 4'b1100;
																assign node29453 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node29457 = (inp[7]) ? node29469 : node29458;
														assign node29458 = (inp[1]) ? node29464 : node29459;
															assign node29459 = (inp[11]) ? 4'b1101 : node29460;
																assign node29460 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node29464 = (inp[11]) ? 4'b1000 : node29465;
																assign node29465 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node29469 = (inp[0]) ? node29475 : node29470;
															assign node29470 = (inp[11]) ? node29472 : 4'b1011;
																assign node29472 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node29475 = (inp[1]) ? 4'b1010 : 4'b1011;
										assign node29478 = (inp[2]) ? node29542 : node29479;
											assign node29479 = (inp[1]) ? node29515 : node29480;
												assign node29480 = (inp[15]) ? node29496 : node29481;
													assign node29481 = (inp[7]) ? node29491 : node29482;
														assign node29482 = (inp[10]) ? node29486 : node29483;
															assign node29483 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node29486 = (inp[0]) ? node29488 : 4'b1001;
																assign node29488 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node29491 = (inp[0]) ? node29493 : 4'b1110;
															assign node29493 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node29496 = (inp[7]) ? node29504 : node29497;
														assign node29497 = (inp[10]) ? node29499 : 4'b1111;
															assign node29499 = (inp[11]) ? 4'b1110 : node29500;
																assign node29500 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node29504 = (inp[10]) ? node29510 : node29505;
															assign node29505 = (inp[0]) ? node29507 : 4'b1100;
																assign node29507 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node29510 = (inp[0]) ? node29512 : 4'b1101;
																assign node29512 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node29515 = (inp[7]) ? node29533 : node29516;
													assign node29516 = (inp[15]) ? node29528 : node29517;
														assign node29517 = (inp[10]) ? node29523 : node29518;
															assign node29518 = (inp[11]) ? node29520 : 4'b1001;
																assign node29520 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node29523 = (inp[0]) ? 4'b1000 : node29524;
																assign node29524 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node29528 = (inp[10]) ? 4'b1010 : node29529;
															assign node29529 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node29533 = (inp[15]) ? node29537 : node29534;
														assign node29534 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node29537 = (inp[10]) ? 4'b1001 : node29538;
															assign node29538 = (inp[11]) ? 4'b1000 : 4'b1001;
											assign node29542 = (inp[1]) ? node29580 : node29543;
												assign node29543 = (inp[7]) ? node29559 : node29544;
													assign node29544 = (inp[15]) ? node29552 : node29545;
														assign node29545 = (inp[10]) ? node29547 : 4'b1101;
															assign node29547 = (inp[0]) ? node29549 : 4'b1100;
																assign node29549 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29552 = (inp[10]) ? node29554 : 4'b1010;
															assign node29554 = (inp[0]) ? 4'b1011 : node29555;
																assign node29555 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node29559 = (inp[15]) ? node29571 : node29560;
														assign node29560 = (inp[10]) ? node29566 : node29561;
															assign node29561 = (inp[11]) ? 4'b1010 : node29562;
																assign node29562 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node29566 = (inp[0]) ? node29568 : 4'b1011;
																assign node29568 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node29571 = (inp[10]) ? node29577 : node29572;
															assign node29572 = (inp[11]) ? node29574 : 4'b1001;
																assign node29574 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node29577 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node29580 = (inp[0]) ? node29596 : node29581;
													assign node29581 = (inp[10]) ? node29587 : node29582;
														assign node29582 = (inp[11]) ? 4'b1101 : node29583;
															assign node29583 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node29587 = (inp[11]) ? node29589 : 4'b1101;
															assign node29589 = (inp[7]) ? node29593 : node29590;
																assign node29590 = (inp[15]) ? 4'b1111 : 4'b1100;
																assign node29593 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node29596 = (inp[10]) ? node29600 : node29597;
														assign node29597 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node29600 = (inp[7]) ? node29604 : node29601;
															assign node29601 = (inp[15]) ? 4'b1110 : 4'b1101;
															assign node29604 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node29607 = (inp[12]) ? node30099 : node29608;
								assign node29608 = (inp[15]) ? node29878 : node29609;
									assign node29609 = (inp[7]) ? node29733 : node29610;
										assign node29610 = (inp[1]) ? node29680 : node29611;
											assign node29611 = (inp[2]) ? node29643 : node29612;
												assign node29612 = (inp[10]) ? node29630 : node29613;
													assign node29613 = (inp[4]) ? node29621 : node29614;
														assign node29614 = (inp[11]) ? node29618 : node29615;
															assign node29615 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node29618 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node29621 = (inp[0]) ? node29623 : 4'b1101;
															assign node29623 = (inp[11]) ? node29627 : node29624;
																assign node29624 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node29627 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node29630 = (inp[0]) ? node29636 : node29631;
														assign node29631 = (inp[9]) ? node29633 : 4'b1100;
															assign node29633 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29636 = (inp[9]) ? node29640 : node29637;
															assign node29637 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node29640 = (inp[11]) ? 4'b1100 : 4'b1101;
												assign node29643 = (inp[4]) ? node29665 : node29644;
													assign node29644 = (inp[10]) ? node29658 : node29645;
														assign node29645 = (inp[0]) ? node29653 : node29646;
															assign node29646 = (inp[9]) ? node29650 : node29647;
																assign node29647 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node29650 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node29653 = (inp[9]) ? node29655 : 4'b1100;
																assign node29655 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29658 = (inp[9]) ? node29660 : 4'b1101;
															assign node29660 = (inp[11]) ? node29662 : 4'b1101;
																assign node29662 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node29665 = (inp[0]) ? node29673 : node29666;
														assign node29666 = (inp[11]) ? node29670 : node29667;
															assign node29667 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node29670 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node29673 = (inp[11]) ? node29677 : node29674;
															assign node29674 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node29677 = (inp[9]) ? 4'b1101 : 4'b1100;
											assign node29680 = (inp[4]) ? node29704 : node29681;
												assign node29681 = (inp[9]) ? node29693 : node29682;
													assign node29682 = (inp[11]) ? node29688 : node29683;
														assign node29683 = (inp[2]) ? 4'b1001 : node29684;
															assign node29684 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node29688 = (inp[2]) ? 4'b1000 : node29689;
															assign node29689 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node29693 = (inp[10]) ? node29695 : 4'b1001;
														assign node29695 = (inp[11]) ? node29701 : node29696;
															assign node29696 = (inp[2]) ? 4'b1000 : node29697;
																assign node29697 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node29701 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node29704 = (inp[0]) ? node29720 : node29705;
													assign node29705 = (inp[2]) ? node29713 : node29706;
														assign node29706 = (inp[11]) ? node29710 : node29707;
															assign node29707 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node29710 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node29713 = (inp[10]) ? node29715 : 4'b1100;
															assign node29715 = (inp[11]) ? 4'b1100 : node29716;
																assign node29716 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node29720 = (inp[2]) ? node29728 : node29721;
														assign node29721 = (inp[11]) ? node29725 : node29722;
															assign node29722 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node29725 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node29728 = (inp[11]) ? 4'b1101 : node29729;
															assign node29729 = (inp[9]) ? 4'b1101 : 4'b1100;
										assign node29733 = (inp[4]) ? node29807 : node29734;
											assign node29734 = (inp[10]) ? node29770 : node29735;
												assign node29735 = (inp[9]) ? node29751 : node29736;
													assign node29736 = (inp[0]) ? node29742 : node29737;
														assign node29737 = (inp[11]) ? node29739 : 4'b1111;
															assign node29739 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node29742 = (inp[11]) ? node29746 : node29743;
															assign node29743 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node29746 = (inp[2]) ? node29748 : 4'b1111;
																assign node29748 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node29751 = (inp[1]) ? node29763 : node29752;
														assign node29752 = (inp[11]) ? node29758 : node29753;
															assign node29753 = (inp[0]) ? 4'b1111 : node29754;
																assign node29754 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node29758 = (inp[2]) ? node29760 : 4'b1110;
																assign node29760 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node29763 = (inp[11]) ? node29765 : 4'b1110;
															assign node29765 = (inp[2]) ? 4'b1111 : node29766;
																assign node29766 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node29770 = (inp[1]) ? node29790 : node29771;
													assign node29771 = (inp[9]) ? node29781 : node29772;
														assign node29772 = (inp[11]) ? node29778 : node29773;
															assign node29773 = (inp[0]) ? 4'b1110 : node29774;
																assign node29774 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node29778 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node29781 = (inp[2]) ? node29785 : node29782;
															assign node29782 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node29785 = (inp[11]) ? node29787 : 4'b1110;
																assign node29787 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node29790 = (inp[0]) ? node29798 : node29791;
														assign node29791 = (inp[11]) ? node29795 : node29792;
															assign node29792 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node29795 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node29798 = (inp[2]) ? node29800 : 4'b1110;
															assign node29800 = (inp[9]) ? node29804 : node29801;
																assign node29801 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node29804 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node29807 = (inp[1]) ? node29845 : node29808;
												assign node29808 = (inp[2]) ? node29828 : node29809;
													assign node29809 = (inp[10]) ? node29821 : node29810;
														assign node29810 = (inp[11]) ? node29816 : node29811;
															assign node29811 = (inp[0]) ? node29813 : 4'b1010;
																assign node29813 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node29816 = (inp[9]) ? 4'b1011 : node29817;
																assign node29817 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node29821 = (inp[9]) ? 4'b1010 : node29822;
															assign node29822 = (inp[0]) ? node29824 : 4'b1010;
																assign node29824 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node29828 = (inp[0]) ? node29836 : node29829;
														assign node29829 = (inp[11]) ? node29833 : node29830;
															assign node29830 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node29833 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node29836 = (inp[10]) ? 4'b1011 : node29837;
															assign node29837 = (inp[9]) ? node29841 : node29838;
																assign node29838 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node29841 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node29845 = (inp[2]) ? node29871 : node29846;
													assign node29846 = (inp[10]) ? node29862 : node29847;
														assign node29847 = (inp[0]) ? node29855 : node29848;
															assign node29848 = (inp[9]) ? node29852 : node29849;
																assign node29849 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node29852 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node29855 = (inp[11]) ? node29859 : node29856;
																assign node29856 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node29859 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node29862 = (inp[11]) ? node29864 : 4'b1110;
															assign node29864 = (inp[0]) ? node29868 : node29865;
																assign node29865 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node29868 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node29871 = (inp[9]) ? node29875 : node29872;
														assign node29872 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node29875 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node29878 = (inp[7]) ? node29964 : node29879;
										assign node29879 = (inp[1]) ? node29921 : node29880;
											assign node29880 = (inp[4]) ? node29898 : node29881;
												assign node29881 = (inp[9]) ? node29893 : node29882;
													assign node29882 = (inp[11]) ? node29888 : node29883;
														assign node29883 = (inp[2]) ? node29885 : 4'b1111;
															assign node29885 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node29888 = (inp[2]) ? node29890 : 4'b1110;
															assign node29890 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node29893 = (inp[11]) ? 4'b1111 : node29894;
														assign node29894 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node29898 = (inp[11]) ? node29910 : node29899;
													assign node29899 = (inp[9]) ? node29905 : node29900;
														assign node29900 = (inp[2]) ? 4'b1011 : node29901;
															assign node29901 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node29905 = (inp[0]) ? 4'b1010 : node29906;
															assign node29906 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node29910 = (inp[9]) ? node29916 : node29911;
														assign node29911 = (inp[0]) ? 4'b1010 : node29912;
															assign node29912 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node29916 = (inp[2]) ? 4'b1011 : node29917;
															assign node29917 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node29921 = (inp[4]) ? node29943 : node29922;
												assign node29922 = (inp[0]) ? node29936 : node29923;
													assign node29923 = (inp[9]) ? node29929 : node29924;
														assign node29924 = (inp[2]) ? 4'b1010 : node29925;
															assign node29925 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node29929 = (inp[11]) ? node29933 : node29930;
															assign node29930 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node29933 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node29936 = (inp[11]) ? node29940 : node29937;
														assign node29937 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node29940 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node29943 = (inp[9]) ? node29953 : node29944;
													assign node29944 = (inp[11]) ? node29950 : node29945;
														assign node29945 = (inp[2]) ? node29947 : 4'b1110;
															assign node29947 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node29950 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node29953 = (inp[11]) ? node29959 : node29954;
														assign node29954 = (inp[2]) ? node29956 : 4'b1111;
															assign node29956 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node29959 = (inp[2]) ? node29961 : 4'b1110;
															assign node29961 = (inp[0]) ? 4'b1111 : 4'b1110;
										assign node29964 = (inp[2]) ? node30056 : node29965;
											assign node29965 = (inp[10]) ? node30011 : node29966;
												assign node29966 = (inp[1]) ? node29986 : node29967;
													assign node29967 = (inp[4]) ? node29981 : node29968;
														assign node29968 = (inp[9]) ? node29976 : node29969;
															assign node29969 = (inp[11]) ? node29973 : node29970;
																assign node29970 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node29973 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node29976 = (inp[0]) ? 4'b1101 : node29977;
																assign node29977 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node29981 = (inp[11]) ? 4'b1001 : node29982;
															assign node29982 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node29986 = (inp[4]) ? node30000 : node29987;
														assign node29987 = (inp[0]) ? node29993 : node29988;
															assign node29988 = (inp[11]) ? 4'b1001 : node29989;
																assign node29989 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node29993 = (inp[9]) ? node29997 : node29994;
																assign node29994 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node29997 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node30000 = (inp[9]) ? node30006 : node30001;
															assign node30001 = (inp[0]) ? 4'b1101 : node30002;
																assign node30002 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node30006 = (inp[11]) ? 4'b1100 : node30007;
																assign node30007 = (inp[0]) ? 4'b1101 : 4'b1100;
												assign node30011 = (inp[4]) ? node30037 : node30012;
													assign node30012 = (inp[1]) ? node30024 : node30013;
														assign node30013 = (inp[11]) ? node30019 : node30014;
															assign node30014 = (inp[0]) ? node30016 : 4'b1100;
																assign node30016 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node30019 = (inp[9]) ? 4'b1101 : node30020;
																assign node30020 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node30024 = (inp[9]) ? node30032 : node30025;
															assign node30025 = (inp[11]) ? node30029 : node30026;
																assign node30026 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node30029 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node30032 = (inp[0]) ? node30034 : 4'b1000;
																assign node30034 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node30037 = (inp[1]) ? node30043 : node30038;
														assign node30038 = (inp[11]) ? node30040 : 4'b1000;
															assign node30040 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node30043 = (inp[11]) ? node30049 : node30044;
															assign node30044 = (inp[9]) ? node30046 : 4'b1100;
																assign node30046 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30049 = (inp[9]) ? node30053 : node30050;
																assign node30050 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node30053 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node30056 = (inp[9]) ? node30076 : node30057;
												assign node30057 = (inp[4]) ? node30065 : node30058;
													assign node30058 = (inp[1]) ? node30062 : node30059;
														assign node30059 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30062 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node30065 = (inp[1]) ? node30073 : node30066;
														assign node30066 = (inp[0]) ? node30070 : node30067;
															assign node30067 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node30070 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node30073 = (inp[11]) ? 4'b1101 : 4'b1100;
												assign node30076 = (inp[11]) ? node30086 : node30077;
													assign node30077 = (inp[1]) ? node30083 : node30078;
														assign node30078 = (inp[4]) ? node30080 : 4'b1101;
															assign node30080 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node30083 = (inp[4]) ? 4'b1101 : 4'b1000;
													assign node30086 = (inp[0]) ? node30094 : node30087;
														assign node30087 = (inp[1]) ? node30091 : node30088;
															assign node30088 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node30091 = (inp[4]) ? 4'b1100 : 4'b1001;
														assign node30094 = (inp[1]) ? node30096 : 4'b1001;
															assign node30096 = (inp[4]) ? 4'b1100 : 4'b1001;
								assign node30099 = (inp[15]) ? node30301 : node30100;
									assign node30100 = (inp[7]) ? node30200 : node30101;
										assign node30101 = (inp[1]) ? node30139 : node30102;
											assign node30102 = (inp[4]) ? node30126 : node30103;
												assign node30103 = (inp[11]) ? node30113 : node30104;
													assign node30104 = (inp[9]) ? node30108 : node30105;
														assign node30105 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node30108 = (inp[2]) ? node30110 : 4'b1101;
															assign node30110 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node30113 = (inp[10]) ? node30121 : node30114;
														assign node30114 = (inp[2]) ? node30116 : 4'b1101;
															assign node30116 = (inp[9]) ? node30118 : 4'b1100;
																assign node30118 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node30121 = (inp[0]) ? node30123 : 4'b1100;
															assign node30123 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node30126 = (inp[11]) ? node30132 : node30127;
													assign node30127 = (inp[9]) ? node30129 : 4'b1100;
														assign node30129 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node30132 = (inp[9]) ? node30134 : 4'b1101;
														assign node30134 = (inp[0]) ? 4'b1100 : node30135;
															assign node30135 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node30139 = (inp[4]) ? node30163 : node30140;
												assign node30140 = (inp[9]) ? node30150 : node30141;
													assign node30141 = (inp[11]) ? node30147 : node30142;
														assign node30142 = (inp[2]) ? 4'b1100 : node30143;
															assign node30143 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node30147 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node30150 = (inp[11]) ? node30158 : node30151;
														assign node30151 = (inp[10]) ? 4'b1101 : node30152;
															assign node30152 = (inp[2]) ? 4'b1101 : node30153;
																assign node30153 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node30158 = (inp[0]) ? node30160 : 4'b1100;
															assign node30160 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node30163 = (inp[10]) ? node30185 : node30164;
													assign node30164 = (inp[0]) ? node30172 : node30165;
														assign node30165 = (inp[9]) ? node30169 : node30166;
															assign node30166 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node30169 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node30172 = (inp[9]) ? node30178 : node30173;
															assign node30173 = (inp[2]) ? 4'b1001 : node30174;
																assign node30174 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node30178 = (inp[11]) ? node30182 : node30179;
																assign node30179 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node30182 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node30185 = (inp[0]) ? node30187 : 4'b1001;
														assign node30187 = (inp[11]) ? node30195 : node30188;
															assign node30188 = (inp[2]) ? node30192 : node30189;
																assign node30189 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node30192 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node30195 = (inp[9]) ? node30197 : 4'b1001;
																assign node30197 = (inp[2]) ? 4'b1001 : 4'b1000;
										assign node30200 = (inp[4]) ? node30242 : node30201;
											assign node30201 = (inp[1]) ? node30219 : node30202;
												assign node30202 = (inp[9]) ? node30214 : node30203;
													assign node30203 = (inp[11]) ? node30209 : node30204;
														assign node30204 = (inp[2]) ? node30206 : 4'b1011;
															assign node30206 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node30209 = (inp[2]) ? node30211 : 4'b1010;
															assign node30211 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node30214 = (inp[11]) ? 4'b1011 : node30215;
														assign node30215 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node30219 = (inp[11]) ? node30231 : node30220;
													assign node30220 = (inp[9]) ? node30226 : node30221;
														assign node30221 = (inp[0]) ? 4'b1110 : node30222;
															assign node30222 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node30226 = (inp[2]) ? node30228 : 4'b1111;
															assign node30228 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node30231 = (inp[9]) ? node30237 : node30232;
														assign node30232 = (inp[2]) ? node30234 : 4'b1111;
															assign node30234 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node30237 = (inp[0]) ? 4'b1110 : node30238;
															assign node30238 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node30242 = (inp[2]) ? node30274 : node30243;
												assign node30243 = (inp[0]) ? node30251 : node30244;
													assign node30244 = (inp[9]) ? node30248 : node30245;
														assign node30245 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node30248 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node30251 = (inp[1]) ? node30259 : node30252;
														assign node30252 = (inp[11]) ? node30256 : node30253;
															assign node30253 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node30256 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node30259 = (inp[10]) ? node30267 : node30260;
															assign node30260 = (inp[11]) ? node30264 : node30261;
																assign node30261 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node30264 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node30267 = (inp[11]) ? node30271 : node30268;
																assign node30268 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node30271 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node30274 = (inp[9]) ? node30286 : node30275;
													assign node30275 = (inp[11]) ? node30281 : node30276;
														assign node30276 = (inp[0]) ? 4'b1110 : node30277;
															assign node30277 = (inp[1]) ? 4'b1110 : 4'b1111;
														assign node30281 = (inp[1]) ? 4'b1111 : node30282;
															assign node30282 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node30286 = (inp[0]) ? 4'b1111 : node30287;
														assign node30287 = (inp[10]) ? node30293 : node30288;
															assign node30288 = (inp[11]) ? 4'b1111 : node30289;
																assign node30289 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node30293 = (inp[1]) ? node30297 : node30294;
																assign node30294 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node30297 = (inp[11]) ? 4'b1110 : 4'b1111;
									assign node30301 = (inp[7]) ? node30423 : node30302;
										assign node30302 = (inp[10]) ? node30348 : node30303;
											assign node30303 = (inp[11]) ? node30331 : node30304;
												assign node30304 = (inp[9]) ? node30314 : node30305;
													assign node30305 = (inp[0]) ? 4'b1111 : node30306;
														assign node30306 = (inp[4]) ? node30310 : node30307;
															assign node30307 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node30310 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node30314 = (inp[0]) ? 4'b1110 : node30315;
														assign node30315 = (inp[1]) ? node30323 : node30316;
															assign node30316 = (inp[2]) ? node30320 : node30317;
																assign node30317 = (inp[4]) ? 4'b1111 : 4'b1110;
																assign node30320 = (inp[4]) ? 4'b1110 : 4'b1111;
															assign node30323 = (inp[4]) ? node30327 : node30324;
																assign node30324 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node30327 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node30331 = (inp[9]) ? node30339 : node30332;
													assign node30332 = (inp[4]) ? 4'b1110 : node30333;
														assign node30333 = (inp[0]) ? 4'b1110 : node30334;
															assign node30334 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node30339 = (inp[0]) ? 4'b1111 : node30340;
														assign node30340 = (inp[4]) ? node30344 : node30341;
															assign node30341 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node30344 = (inp[2]) ? 4'b1111 : 4'b1110;
											assign node30348 = (inp[4]) ? node30386 : node30349;
												assign node30349 = (inp[2]) ? node30363 : node30350;
													assign node30350 = (inp[0]) ? node30356 : node30351;
														assign node30351 = (inp[9]) ? node30353 : 4'b1111;
															assign node30353 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node30356 = (inp[1]) ? node30358 : 4'b1110;
															assign node30358 = (inp[11]) ? node30360 : 4'b1111;
																assign node30360 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node30363 = (inp[11]) ? node30377 : node30364;
														assign node30364 = (inp[1]) ? node30372 : node30365;
															assign node30365 = (inp[9]) ? node30369 : node30366;
																assign node30366 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node30369 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node30372 = (inp[0]) ? 4'b1111 : node30373;
																assign node30373 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node30377 = (inp[1]) ? 4'b1110 : node30378;
															assign node30378 = (inp[9]) ? node30382 : node30379;
																assign node30379 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node30382 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node30386 = (inp[2]) ? node30416 : node30387;
													assign node30387 = (inp[9]) ? node30401 : node30388;
														assign node30388 = (inp[1]) ? node30394 : node30389;
															assign node30389 = (inp[0]) ? node30391 : 4'b1110;
																assign node30391 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node30394 = (inp[11]) ? node30398 : node30395;
																assign node30395 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node30398 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node30401 = (inp[1]) ? node30409 : node30402;
															assign node30402 = (inp[11]) ? node30406 : node30403;
																assign node30403 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node30406 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node30409 = (inp[0]) ? node30413 : node30410;
																assign node30410 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node30413 = (inp[11]) ? 4'b1111 : 4'b1110;
													assign node30416 = (inp[9]) ? node30420 : node30417;
														assign node30417 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node30420 = (inp[11]) ? 4'b1111 : 4'b1110;
										assign node30423 = (inp[2]) ? node30475 : node30424;
											assign node30424 = (inp[0]) ? node30446 : node30425;
												assign node30425 = (inp[11]) ? node30441 : node30426;
													assign node30426 = (inp[10]) ? node30434 : node30427;
														assign node30427 = (inp[4]) ? node30431 : node30428;
															assign node30428 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node30431 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node30434 = (inp[9]) ? node30438 : node30435;
															assign node30435 = (inp[4]) ? 4'b1101 : 4'b1100;
															assign node30438 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node30441 = (inp[4]) ? node30443 : 4'b1100;
														assign node30443 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node30446 = (inp[1]) ? node30468 : node30447;
													assign node30447 = (inp[10]) ? node30459 : node30448;
														assign node30448 = (inp[4]) ? node30454 : node30449;
															assign node30449 = (inp[11]) ? node30451 : 4'b1101;
																assign node30451 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node30454 = (inp[9]) ? node30456 : 4'b1100;
																assign node30456 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node30459 = (inp[4]) ? node30465 : node30460;
															assign node30460 = (inp[9]) ? node30462 : 4'b1100;
																assign node30462 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node30465 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node30468 = (inp[11]) ? node30472 : node30469;
														assign node30469 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node30472 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node30475 = (inp[4]) ? node30505 : node30476;
												assign node30476 = (inp[10]) ? node30490 : node30477;
													assign node30477 = (inp[9]) ? node30485 : node30478;
														assign node30478 = (inp[0]) ? node30482 : node30479;
															assign node30479 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node30482 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30485 = (inp[11]) ? 4'b1101 : node30486;
															assign node30486 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node30490 = (inp[1]) ? node30492 : 4'b1101;
														assign node30492 = (inp[11]) ? node30500 : node30493;
															assign node30493 = (inp[9]) ? node30497 : node30494;
																assign node30494 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node30497 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node30500 = (inp[9]) ? node30502 : 4'b1101;
																assign node30502 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node30505 = (inp[1]) ? node30513 : node30506;
													assign node30506 = (inp[9]) ? node30510 : node30507;
														assign node30507 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30510 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node30513 = (inp[9]) ? node30517 : node30514;
														assign node30514 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node30517 = (inp[11]) ? 4'b1100 : 4'b1101;
					assign node30520 = (inp[13]) ? node32538 : node30521;
						assign node30521 = (inp[6]) ? node31731 : node30522;
							assign node30522 = (inp[2]) ? node31146 : node30523;
								assign node30523 = (inp[12]) ? node30837 : node30524;
									assign node30524 = (inp[7]) ? node30684 : node30525;
										assign node30525 = (inp[4]) ? node30613 : node30526;
											assign node30526 = (inp[0]) ? node30570 : node30527;
												assign node30527 = (inp[15]) ? node30551 : node30528;
													assign node30528 = (inp[1]) ? node30536 : node30529;
														assign node30529 = (inp[11]) ? node30531 : 4'b1000;
															assign node30531 = (inp[9]) ? node30533 : 4'b1000;
																assign node30533 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node30536 = (inp[9]) ? node30544 : node30537;
															assign node30537 = (inp[11]) ? node30541 : node30538;
																assign node30538 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node30541 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node30544 = (inp[11]) ? node30548 : node30545;
																assign node30545 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node30548 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node30551 = (inp[1]) ? node30563 : node30552;
														assign node30552 = (inp[11]) ? node30558 : node30553;
															assign node30553 = (inp[9]) ? node30555 : 4'b1001;
																assign node30555 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node30558 = (inp[10]) ? 4'b1001 : node30559;
																assign node30559 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node30563 = (inp[9]) ? node30567 : node30564;
															assign node30564 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node30567 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node30570 = (inp[15]) ? node30588 : node30571;
													assign node30571 = (inp[10]) ? node30577 : node30572;
														assign node30572 = (inp[11]) ? node30574 : 4'b1001;
															assign node30574 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node30577 = (inp[9]) ? node30583 : node30578;
															assign node30578 = (inp[11]) ? 4'b1001 : node30579;
																assign node30579 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node30583 = (inp[11]) ? 4'b1000 : node30584;
																assign node30584 = (inp[1]) ? 4'b1000 : 4'b1001;
													assign node30588 = (inp[10]) ? node30598 : node30589;
														assign node30589 = (inp[11]) ? node30591 : 4'b1000;
															assign node30591 = (inp[1]) ? node30595 : node30592;
																assign node30592 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node30595 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node30598 = (inp[11]) ? node30606 : node30599;
															assign node30599 = (inp[1]) ? node30603 : node30600;
																assign node30600 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node30603 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node30606 = (inp[9]) ? node30610 : node30607;
																assign node30607 = (inp[1]) ? 4'b1000 : 4'b1001;
																assign node30610 = (inp[1]) ? 4'b1001 : 4'b1000;
											assign node30613 = (inp[15]) ? node30643 : node30614;
												assign node30614 = (inp[9]) ? node30634 : node30615;
													assign node30615 = (inp[1]) ? node30623 : node30616;
														assign node30616 = (inp[10]) ? 4'b1011 : node30617;
															assign node30617 = (inp[0]) ? 4'b1010 : node30618;
																assign node30618 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node30623 = (inp[10]) ? node30629 : node30624;
															assign node30624 = (inp[11]) ? 4'b1011 : node30625;
																assign node30625 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node30629 = (inp[0]) ? node30631 : 4'b1010;
																assign node30631 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node30634 = (inp[10]) ? node30640 : node30635;
														assign node30635 = (inp[11]) ? 4'b1010 : node30636;
															assign node30636 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node30640 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node30643 = (inp[11]) ? node30659 : node30644;
													assign node30644 = (inp[10]) ? node30652 : node30645;
														assign node30645 = (inp[9]) ? node30649 : node30646;
															assign node30646 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node30649 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node30652 = (inp[1]) ? node30656 : node30653;
															assign node30653 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node30656 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node30659 = (inp[0]) ? node30675 : node30660;
														assign node30660 = (inp[9]) ? node30668 : node30661;
															assign node30661 = (inp[10]) ? node30665 : node30662;
																assign node30662 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node30665 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node30668 = (inp[10]) ? node30672 : node30669;
																assign node30669 = (inp[1]) ? 4'b1101 : 4'b1100;
																assign node30672 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node30675 = (inp[9]) ? node30677 : 4'b1100;
															assign node30677 = (inp[10]) ? node30681 : node30678;
																assign node30678 = (inp[1]) ? 4'b1100 : 4'b1101;
																assign node30681 = (inp[1]) ? 4'b1101 : 4'b1100;
										assign node30684 = (inp[4]) ? node30762 : node30685;
											assign node30685 = (inp[10]) ? node30717 : node30686;
												assign node30686 = (inp[9]) ? node30706 : node30687;
													assign node30687 = (inp[0]) ? node30697 : node30688;
														assign node30688 = (inp[1]) ? node30694 : node30689;
															assign node30689 = (inp[15]) ? node30691 : 4'b1111;
																assign node30691 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node30694 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node30697 = (inp[1]) ? node30703 : node30698;
															assign node30698 = (inp[15]) ? 4'b1011 : node30699;
																assign node30699 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node30703 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node30706 = (inp[1]) ? node30712 : node30707;
														assign node30707 = (inp[15]) ? 4'b1010 : node30708;
															assign node30708 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node30712 = (inp[15]) ? 4'b1111 : node30713;
															assign node30713 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node30717 = (inp[9]) ? node30743 : node30718;
													assign node30718 = (inp[0]) ? node30730 : node30719;
														assign node30719 = (inp[11]) ? node30725 : node30720;
															assign node30720 = (inp[1]) ? node30722 : 4'b1010;
																assign node30722 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node30725 = (inp[1]) ? node30727 : 4'b1011;
																assign node30727 = (inp[15]) ? 4'b1111 : 4'b1011;
														assign node30730 = (inp[11]) ? node30736 : node30731;
															assign node30731 = (inp[15]) ? 4'b1010 : node30732;
																assign node30732 = (inp[1]) ? 4'b1010 : 4'b1111;
															assign node30736 = (inp[1]) ? node30740 : node30737;
																assign node30737 = (inp[15]) ? 4'b1010 : 4'b1110;
																assign node30740 = (inp[15]) ? 4'b1111 : 4'b1010;
													assign node30743 = (inp[0]) ? node30753 : node30744;
														assign node30744 = (inp[1]) ? node30750 : node30745;
															assign node30745 = (inp[15]) ? node30747 : 4'b1111;
																assign node30747 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node30750 = (inp[15]) ? 4'b1110 : 4'b1010;
														assign node30753 = (inp[11]) ? 4'b1011 : node30754;
															assign node30754 = (inp[1]) ? node30758 : node30755;
																assign node30755 = (inp[15]) ? 4'b1011 : 4'b1110;
																assign node30758 = (inp[15]) ? 4'b1111 : 4'b1011;
											assign node30762 = (inp[15]) ? node30806 : node30763;
												assign node30763 = (inp[0]) ? node30781 : node30764;
													assign node30764 = (inp[9]) ? node30776 : node30765;
														assign node30765 = (inp[10]) ? node30771 : node30766;
															assign node30766 = (inp[1]) ? 4'b1100 : node30767;
																assign node30767 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node30771 = (inp[11]) ? 4'b1101 : node30772;
																assign node30772 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node30776 = (inp[10]) ? 4'b1100 : node30777;
															assign node30777 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node30781 = (inp[11]) ? node30797 : node30782;
														assign node30782 = (inp[1]) ? node30790 : node30783;
															assign node30783 = (inp[10]) ? node30787 : node30784;
																assign node30784 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node30787 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node30790 = (inp[10]) ? node30794 : node30791;
																assign node30791 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node30794 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node30797 = (inp[1]) ? 4'b1101 : node30798;
															assign node30798 = (inp[10]) ? node30802 : node30799;
																assign node30799 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node30802 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node30806 = (inp[1]) ? node30822 : node30807;
													assign node30807 = (inp[9]) ? node30813 : node30808;
														assign node30808 = (inp[10]) ? 4'b1111 : node30809;
															assign node30809 = (inp[11]) ? 4'b1110 : 4'b1111;
														assign node30813 = (inp[11]) ? 4'b1110 : node30814;
															assign node30814 = (inp[10]) ? node30818 : node30815;
																assign node30815 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node30818 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node30822 = (inp[10]) ? node30828 : node30823;
														assign node30823 = (inp[11]) ? node30825 : 4'b1011;
															assign node30825 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node30828 = (inp[11]) ? 4'b1011 : node30829;
															assign node30829 = (inp[9]) ? node30833 : node30830;
																assign node30830 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node30833 = (inp[0]) ? 4'b1010 : 4'b1011;
									assign node30837 = (inp[7]) ? node30995 : node30838;
										assign node30838 = (inp[15]) ? node30910 : node30839;
											assign node30839 = (inp[4]) ? node30873 : node30840;
												assign node30840 = (inp[1]) ? node30860 : node30841;
													assign node30841 = (inp[10]) ? node30851 : node30842;
														assign node30842 = (inp[9]) ? node30848 : node30843;
															assign node30843 = (inp[0]) ? node30845 : 4'b1010;
																assign node30845 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node30848 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node30851 = (inp[11]) ? node30857 : node30852;
															assign node30852 = (inp[0]) ? node30854 : 4'b1010;
																assign node30854 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node30857 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node30860 = (inp[0]) ? node30868 : node30861;
														assign node30861 = (inp[9]) ? 4'b1010 : node30862;
															assign node30862 = (inp[10]) ? node30864 : 4'b1011;
																assign node30864 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node30868 = (inp[10]) ? 4'b1011 : node30869;
															assign node30869 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node30873 = (inp[1]) ? node30889 : node30874;
													assign node30874 = (inp[11]) ? node30884 : node30875;
														assign node30875 = (inp[0]) ? 4'b1000 : node30876;
															assign node30876 = (inp[9]) ? node30880 : node30877;
																assign node30877 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node30880 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node30884 = (inp[9]) ? 4'b1000 : node30885;
															assign node30885 = (inp[10]) ? 4'b1000 : 4'b1001;
													assign node30889 = (inp[11]) ? node30903 : node30890;
														assign node30890 = (inp[10]) ? node30898 : node30891;
															assign node30891 = (inp[9]) ? node30895 : node30892;
																assign node30892 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node30895 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node30898 = (inp[0]) ? 4'b1100 : node30899;
																assign node30899 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node30903 = (inp[10]) ? node30907 : node30904;
															assign node30904 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node30907 = (inp[9]) ? 4'b1100 : 4'b1101;
											assign node30910 = (inp[1]) ? node30950 : node30911;
												assign node30911 = (inp[10]) ? node30937 : node30912;
													assign node30912 = (inp[0]) ? node30924 : node30913;
														assign node30913 = (inp[11]) ? node30919 : node30914;
															assign node30914 = (inp[4]) ? 4'b1011 : node30915;
																assign node30915 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node30919 = (inp[9]) ? node30921 : 4'b1011;
																assign node30921 = (inp[4]) ? 4'b1010 : 4'b1011;
														assign node30924 = (inp[9]) ? node30932 : node30925;
															assign node30925 = (inp[11]) ? node30929 : node30926;
																assign node30926 = (inp[4]) ? 4'b1010 : 4'b1011;
																assign node30929 = (inp[4]) ? 4'b1011 : 4'b1010;
															assign node30932 = (inp[11]) ? 4'b1010 : node30933;
																assign node30933 = (inp[4]) ? 4'b1011 : 4'b1010;
													assign node30937 = (inp[4]) ? node30945 : node30938;
														assign node30938 = (inp[9]) ? 4'b1010 : node30939;
															assign node30939 = (inp[11]) ? 4'b1011 : node30940;
																assign node30940 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node30945 = (inp[9]) ? node30947 : 4'b1010;
															assign node30947 = (inp[11]) ? 4'b1011 : 4'b1010;
												assign node30950 = (inp[9]) ? node30976 : node30951;
													assign node30951 = (inp[11]) ? node30961 : node30952;
														assign node30952 = (inp[10]) ? node30954 : 4'b1010;
															assign node30954 = (inp[4]) ? node30958 : node30955;
																assign node30955 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node30958 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node30961 = (inp[0]) ? node30969 : node30962;
															assign node30962 = (inp[10]) ? node30966 : node30963;
																assign node30963 = (inp[4]) ? 4'b1011 : 4'b1010;
																assign node30966 = (inp[4]) ? 4'b1010 : 4'b1011;
															assign node30969 = (inp[10]) ? node30973 : node30970;
																assign node30970 = (inp[4]) ? 4'b1011 : 4'b1010;
																assign node30973 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node30976 = (inp[10]) ? node30986 : node30977;
														assign node30977 = (inp[4]) ? node30983 : node30978;
															assign node30978 = (inp[11]) ? 4'b1011 : node30979;
																assign node30979 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node30983 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node30986 = (inp[4]) ? node30990 : node30987;
															assign node30987 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node30990 = (inp[0]) ? node30992 : 4'b1011;
																assign node30992 = (inp[11]) ? 4'b1011 : 4'b1010;
										assign node30995 = (inp[15]) ? node31073 : node30996;
											assign node30996 = (inp[4]) ? node31032 : node30997;
												assign node30997 = (inp[11]) ? node31013 : node30998;
													assign node30998 = (inp[0]) ? node31006 : node30999;
														assign node30999 = (inp[10]) ? node31003 : node31000;
															assign node31000 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node31003 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node31006 = (inp[9]) ? node31008 : 4'b1101;
															assign node31008 = (inp[1]) ? node31010 : 4'b1101;
																assign node31010 = (inp[10]) ? 4'b1100 : 4'b1101;
													assign node31013 = (inp[1]) ? node31027 : node31014;
														assign node31014 = (inp[0]) ? node31022 : node31015;
															assign node31015 = (inp[10]) ? node31019 : node31016;
																assign node31016 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node31019 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node31022 = (inp[10]) ? node31024 : 4'b1100;
																assign node31024 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node31027 = (inp[0]) ? node31029 : 4'b1100;
															assign node31029 = (inp[10]) ? 4'b1100 : 4'b1101;
												assign node31032 = (inp[11]) ? node31056 : node31033;
													assign node31033 = (inp[0]) ? node31045 : node31034;
														assign node31034 = (inp[1]) ? node31040 : node31035;
															assign node31035 = (inp[10]) ? 4'b1011 : node31036;
																assign node31036 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node31040 = (inp[9]) ? node31042 : 4'b1011;
																assign node31042 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node31045 = (inp[1]) ? node31051 : node31046;
															assign node31046 = (inp[9]) ? 4'b1011 : node31047;
																assign node31047 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node31051 = (inp[9]) ? 4'b1010 : node31052;
																assign node31052 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node31056 = (inp[9]) ? node31066 : node31057;
														assign node31057 = (inp[10]) ? node31063 : node31058;
															assign node31058 = (inp[0]) ? 4'b1010 : node31059;
																assign node31059 = (inp[1]) ? 4'b1010 : 4'b1011;
															assign node31063 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node31066 = (inp[1]) ? 4'b1010 : node31067;
															assign node31067 = (inp[10]) ? node31069 : 4'b1010;
																assign node31069 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node31073 = (inp[4]) ? node31117 : node31074;
												assign node31074 = (inp[1]) ? node31096 : node31075;
													assign node31075 = (inp[10]) ? node31087 : node31076;
														assign node31076 = (inp[9]) ? node31082 : node31077;
															assign node31077 = (inp[11]) ? 4'b1000 : node31078;
																assign node31078 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node31082 = (inp[11]) ? 4'b1001 : node31083;
																assign node31083 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node31087 = (inp[9]) ? node31091 : node31088;
															assign node31088 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node31091 = (inp[0]) ? node31093 : 4'b1000;
																assign node31093 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node31096 = (inp[10]) ? node31106 : node31097;
														assign node31097 = (inp[9]) ? node31103 : node31098;
															assign node31098 = (inp[0]) ? node31100 : 4'b1000;
																assign node31100 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node31103 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node31106 = (inp[9]) ? node31112 : node31107;
															assign node31107 = (inp[11]) ? 4'b1001 : node31108;
																assign node31108 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node31112 = (inp[11]) ? 4'b1000 : node31113;
																assign node31113 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node31117 = (inp[11]) ? node31131 : node31118;
													assign node31118 = (inp[0]) ? node31124 : node31119;
														assign node31119 = (inp[9]) ? node31121 : 4'b1001;
															assign node31121 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node31124 = (inp[10]) ? node31128 : node31125;
															assign node31125 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node31128 = (inp[9]) ? 4'b1000 : 4'b1001;
													assign node31131 = (inp[1]) ? node31139 : node31132;
														assign node31132 = (inp[10]) ? node31136 : node31133;
															assign node31133 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node31136 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node31139 = (inp[9]) ? node31143 : node31140;
															assign node31140 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node31143 = (inp[10]) ? 4'b1001 : 4'b1000;
								assign node31146 = (inp[12]) ? node31486 : node31147;
									assign node31147 = (inp[7]) ? node31323 : node31148;
										assign node31148 = (inp[15]) ? node31240 : node31149;
											assign node31149 = (inp[4]) ? node31193 : node31150;
												assign node31150 = (inp[1]) ? node31174 : node31151;
													assign node31151 = (inp[11]) ? node31161 : node31152;
														assign node31152 = (inp[0]) ? 4'b1101 : node31153;
															assign node31153 = (inp[10]) ? node31157 : node31154;
																assign node31154 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node31157 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node31161 = (inp[0]) ? node31167 : node31162;
															assign node31162 = (inp[10]) ? node31164 : 4'b1101;
																assign node31164 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node31167 = (inp[10]) ? node31171 : node31168;
																assign node31168 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node31171 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node31174 = (inp[0]) ? node31186 : node31175;
														assign node31175 = (inp[9]) ? node31181 : node31176;
															assign node31176 = (inp[11]) ? node31178 : 4'b1101;
																assign node31178 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node31181 = (inp[11]) ? node31183 : 4'b1100;
																assign node31183 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node31186 = (inp[10]) ? node31190 : node31187;
															assign node31187 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node31190 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node31193 = (inp[1]) ? node31213 : node31194;
													assign node31194 = (inp[10]) ? node31206 : node31195;
														assign node31195 = (inp[9]) ? node31201 : node31196;
															assign node31196 = (inp[0]) ? 4'b1111 : node31197;
																assign node31197 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node31201 = (inp[11]) ? node31203 : 4'b1110;
																assign node31203 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31206 = (inp[9]) ? node31208 : 4'b1110;
															assign node31208 = (inp[0]) ? 4'b1111 : node31209;
																assign node31209 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node31213 = (inp[0]) ? node31227 : node31214;
														assign node31214 = (inp[11]) ? node31220 : node31215;
															assign node31215 = (inp[10]) ? node31217 : 4'b1111;
																assign node31217 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node31220 = (inp[10]) ? node31224 : node31221;
																assign node31221 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node31224 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node31227 = (inp[10]) ? node31233 : node31228;
															assign node31228 = (inp[9]) ? node31230 : 4'b1110;
																assign node31230 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node31233 = (inp[9]) ? node31237 : node31234;
																assign node31234 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node31237 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node31240 = (inp[4]) ? node31282 : node31241;
												assign node31241 = (inp[1]) ? node31259 : node31242;
													assign node31242 = (inp[0]) ? node31248 : node31243;
														assign node31243 = (inp[10]) ? node31245 : 4'b1101;
															assign node31245 = (inp[9]) ? 4'b1100 : 4'b1101;
														assign node31248 = (inp[10]) ? node31254 : node31249;
															assign node31249 = (inp[11]) ? node31251 : 4'b1100;
																assign node31251 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node31254 = (inp[11]) ? node31256 : 4'b1101;
																assign node31256 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node31259 = (inp[11]) ? node31275 : node31260;
														assign node31260 = (inp[10]) ? node31268 : node31261;
															assign node31261 = (inp[9]) ? node31265 : node31262;
																assign node31262 = (inp[0]) ? 4'b1100 : 4'b1101;
																assign node31265 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node31268 = (inp[9]) ? node31272 : node31269;
																assign node31269 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node31272 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node31275 = (inp[10]) ? node31279 : node31276;
															assign node31276 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node31279 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node31282 = (inp[10]) ? node31302 : node31283;
													assign node31283 = (inp[1]) ? node31293 : node31284;
														assign node31284 = (inp[9]) ? node31290 : node31285;
															assign node31285 = (inp[11]) ? 4'b1000 : node31286;
																assign node31286 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node31290 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node31293 = (inp[9]) ? node31297 : node31294;
															assign node31294 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node31297 = (inp[0]) ? node31299 : 4'b1000;
																assign node31299 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node31302 = (inp[1]) ? node31314 : node31303;
														assign node31303 = (inp[9]) ? node31309 : node31304;
															assign node31304 = (inp[11]) ? 4'b1001 : node31305;
																assign node31305 = (inp[0]) ? 4'b1000 : 4'b1001;
															assign node31309 = (inp[0]) ? node31311 : 4'b1000;
																assign node31311 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node31314 = (inp[9]) ? node31318 : node31315;
															assign node31315 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node31318 = (inp[11]) ? 4'b1001 : node31319;
																assign node31319 = (inp[0]) ? 4'b1000 : 4'b1001;
										assign node31323 = (inp[15]) ? node31401 : node31324;
											assign node31324 = (inp[4]) ? node31368 : node31325;
												assign node31325 = (inp[1]) ? node31345 : node31326;
													assign node31326 = (inp[10]) ? node31336 : node31327;
														assign node31327 = (inp[11]) ? node31331 : node31328;
															assign node31328 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node31331 = (inp[9]) ? 4'b1011 : node31332;
																assign node31332 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node31336 = (inp[11]) ? node31338 : 4'b1011;
															assign node31338 = (inp[9]) ? node31342 : node31339;
																assign node31339 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node31342 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node31345 = (inp[0]) ? node31353 : node31346;
														assign node31346 = (inp[11]) ? node31348 : 4'b1111;
															assign node31348 = (inp[10]) ? 4'b1111 : node31349;
																assign node31349 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node31353 = (inp[11]) ? node31361 : node31354;
															assign node31354 = (inp[9]) ? node31358 : node31355;
																assign node31355 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node31358 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node31361 = (inp[10]) ? node31365 : node31362;
																assign node31362 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node31365 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node31368 = (inp[11]) ? node31384 : node31369;
													assign node31369 = (inp[9]) ? node31377 : node31370;
														assign node31370 = (inp[10]) ? 4'b1000 : node31371;
															assign node31371 = (inp[0]) ? node31373 : 4'b1001;
																assign node31373 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node31377 = (inp[10]) ? node31379 : 4'b1000;
															assign node31379 = (inp[0]) ? node31381 : 4'b1001;
																assign node31381 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node31384 = (inp[1]) ? node31390 : node31385;
														assign node31385 = (inp[10]) ? 4'b1001 : node31386;
															assign node31386 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node31390 = (inp[10]) ? node31396 : node31391;
															assign node31391 = (inp[0]) ? 4'b1001 : node31392;
																assign node31392 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node31396 = (inp[0]) ? 4'b1000 : node31397;
																assign node31397 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node31401 = (inp[11]) ? node31445 : node31402;
												assign node31402 = (inp[10]) ? node31422 : node31403;
													assign node31403 = (inp[9]) ? node31413 : node31404;
														assign node31404 = (inp[1]) ? node31408 : node31405;
															assign node31405 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node31408 = (inp[4]) ? node31410 : 4'b1010;
																assign node31410 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node31413 = (inp[1]) ? node31417 : node31414;
															assign node31414 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node31417 = (inp[4]) ? node31419 : 4'b1011;
																assign node31419 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node31422 = (inp[0]) ? node31430 : node31423;
														assign node31423 = (inp[1]) ? node31425 : 4'b1110;
															assign node31425 = (inp[4]) ? node31427 : 4'b1011;
																assign node31427 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node31430 = (inp[9]) ? node31438 : node31431;
															assign node31431 = (inp[1]) ? node31435 : node31432;
																assign node31432 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node31435 = (inp[4]) ? 4'b1110 : 4'b1011;
															assign node31438 = (inp[4]) ? node31442 : node31439;
																assign node31439 = (inp[1]) ? 4'b1010 : 4'b1111;
																assign node31442 = (inp[1]) ? 4'b1111 : 4'b1011;
												assign node31445 = (inp[0]) ? node31471 : node31446;
													assign node31446 = (inp[1]) ? node31460 : node31447;
														assign node31447 = (inp[4]) ? node31453 : node31448;
															assign node31448 = (inp[9]) ? 4'b1110 : node31449;
																assign node31449 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node31453 = (inp[9]) ? node31457 : node31454;
																assign node31454 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node31457 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node31460 = (inp[4]) ? node31466 : node31461;
															assign node31461 = (inp[9]) ? node31463 : 4'b1010;
																assign node31463 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node31466 = (inp[10]) ? 4'b1110 : node31467;
																assign node31467 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node31471 = (inp[4]) ? node31481 : node31472;
														assign node31472 = (inp[1]) ? node31478 : node31473;
															assign node31473 = (inp[10]) ? 4'b1111 : node31474;
																assign node31474 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node31478 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node31481 = (inp[1]) ? node31483 : 4'b1010;
															assign node31483 = (inp[9]) ? 4'b1110 : 4'b1111;
									assign node31486 = (inp[7]) ? node31596 : node31487;
										assign node31487 = (inp[4]) ? node31539 : node31488;
											assign node31488 = (inp[1]) ? node31514 : node31489;
												assign node31489 = (inp[11]) ? node31507 : node31490;
													assign node31490 = (inp[9]) ? node31498 : node31491;
														assign node31491 = (inp[10]) ? node31495 : node31492;
															assign node31492 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node31495 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31498 = (inp[15]) ? 4'b1110 : node31499;
															assign node31499 = (inp[0]) ? node31503 : node31500;
																assign node31500 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node31503 = (inp[10]) ? 4'b1111 : 4'b1110;
													assign node31507 = (inp[10]) ? node31511 : node31508;
														assign node31508 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node31511 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node31514 = (inp[9]) ? node31530 : node31515;
													assign node31515 = (inp[10]) ? node31527 : node31516;
														assign node31516 = (inp[11]) ? node31522 : node31517;
															assign node31517 = (inp[15]) ? node31519 : 4'b1111;
																assign node31519 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node31522 = (inp[0]) ? node31524 : 4'b1110;
																assign node31524 = (inp[15]) ? 4'b1110 : 4'b1111;
														assign node31527 = (inp[15]) ? 4'b1111 : 4'b1110;
													assign node31530 = (inp[10]) ? node31534 : node31531;
														assign node31531 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node31534 = (inp[15]) ? 4'b1110 : node31535;
															assign node31535 = (inp[11]) ? 4'b1110 : 4'b1111;
											assign node31539 = (inp[15]) ? node31577 : node31540;
												assign node31540 = (inp[1]) ? node31556 : node31541;
													assign node31541 = (inp[0]) ? node31543 : 4'b1100;
														assign node31543 = (inp[10]) ? node31549 : node31544;
															assign node31544 = (inp[9]) ? node31546 : 4'b1101;
																assign node31546 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node31549 = (inp[11]) ? node31553 : node31550;
																assign node31550 = (inp[9]) ? 4'b1101 : 4'b1100;
																assign node31553 = (inp[9]) ? 4'b1100 : 4'b1101;
													assign node31556 = (inp[11]) ? node31564 : node31557;
														assign node31557 = (inp[9]) ? node31561 : node31558;
															assign node31558 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node31561 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node31564 = (inp[9]) ? node31572 : node31565;
															assign node31565 = (inp[0]) ? node31569 : node31566;
																assign node31566 = (inp[10]) ? 4'b1001 : 4'b1000;
																assign node31569 = (inp[10]) ? 4'b1000 : 4'b1001;
															assign node31572 = (inp[10]) ? node31574 : 4'b1000;
																assign node31574 = (inp[0]) ? 4'b1001 : 4'b1000;
												assign node31577 = (inp[9]) ? node31585 : node31578;
													assign node31578 = (inp[10]) ? 4'b1111 : node31579;
														assign node31579 = (inp[11]) ? 4'b1110 : node31580;
															assign node31580 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node31585 = (inp[10]) ? node31591 : node31586;
														assign node31586 = (inp[11]) ? 4'b1111 : node31587;
															assign node31587 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31591 = (inp[0]) ? node31593 : 4'b1110;
															assign node31593 = (inp[11]) ? 4'b1110 : 4'b1111;
										assign node31596 = (inp[4]) ? node31672 : node31597;
											assign node31597 = (inp[15]) ? node31635 : node31598;
												assign node31598 = (inp[9]) ? node31614 : node31599;
													assign node31599 = (inp[11]) ? node31609 : node31600;
														assign node31600 = (inp[10]) ? node31606 : node31601;
															assign node31601 = (inp[0]) ? 4'b1001 : node31602;
																assign node31602 = (inp[1]) ? 4'b1001 : 4'b1000;
															assign node31606 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node31609 = (inp[10]) ? 4'b1001 : node31610;
															assign node31610 = (inp[1]) ? 4'b1001 : 4'b1000;
													assign node31614 = (inp[11]) ? node31624 : node31615;
														assign node31615 = (inp[1]) ? 4'b1000 : node31616;
															assign node31616 = (inp[10]) ? node31620 : node31617;
																assign node31617 = (inp[0]) ? 4'b1000 : 4'b1001;
																assign node31620 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node31624 = (inp[10]) ? node31630 : node31625;
															assign node31625 = (inp[0]) ? node31627 : 4'b1001;
																assign node31627 = (inp[1]) ? 4'b1000 : 4'b1001;
															assign node31630 = (inp[0]) ? node31632 : 4'b1000;
																assign node31632 = (inp[1]) ? 4'b1001 : 4'b1000;
												assign node31635 = (inp[1]) ? node31653 : node31636;
													assign node31636 = (inp[9]) ? node31642 : node31637;
														assign node31637 = (inp[10]) ? node31639 : 4'b1100;
															assign node31639 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node31642 = (inp[10]) ? node31648 : node31643;
															assign node31643 = (inp[11]) ? 4'b1101 : node31644;
																assign node31644 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node31648 = (inp[0]) ? node31650 : 4'b1100;
																assign node31650 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node31653 = (inp[9]) ? node31663 : node31654;
														assign node31654 = (inp[0]) ? node31656 : 4'b1101;
															assign node31656 = (inp[11]) ? node31660 : node31657;
																assign node31657 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node31660 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node31663 = (inp[10]) ? node31667 : node31664;
															assign node31664 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node31667 = (inp[11]) ? 4'b1100 : node31668;
																assign node31668 = (inp[0]) ? 4'b1101 : 4'b1100;
											assign node31672 = (inp[15]) ? node31710 : node31673;
												assign node31673 = (inp[9]) ? node31691 : node31674;
													assign node31674 = (inp[10]) ? node31684 : node31675;
														assign node31675 = (inp[11]) ? node31679 : node31676;
															assign node31676 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node31679 = (inp[1]) ? 4'b1111 : node31680;
																assign node31680 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node31684 = (inp[11]) ? node31688 : node31685;
															assign node31685 = (inp[1]) ? 4'b1111 : 4'b1110;
															assign node31688 = (inp[1]) ? 4'b1110 : 4'b1111;
													assign node31691 = (inp[10]) ? node31701 : node31692;
														assign node31692 = (inp[11]) ? node31698 : node31693;
															assign node31693 = (inp[1]) ? node31695 : 4'b1110;
																assign node31695 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node31698 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31701 = (inp[1]) ? node31707 : node31702;
															assign node31702 = (inp[11]) ? node31704 : 4'b1111;
																assign node31704 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node31707 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node31710 = (inp[9]) ? node31722 : node31711;
													assign node31711 = (inp[10]) ? node31717 : node31712;
														assign node31712 = (inp[11]) ? 4'b1100 : node31713;
															assign node31713 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node31717 = (inp[11]) ? 4'b1101 : node31718;
															assign node31718 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node31722 = (inp[10]) ? node31728 : node31723;
														assign node31723 = (inp[11]) ? 4'b1101 : node31724;
															assign node31724 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node31728 = (inp[11]) ? 4'b1100 : 4'b1101;
							assign node31731 = (inp[12]) ? node32167 : node31732;
								assign node31732 = (inp[15]) ? node31942 : node31733;
									assign node31733 = (inp[7]) ? node31857 : node31734;
										assign node31734 = (inp[1]) ? node31796 : node31735;
											assign node31735 = (inp[10]) ? node31769 : node31736;
												assign node31736 = (inp[4]) ? node31756 : node31737;
													assign node31737 = (inp[2]) ? node31745 : node31738;
														assign node31738 = (inp[0]) ? node31740 : 4'b1101;
															assign node31740 = (inp[9]) ? 4'b1100 : node31741;
																assign node31741 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node31745 = (inp[0]) ? node31751 : node31746;
															assign node31746 = (inp[9]) ? 4'b1100 : node31747;
																assign node31747 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node31751 = (inp[11]) ? 4'b1101 : node31752;
																assign node31752 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node31756 = (inp[0]) ? 4'b1101 : node31757;
														assign node31757 = (inp[2]) ? node31763 : node31758;
															assign node31758 = (inp[9]) ? node31760 : 4'b1101;
																assign node31760 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node31763 = (inp[11]) ? 4'b1100 : node31764;
																assign node31764 = (inp[9]) ? 4'b1101 : 4'b1100;
												assign node31769 = (inp[0]) ? node31777 : node31770;
													assign node31770 = (inp[9]) ? node31774 : node31771;
														assign node31771 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node31774 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node31777 = (inp[11]) ? node31787 : node31778;
														assign node31778 = (inp[9]) ? node31780 : 4'b1100;
															assign node31780 = (inp[4]) ? node31784 : node31781;
																assign node31781 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node31784 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node31787 = (inp[4]) ? node31789 : 4'b1101;
															assign node31789 = (inp[9]) ? node31793 : node31790;
																assign node31790 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node31793 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node31796 = (inp[4]) ? node31836 : node31797;
												assign node31797 = (inp[0]) ? node31821 : node31798;
													assign node31798 = (inp[10]) ? node31812 : node31799;
														assign node31799 = (inp[2]) ? node31805 : node31800;
															assign node31800 = (inp[9]) ? node31802 : 4'b1000;
																assign node31802 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node31805 = (inp[9]) ? node31809 : node31806;
																assign node31806 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node31809 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node31812 = (inp[9]) ? 4'b1000 : node31813;
															assign node31813 = (inp[2]) ? node31817 : node31814;
																assign node31814 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node31817 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node31821 = (inp[2]) ? node31829 : node31822;
														assign node31822 = (inp[9]) ? node31826 : node31823;
															assign node31823 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node31826 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node31829 = (inp[11]) ? node31833 : node31830;
															assign node31830 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node31833 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node31836 = (inp[9]) ? node31846 : node31837;
													assign node31837 = (inp[11]) ? node31841 : node31838;
														assign node31838 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node31841 = (inp[0]) ? 4'b1101 : node31842;
															assign node31842 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node31846 = (inp[11]) ? node31852 : node31847;
														assign node31847 = (inp[0]) ? 4'b1101 : node31848;
															assign node31848 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node31852 = (inp[0]) ? 4'b1100 : node31853;
															assign node31853 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node31857 = (inp[1]) ? node31897 : node31858;
											assign node31858 = (inp[4]) ? node31880 : node31859;
												assign node31859 = (inp[11]) ? node31871 : node31860;
													assign node31860 = (inp[9]) ? node31866 : node31861;
														assign node31861 = (inp[2]) ? 4'b1111 : node31862;
															assign node31862 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31866 = (inp[0]) ? node31868 : 4'b1110;
															assign node31868 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node31871 = (inp[2]) ? node31877 : node31872;
														assign node31872 = (inp[9]) ? node31874 : 4'b1111;
															assign node31874 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31877 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node31880 = (inp[9]) ? node31886 : node31881;
													assign node31881 = (inp[11]) ? 4'b1010 : node31882;
														assign node31882 = (inp[0]) ? 4'b1011 : 4'b1010;
													assign node31886 = (inp[11]) ? node31892 : node31887;
														assign node31887 = (inp[0]) ? 4'b1010 : node31888;
															assign node31888 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node31892 = (inp[0]) ? 4'b1011 : node31893;
															assign node31893 = (inp[2]) ? 4'b1011 : 4'b1010;
											assign node31897 = (inp[2]) ? node31919 : node31898;
												assign node31898 = (inp[9]) ? node31910 : node31899;
													assign node31899 = (inp[11]) ? node31905 : node31900;
														assign node31900 = (inp[0]) ? 4'b1111 : node31901;
															assign node31901 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node31905 = (inp[0]) ? 4'b1110 : node31906;
															assign node31906 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node31910 = (inp[11]) ? node31916 : node31911;
														assign node31911 = (inp[0]) ? 4'b1110 : node31912;
															assign node31912 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node31916 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node31919 = (inp[11]) ? node31931 : node31920;
													assign node31920 = (inp[9]) ? node31926 : node31921;
														assign node31921 = (inp[0]) ? 4'b1111 : node31922;
															assign node31922 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node31926 = (inp[4]) ? 4'b1110 : node31927;
															assign node31927 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node31931 = (inp[9]) ? node31937 : node31932;
														assign node31932 = (inp[4]) ? 4'b1110 : node31933;
															assign node31933 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31937 = (inp[4]) ? 4'b1111 : node31938;
															assign node31938 = (inp[0]) ? 4'b1111 : 4'b1110;
									assign node31942 = (inp[7]) ? node32032 : node31943;
										assign node31943 = (inp[9]) ? node31989 : node31944;
											assign node31944 = (inp[0]) ? node31962 : node31945;
												assign node31945 = (inp[11]) ? node31953 : node31946;
													assign node31946 = (inp[4]) ? node31950 : node31947;
														assign node31947 = (inp[1]) ? 4'b1011 : 4'b1110;
														assign node31950 = (inp[1]) ? 4'b1111 : 4'b1011;
													assign node31953 = (inp[1]) ? node31959 : node31954;
														assign node31954 = (inp[4]) ? node31956 : 4'b1111;
															assign node31956 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node31959 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node31962 = (inp[11]) ? node31976 : node31963;
													assign node31963 = (inp[1]) ? node31969 : node31964;
														assign node31964 = (inp[4]) ? 4'b1010 : node31965;
															assign node31965 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node31969 = (inp[4]) ? node31973 : node31970;
															assign node31970 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node31973 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node31976 = (inp[2]) ? node31984 : node31977;
														assign node31977 = (inp[1]) ? node31981 : node31978;
															assign node31978 = (inp[4]) ? 4'b1011 : 4'b1110;
															assign node31981 = (inp[4]) ? 4'b1110 : 4'b1011;
														assign node31984 = (inp[4]) ? node31986 : 4'b1111;
															assign node31986 = (inp[1]) ? 4'b1111 : 4'b1011;
											assign node31989 = (inp[11]) ? node32013 : node31990;
												assign node31990 = (inp[1]) ? node32002 : node31991;
													assign node31991 = (inp[4]) ? node31997 : node31992;
														assign node31992 = (inp[2]) ? 4'b1111 : node31993;
															assign node31993 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node31997 = (inp[0]) ? 4'b1011 : node31998;
															assign node31998 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node32002 = (inp[4]) ? node32008 : node32003;
														assign node32003 = (inp[2]) ? 4'b1010 : node32004;
															assign node32004 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node32008 = (inp[2]) ? node32010 : 4'b1110;
															assign node32010 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node32013 = (inp[1]) ? node32021 : node32014;
													assign node32014 = (inp[4]) ? node32016 : 4'b1110;
														assign node32016 = (inp[2]) ? 4'b1010 : node32017;
															assign node32017 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node32021 = (inp[4]) ? node32027 : node32022;
														assign node32022 = (inp[2]) ? 4'b1011 : node32023;
															assign node32023 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node32027 = (inp[2]) ? node32029 : 4'b1111;
															assign node32029 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node32032 = (inp[0]) ? node32096 : node32033;
											assign node32033 = (inp[11]) ? node32061 : node32034;
												assign node32034 = (inp[9]) ? node32048 : node32035;
													assign node32035 = (inp[2]) ? node32043 : node32036;
														assign node32036 = (inp[1]) ? node32040 : node32037;
															assign node32037 = (inp[4]) ? 4'b1000 : 4'b1101;
															assign node32040 = (inp[4]) ? 4'b1101 : 4'b1000;
														assign node32043 = (inp[10]) ? node32045 : 4'b1100;
															assign node32045 = (inp[1]) ? 4'b1100 : 4'b1000;
													assign node32048 = (inp[1]) ? node32054 : node32049;
														assign node32049 = (inp[4]) ? 4'b1001 : node32050;
															assign node32050 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node32054 = (inp[4]) ? node32058 : node32055;
															assign node32055 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node32058 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node32061 = (inp[10]) ? node32081 : node32062;
													assign node32062 = (inp[2]) ? node32074 : node32063;
														assign node32063 = (inp[1]) ? node32069 : node32064;
															assign node32064 = (inp[4]) ? node32066 : 4'b1101;
																assign node32066 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node32069 = (inp[4]) ? 4'b1100 : node32070;
																assign node32070 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node32074 = (inp[9]) ? 4'b1100 : node32075;
															assign node32075 = (inp[1]) ? node32077 : 4'b1101;
																assign node32077 = (inp[4]) ? 4'b1101 : 4'b1000;
													assign node32081 = (inp[1]) ? node32087 : node32082;
														assign node32082 = (inp[2]) ? 4'b1100 : node32083;
															assign node32083 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node32087 = (inp[4]) ? node32089 : 4'b1001;
															assign node32089 = (inp[9]) ? node32093 : node32090;
																assign node32090 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node32093 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node32096 = (inp[10]) ? node32134 : node32097;
												assign node32097 = (inp[9]) ? node32115 : node32098;
													assign node32098 = (inp[11]) ? node32108 : node32099;
														assign node32099 = (inp[1]) ? node32105 : node32100;
															assign node32100 = (inp[4]) ? node32102 : 4'b1101;
																assign node32102 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node32105 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node32108 = (inp[1]) ? node32112 : node32109;
															assign node32109 = (inp[4]) ? 4'b1001 : 4'b1100;
															assign node32112 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node32115 = (inp[11]) ? node32125 : node32116;
														assign node32116 = (inp[1]) ? node32122 : node32117;
															assign node32117 = (inp[2]) ? node32119 : 4'b1001;
																assign node32119 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node32122 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node32125 = (inp[1]) ? node32131 : node32126;
															assign node32126 = (inp[4]) ? node32128 : 4'b1101;
																assign node32128 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node32131 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node32134 = (inp[4]) ? node32150 : node32135;
													assign node32135 = (inp[1]) ? node32143 : node32136;
														assign node32136 = (inp[9]) ? node32140 : node32137;
															assign node32137 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node32140 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node32143 = (inp[9]) ? node32147 : node32144;
															assign node32144 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node32147 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node32150 = (inp[1]) ? node32164 : node32151;
														assign node32151 = (inp[9]) ? node32159 : node32152;
															assign node32152 = (inp[2]) ? node32156 : node32153;
																assign node32153 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node32156 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node32159 = (inp[11]) ? 4'b1000 : node32160;
																assign node32160 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node32164 = (inp[9]) ? 4'b1101 : 4'b1100;
								assign node32167 = (inp[15]) ? node32393 : node32168;
									assign node32168 = (inp[7]) ? node32264 : node32169;
										assign node32169 = (inp[4]) ? node32215 : node32170;
											assign node32170 = (inp[11]) ? node32194 : node32171;
												assign node32171 = (inp[2]) ? node32183 : node32172;
													assign node32172 = (inp[9]) ? node32178 : node32173;
														assign node32173 = (inp[1]) ? 4'b1101 : node32174;
															assign node32174 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node32178 = (inp[1]) ? 4'b1100 : node32179;
															assign node32179 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node32183 = (inp[9]) ? node32189 : node32184;
														assign node32184 = (inp[1]) ? node32186 : 4'b1100;
															assign node32186 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node32189 = (inp[1]) ? node32191 : 4'b1101;
															assign node32191 = (inp[0]) ? 4'b1100 : 4'b1101;
												assign node32194 = (inp[0]) ? node32204 : node32195;
													assign node32195 = (inp[9]) ? node32199 : node32196;
														assign node32196 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node32199 = (inp[2]) ? 4'b1100 : node32200;
															assign node32200 = (inp[1]) ? 4'b1101 : 4'b1100;
													assign node32204 = (inp[9]) ? node32210 : node32205;
														assign node32205 = (inp[2]) ? node32207 : 4'b1100;
															assign node32207 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node32210 = (inp[1]) ? 4'b1101 : node32211;
															assign node32211 = (inp[10]) ? 4'b1101 : 4'b1100;
											assign node32215 = (inp[1]) ? node32247 : node32216;
												assign node32216 = (inp[0]) ? node32240 : node32217;
													assign node32217 = (inp[9]) ? node32225 : node32218;
														assign node32218 = (inp[11]) ? node32222 : node32219;
															assign node32219 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node32222 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node32225 = (inp[10]) ? node32233 : node32226;
															assign node32226 = (inp[11]) ? node32230 : node32227;
																assign node32227 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node32230 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node32233 = (inp[2]) ? node32237 : node32234;
																assign node32234 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node32237 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node32240 = (inp[11]) ? node32244 : node32241;
														assign node32241 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node32244 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node32247 = (inp[2]) ? node32255 : node32248;
													assign node32248 = (inp[9]) ? node32252 : node32249;
														assign node32249 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node32252 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node32255 = (inp[11]) ? 4'b1000 : node32256;
														assign node32256 = (inp[0]) ? node32260 : node32257;
															assign node32257 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node32260 = (inp[9]) ? 4'b1000 : 4'b1001;
										assign node32264 = (inp[1]) ? node32328 : node32265;
											assign node32265 = (inp[4]) ? node32307 : node32266;
												assign node32266 = (inp[2]) ? node32288 : node32267;
													assign node32267 = (inp[10]) ? node32281 : node32268;
														assign node32268 = (inp[9]) ? node32276 : node32269;
															assign node32269 = (inp[11]) ? node32273 : node32270;
																assign node32270 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node32273 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node32276 = (inp[0]) ? 4'b1010 : node32277;
																assign node32277 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node32281 = (inp[11]) ? node32283 : 4'b1010;
															assign node32283 = (inp[0]) ? 4'b1010 : node32284;
																assign node32284 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node32288 = (inp[10]) ? node32294 : node32289;
														assign node32289 = (inp[0]) ? 4'b1010 : node32290;
															assign node32290 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node32294 = (inp[0]) ? node32302 : node32295;
															assign node32295 = (inp[11]) ? node32299 : node32296;
																assign node32296 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node32299 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node32302 = (inp[9]) ? node32304 : 4'b1011;
																assign node32304 = (inp[11]) ? 4'b1010 : 4'b1011;
												assign node32307 = (inp[2]) ? node32313 : node32308;
													assign node32308 = (inp[11]) ? 4'b1111 : node32309;
														assign node32309 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node32313 = (inp[0]) ? node32321 : node32314;
														assign node32314 = (inp[11]) ? node32318 : node32315;
															assign node32315 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node32318 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node32321 = (inp[11]) ? node32325 : node32322;
															assign node32322 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node32325 = (inp[9]) ? 4'b1111 : 4'b1110;
											assign node32328 = (inp[10]) ? node32360 : node32329;
												assign node32329 = (inp[11]) ? node32347 : node32330;
													assign node32330 = (inp[9]) ? node32338 : node32331;
														assign node32331 = (inp[2]) ? 4'b1111 : node32332;
															assign node32332 = (inp[4]) ? node32334 : 4'b1110;
																assign node32334 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node32338 = (inp[2]) ? 4'b1110 : node32339;
															assign node32339 = (inp[0]) ? node32343 : node32340;
																assign node32340 = (inp[4]) ? 4'b1111 : 4'b1110;
																assign node32343 = (inp[4]) ? 4'b1110 : 4'b1111;
													assign node32347 = (inp[0]) ? node32353 : node32348;
														assign node32348 = (inp[4]) ? 4'b1111 : node32349;
															assign node32349 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node32353 = (inp[4]) ? 4'b1110 : node32354;
															assign node32354 = (inp[2]) ? 4'b1110 : node32355;
																assign node32355 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node32360 = (inp[11]) ? node32376 : node32361;
													assign node32361 = (inp[9]) ? node32369 : node32362;
														assign node32362 = (inp[2]) ? 4'b1111 : node32363;
															assign node32363 = (inp[0]) ? 4'b1110 : node32364;
																assign node32364 = (inp[4]) ? 4'b1110 : 4'b1111;
														assign node32369 = (inp[2]) ? 4'b1110 : node32370;
															assign node32370 = (inp[4]) ? node32372 : 4'b1110;
																assign node32372 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node32376 = (inp[9]) ? node32384 : node32377;
														assign node32377 = (inp[2]) ? 4'b1110 : node32378;
															assign node32378 = (inp[0]) ? 4'b1111 : node32379;
																assign node32379 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node32384 = (inp[2]) ? 4'b1111 : node32385;
															assign node32385 = (inp[4]) ? node32389 : node32386;
																assign node32386 = (inp[0]) ? 4'b1110 : 4'b1111;
																assign node32389 = (inp[0]) ? 4'b1111 : 4'b1110;
									assign node32393 = (inp[7]) ? node32491 : node32394;
										assign node32394 = (inp[2]) ? node32458 : node32395;
											assign node32395 = (inp[0]) ? node32437 : node32396;
												assign node32396 = (inp[4]) ? node32422 : node32397;
													assign node32397 = (inp[1]) ? node32413 : node32398;
														assign node32398 = (inp[10]) ? node32406 : node32399;
															assign node32399 = (inp[11]) ? node32403 : node32400;
																assign node32400 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node32403 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node32406 = (inp[11]) ? node32410 : node32407;
																assign node32407 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node32410 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node32413 = (inp[10]) ? node32417 : node32414;
															assign node32414 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node32417 = (inp[11]) ? node32419 : 4'b1111;
																assign node32419 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node32422 = (inp[1]) ? node32430 : node32423;
														assign node32423 = (inp[11]) ? node32427 : node32424;
															assign node32424 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node32427 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node32430 = (inp[10]) ? node32434 : node32431;
															assign node32431 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node32434 = (inp[11]) ? 4'b1111 : 4'b1110;
												assign node32437 = (inp[11]) ? node32451 : node32438;
													assign node32438 = (inp[1]) ? node32446 : node32439;
														assign node32439 = (inp[4]) ? node32443 : node32440;
															assign node32440 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node32443 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node32446 = (inp[9]) ? node32448 : 4'b1111;
															assign node32448 = (inp[4]) ? 4'b1111 : 4'b1110;
													assign node32451 = (inp[9]) ? node32455 : node32452;
														assign node32452 = (inp[4]) ? 4'b1111 : 4'b1110;
														assign node32455 = (inp[4]) ? 4'b1110 : 4'b1111;
											assign node32458 = (inp[4]) ? node32466 : node32459;
												assign node32459 = (inp[11]) ? node32463 : node32460;
													assign node32460 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node32463 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node32466 = (inp[1]) ? node32476 : node32467;
													assign node32467 = (inp[10]) ? 4'b1110 : node32468;
														assign node32468 = (inp[9]) ? node32472 : node32469;
															assign node32469 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node32472 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node32476 = (inp[10]) ? node32484 : node32477;
														assign node32477 = (inp[11]) ? node32481 : node32478;
															assign node32478 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node32481 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node32484 = (inp[11]) ? node32488 : node32485;
															assign node32485 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node32488 = (inp[9]) ? 4'b1110 : 4'b1111;
										assign node32491 = (inp[0]) ? node32515 : node32492;
											assign node32492 = (inp[11]) ? node32504 : node32493;
												assign node32493 = (inp[9]) ? node32499 : node32494;
													assign node32494 = (inp[4]) ? node32496 : 4'b1100;
														assign node32496 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node32499 = (inp[4]) ? node32501 : 4'b1101;
														assign node32501 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node32504 = (inp[9]) ? node32510 : node32505;
													assign node32505 = (inp[4]) ? node32507 : 4'b1101;
														assign node32507 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node32510 = (inp[4]) ? node32512 : 4'b1100;
														assign node32512 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node32515 = (inp[9]) ? node32527 : node32516;
												assign node32516 = (inp[11]) ? node32522 : node32517;
													assign node32517 = (inp[2]) ? 4'b1100 : node32518;
														assign node32518 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node32522 = (inp[2]) ? 4'b1101 : node32523;
														assign node32523 = (inp[4]) ? 4'b1101 : 4'b1100;
												assign node32527 = (inp[11]) ? node32533 : node32528;
													assign node32528 = (inp[2]) ? 4'b1101 : node32529;
														assign node32529 = (inp[4]) ? 4'b1101 : 4'b1100;
													assign node32533 = (inp[2]) ? 4'b1100 : node32534;
														assign node32534 = (inp[4]) ? 4'b1100 : 4'b1101;
						assign node32538 = (inp[6]) ? node33626 : node32539;
							assign node32539 = (inp[2]) ? node33095 : node32540;
								assign node32540 = (inp[12]) ? node32816 : node32541;
									assign node32541 = (inp[7]) ? node32673 : node32542;
										assign node32542 = (inp[4]) ? node32618 : node32543;
											assign node32543 = (inp[10]) ? node32579 : node32544;
												assign node32544 = (inp[1]) ? node32558 : node32545;
													assign node32545 = (inp[9]) ? node32551 : node32546;
														assign node32546 = (inp[15]) ? 4'b1101 : node32547;
															assign node32547 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node32551 = (inp[15]) ? 4'b1100 : node32552;
															assign node32552 = (inp[11]) ? node32554 : 4'b1101;
																assign node32554 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node32558 = (inp[11]) ? node32570 : node32559;
														assign node32559 = (inp[9]) ? node32565 : node32560;
															assign node32560 = (inp[0]) ? 4'b1100 : node32561;
																assign node32561 = (inp[15]) ? 4'b1100 : 4'b1101;
															assign node32565 = (inp[0]) ? 4'b1101 : node32566;
																assign node32566 = (inp[15]) ? 4'b1101 : 4'b1100;
														assign node32570 = (inp[9]) ? node32574 : node32571;
															assign node32571 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node32574 = (inp[0]) ? node32576 : 4'b1100;
																assign node32576 = (inp[15]) ? 4'b1101 : 4'b1100;
												assign node32579 = (inp[15]) ? node32601 : node32580;
													assign node32580 = (inp[11]) ? node32590 : node32581;
														assign node32581 = (inp[9]) ? node32587 : node32582;
															assign node32582 = (inp[0]) ? 4'b1101 : node32583;
																assign node32583 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node32587 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node32590 = (inp[9]) ? node32596 : node32591;
															assign node32591 = (inp[1]) ? 4'b1100 : node32592;
																assign node32592 = (inp[0]) ? 4'b1101 : 4'b1100;
															assign node32596 = (inp[1]) ? 4'b1101 : node32597;
																assign node32597 = (inp[0]) ? 4'b1100 : 4'b1101;
													assign node32601 = (inp[9]) ? node32607 : node32602;
														assign node32602 = (inp[1]) ? 4'b1101 : node32603;
															assign node32603 = (inp[11]) ? 4'b1101 : 4'b1100;
														assign node32607 = (inp[1]) ? node32613 : node32608;
															assign node32608 = (inp[0]) ? 4'b1101 : node32609;
																assign node32609 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node32613 = (inp[11]) ? node32615 : 4'b1100;
																assign node32615 = (inp[0]) ? 4'b1100 : 4'b1101;
											assign node32618 = (inp[15]) ? node32638 : node32619;
												assign node32619 = (inp[10]) ? node32629 : node32620;
													assign node32620 = (inp[9]) ? node32624 : node32621;
														assign node32621 = (inp[1]) ? 4'b1111 : 4'b1110;
														assign node32624 = (inp[0]) ? node32626 : 4'b1110;
															assign node32626 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node32629 = (inp[11]) ? 4'b1111 : node32630;
														assign node32630 = (inp[9]) ? node32632 : 4'b1110;
															assign node32632 = (inp[1]) ? 4'b1111 : node32633;
																assign node32633 = (inp[0]) ? 4'b1110 : 4'b1111;
												assign node32638 = (inp[0]) ? node32662 : node32639;
													assign node32639 = (inp[10]) ? node32655 : node32640;
														assign node32640 = (inp[1]) ? node32648 : node32641;
															assign node32641 = (inp[9]) ? node32645 : node32642;
																assign node32642 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node32645 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node32648 = (inp[9]) ? node32652 : node32649;
																assign node32649 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node32652 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node32655 = (inp[1]) ? 4'b1001 : node32656;
															assign node32656 = (inp[9]) ? 4'b1001 : node32657;
																assign node32657 = (inp[11]) ? 4'b1000 : 4'b1001;
													assign node32662 = (inp[10]) ? 4'b1000 : node32663;
														assign node32663 = (inp[11]) ? 4'b1001 : node32664;
															assign node32664 = (inp[1]) ? node32668 : node32665;
																assign node32665 = (inp[9]) ? 4'b1001 : 4'b1000;
																assign node32668 = (inp[9]) ? 4'b1000 : 4'b1001;
										assign node32673 = (inp[4]) ? node32745 : node32674;
											assign node32674 = (inp[15]) ? node32714 : node32675;
												assign node32675 = (inp[1]) ? node32693 : node32676;
													assign node32676 = (inp[0]) ? node32684 : node32677;
														assign node32677 = (inp[9]) ? node32681 : node32678;
															assign node32678 = (inp[10]) ? 4'b1011 : 4'b1010;
															assign node32681 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node32684 = (inp[11]) ? node32686 : 4'b1010;
															assign node32686 = (inp[9]) ? node32690 : node32687;
																assign node32687 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node32690 = (inp[10]) ? 4'b1010 : 4'b1011;
													assign node32693 = (inp[0]) ? node32701 : node32694;
														assign node32694 = (inp[9]) ? node32698 : node32695;
															assign node32695 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node32698 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node32701 = (inp[10]) ? node32709 : node32702;
															assign node32702 = (inp[9]) ? node32706 : node32703;
																assign node32703 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node32706 = (inp[11]) ? 4'b1111 : 4'b1110;
															assign node32709 = (inp[11]) ? node32711 : 4'b1111;
																assign node32711 = (inp[9]) ? 4'b1110 : 4'b1111;
												assign node32714 = (inp[1]) ? node32730 : node32715;
													assign node32715 = (inp[10]) ? node32725 : node32716;
														assign node32716 = (inp[9]) ? node32720 : node32717;
															assign node32717 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node32720 = (inp[11]) ? 4'b1110 : node32721;
																assign node32721 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node32725 = (inp[9]) ? 4'b1111 : node32726;
															assign node32726 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node32730 = (inp[11]) ? node32740 : node32731;
														assign node32731 = (inp[0]) ? node32733 : 4'b1010;
															assign node32733 = (inp[10]) ? node32737 : node32734;
																assign node32734 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node32737 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node32740 = (inp[10]) ? node32742 : 4'b1011;
															assign node32742 = (inp[9]) ? 4'b1010 : 4'b1011;
											assign node32745 = (inp[15]) ? node32785 : node32746;
												assign node32746 = (inp[1]) ? node32762 : node32747;
													assign node32747 = (inp[11]) ? node32755 : node32748;
														assign node32748 = (inp[10]) ? node32752 : node32749;
															assign node32749 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node32752 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node32755 = (inp[0]) ? node32757 : 4'b1000;
															assign node32757 = (inp[10]) ? 4'b1000 : node32758;
																assign node32758 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node32762 = (inp[0]) ? node32778 : node32763;
														assign node32763 = (inp[11]) ? node32771 : node32764;
															assign node32764 = (inp[9]) ? node32768 : node32765;
																assign node32765 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node32768 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node32771 = (inp[9]) ? node32775 : node32772;
																assign node32772 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node32775 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node32778 = (inp[11]) ? 4'b1001 : node32779;
															assign node32779 = (inp[9]) ? node32781 : 4'b1001;
																assign node32781 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node32785 = (inp[1]) ? node32799 : node32786;
													assign node32786 = (inp[9]) ? node32794 : node32787;
														assign node32787 = (inp[10]) ? node32789 : 4'b1010;
															assign node32789 = (inp[0]) ? node32791 : 4'b1011;
																assign node32791 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node32794 = (inp[10]) ? 4'b1010 : node32795;
															assign node32795 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node32799 = (inp[11]) ? node32807 : node32800;
														assign node32800 = (inp[9]) ? node32804 : node32801;
															assign node32801 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node32804 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node32807 = (inp[9]) ? node32809 : 4'b1111;
															assign node32809 = (inp[10]) ? node32813 : node32810;
																assign node32810 = (inp[0]) ? 4'b1111 : 4'b1110;
																assign node32813 = (inp[0]) ? 4'b1110 : 4'b1111;
									assign node32816 = (inp[7]) ? node32952 : node32817;
										assign node32817 = (inp[4]) ? node32887 : node32818;
											assign node32818 = (inp[11]) ? node32840 : node32819;
												assign node32819 = (inp[15]) ? node32833 : node32820;
													assign node32820 = (inp[1]) ? node32828 : node32821;
														assign node32821 = (inp[9]) ? node32825 : node32822;
															assign node32822 = (inp[10]) ? 4'b1111 : 4'b1110;
															assign node32825 = (inp[10]) ? 4'b1110 : 4'b1111;
														assign node32828 = (inp[0]) ? 4'b1111 : node32829;
															assign node32829 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node32833 = (inp[10]) ? node32837 : node32834;
														assign node32834 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node32837 = (inp[9]) ? 4'b1111 : 4'b1110;
												assign node32840 = (inp[9]) ? node32862 : node32841;
													assign node32841 = (inp[10]) ? node32851 : node32842;
														assign node32842 = (inp[15]) ? node32848 : node32843;
															assign node32843 = (inp[0]) ? 4'b1110 : node32844;
																assign node32844 = (inp[1]) ? 4'b1110 : 4'b1111;
															assign node32848 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node32851 = (inp[1]) ? node32857 : node32852;
															assign node32852 = (inp[15]) ? 4'b1111 : node32853;
																assign node32853 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node32857 = (inp[15]) ? node32859 : 4'b1111;
																assign node32859 = (inp[0]) ? 4'b1110 : 4'b1111;
													assign node32862 = (inp[1]) ? node32878 : node32863;
														assign node32863 = (inp[15]) ? node32871 : node32864;
															assign node32864 = (inp[0]) ? node32868 : node32865;
																assign node32865 = (inp[10]) ? 4'b1111 : 4'b1110;
																assign node32868 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node32871 = (inp[0]) ? node32875 : node32872;
																assign node32872 = (inp[10]) ? 4'b1110 : 4'b1111;
																assign node32875 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node32878 = (inp[10]) ? node32882 : node32879;
															assign node32879 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node32882 = (inp[15]) ? node32884 : 4'b1110;
																assign node32884 = (inp[0]) ? 4'b1111 : 4'b1110;
											assign node32887 = (inp[15]) ? node32923 : node32888;
												assign node32888 = (inp[1]) ? node32904 : node32889;
													assign node32889 = (inp[11]) ? node32895 : node32890;
														assign node32890 = (inp[9]) ? 4'b1101 : node32891;
															assign node32891 = (inp[10]) ? 4'b1100 : 4'b1101;
														assign node32895 = (inp[0]) ? node32897 : 4'b1100;
															assign node32897 = (inp[9]) ? node32901 : node32898;
																assign node32898 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node32901 = (inp[10]) ? 4'b1101 : 4'b1100;
													assign node32904 = (inp[11]) ? node32912 : node32905;
														assign node32905 = (inp[9]) ? 4'b1000 : node32906;
															assign node32906 = (inp[0]) ? 4'b1000 : node32907;
																assign node32907 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node32912 = (inp[0]) ? node32918 : node32913;
															assign node32913 = (inp[10]) ? node32915 : 4'b1001;
																assign node32915 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node32918 = (inp[9]) ? 4'b1000 : node32919;
																assign node32919 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node32923 = (inp[11]) ? node32933 : node32924;
													assign node32924 = (inp[0]) ? 4'b1111 : node32925;
														assign node32925 = (inp[10]) ? node32929 : node32926;
															assign node32926 = (inp[9]) ? 4'b1111 : 4'b1110;
															assign node32929 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node32933 = (inp[9]) ? node32941 : node32934;
														assign node32934 = (inp[10]) ? node32938 : node32935;
															assign node32935 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node32938 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node32941 = (inp[1]) ? node32947 : node32942;
															assign node32942 = (inp[0]) ? node32944 : 4'b1111;
																assign node32944 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node32947 = (inp[10]) ? node32949 : 4'b1110;
																assign node32949 = (inp[0]) ? 4'b1110 : 4'b1111;
										assign node32952 = (inp[15]) ? node33006 : node32953;
											assign node32953 = (inp[4]) ? node32979 : node32954;
												assign node32954 = (inp[9]) ? node32962 : node32955;
													assign node32955 = (inp[10]) ? 4'b1001 : node32956;
														assign node32956 = (inp[1]) ? node32958 : 4'b1000;
															assign node32958 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node32962 = (inp[10]) ? node32972 : node32963;
														assign node32963 = (inp[0]) ? node32967 : node32964;
															assign node32964 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node32967 = (inp[1]) ? node32969 : 4'b1001;
																assign node32969 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node32972 = (inp[1]) ? 4'b1000 : node32973;
															assign node32973 = (inp[0]) ? 4'b1000 : node32974;
																assign node32974 = (inp[11]) ? 4'b1001 : 4'b1000;
												assign node32979 = (inp[11]) ? node32993 : node32980;
													assign node32980 = (inp[9]) ? node32988 : node32981;
														assign node32981 = (inp[10]) ? 4'b1111 : node32982;
															assign node32982 = (inp[1]) ? 4'b1110 : node32983;
																assign node32983 = (inp[0]) ? 4'b1110 : 4'b1111;
														assign node32988 = (inp[10]) ? 4'b1110 : node32989;
															assign node32989 = (inp[1]) ? 4'b1111 : 4'b1110;
													assign node32993 = (inp[9]) ? node33001 : node32994;
														assign node32994 = (inp[1]) ? node32998 : node32995;
															assign node32995 = (inp[10]) ? 4'b1110 : 4'b1111;
															assign node32998 = (inp[10]) ? 4'b1111 : 4'b1110;
														assign node33001 = (inp[10]) ? 4'b1111 : node33002;
															assign node33002 = (inp[1]) ? 4'b1111 : 4'b1110;
											assign node33006 = (inp[1]) ? node33048 : node33007;
												assign node33007 = (inp[10]) ? node33027 : node33008;
													assign node33008 = (inp[4]) ? node33018 : node33009;
														assign node33009 = (inp[11]) ? node33011 : 4'b1100;
															assign node33011 = (inp[9]) ? node33015 : node33012;
																assign node33012 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node33015 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node33018 = (inp[9]) ? node33024 : node33019;
															assign node33019 = (inp[0]) ? 4'b1100 : node33020;
																assign node33020 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node33024 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node33027 = (inp[0]) ? node33041 : node33028;
														assign node33028 = (inp[4]) ? node33034 : node33029;
															assign node33029 = (inp[9]) ? node33031 : 4'b1101;
																assign node33031 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node33034 = (inp[11]) ? node33038 : node33035;
																assign node33035 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node33038 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node33041 = (inp[4]) ? node33045 : node33042;
															assign node33042 = (inp[9]) ? 4'b1101 : 4'b1100;
															assign node33045 = (inp[9]) ? 4'b1100 : 4'b1101;
												assign node33048 = (inp[9]) ? node33078 : node33049;
													assign node33049 = (inp[11]) ? node33065 : node33050;
														assign node33050 = (inp[0]) ? node33058 : node33051;
															assign node33051 = (inp[4]) ? node33055 : node33052;
																assign node33052 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node33055 = (inp[10]) ? 4'b1101 : 4'b1100;
															assign node33058 = (inp[4]) ? node33062 : node33059;
																assign node33059 = (inp[10]) ? 4'b1100 : 4'b1101;
																assign node33062 = (inp[10]) ? 4'b1101 : 4'b1100;
														assign node33065 = (inp[10]) ? node33073 : node33066;
															assign node33066 = (inp[4]) ? node33070 : node33067;
																assign node33067 = (inp[0]) ? 4'b1101 : 4'b1100;
																assign node33070 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node33073 = (inp[0]) ? 4'b1100 : node33074;
																assign node33074 = (inp[4]) ? 4'b1100 : 4'b1101;
													assign node33078 = (inp[10]) ? node33084 : node33079;
														assign node33079 = (inp[4]) ? 4'b1101 : node33080;
															assign node33080 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node33084 = (inp[4]) ? node33090 : node33085;
															assign node33085 = (inp[0]) ? 4'b1101 : node33086;
																assign node33086 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node33090 = (inp[0]) ? 4'b1100 : node33091;
																assign node33091 = (inp[11]) ? 4'b1101 : 4'b1100;
								assign node33095 = (inp[7]) ? node33339 : node33096;
									assign node33096 = (inp[12]) ? node33240 : node33097;
										assign node33097 = (inp[4]) ? node33169 : node33098;
											assign node33098 = (inp[0]) ? node33128 : node33099;
												assign node33099 = (inp[10]) ? node33115 : node33100;
													assign node33100 = (inp[9]) ? node33108 : node33101;
														assign node33101 = (inp[11]) ? node33103 : 4'b1001;
															assign node33103 = (inp[1]) ? node33105 : 4'b1001;
																assign node33105 = (inp[15]) ? 4'b1001 : 4'b1000;
														assign node33108 = (inp[1]) ? node33112 : node33109;
															assign node33109 = (inp[15]) ? 4'b1001 : 4'b1000;
															assign node33112 = (inp[15]) ? 4'b1000 : 4'b1001;
													assign node33115 = (inp[15]) ? node33121 : node33116;
														assign node33116 = (inp[9]) ? 4'b1001 : node33117;
															assign node33117 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node33121 = (inp[1]) ? node33125 : node33122;
															assign node33122 = (inp[9]) ? 4'b1000 : 4'b1001;
															assign node33125 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node33128 = (inp[11]) ? node33150 : node33129;
													assign node33129 = (inp[15]) ? node33141 : node33130;
														assign node33130 = (inp[10]) ? node33136 : node33131;
															assign node33131 = (inp[1]) ? 4'b1000 : node33132;
																assign node33132 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node33136 = (inp[9]) ? node33138 : 4'b1001;
																assign node33138 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node33141 = (inp[10]) ? 4'b1000 : node33142;
															assign node33142 = (inp[1]) ? node33146 : node33143;
																assign node33143 = (inp[9]) ? 4'b1000 : 4'b1001;
																assign node33146 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node33150 = (inp[15]) ? node33162 : node33151;
														assign node33151 = (inp[1]) ? node33157 : node33152;
															assign node33152 = (inp[10]) ? node33154 : 4'b1000;
																assign node33154 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node33157 = (inp[10]) ? node33159 : 4'b1001;
																assign node33159 = (inp[9]) ? 4'b1001 : 4'b1000;
														assign node33162 = (inp[1]) ? node33164 : 4'b1001;
															assign node33164 = (inp[10]) ? 4'b1000 : node33165;
																assign node33165 = (inp[9]) ? 4'b1000 : 4'b1001;
											assign node33169 = (inp[15]) ? node33205 : node33170;
												assign node33170 = (inp[0]) ? node33186 : node33171;
													assign node33171 = (inp[11]) ? node33179 : node33172;
														assign node33172 = (inp[1]) ? 4'b1011 : node33173;
															assign node33173 = (inp[10]) ? node33175 : 4'b1011;
																assign node33175 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node33179 = (inp[9]) ? node33183 : node33180;
															assign node33180 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node33183 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node33186 = (inp[11]) ? node33194 : node33187;
														assign node33187 = (inp[10]) ? node33191 : node33188;
															assign node33188 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node33191 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node33194 = (inp[10]) ? node33200 : node33195;
															assign node33195 = (inp[1]) ? 4'b1011 : node33196;
																assign node33196 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node33200 = (inp[1]) ? 4'b1010 : node33201;
																assign node33201 = (inp[9]) ? 4'b1010 : 4'b1011;
												assign node33205 = (inp[9]) ? node33221 : node33206;
													assign node33206 = (inp[10]) ? node33214 : node33207;
														assign node33207 = (inp[1]) ? 4'b1100 : node33208;
															assign node33208 = (inp[11]) ? node33210 : 4'b1101;
																assign node33210 = (inp[0]) ? 4'b1101 : 4'b1100;
														assign node33214 = (inp[1]) ? 4'b1101 : node33215;
															assign node33215 = (inp[0]) ? 4'b1100 : node33216;
																assign node33216 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node33221 = (inp[0]) ? node33229 : node33222;
														assign node33222 = (inp[11]) ? node33224 : 4'b1101;
															assign node33224 = (inp[10]) ? node33226 : 4'b1101;
																assign node33226 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node33229 = (inp[11]) ? node33235 : node33230;
															assign node33230 = (inp[1]) ? node33232 : 4'b1101;
																assign node33232 = (inp[10]) ? 4'b1100 : 4'b1101;
															assign node33235 = (inp[1]) ? 4'b1100 : node33236;
																assign node33236 = (inp[10]) ? 4'b1101 : 4'b1100;
										assign node33240 = (inp[15]) ? node33300 : node33241;
											assign node33241 = (inp[4]) ? node33269 : node33242;
												assign node33242 = (inp[11]) ? node33250 : node33243;
													assign node33243 = (inp[0]) ? node33245 : 4'b1011;
														assign node33245 = (inp[10]) ? 4'b1011 : node33246;
															assign node33246 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node33250 = (inp[10]) ? node33260 : node33251;
														assign node33251 = (inp[9]) ? node33257 : node33252;
															assign node33252 = (inp[1]) ? node33254 : 4'b1011;
																assign node33254 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node33257 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node33260 = (inp[9]) ? node33266 : node33261;
															assign node33261 = (inp[0]) ? node33263 : 4'b1010;
																assign node33263 = (inp[1]) ? 4'b1011 : 4'b1010;
															assign node33266 = (inp[0]) ? 4'b1010 : 4'b1011;
												assign node33269 = (inp[1]) ? node33285 : node33270;
													assign node33270 = (inp[0]) ? node33276 : node33271;
														assign node33271 = (inp[9]) ? 4'b1001 : node33272;
															assign node33272 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node33276 = (inp[10]) ? node33278 : 4'b1000;
															assign node33278 = (inp[9]) ? node33282 : node33279;
																assign node33279 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node33282 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node33285 = (inp[9]) ? node33289 : node33286;
														assign node33286 = (inp[0]) ? 4'b1100 : 4'b1101;
														assign node33289 = (inp[10]) ? node33295 : node33290;
															assign node33290 = (inp[11]) ? 4'b1101 : node33291;
																assign node33291 = (inp[0]) ? 4'b1100 : 4'b1101;
															assign node33295 = (inp[0]) ? node33297 : 4'b1100;
																assign node33297 = (inp[11]) ? 4'b1100 : 4'b1101;
											assign node33300 = (inp[0]) ? node33308 : node33301;
												assign node33301 = (inp[9]) ? node33305 : node33302;
													assign node33302 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node33305 = (inp[10]) ? 4'b1010 : 4'b1011;
												assign node33308 = (inp[9]) ? node33316 : node33309;
													assign node33309 = (inp[10]) ? node33313 : node33310;
														assign node33310 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node33313 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node33316 = (inp[4]) ? node33324 : node33317;
														assign node33317 = (inp[10]) ? node33321 : node33318;
															assign node33318 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node33321 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node33324 = (inp[1]) ? node33332 : node33325;
															assign node33325 = (inp[11]) ? node33329 : node33326;
																assign node33326 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node33329 = (inp[10]) ? 4'b1010 : 4'b1011;
															assign node33332 = (inp[10]) ? node33336 : node33333;
																assign node33333 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node33336 = (inp[11]) ? 4'b1010 : 4'b1011;
									assign node33339 = (inp[12]) ? node33507 : node33340;
										assign node33340 = (inp[4]) ? node33432 : node33341;
											assign node33341 = (inp[11]) ? node33389 : node33342;
												assign node33342 = (inp[15]) ? node33362 : node33343;
													assign node33343 = (inp[1]) ? node33357 : node33344;
														assign node33344 = (inp[0]) ? node33350 : node33345;
															assign node33345 = (inp[10]) ? node33347 : 4'b1111;
																assign node33347 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node33350 = (inp[10]) ? node33354 : node33351;
																assign node33351 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node33354 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node33357 = (inp[10]) ? node33359 : 4'b1011;
															assign node33359 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node33362 = (inp[1]) ? node33378 : node33363;
														assign node33363 = (inp[0]) ? node33371 : node33364;
															assign node33364 = (inp[10]) ? node33368 : node33365;
																assign node33365 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node33368 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node33371 = (inp[9]) ? node33375 : node33372;
																assign node33372 = (inp[10]) ? 4'b1010 : 4'b1011;
																assign node33375 = (inp[10]) ? 4'b1011 : 4'b1010;
														assign node33378 = (inp[0]) ? node33384 : node33379;
															assign node33379 = (inp[10]) ? node33381 : 4'b1110;
																assign node33381 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node33384 = (inp[9]) ? node33386 : 4'b1111;
																assign node33386 = (inp[10]) ? 4'b1111 : 4'b1110;
												assign node33389 = (inp[10]) ? node33415 : node33390;
													assign node33390 = (inp[9]) ? node33402 : node33391;
														assign node33391 = (inp[15]) ? node33397 : node33392;
															assign node33392 = (inp[1]) ? node33394 : 4'b1110;
																assign node33394 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node33397 = (inp[1]) ? 4'b1110 : node33398;
																assign node33398 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node33402 = (inp[0]) ? node33410 : node33403;
															assign node33403 = (inp[1]) ? node33407 : node33404;
																assign node33404 = (inp[15]) ? 4'b1011 : 4'b1111;
																assign node33407 = (inp[15]) ? 4'b1111 : 4'b1010;
															assign node33410 = (inp[1]) ? node33412 : 4'b1010;
																assign node33412 = (inp[15]) ? 4'b1111 : 4'b1011;
													assign node33415 = (inp[9]) ? node33425 : node33416;
														assign node33416 = (inp[1]) ? node33420 : node33417;
															assign node33417 = (inp[0]) ? 4'b1010 : 4'b1111;
															assign node33420 = (inp[15]) ? 4'b1111 : node33421;
																assign node33421 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node33425 = (inp[15]) ? 4'b1110 : node33426;
															assign node33426 = (inp[1]) ? node33428 : 4'b1110;
																assign node33428 = (inp[0]) ? 4'b1010 : 4'b1011;
											assign node33432 = (inp[15]) ? node33470 : node33433;
												assign node33433 = (inp[0]) ? node33447 : node33434;
													assign node33434 = (inp[9]) ? node33442 : node33435;
														assign node33435 = (inp[10]) ? node33437 : 4'b1100;
															assign node33437 = (inp[11]) ? 4'b1101 : node33438;
																assign node33438 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node33442 = (inp[10]) ? node33444 : 4'b1101;
															assign node33444 = (inp[11]) ? 4'b1100 : 4'b1101;
													assign node33447 = (inp[9]) ? node33459 : node33448;
														assign node33448 = (inp[10]) ? node33454 : node33449;
															assign node33449 = (inp[1]) ? node33451 : 4'b1101;
																assign node33451 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node33454 = (inp[11]) ? node33456 : 4'b1100;
																assign node33456 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node33459 = (inp[10]) ? node33465 : node33460;
															assign node33460 = (inp[1]) ? node33462 : 4'b1100;
																assign node33462 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node33465 = (inp[11]) ? node33467 : 4'b1101;
																assign node33467 = (inp[1]) ? 4'b1100 : 4'b1101;
												assign node33470 = (inp[1]) ? node33492 : node33471;
													assign node33471 = (inp[11]) ? node33485 : node33472;
														assign node33472 = (inp[10]) ? node33478 : node33473;
															assign node33473 = (inp[9]) ? node33475 : 4'b1110;
																assign node33475 = (inp[0]) ? 4'b1111 : 4'b1110;
															assign node33478 = (inp[0]) ? node33482 : node33479;
																assign node33479 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node33482 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node33485 = (inp[10]) ? node33489 : node33486;
															assign node33486 = (inp[9]) ? 4'b1110 : 4'b1111;
															assign node33489 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node33492 = (inp[10]) ? node33502 : node33493;
														assign node33493 = (inp[0]) ? node33495 : 4'b1010;
															assign node33495 = (inp[11]) ? node33499 : node33496;
																assign node33496 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node33499 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node33502 = (inp[9]) ? node33504 : 4'b1011;
															assign node33504 = (inp[11]) ? 4'b1010 : 4'b1011;
										assign node33507 = (inp[15]) ? node33581 : node33508;
											assign node33508 = (inp[4]) ? node33546 : node33509;
												assign node33509 = (inp[10]) ? node33529 : node33510;
													assign node33510 = (inp[9]) ? node33522 : node33511;
														assign node33511 = (inp[11]) ? node33517 : node33512;
															assign node33512 = (inp[0]) ? node33514 : 4'b1100;
																assign node33514 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node33517 = (inp[0]) ? 4'b1100 : node33518;
																assign node33518 = (inp[1]) ? 4'b1100 : 4'b1101;
														assign node33522 = (inp[0]) ? node33526 : node33523;
															assign node33523 = (inp[1]) ? 4'b1101 : 4'b1100;
															assign node33526 = (inp[1]) ? 4'b1100 : 4'b1101;
													assign node33529 = (inp[9]) ? node33537 : node33530;
														assign node33530 = (inp[11]) ? node33532 : 4'b1101;
															assign node33532 = (inp[0]) ? 4'b1101 : node33533;
																assign node33533 = (inp[1]) ? 4'b1101 : 4'b1100;
														assign node33537 = (inp[0]) ? node33543 : node33538;
															assign node33538 = (inp[11]) ? node33540 : 4'b1100;
																assign node33540 = (inp[1]) ? 4'b1100 : 4'b1101;
															assign node33543 = (inp[1]) ? 4'b1101 : 4'b1100;
												assign node33546 = (inp[1]) ? node33562 : node33547;
													assign node33547 = (inp[9]) ? node33557 : node33548;
														assign node33548 = (inp[10]) ? node33554 : node33549;
															assign node33549 = (inp[11]) ? node33551 : 4'b1010;
																assign node33551 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node33554 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node33557 = (inp[10]) ? 4'b1010 : node33558;
															assign node33558 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node33562 = (inp[9]) ? node33572 : node33563;
														assign node33563 = (inp[11]) ? 4'b1010 : node33564;
															assign node33564 = (inp[0]) ? node33568 : node33565;
																assign node33565 = (inp[10]) ? 4'b1011 : 4'b1010;
																assign node33568 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node33572 = (inp[0]) ? node33574 : 4'b1011;
															assign node33574 = (inp[10]) ? node33578 : node33575;
																assign node33575 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node33578 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node33581 = (inp[11]) ? node33619 : node33582;
												assign node33582 = (inp[4]) ? node33596 : node33583;
													assign node33583 = (inp[0]) ? node33591 : node33584;
														assign node33584 = (inp[9]) ? node33588 : node33585;
															assign node33585 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node33588 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node33591 = (inp[9]) ? node33593 : 4'b1001;
															assign node33593 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node33596 = (inp[1]) ? node33606 : node33597;
														assign node33597 = (inp[9]) ? node33599 : 4'b1001;
															assign node33599 = (inp[0]) ? node33603 : node33600;
																assign node33600 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node33603 = (inp[10]) ? 4'b1001 : 4'b1000;
														assign node33606 = (inp[9]) ? node33612 : node33607;
															assign node33607 = (inp[0]) ? 4'b1000 : node33608;
																assign node33608 = (inp[10]) ? 4'b1001 : 4'b1000;
															assign node33612 = (inp[0]) ? node33616 : node33613;
																assign node33613 = (inp[10]) ? 4'b1000 : 4'b1001;
																assign node33616 = (inp[10]) ? 4'b1001 : 4'b1000;
												assign node33619 = (inp[10]) ? node33623 : node33620;
													assign node33620 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node33623 = (inp[9]) ? 4'b1000 : 4'b1001;
							assign node33626 = (inp[12]) ? node34080 : node33627;
								assign node33627 = (inp[15]) ? node33835 : node33628;
									assign node33628 = (inp[7]) ? node33732 : node33629;
										assign node33629 = (inp[1]) ? node33669 : node33630;
											assign node33630 = (inp[9]) ? node33650 : node33631;
												assign node33631 = (inp[11]) ? node33641 : node33632;
													assign node33632 = (inp[0]) ? node33634 : 4'b1001;
														assign node33634 = (inp[2]) ? node33638 : node33635;
															assign node33635 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node33638 = (inp[4]) ? 4'b1000 : 4'b1001;
													assign node33641 = (inp[0]) ? node33643 : 4'b1000;
														assign node33643 = (inp[4]) ? node33647 : node33644;
															assign node33644 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node33647 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node33650 = (inp[11]) ? node33658 : node33651;
													assign node33651 = (inp[2]) ? 4'b1000 : node33652;
														assign node33652 = (inp[4]) ? 4'b1000 : node33653;
															assign node33653 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node33658 = (inp[0]) ? node33660 : 4'b1001;
														assign node33660 = (inp[10]) ? node33662 : 4'b1001;
															assign node33662 = (inp[2]) ? node33666 : node33663;
																assign node33663 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node33666 = (inp[4]) ? 4'b1000 : 4'b1001;
											assign node33669 = (inp[4]) ? node33709 : node33670;
												assign node33670 = (inp[0]) ? node33690 : node33671;
													assign node33671 = (inp[10]) ? node33679 : node33672;
														assign node33672 = (inp[11]) ? node33676 : node33673;
															assign node33673 = (inp[9]) ? 4'b1100 : 4'b1101;
															assign node33676 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node33679 = (inp[2]) ? node33685 : node33680;
															assign node33680 = (inp[9]) ? node33682 : 4'b1100;
																assign node33682 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node33685 = (inp[9]) ? node33687 : 4'b1101;
																assign node33687 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node33690 = (inp[10]) ? node33698 : node33691;
														assign node33691 = (inp[2]) ? 4'b1101 : node33692;
															assign node33692 = (inp[11]) ? 4'b1101 : node33693;
																assign node33693 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node33698 = (inp[9]) ? node33704 : node33699;
															assign node33699 = (inp[2]) ? node33701 : 4'b1101;
																assign node33701 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node33704 = (inp[11]) ? node33706 : 4'b1100;
																assign node33706 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node33709 = (inp[2]) ? node33725 : node33710;
													assign node33710 = (inp[11]) ? node33720 : node33711;
														assign node33711 = (inp[10]) ? node33717 : node33712;
															assign node33712 = (inp[0]) ? 4'b1001 : node33713;
																assign node33713 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node33717 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node33720 = (inp[9]) ? node33722 : 4'b1001;
															assign node33722 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node33725 = (inp[11]) ? node33729 : node33726;
														assign node33726 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node33729 = (inp[9]) ? 4'b1001 : 4'b1000;
										assign node33732 = (inp[1]) ? node33784 : node33733;
											assign node33733 = (inp[4]) ? node33755 : node33734;
												assign node33734 = (inp[9]) ? node33746 : node33735;
													assign node33735 = (inp[11]) ? node33741 : node33736;
														assign node33736 = (inp[2]) ? 4'b1010 : node33737;
															assign node33737 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node33741 = (inp[2]) ? 4'b1011 : node33742;
															assign node33742 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node33746 = (inp[11]) ? node33750 : node33747;
														assign node33747 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node33750 = (inp[0]) ? node33752 : 4'b1010;
															assign node33752 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node33755 = (inp[0]) ? node33763 : node33756;
													assign node33756 = (inp[9]) ? node33760 : node33757;
														assign node33757 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node33760 = (inp[11]) ? 4'b1110 : 4'b1111;
													assign node33763 = (inp[10]) ? node33773 : node33764;
														assign node33764 = (inp[2]) ? 4'b1111 : node33765;
															assign node33765 = (inp[11]) ? node33769 : node33766;
																assign node33766 = (inp[9]) ? 4'b1111 : 4'b1110;
																assign node33769 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node33773 = (inp[9]) ? node33779 : node33774;
															assign node33774 = (inp[11]) ? 4'b1110 : node33775;
																assign node33775 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node33779 = (inp[2]) ? node33781 : 4'b1111;
																assign node33781 = (inp[11]) ? 4'b1111 : 4'b1110;
											assign node33784 = (inp[0]) ? node33828 : node33785;
												assign node33785 = (inp[10]) ? node33803 : node33786;
													assign node33786 = (inp[2]) ? node33794 : node33787;
														assign node33787 = (inp[4]) ? node33791 : node33788;
															assign node33788 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node33791 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node33794 = (inp[9]) ? node33796 : 4'b1011;
															assign node33796 = (inp[11]) ? node33800 : node33797;
																assign node33797 = (inp[4]) ? 4'b1011 : 4'b1010;
																assign node33800 = (inp[4]) ? 4'b1010 : 4'b1011;
													assign node33803 = (inp[4]) ? node33813 : node33804;
														assign node33804 = (inp[11]) ? node33806 : 4'b1010;
															assign node33806 = (inp[9]) ? node33810 : node33807;
																assign node33807 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node33810 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node33813 = (inp[11]) ? node33821 : node33814;
															assign node33814 = (inp[2]) ? node33818 : node33815;
																assign node33815 = (inp[9]) ? 4'b1010 : 4'b1011;
																assign node33818 = (inp[9]) ? 4'b1011 : 4'b1010;
															assign node33821 = (inp[9]) ? node33825 : node33822;
																assign node33822 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node33825 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node33828 = (inp[11]) ? node33832 : node33829;
													assign node33829 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node33832 = (inp[9]) ? 4'b1010 : 4'b1011;
									assign node33835 = (inp[7]) ? node33939 : node33836;
										assign node33836 = (inp[4]) ? node33886 : node33837;
											assign node33837 = (inp[1]) ? node33861 : node33838;
												assign node33838 = (inp[11]) ? node33850 : node33839;
													assign node33839 = (inp[9]) ? node33845 : node33840;
														assign node33840 = (inp[2]) ? 4'b1010 : node33841;
															assign node33841 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node33845 = (inp[2]) ? 4'b1011 : node33846;
															assign node33846 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node33850 = (inp[9]) ? node33856 : node33851;
														assign node33851 = (inp[2]) ? 4'b1011 : node33852;
															assign node33852 = (inp[0]) ? 4'b1010 : 4'b1011;
														assign node33856 = (inp[0]) ? node33858 : 4'b1010;
															assign node33858 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node33861 = (inp[10]) ? node33881 : node33862;
													assign node33862 = (inp[9]) ? node33874 : node33863;
														assign node33863 = (inp[11]) ? node33869 : node33864;
															assign node33864 = (inp[2]) ? node33866 : 4'b1110;
																assign node33866 = (inp[0]) ? 4'b1110 : 4'b1111;
															assign node33869 = (inp[2]) ? node33871 : 4'b1111;
																assign node33871 = (inp[0]) ? 4'b1111 : 4'b1110;
														assign node33874 = (inp[11]) ? 4'b1110 : node33875;
															assign node33875 = (inp[2]) ? node33877 : 4'b1111;
																assign node33877 = (inp[0]) ? 4'b1111 : 4'b1110;
													assign node33881 = (inp[0]) ? 4'b1110 : node33882;
														assign node33882 = (inp[9]) ? 4'b1110 : 4'b1111;
											assign node33886 = (inp[1]) ? node33918 : node33887;
												assign node33887 = (inp[2]) ? node33895 : node33888;
													assign node33888 = (inp[11]) ? node33892 : node33889;
														assign node33889 = (inp[9]) ? 4'b1111 : 4'b1110;
														assign node33892 = (inp[9]) ? 4'b1110 : 4'b1111;
													assign node33895 = (inp[10]) ? node33905 : node33896;
														assign node33896 = (inp[0]) ? node33898 : 4'b1111;
															assign node33898 = (inp[9]) ? node33902 : node33899;
																assign node33899 = (inp[11]) ? 4'b1110 : 4'b1111;
																assign node33902 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node33905 = (inp[9]) ? node33913 : node33906;
															assign node33906 = (inp[0]) ? node33910 : node33907;
																assign node33907 = (inp[11]) ? 4'b1111 : 4'b1110;
																assign node33910 = (inp[11]) ? 4'b1110 : 4'b1111;
															assign node33913 = (inp[11]) ? node33915 : 4'b1111;
																assign node33915 = (inp[0]) ? 4'b1111 : 4'b1110;
												assign node33918 = (inp[11]) ? node33930 : node33919;
													assign node33919 = (inp[9]) ? node33925 : node33920;
														assign node33920 = (inp[0]) ? node33922 : 4'b1011;
															assign node33922 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node33925 = (inp[0]) ? node33927 : 4'b1010;
															assign node33927 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node33930 = (inp[2]) ? node33932 : 4'b1011;
														assign node33932 = (inp[9]) ? node33936 : node33933;
															assign node33933 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node33936 = (inp[0]) ? 4'b1010 : 4'b1011;
										assign node33939 = (inp[0]) ? node34005 : node33940;
											assign node33940 = (inp[9]) ? node33968 : node33941;
												assign node33941 = (inp[11]) ? node33955 : node33942;
													assign node33942 = (inp[2]) ? node33950 : node33943;
														assign node33943 = (inp[1]) ? node33947 : node33944;
															assign node33944 = (inp[4]) ? 4'b1100 : 4'b1001;
															assign node33947 = (inp[4]) ? 4'b1001 : 4'b1100;
														assign node33950 = (inp[1]) ? 4'b1000 : node33951;
															assign node33951 = (inp[4]) ? 4'b1101 : 4'b1000;
													assign node33955 = (inp[1]) ? node33963 : node33956;
														assign node33956 = (inp[4]) ? node33960 : node33957;
															assign node33957 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node33960 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node33963 = (inp[4]) ? node33965 : 4'b1101;
															assign node33965 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node33968 = (inp[10]) ? node33984 : node33969;
													assign node33969 = (inp[4]) ? node33977 : node33970;
														assign node33970 = (inp[1]) ? 4'b1100 : node33971;
															assign node33971 = (inp[2]) ? 4'b1000 : node33972;
																assign node33972 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node33977 = (inp[1]) ? node33979 : 4'b1100;
															assign node33979 = (inp[11]) ? node33981 : 4'b1001;
																assign node33981 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node33984 = (inp[11]) ? node33996 : node33985;
														assign node33985 = (inp[1]) ? node33991 : node33986;
															assign node33986 = (inp[4]) ? 4'b1100 : node33987;
																assign node33987 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node33991 = (inp[4]) ? node33993 : 4'b1101;
																assign node33993 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node33996 = (inp[1]) ? node34002 : node33997;
															assign node33997 = (inp[4]) ? 4'b1101 : node33998;
																assign node33998 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node34002 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node34005 = (inp[10]) ? node34041 : node34006;
												assign node34006 = (inp[1]) ? node34024 : node34007;
													assign node34007 = (inp[4]) ? node34015 : node34008;
														assign node34008 = (inp[9]) ? node34012 : node34009;
															assign node34009 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node34012 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node34015 = (inp[2]) ? 4'b1100 : node34016;
															assign node34016 = (inp[9]) ? node34020 : node34017;
																assign node34017 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node34020 = (inp[11]) ? 4'b1101 : 4'b1100;
													assign node34024 = (inp[4]) ? node34038 : node34025;
														assign node34025 = (inp[9]) ? node34031 : node34026;
															assign node34026 = (inp[2]) ? 4'b1100 : node34027;
																assign node34027 = (inp[11]) ? 4'b1100 : 4'b1101;
															assign node34031 = (inp[2]) ? node34035 : node34032;
																assign node34032 = (inp[11]) ? 4'b1101 : 4'b1100;
																assign node34035 = (inp[11]) ? 4'b1100 : 4'b1101;
														assign node34038 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node34041 = (inp[4]) ? node34057 : node34042;
													assign node34042 = (inp[1]) ? node34050 : node34043;
														assign node34043 = (inp[9]) ? node34047 : node34044;
															assign node34044 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node34047 = (inp[11]) ? 4'b1001 : 4'b1000;
														assign node34050 = (inp[2]) ? node34052 : 4'b1101;
															assign node34052 = (inp[11]) ? 4'b1100 : node34053;
																assign node34053 = (inp[9]) ? 4'b1101 : 4'b1100;
													assign node34057 = (inp[1]) ? node34073 : node34058;
														assign node34058 = (inp[2]) ? node34066 : node34059;
															assign node34059 = (inp[9]) ? node34063 : node34060;
																assign node34060 = (inp[11]) ? 4'b1100 : 4'b1101;
																assign node34063 = (inp[11]) ? 4'b1101 : 4'b1100;
															assign node34066 = (inp[11]) ? node34070 : node34067;
																assign node34067 = (inp[9]) ? 4'b1100 : 4'b1101;
																assign node34070 = (inp[9]) ? 4'b1101 : 4'b1100;
														assign node34073 = (inp[11]) ? node34077 : node34074;
															assign node34074 = (inp[9]) ? 4'b1001 : 4'b1000;
															assign node34077 = (inp[9]) ? 4'b1000 : 4'b1001;
								assign node34080 = (inp[15]) ? node34322 : node34081;
									assign node34081 = (inp[7]) ? node34183 : node34082;
										assign node34082 = (inp[4]) ? node34130 : node34083;
											assign node34083 = (inp[2]) ? node34107 : node34084;
												assign node34084 = (inp[9]) ? node34096 : node34085;
													assign node34085 = (inp[11]) ? node34091 : node34086;
														assign node34086 = (inp[1]) ? 4'b1000 : node34087;
															assign node34087 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node34091 = (inp[1]) ? 4'b1001 : node34092;
															assign node34092 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node34096 = (inp[11]) ? node34102 : node34097;
														assign node34097 = (inp[1]) ? 4'b1001 : node34098;
															assign node34098 = (inp[0]) ? 4'b1001 : 4'b1000;
														assign node34102 = (inp[1]) ? 4'b1000 : node34103;
															assign node34103 = (inp[0]) ? 4'b1000 : 4'b1001;
												assign node34107 = (inp[9]) ? node34119 : node34108;
													assign node34108 = (inp[11]) ? node34114 : node34109;
														assign node34109 = (inp[1]) ? node34111 : 4'b1001;
															assign node34111 = (inp[0]) ? 4'b1000 : 4'b1001;
														assign node34114 = (inp[1]) ? node34116 : 4'b1000;
															assign node34116 = (inp[0]) ? 4'b1001 : 4'b1000;
													assign node34119 = (inp[11]) ? node34125 : node34120;
														assign node34120 = (inp[0]) ? node34122 : 4'b1000;
															assign node34122 = (inp[1]) ? 4'b1001 : 4'b1000;
														assign node34125 = (inp[0]) ? node34127 : 4'b1001;
															assign node34127 = (inp[1]) ? 4'b1000 : 4'b1001;
											assign node34130 = (inp[1]) ? node34160 : node34131;
												assign node34131 = (inp[2]) ? node34153 : node34132;
													assign node34132 = (inp[10]) ? node34144 : node34133;
														assign node34133 = (inp[11]) ? node34139 : node34134;
															assign node34134 = (inp[9]) ? 4'b1001 : node34135;
																assign node34135 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node34139 = (inp[0]) ? 4'b1000 : node34140;
																assign node34140 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node34144 = (inp[11]) ? 4'b1001 : node34145;
															assign node34145 = (inp[9]) ? node34149 : node34146;
																assign node34146 = (inp[0]) ? 4'b1001 : 4'b1000;
																assign node34149 = (inp[0]) ? 4'b1000 : 4'b1001;
													assign node34153 = (inp[11]) ? node34157 : node34154;
														assign node34154 = (inp[9]) ? 4'b1000 : 4'b1001;
														assign node34157 = (inp[9]) ? 4'b1001 : 4'b1000;
												assign node34160 = (inp[10]) ? node34176 : node34161;
													assign node34161 = (inp[9]) ? node34171 : node34162;
														assign node34162 = (inp[11]) ? node34166 : node34163;
															assign node34163 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node34166 = (inp[0]) ? 4'b1101 : node34167;
																assign node34167 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node34171 = (inp[11]) ? 4'b1100 : node34172;
															assign node34172 = (inp[0]) ? 4'b1101 : 4'b1100;
													assign node34176 = (inp[11]) ? node34178 : 4'b1101;
														assign node34178 = (inp[0]) ? 4'b1101 : node34179;
															assign node34179 = (inp[9]) ? 4'b1101 : 4'b1100;
										assign node34183 = (inp[1]) ? node34239 : node34184;
											assign node34184 = (inp[4]) ? node34214 : node34185;
												assign node34185 = (inp[0]) ? node34207 : node34186;
													assign node34186 = (inp[11]) ? node34198 : node34187;
														assign node34187 = (inp[10]) ? node34193 : node34188;
															assign node34188 = (inp[9]) ? 4'b1111 : node34189;
																assign node34189 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node34193 = (inp[2]) ? node34195 : 4'b1111;
																assign node34195 = (inp[9]) ? 4'b1110 : 4'b1111;
														assign node34198 = (inp[10]) ? node34200 : 4'b1110;
															assign node34200 = (inp[2]) ? node34204 : node34201;
																assign node34201 = (inp[9]) ? 4'b1110 : 4'b1111;
																assign node34204 = (inp[9]) ? 4'b1111 : 4'b1110;
													assign node34207 = (inp[9]) ? node34211 : node34208;
														assign node34208 = (inp[11]) ? 4'b1111 : 4'b1110;
														assign node34211 = (inp[11]) ? 4'b1110 : 4'b1111;
												assign node34214 = (inp[2]) ? node34222 : node34215;
													assign node34215 = (inp[11]) ? node34219 : node34216;
														assign node34216 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node34219 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node34222 = (inp[10]) ? node34228 : node34223;
														assign node34223 = (inp[9]) ? node34225 : 4'b1010;
															assign node34225 = (inp[0]) ? 4'b1011 : 4'b1010;
														assign node34228 = (inp[9]) ? node34234 : node34229;
															assign node34229 = (inp[11]) ? 4'b1011 : node34230;
																assign node34230 = (inp[0]) ? 4'b1010 : 4'b1011;
															assign node34234 = (inp[11]) ? 4'b1010 : node34235;
																assign node34235 = (inp[0]) ? 4'b1011 : 4'b1010;
											assign node34239 = (inp[10]) ? node34279 : node34240;
												assign node34240 = (inp[0]) ? node34260 : node34241;
													assign node34241 = (inp[2]) ? node34255 : node34242;
														assign node34242 = (inp[11]) ? node34250 : node34243;
															assign node34243 = (inp[4]) ? node34247 : node34244;
																assign node34244 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node34247 = (inp[9]) ? 4'b1010 : 4'b1011;
															assign node34250 = (inp[9]) ? node34252 : 4'b1011;
																assign node34252 = (inp[4]) ? 4'b1011 : 4'b1010;
														assign node34255 = (inp[9]) ? 4'b1011 : node34256;
															assign node34256 = (inp[11]) ? 4'b1011 : 4'b1010;
													assign node34260 = (inp[11]) ? node34270 : node34261;
														assign node34261 = (inp[4]) ? 4'b1011 : node34262;
															assign node34262 = (inp[9]) ? node34266 : node34263;
																assign node34263 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node34266 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node34270 = (inp[9]) ? node34274 : node34271;
															assign node34271 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node34274 = (inp[2]) ? 4'b1010 : node34275;
																assign node34275 = (inp[4]) ? 4'b1010 : 4'b1011;
												assign node34279 = (inp[2]) ? node34305 : node34280;
													assign node34280 = (inp[4]) ? node34290 : node34281;
														assign node34281 = (inp[0]) ? 4'b1011 : node34282;
															assign node34282 = (inp[11]) ? node34286 : node34283;
																assign node34283 = (inp[9]) ? 4'b1011 : 4'b1010;
																assign node34286 = (inp[9]) ? 4'b1010 : 4'b1011;
														assign node34290 = (inp[9]) ? node34298 : node34291;
															assign node34291 = (inp[11]) ? node34295 : node34292;
																assign node34292 = (inp[0]) ? 4'b1010 : 4'b1011;
																assign node34295 = (inp[0]) ? 4'b1011 : 4'b1010;
															assign node34298 = (inp[11]) ? node34302 : node34299;
																assign node34299 = (inp[0]) ? 4'b1011 : 4'b1010;
																assign node34302 = (inp[0]) ? 4'b1010 : 4'b1011;
													assign node34305 = (inp[0]) ? node34313 : node34306;
														assign node34306 = (inp[9]) ? node34310 : node34307;
															assign node34307 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node34310 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node34313 = (inp[4]) ? node34315 : 4'b1010;
															assign node34315 = (inp[9]) ? node34319 : node34316;
																assign node34316 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node34319 = (inp[11]) ? 4'b1010 : 4'b1011;
									assign node34322 = (inp[7]) ? node34406 : node34323;
										assign node34323 = (inp[0]) ? node34361 : node34324;
											assign node34324 = (inp[2]) ? node34346 : node34325;
												assign node34325 = (inp[9]) ? node34339 : node34326;
													assign node34326 = (inp[1]) ? node34332 : node34327;
														assign node34327 = (inp[4]) ? node34329 : 4'b1010;
															assign node34329 = (inp[11]) ? 4'b1010 : 4'b1011;
														assign node34332 = (inp[4]) ? node34336 : node34333;
															assign node34333 = (inp[11]) ? 4'b1011 : 4'b1010;
															assign node34336 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node34339 = (inp[11]) ? node34343 : node34340;
														assign node34340 = (inp[4]) ? 4'b1010 : 4'b1011;
														assign node34343 = (inp[4]) ? 4'b1011 : 4'b1010;
												assign node34346 = (inp[1]) ? node34354 : node34347;
													assign node34347 = (inp[11]) ? node34351 : node34348;
														assign node34348 = (inp[9]) ? 4'b1011 : 4'b1010;
														assign node34351 = (inp[9]) ? 4'b1010 : 4'b1011;
													assign node34354 = (inp[9]) ? node34358 : node34355;
														assign node34355 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node34358 = (inp[11]) ? 4'b1010 : 4'b1011;
											assign node34361 = (inp[4]) ? node34399 : node34362;
												assign node34362 = (inp[1]) ? node34386 : node34363;
													assign node34363 = (inp[9]) ? node34373 : node34364;
														assign node34364 = (inp[10]) ? 4'b1011 : node34365;
															assign node34365 = (inp[2]) ? node34369 : node34366;
																assign node34366 = (inp[11]) ? 4'b1010 : 4'b1011;
																assign node34369 = (inp[11]) ? 4'b1011 : 4'b1010;
														assign node34373 = (inp[10]) ? node34381 : node34374;
															assign node34374 = (inp[2]) ? node34378 : node34375;
																assign node34375 = (inp[11]) ? 4'b1011 : 4'b1010;
																assign node34378 = (inp[11]) ? 4'b1010 : 4'b1011;
															assign node34381 = (inp[2]) ? node34383 : 4'b1010;
																assign node34383 = (inp[11]) ? 4'b1010 : 4'b1011;
													assign node34386 = (inp[11]) ? node34392 : node34387;
														assign node34387 = (inp[9]) ? 4'b1010 : node34388;
															assign node34388 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node34392 = (inp[9]) ? node34396 : node34393;
															assign node34393 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node34396 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node34399 = (inp[11]) ? node34403 : node34400;
													assign node34400 = (inp[9]) ? 4'b1011 : 4'b1010;
													assign node34403 = (inp[9]) ? 4'b1010 : 4'b1011;
										assign node34406 = (inp[2]) ? node34494 : node34407;
											assign node34407 = (inp[10]) ? node34453 : node34408;
												assign node34408 = (inp[9]) ? node34426 : node34409;
													assign node34409 = (inp[0]) ? node34419 : node34410;
														assign node34410 = (inp[1]) ? node34412 : 4'b1000;
															assign node34412 = (inp[11]) ? node34416 : node34413;
																assign node34413 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node34416 = (inp[4]) ? 4'b1000 : 4'b1001;
														assign node34419 = (inp[4]) ? node34423 : node34420;
															assign node34420 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node34423 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node34426 = (inp[11]) ? node34438 : node34427;
														assign node34427 = (inp[1]) ? node34433 : node34428;
															assign node34428 = (inp[4]) ? node34430 : 4'b1001;
																assign node34430 = (inp[0]) ? 4'b1001 : 4'b1000;
															assign node34433 = (inp[0]) ? node34435 : 4'b1001;
																assign node34435 = (inp[4]) ? 4'b1001 : 4'b1000;
														assign node34438 = (inp[1]) ? node34446 : node34439;
															assign node34439 = (inp[0]) ? node34443 : node34440;
																assign node34440 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node34443 = (inp[4]) ? 4'b1000 : 4'b1001;
															assign node34446 = (inp[0]) ? node34450 : node34447;
																assign node34447 = (inp[4]) ? 4'b1001 : 4'b1000;
																assign node34450 = (inp[4]) ? 4'b1000 : 4'b1001;
												assign node34453 = (inp[9]) ? node34479 : node34454;
													assign node34454 = (inp[0]) ? node34470 : node34455;
														assign node34455 = (inp[1]) ? node34463 : node34456;
															assign node34456 = (inp[4]) ? node34460 : node34457;
																assign node34457 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node34460 = (inp[11]) ? 4'b1000 : 4'b1001;
															assign node34463 = (inp[4]) ? node34467 : node34464;
																assign node34464 = (inp[11]) ? 4'b1001 : 4'b1000;
																assign node34467 = (inp[11]) ? 4'b1000 : 4'b1001;
														assign node34470 = (inp[1]) ? node34476 : node34471;
															assign node34471 = (inp[11]) ? node34473 : 4'b1001;
																assign node34473 = (inp[4]) ? 4'b1001 : 4'b1000;
															assign node34476 = (inp[11]) ? 4'b1001 : 4'b1000;
													assign node34479 = (inp[0]) ? 4'b1000 : node34480;
														assign node34480 = (inp[1]) ? node34488 : node34481;
															assign node34481 = (inp[4]) ? node34485 : node34482;
																assign node34482 = (inp[11]) ? 4'b1000 : 4'b1001;
																assign node34485 = (inp[11]) ? 4'b1001 : 4'b1000;
															assign node34488 = (inp[11]) ? node34490 : 4'b1000;
																assign node34490 = (inp[4]) ? 4'b1001 : 4'b1000;
											assign node34494 = (inp[10]) ? node34502 : node34495;
												assign node34495 = (inp[11]) ? node34499 : node34496;
													assign node34496 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node34499 = (inp[9]) ? 4'b1000 : 4'b1001;
												assign node34502 = (inp[11]) ? node34506 : node34503;
													assign node34503 = (inp[9]) ? 4'b1001 : 4'b1000;
													assign node34506 = (inp[9]) ? 4'b1000 : 4'b1001;
				assign node34509 = (inp[7]) ? node37751 : node34510;
					assign node34510 = (inp[6]) ? node36932 : node34511;
						assign node34511 = (inp[12]) ? node35723 : node34512;
							assign node34512 = (inp[15]) ? node35090 : node34513;
								assign node34513 = (inp[4]) ? node34811 : node34514;
									assign node34514 = (inp[1]) ? node34672 : node34515;
										assign node34515 = (inp[13]) ? node34593 : node34516;
											assign node34516 = (inp[9]) ? node34556 : node34517;
												assign node34517 = (inp[0]) ? node34537 : node34518;
													assign node34518 = (inp[10]) ? node34530 : node34519;
														assign node34519 = (inp[11]) ? node34523 : node34520;
															assign node34520 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node34523 = (inp[2]) ? node34527 : node34524;
																assign node34524 = (inp[5]) ? 4'b0111 : 4'b0011;
																assign node34527 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node34530 = (inp[2]) ? 4'b0111 : node34531;
															assign node34531 = (inp[11]) ? 4'b0010 : node34532;
																assign node34532 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node34537 = (inp[10]) ? node34547 : node34538;
														assign node34538 = (inp[2]) ? node34542 : node34539;
															assign node34539 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node34542 = (inp[5]) ? 4'b0010 : node34543;
																assign node34543 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node34547 = (inp[2]) ? node34551 : node34548;
															assign node34548 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node34551 = (inp[5]) ? 4'b0011 : node34552;
																assign node34552 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node34556 = (inp[0]) ? node34574 : node34557;
													assign node34557 = (inp[10]) ? node34567 : node34558;
														assign node34558 = (inp[2]) ? node34564 : node34559;
															assign node34559 = (inp[5]) ? node34561 : 4'b0010;
																assign node34561 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node34564 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node34567 = (inp[11]) ? 4'b0010 : node34568;
															assign node34568 = (inp[5]) ? 4'b0110 : node34569;
																assign node34569 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node34574 = (inp[10]) ? node34584 : node34575;
														assign node34575 = (inp[2]) ? node34579 : node34576;
															assign node34576 = (inp[5]) ? 4'b0110 : 4'b0010;
															assign node34579 = (inp[5]) ? 4'b0011 : node34580;
																assign node34580 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node34584 = (inp[2]) ? node34588 : node34585;
															assign node34585 = (inp[5]) ? 4'b0111 : 4'b0011;
															assign node34588 = (inp[5]) ? 4'b0010 : node34589;
																assign node34589 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node34593 = (inp[11]) ? node34629 : node34594;
												assign node34594 = (inp[9]) ? node34614 : node34595;
													assign node34595 = (inp[10]) ? node34605 : node34596;
														assign node34596 = (inp[2]) ? node34602 : node34597;
															assign node34597 = (inp[5]) ? node34599 : 4'b0110;
																assign node34599 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node34602 = (inp[5]) ? 4'b0111 : 4'b0011;
														assign node34605 = (inp[2]) ? node34611 : node34606;
															assign node34606 = (inp[5]) ? node34608 : 4'b0111;
																assign node34608 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node34611 = (inp[5]) ? 4'b0110 : 4'b0010;
													assign node34614 = (inp[10]) ? node34622 : node34615;
														assign node34615 = (inp[2]) ? node34619 : node34616;
															assign node34616 = (inp[0]) ? 4'b0011 : 4'b0111;
															assign node34619 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node34622 = (inp[2]) ? node34626 : node34623;
															assign node34623 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node34626 = (inp[5]) ? 4'b0111 : 4'b0011;
												assign node34629 = (inp[9]) ? node34651 : node34630;
													assign node34630 = (inp[10]) ? node34640 : node34631;
														assign node34631 = (inp[2]) ? node34635 : node34632;
															assign node34632 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node34635 = (inp[0]) ? node34637 : 4'b0111;
																assign node34637 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node34640 = (inp[5]) ? node34648 : node34641;
															assign node34641 = (inp[2]) ? node34645 : node34642;
																assign node34642 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node34645 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node34648 = (inp[0]) ? 4'b0111 : 4'b0011;
													assign node34651 = (inp[10]) ? node34661 : node34652;
														assign node34652 = (inp[2]) ? node34656 : node34653;
															assign node34653 = (inp[5]) ? 4'b0011 : 4'b0111;
															assign node34656 = (inp[5]) ? 4'b0110 : node34657;
																assign node34657 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node34661 = (inp[5]) ? node34669 : node34662;
															assign node34662 = (inp[2]) ? node34666 : node34663;
																assign node34663 = (inp[0]) ? 4'b0111 : 4'b0110;
																assign node34666 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node34669 = (inp[2]) ? 4'b0110 : 4'b0010;
										assign node34672 = (inp[5]) ? node34754 : node34673;
											assign node34673 = (inp[10]) ? node34711 : node34674;
												assign node34674 = (inp[0]) ? node34692 : node34675;
													assign node34675 = (inp[9]) ? node34683 : node34676;
														assign node34676 = (inp[11]) ? 4'b0111 : node34677;
															assign node34677 = (inp[2]) ? 4'b0011 : node34678;
																assign node34678 = (inp[13]) ? 4'b0011 : 4'b0110;
														assign node34683 = (inp[13]) ? node34689 : node34684;
															assign node34684 = (inp[2]) ? 4'b0011 : node34685;
																assign node34685 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node34689 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node34692 = (inp[2]) ? node34700 : node34693;
														assign node34693 = (inp[13]) ? node34697 : node34694;
															assign node34694 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node34697 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node34700 = (inp[13]) ? node34704 : node34701;
															assign node34701 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node34704 = (inp[9]) ? node34708 : node34705;
																assign node34705 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node34708 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node34711 = (inp[0]) ? node34733 : node34712;
													assign node34712 = (inp[11]) ? node34726 : node34713;
														assign node34713 = (inp[9]) ? node34721 : node34714;
															assign node34714 = (inp[2]) ? node34718 : node34715;
																assign node34715 = (inp[13]) ? 4'b0010 : 4'b0111;
																assign node34718 = (inp[13]) ? 4'b0110 : 4'b0010;
															assign node34721 = (inp[13]) ? node34723 : 4'b0011;
																assign node34723 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node34726 = (inp[9]) ? node34728 : 4'b0011;
															assign node34728 = (inp[2]) ? 4'b0010 : node34729;
																assign node34729 = (inp[13]) ? 4'b0010 : 4'b0111;
													assign node34733 = (inp[11]) ? node34743 : node34734;
														assign node34734 = (inp[13]) ? node34740 : node34735;
															assign node34735 = (inp[2]) ? 4'b0010 : node34736;
																assign node34736 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node34740 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node34743 = (inp[13]) ? node34749 : node34744;
															assign node34744 = (inp[2]) ? 4'b0011 : node34745;
																assign node34745 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node34749 = (inp[9]) ? node34751 : 4'b0111;
																assign node34751 = (inp[2]) ? 4'b0110 : 4'b0010;
											assign node34754 = (inp[13]) ? node34786 : node34755;
												assign node34755 = (inp[2]) ? node34767 : node34756;
													assign node34756 = (inp[10]) ? node34760 : node34757;
														assign node34757 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node34760 = (inp[9]) ? 4'b0110 : node34761;
															assign node34761 = (inp[11]) ? node34763 : 4'b0111;
																assign node34763 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node34767 = (inp[10]) ? node34775 : node34768;
														assign node34768 = (inp[9]) ? node34770 : 4'b0011;
															assign node34770 = (inp[0]) ? node34772 : 4'b0010;
																assign node34772 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node34775 = (inp[9]) ? node34781 : node34776;
															assign node34776 = (inp[0]) ? node34778 : 4'b0010;
																assign node34778 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node34781 = (inp[0]) ? node34783 : 4'b0011;
																assign node34783 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node34786 = (inp[2]) ? node34802 : node34787;
													assign node34787 = (inp[0]) ? node34789 : 4'b0011;
														assign node34789 = (inp[11]) ? node34795 : node34790;
															assign node34790 = (inp[9]) ? node34792 : 4'b0011;
																assign node34792 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node34795 = (inp[10]) ? node34799 : node34796;
																assign node34796 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node34799 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node34802 = (inp[9]) ? 4'b0111 : node34803;
														assign node34803 = (inp[10]) ? node34805 : 4'b0111;
															assign node34805 = (inp[0]) ? 4'b0110 : node34806;
																assign node34806 = (inp[11]) ? 4'b0110 : 4'b0111;
									assign node34811 = (inp[5]) ? node34943 : node34812;
										assign node34812 = (inp[2]) ? node34868 : node34813;
											assign node34813 = (inp[13]) ? node34841 : node34814;
												assign node34814 = (inp[0]) ? node34826 : node34815;
													assign node34815 = (inp[11]) ? node34817 : 4'b0000;
														assign node34817 = (inp[1]) ? node34819 : 4'b0000;
															assign node34819 = (inp[10]) ? node34823 : node34820;
																assign node34820 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node34823 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node34826 = (inp[10]) ? node34832 : node34827;
														assign node34827 = (inp[9]) ? node34829 : 4'b0001;
															assign node34829 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node34832 = (inp[9]) ? node34838 : node34833;
															assign node34833 = (inp[1]) ? node34835 : 4'b0000;
																assign node34835 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node34838 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node34841 = (inp[9]) ? node34861 : node34842;
													assign node34842 = (inp[10]) ? node34850 : node34843;
														assign node34843 = (inp[1]) ? node34845 : 4'b0100;
															assign node34845 = (inp[0]) ? 4'b0100 : node34846;
																assign node34846 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node34850 = (inp[0]) ? node34856 : node34851;
															assign node34851 = (inp[11]) ? 4'b0101 : node34852;
																assign node34852 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node34856 = (inp[11]) ? node34858 : 4'b0101;
																assign node34858 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node34861 = (inp[10]) ? 4'b0100 : node34862;
														assign node34862 = (inp[11]) ? 4'b0101 : node34863;
															assign node34863 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node34868 = (inp[13]) ? node34904 : node34869;
												assign node34869 = (inp[9]) ? node34887 : node34870;
													assign node34870 = (inp[10]) ? node34878 : node34871;
														assign node34871 = (inp[1]) ? 4'b0101 : node34872;
															assign node34872 = (inp[11]) ? node34874 : 4'b0101;
																assign node34874 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node34878 = (inp[0]) ? node34884 : node34879;
															assign node34879 = (inp[1]) ? node34881 : 4'b0100;
																assign node34881 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node34884 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node34887 = (inp[10]) ? node34893 : node34888;
														assign node34888 = (inp[1]) ? 4'b0100 : node34889;
															assign node34889 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node34893 = (inp[0]) ? node34899 : node34894;
															assign node34894 = (inp[1]) ? node34896 : 4'b0101;
																assign node34896 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node34899 = (inp[1]) ? 4'b0101 : node34900;
																assign node34900 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node34904 = (inp[1]) ? node34922 : node34905;
													assign node34905 = (inp[10]) ? node34911 : node34906;
														assign node34906 = (inp[9]) ? node34908 : 4'b0000;
															assign node34908 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node34911 = (inp[9]) ? node34917 : node34912;
															assign node34912 = (inp[0]) ? node34914 : 4'b0001;
																assign node34914 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node34917 = (inp[11]) ? node34919 : 4'b0000;
																assign node34919 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node34922 = (inp[0]) ? node34930 : node34923;
														assign node34923 = (inp[11]) ? 4'b0001 : node34924;
															assign node34924 = (inp[9]) ? 4'b0001 : node34925;
																assign node34925 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node34930 = (inp[11]) ? node34936 : node34931;
															assign node34931 = (inp[10]) ? node34933 : 4'b0000;
																assign node34933 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node34936 = (inp[10]) ? node34940 : node34937;
																assign node34937 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node34940 = (inp[9]) ? 4'b0000 : 4'b0001;
										assign node34943 = (inp[9]) ? node35019 : node34944;
											assign node34944 = (inp[0]) ? node34984 : node34945;
												assign node34945 = (inp[2]) ? node34969 : node34946;
													assign node34946 = (inp[13]) ? node34958 : node34947;
														assign node34947 = (inp[1]) ? node34955 : node34948;
															assign node34948 = (inp[11]) ? node34952 : node34949;
																assign node34949 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node34952 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node34955 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node34958 = (inp[1]) ? node34962 : node34959;
															assign node34959 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node34962 = (inp[10]) ? node34966 : node34963;
																assign node34963 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node34966 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node34969 = (inp[1]) ? node34975 : node34970;
														assign node34970 = (inp[13]) ? 4'b0001 : node34971;
															assign node34971 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node34975 = (inp[13]) ? node34981 : node34976;
															assign node34976 = (inp[11]) ? node34978 : 4'b0000;
																assign node34978 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node34981 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node34984 = (inp[10]) ? node35000 : node34985;
													assign node34985 = (inp[13]) ? node34987 : 4'b0100;
														assign node34987 = (inp[11]) ? node34995 : node34988;
															assign node34988 = (inp[2]) ? node34992 : node34989;
																assign node34989 = (inp[1]) ? 4'b0001 : 4'b0101;
																assign node34992 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node34995 = (inp[1]) ? node34997 : 4'b0100;
																assign node34997 = (inp[2]) ? 4'b0100 : 4'b0001;
													assign node35000 = (inp[11]) ? node35010 : node35001;
														assign node35001 = (inp[13]) ? node35005 : node35002;
															assign node35002 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node35005 = (inp[2]) ? node35007 : 4'b0000;
																assign node35007 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node35010 = (inp[13]) ? 4'b0101 : node35011;
															assign node35011 = (inp[2]) ? node35015 : node35012;
																assign node35012 = (inp[1]) ? 4'b0101 : 4'b0001;
																assign node35015 = (inp[1]) ? 4'b0001 : 4'b0100;
											assign node35019 = (inp[0]) ? node35065 : node35020;
												assign node35020 = (inp[10]) ? node35042 : node35021;
													assign node35021 = (inp[13]) ? node35035 : node35022;
														assign node35022 = (inp[11]) ? node35030 : node35023;
															assign node35023 = (inp[2]) ? node35027 : node35024;
																assign node35024 = (inp[1]) ? 4'b0100 : 4'b0000;
																assign node35027 = (inp[1]) ? 4'b0000 : 4'b0101;
															assign node35030 = (inp[2]) ? node35032 : 4'b0101;
																assign node35032 = (inp[1]) ? 4'b0001 : 4'b0101;
														assign node35035 = (inp[1]) ? node35039 : node35036;
															assign node35036 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node35039 = (inp[2]) ? 4'b0100 : 4'b0001;
													assign node35042 = (inp[13]) ? node35056 : node35043;
														assign node35043 = (inp[11]) ? node35049 : node35044;
															assign node35044 = (inp[2]) ? 4'b0100 : node35045;
																assign node35045 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node35049 = (inp[2]) ? node35053 : node35050;
																assign node35050 = (inp[1]) ? 4'b0100 : 4'b0000;
																assign node35053 = (inp[1]) ? 4'b0000 : 4'b0100;
														assign node35056 = (inp[1]) ? node35060 : node35057;
															assign node35057 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node35060 = (inp[2]) ? 4'b0101 : node35061;
																assign node35061 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node35065 = (inp[10]) ? node35073 : node35066;
													assign node35066 = (inp[1]) ? node35068 : 4'b0001;
														assign node35068 = (inp[13]) ? 4'b0100 : node35069;
															assign node35069 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node35073 = (inp[11]) ? node35083 : node35074;
														assign node35074 = (inp[13]) ? node35076 : 4'b0000;
															assign node35076 = (inp[1]) ? node35080 : node35077;
																assign node35077 = (inp[2]) ? 4'b0001 : 4'b0101;
																assign node35080 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node35083 = (inp[1]) ? 4'b0100 : node35084;
															assign node35084 = (inp[13]) ? 4'b0000 : node35085;
																assign node35085 = (inp[2]) ? 4'b0101 : 4'b0000;
								assign node35090 = (inp[9]) ? node35418 : node35091;
									assign node35091 = (inp[1]) ? node35253 : node35092;
										assign node35092 = (inp[0]) ? node35180 : node35093;
											assign node35093 = (inp[10]) ? node35139 : node35094;
												assign node35094 = (inp[13]) ? node35116 : node35095;
													assign node35095 = (inp[11]) ? node35107 : node35096;
														assign node35096 = (inp[5]) ? node35102 : node35097;
															assign node35097 = (inp[4]) ? node35099 : 4'b0100;
																assign node35099 = (inp[2]) ? 4'b0000 : 4'b0100;
															assign node35102 = (inp[4]) ? node35104 : 4'b0101;
																assign node35104 = (inp[2]) ? 4'b0001 : 4'b0101;
														assign node35107 = (inp[2]) ? node35113 : node35108;
															assign node35108 = (inp[4]) ? 4'b0100 : node35109;
																assign node35109 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node35113 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node35116 = (inp[2]) ? node35130 : node35117;
														assign node35117 = (inp[4]) ? node35123 : node35118;
															assign node35118 = (inp[11]) ? 4'b0101 : node35119;
																assign node35119 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node35123 = (inp[11]) ? node35127 : node35124;
																assign node35124 = (inp[5]) ? 4'b0001 : 4'b0000;
																assign node35127 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node35130 = (inp[4]) ? node35136 : node35131;
															assign node35131 = (inp[11]) ? 4'b0000 : node35132;
																assign node35132 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node35136 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node35139 = (inp[4]) ? node35153 : node35140;
													assign node35140 = (inp[2]) ? node35146 : node35141;
														assign node35141 = (inp[11]) ? 4'b0100 : node35142;
															assign node35142 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node35146 = (inp[13]) ? 4'b0001 : node35147;
															assign node35147 = (inp[5]) ? node35149 : 4'b0101;
																assign node35149 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node35153 = (inp[5]) ? node35165 : node35154;
														assign node35154 = (inp[11]) ? node35160 : node35155;
															assign node35155 = (inp[13]) ? 4'b0100 : node35156;
																assign node35156 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node35160 = (inp[13]) ? 4'b0100 : node35161;
																assign node35161 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node35165 = (inp[11]) ? node35173 : node35166;
															assign node35166 = (inp[2]) ? node35170 : node35167;
																assign node35167 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node35170 = (inp[13]) ? 4'b0101 : 4'b0000;
															assign node35173 = (inp[2]) ? node35177 : node35174;
																assign node35174 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node35177 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node35180 = (inp[5]) ? node35222 : node35181;
												assign node35181 = (inp[10]) ? node35207 : node35182;
													assign node35182 = (inp[13]) ? node35196 : node35183;
														assign node35183 = (inp[11]) ? node35189 : node35184;
															assign node35184 = (inp[2]) ? 4'b0001 : node35185;
																assign node35185 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node35189 = (inp[2]) ? node35193 : node35190;
																assign node35190 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node35193 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node35196 = (inp[2]) ? node35200 : node35197;
															assign node35197 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node35200 = (inp[4]) ? node35204 : node35201;
																assign node35201 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node35204 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node35207 = (inp[2]) ? node35213 : node35208;
														assign node35208 = (inp[4]) ? 4'b0100 : node35209;
															assign node35209 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node35213 = (inp[4]) ? node35219 : node35214;
															assign node35214 = (inp[11]) ? 4'b0000 : node35215;
																assign node35215 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node35219 = (inp[13]) ? 4'b0101 : 4'b0000;
												assign node35222 = (inp[10]) ? node35238 : node35223;
													assign node35223 = (inp[13]) ? node35233 : node35224;
														assign node35224 = (inp[2]) ? node35230 : node35225;
															assign node35225 = (inp[4]) ? 4'b0100 : node35226;
																assign node35226 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node35230 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node35233 = (inp[4]) ? node35235 : 4'b0101;
															assign node35235 = (inp[2]) ? 4'b0101 : 4'b0000;
													assign node35238 = (inp[2]) ? node35246 : node35239;
														assign node35239 = (inp[13]) ? node35243 : node35240;
															assign node35240 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node35243 = (inp[4]) ? 4'b0001 : 4'b0100;
														assign node35246 = (inp[13]) ? node35250 : node35247;
															assign node35247 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node35250 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node35253 = (inp[5]) ? node35335 : node35254;
											assign node35254 = (inp[10]) ? node35302 : node35255;
												assign node35255 = (inp[4]) ? node35275 : node35256;
													assign node35256 = (inp[2]) ? node35268 : node35257;
														assign node35257 = (inp[13]) ? node35263 : node35258;
															assign node35258 = (inp[0]) ? 4'b0000 : node35259;
																assign node35259 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node35263 = (inp[11]) ? node35265 : 4'b0100;
																assign node35265 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node35268 = (inp[13]) ? 4'b0001 : node35269;
															assign node35269 = (inp[0]) ? node35271 : 4'b0101;
																assign node35271 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node35275 = (inp[11]) ? node35289 : node35276;
														assign node35276 = (inp[0]) ? node35282 : node35277;
															assign node35277 = (inp[13]) ? node35279 : 4'b0001;
																assign node35279 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node35282 = (inp[13]) ? node35286 : node35283;
																assign node35283 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node35286 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node35289 = (inp[0]) ? node35297 : node35290;
															assign node35290 = (inp[2]) ? node35294 : node35291;
																assign node35291 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node35294 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node35297 = (inp[2]) ? 4'b0000 : node35298;
																assign node35298 = (inp[13]) ? 4'b0000 : 4'b0100;
												assign node35302 = (inp[0]) ? node35318 : node35303;
													assign node35303 = (inp[2]) ? node35311 : node35304;
														assign node35304 = (inp[11]) ? 4'b0101 : node35305;
															assign node35305 = (inp[4]) ? node35307 : 4'b0101;
																assign node35307 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node35311 = (inp[4]) ? node35315 : node35312;
															assign node35312 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node35315 = (inp[13]) ? 4'b0101 : 4'b0000;
													assign node35318 = (inp[13]) ? node35324 : node35319;
														assign node35319 = (inp[2]) ? node35321 : 4'b0101;
															assign node35321 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node35324 = (inp[4]) ? node35330 : node35325;
															assign node35325 = (inp[2]) ? node35327 : 4'b0100;
																assign node35327 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node35330 = (inp[2]) ? node35332 : 4'b0001;
																assign node35332 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node35335 = (inp[10]) ? node35379 : node35336;
												assign node35336 = (inp[2]) ? node35358 : node35337;
													assign node35337 = (inp[11]) ? node35349 : node35338;
														assign node35338 = (inp[4]) ? node35344 : node35339;
															assign node35339 = (inp[13]) ? node35341 : 4'b0101;
																assign node35341 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node35344 = (inp[13]) ? 4'b0101 : node35345;
																assign node35345 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node35349 = (inp[4]) ? node35353 : node35350;
															assign node35350 = (inp[13]) ? 4'b0000 : 4'b0100;
															assign node35353 = (inp[0]) ? 4'b0100 : node35354;
																assign node35354 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node35358 = (inp[11]) ? node35370 : node35359;
														assign node35359 = (inp[0]) ? node35365 : node35360;
															assign node35360 = (inp[13]) ? node35362 : 4'b0101;
																assign node35362 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node35365 = (inp[4]) ? 4'b0101 : node35366;
																assign node35366 = (inp[13]) ? 4'b0101 : 4'b0001;
														assign node35370 = (inp[0]) ? node35376 : node35371;
															assign node35371 = (inp[13]) ? node35373 : 4'b0001;
																assign node35373 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node35376 = (inp[4]) ? 4'b0100 : 4'b0001;
												assign node35379 = (inp[0]) ? node35395 : node35380;
													assign node35380 = (inp[2]) ? node35388 : node35381;
														assign node35381 = (inp[4]) ? node35385 : node35382;
															assign node35382 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node35385 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node35388 = (inp[4]) ? node35392 : node35389;
															assign node35389 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node35392 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node35395 = (inp[11]) ? node35407 : node35396;
														assign node35396 = (inp[2]) ? node35402 : node35397;
															assign node35397 = (inp[4]) ? 4'b0000 : node35398;
																assign node35398 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node35402 = (inp[4]) ? node35404 : 4'b0100;
																assign node35404 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node35407 = (inp[13]) ? node35413 : node35408;
															assign node35408 = (inp[4]) ? 4'b0101 : node35409;
																assign node35409 = (inp[2]) ? 4'b0000 : 4'b0101;
															assign node35413 = (inp[2]) ? node35415 : 4'b0001;
																assign node35415 = (inp[4]) ? 4'b0001 : 4'b0101;
									assign node35418 = (inp[11]) ? node35578 : node35419;
										assign node35419 = (inp[2]) ? node35503 : node35420;
											assign node35420 = (inp[0]) ? node35452 : node35421;
												assign node35421 = (inp[1]) ? node35435 : node35422;
													assign node35422 = (inp[10]) ? node35426 : node35423;
														assign node35423 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node35426 = (inp[5]) ? node35428 : 4'b0000;
															assign node35428 = (inp[4]) ? node35432 : node35429;
																assign node35429 = (inp[13]) ? 4'b0100 : 4'b0000;
																assign node35432 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node35435 = (inp[10]) ? node35447 : node35436;
														assign node35436 = (inp[5]) ? node35444 : node35437;
															assign node35437 = (inp[13]) ? node35441 : node35438;
																assign node35438 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node35441 = (inp[4]) ? 4'b0000 : 4'b0101;
															assign node35444 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node35447 = (inp[5]) ? node35449 : 4'b0001;
															assign node35449 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node35452 = (inp[1]) ? node35480 : node35453;
													assign node35453 = (inp[10]) ? node35467 : node35454;
														assign node35454 = (inp[5]) ? node35460 : node35455;
															assign node35455 = (inp[13]) ? node35457 : 4'b0100;
																assign node35457 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node35460 = (inp[13]) ? node35464 : node35461;
																assign node35461 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node35464 = (inp[4]) ? 4'b0001 : 4'b0100;
														assign node35467 = (inp[5]) ? node35475 : node35468;
															assign node35468 = (inp[13]) ? node35472 : node35469;
																assign node35469 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node35472 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node35475 = (inp[4]) ? node35477 : 4'b0101;
																assign node35477 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node35480 = (inp[10]) ? node35494 : node35481;
														assign node35481 = (inp[4]) ? node35489 : node35482;
															assign node35482 = (inp[13]) ? node35486 : node35483;
																assign node35483 = (inp[5]) ? 4'b0101 : 4'b0001;
																assign node35486 = (inp[5]) ? 4'b0001 : 4'b0101;
															assign node35489 = (inp[5]) ? node35491 : 4'b0001;
																assign node35491 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node35494 = (inp[5]) ? node35496 : 4'b0000;
															assign node35496 = (inp[4]) ? node35500 : node35497;
																assign node35497 = (inp[13]) ? 4'b0000 : 4'b0100;
																assign node35500 = (inp[13]) ? 4'b0101 : 4'b0001;
											assign node35503 = (inp[13]) ? node35549 : node35504;
												assign node35504 = (inp[4]) ? node35528 : node35505;
													assign node35505 = (inp[1]) ? node35517 : node35506;
														assign node35506 = (inp[10]) ? node35512 : node35507;
															assign node35507 = (inp[0]) ? 4'b0101 : node35508;
																assign node35508 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node35512 = (inp[0]) ? 4'b0100 : node35513;
																assign node35513 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node35517 = (inp[5]) ? node35521 : node35518;
															assign node35518 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node35521 = (inp[10]) ? node35525 : node35522;
																assign node35522 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node35525 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node35528 = (inp[1]) ? node35540 : node35529;
														assign node35529 = (inp[5]) ? node35535 : node35530;
															assign node35530 = (inp[0]) ? node35532 : 4'b0000;
																assign node35532 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node35535 = (inp[10]) ? node35537 : 4'b0001;
																assign node35537 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node35540 = (inp[5]) ? node35546 : node35541;
															assign node35541 = (inp[10]) ? node35543 : 4'b0001;
																assign node35543 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node35546 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node35549 = (inp[4]) ? node35565 : node35550;
													assign node35550 = (inp[5]) ? node35556 : node35551;
														assign node35551 = (inp[1]) ? node35553 : 4'b0000;
															assign node35553 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node35556 = (inp[1]) ? node35562 : node35557;
															assign node35557 = (inp[0]) ? 4'b0001 : node35558;
																assign node35558 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node35562 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node35565 = (inp[5]) ? node35573 : node35566;
														assign node35566 = (inp[10]) ? node35570 : node35567;
															assign node35567 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node35570 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node35573 = (inp[1]) ? 4'b0000 : node35574;
															assign node35574 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node35578 = (inp[2]) ? node35646 : node35579;
											assign node35579 = (inp[10]) ? node35613 : node35580;
												assign node35580 = (inp[1]) ? node35598 : node35581;
													assign node35581 = (inp[5]) ? node35589 : node35582;
														assign node35582 = (inp[0]) ? node35584 : 4'b0100;
															assign node35584 = (inp[13]) ? 4'b0000 : node35585;
																assign node35585 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node35589 = (inp[4]) ? node35595 : node35590;
															assign node35590 = (inp[13]) ? 4'b0100 : node35591;
																assign node35591 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node35595 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node35598 = (inp[4]) ? node35604 : node35599;
														assign node35599 = (inp[5]) ? 4'b0101 : node35600;
															assign node35600 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node35604 = (inp[5]) ? node35608 : node35605;
															assign node35605 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node35608 = (inp[13]) ? node35610 : 4'b0000;
																assign node35610 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node35613 = (inp[5]) ? node35627 : node35614;
													assign node35614 = (inp[1]) ? node35624 : node35615;
														assign node35615 = (inp[0]) ? node35619 : node35616;
															assign node35616 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node35619 = (inp[4]) ? node35621 : 4'b0001;
																assign node35621 = (inp[13]) ? 4'b0001 : 4'b0101;
														assign node35624 = (inp[13]) ? 4'b0101 : 4'b0000;
													assign node35627 = (inp[4]) ? node35637 : node35628;
														assign node35628 = (inp[1]) ? node35634 : node35629;
															assign node35629 = (inp[13]) ? 4'b0101 : node35630;
																assign node35630 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node35634 = (inp[13]) ? 4'b0000 : 4'b0100;
														assign node35637 = (inp[0]) ? node35641 : node35638;
															assign node35638 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node35641 = (inp[1]) ? 4'b0100 : node35642;
																assign node35642 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node35646 = (inp[10]) ? node35682 : node35647;
												assign node35647 = (inp[5]) ? node35669 : node35648;
													assign node35648 = (inp[4]) ? node35658 : node35649;
														assign node35649 = (inp[13]) ? node35651 : 4'b0100;
															assign node35651 = (inp[1]) ? node35655 : node35652;
																assign node35652 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node35655 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node35658 = (inp[13]) ? node35662 : node35659;
															assign node35659 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node35662 = (inp[0]) ? node35666 : node35663;
																assign node35663 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node35666 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node35669 = (inp[1]) ? node35679 : node35670;
														assign node35670 = (inp[13]) ? node35674 : node35671;
															assign node35671 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node35674 = (inp[4]) ? node35676 : 4'b0001;
																assign node35676 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node35679 = (inp[0]) ? 4'b0101 : 4'b0000;
												assign node35682 = (inp[5]) ? node35702 : node35683;
													assign node35683 = (inp[4]) ? node35693 : node35684;
														assign node35684 = (inp[13]) ? node35686 : 4'b0101;
															assign node35686 = (inp[0]) ? node35690 : node35687;
																assign node35687 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node35690 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node35693 = (inp[13]) ? node35697 : node35694;
															assign node35694 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node35697 = (inp[0]) ? 4'b0100 : node35698;
																assign node35698 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node35702 = (inp[1]) ? node35716 : node35703;
														assign node35703 = (inp[0]) ? node35711 : node35704;
															assign node35704 = (inp[13]) ? node35708 : node35705;
																assign node35705 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node35708 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node35711 = (inp[4]) ? node35713 : 4'b0000;
																assign node35713 = (inp[13]) ? 4'b0101 : 4'b0000;
														assign node35716 = (inp[0]) ? 4'b0100 : node35717;
															assign node35717 = (inp[13]) ? node35719 : 4'b0101;
																assign node35719 = (inp[4]) ? 4'b0001 : 4'b0101;
							assign node35723 = (inp[4]) ? node36283 : node35724;
								assign node35724 = (inp[15]) ? node36024 : node35725;
									assign node35725 = (inp[0]) ? node35901 : node35726;
										assign node35726 = (inp[1]) ? node35816 : node35727;
											assign node35727 = (inp[10]) ? node35775 : node35728;
												assign node35728 = (inp[5]) ? node35750 : node35729;
													assign node35729 = (inp[11]) ? node35739 : node35730;
														assign node35730 = (inp[9]) ? 4'b0101 : node35731;
															assign node35731 = (inp[13]) ? node35735 : node35732;
																assign node35732 = (inp[2]) ? 4'b0001 : 4'b0100;
																assign node35735 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node35739 = (inp[2]) ? node35745 : node35740;
															assign node35740 = (inp[13]) ? node35742 : 4'b0100;
																assign node35742 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node35745 = (inp[13]) ? node35747 : 4'b0001;
																assign node35747 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node35750 = (inp[2]) ? node35762 : node35751;
														assign node35751 = (inp[13]) ? node35755 : node35752;
															assign node35752 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node35755 = (inp[11]) ? node35759 : node35756;
																assign node35756 = (inp[9]) ? 4'b0100 : 4'b0101;
																assign node35759 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node35762 = (inp[13]) ? node35770 : node35763;
															assign node35763 = (inp[9]) ? node35767 : node35764;
																assign node35764 = (inp[11]) ? 4'b0100 : 4'b0101;
																assign node35767 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node35770 = (inp[9]) ? 4'b0000 : node35771;
																assign node35771 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node35775 = (inp[5]) ? node35793 : node35776;
													assign node35776 = (inp[9]) ? node35786 : node35777;
														assign node35777 = (inp[11]) ? 4'b0100 : node35778;
															assign node35778 = (inp[2]) ? node35782 : node35779;
																assign node35779 = (inp[13]) ? 4'b0000 : 4'b0101;
																assign node35782 = (inp[13]) ? 4'b0100 : 4'b0000;
														assign node35786 = (inp[13]) ? 4'b0101 : node35787;
															assign node35787 = (inp[2]) ? 4'b0000 : node35788;
																assign node35788 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node35793 = (inp[13]) ? node35805 : node35794;
														assign node35794 = (inp[2]) ? node35798 : node35795;
															assign node35795 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node35798 = (inp[11]) ? node35802 : node35799;
																assign node35799 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node35802 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node35805 = (inp[2]) ? node35811 : node35806;
															assign node35806 = (inp[9]) ? 4'b0100 : node35807;
																assign node35807 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node35811 = (inp[9]) ? node35813 : 4'b0000;
																assign node35813 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node35816 = (inp[13]) ? node35860 : node35817;
												assign node35817 = (inp[2]) ? node35835 : node35818;
													assign node35818 = (inp[9]) ? node35828 : node35819;
														assign node35819 = (inp[5]) ? node35823 : node35820;
															assign node35820 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node35823 = (inp[11]) ? 4'b0001 : node35824;
																assign node35824 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node35828 = (inp[10]) ? node35832 : node35829;
															assign node35829 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node35832 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node35835 = (inp[11]) ? node35851 : node35836;
														assign node35836 = (inp[5]) ? node35844 : node35837;
															assign node35837 = (inp[10]) ? node35841 : node35838;
																assign node35838 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node35841 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node35844 = (inp[9]) ? node35848 : node35845;
																assign node35845 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node35848 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node35851 = (inp[10]) ? 4'b0101 : node35852;
															assign node35852 = (inp[9]) ? node35856 : node35853;
																assign node35853 = (inp[5]) ? 4'b0100 : 4'b0101;
																assign node35856 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node35860 = (inp[2]) ? node35878 : node35861;
													assign node35861 = (inp[10]) ? node35873 : node35862;
														assign node35862 = (inp[9]) ? node35868 : node35863;
															assign node35863 = (inp[11]) ? node35865 : 4'b0100;
																assign node35865 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node35868 = (inp[11]) ? node35870 : 4'b0101;
																assign node35870 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node35873 = (inp[9]) ? node35875 : 4'b0101;
															assign node35875 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node35878 = (inp[11]) ? node35886 : node35879;
														assign node35879 = (inp[10]) ? node35883 : node35880;
															assign node35880 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node35883 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node35886 = (inp[5]) ? node35894 : node35887;
															assign node35887 = (inp[10]) ? node35891 : node35888;
																assign node35888 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node35891 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node35894 = (inp[10]) ? node35898 : node35895;
																assign node35895 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node35898 = (inp[9]) ? 4'b0001 : 4'b0000;
										assign node35901 = (inp[9]) ? node35965 : node35902;
											assign node35902 = (inp[5]) ? node35934 : node35903;
												assign node35903 = (inp[13]) ? node35925 : node35904;
													assign node35904 = (inp[10]) ? node35916 : node35905;
														assign node35905 = (inp[11]) ? node35911 : node35906;
															assign node35906 = (inp[1]) ? node35908 : 4'b0101;
																assign node35908 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node35911 = (inp[1]) ? node35913 : 4'b0000;
																assign node35913 = (inp[2]) ? 4'b0101 : 4'b0000;
														assign node35916 = (inp[2]) ? node35922 : node35917;
															assign node35917 = (inp[1]) ? node35919 : 4'b0100;
																assign node35919 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node35922 = (inp[1]) ? 4'b0100 : 4'b0001;
													assign node35925 = (inp[10]) ? node35927 : 4'b0000;
														assign node35927 = (inp[1]) ? node35931 : node35928;
															assign node35928 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node35931 = (inp[2]) ? 4'b0001 : 4'b0100;
												assign node35934 = (inp[11]) ? node35946 : node35935;
													assign node35935 = (inp[10]) ? node35937 : 4'b0001;
														assign node35937 = (inp[1]) ? node35939 : 4'b0101;
															assign node35939 = (inp[13]) ? node35943 : node35940;
																assign node35940 = (inp[2]) ? 4'b0101 : 4'b0000;
																assign node35943 = (inp[2]) ? 4'b0000 : 4'b0101;
													assign node35946 = (inp[1]) ? node35954 : node35947;
														assign node35947 = (inp[10]) ? 4'b0101 : node35948;
															assign node35948 = (inp[2]) ? 4'b0100 : node35949;
																assign node35949 = (inp[13]) ? 4'b0100 : 4'b0001;
														assign node35954 = (inp[2]) ? node35958 : node35955;
															assign node35955 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node35958 = (inp[13]) ? node35962 : node35959;
																assign node35959 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node35962 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node35965 = (inp[13]) ? node35997 : node35966;
												assign node35966 = (inp[2]) ? node35986 : node35967;
													assign node35967 = (inp[10]) ? node35977 : node35968;
														assign node35968 = (inp[1]) ? node35972 : node35969;
															assign node35969 = (inp[5]) ? 4'b0000 : 4'b0100;
															assign node35972 = (inp[11]) ? node35974 : 4'b0000;
																assign node35974 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node35977 = (inp[5]) ? node35981 : node35978;
															assign node35978 = (inp[1]) ? 4'b0000 : 4'b0101;
															assign node35981 = (inp[1]) ? 4'b0001 : node35982;
																assign node35982 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node35986 = (inp[1]) ? node35992 : node35987;
														assign node35987 = (inp[10]) ? 4'b0000 : node35988;
															assign node35988 = (inp[5]) ? 4'b0101 : 4'b0001;
														assign node35992 = (inp[5]) ? 4'b0100 : node35993;
															assign node35993 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node35997 = (inp[2]) ? node36009 : node35998;
													assign node35998 = (inp[5]) ? node36006 : node35999;
														assign node35999 = (inp[1]) ? node36003 : node36000;
															assign node36000 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node36003 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node36006 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node36009 = (inp[1]) ? node36017 : node36010;
														assign node36010 = (inp[5]) ? 4'b0000 : node36011;
															assign node36011 = (inp[10]) ? node36013 : 4'b0100;
																assign node36013 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node36017 = (inp[10]) ? node36019 : 4'b0001;
															assign node36019 = (inp[11]) ? 4'b0000 : node36020;
																assign node36020 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node36024 = (inp[9]) ? node36150 : node36025;
										assign node36025 = (inp[13]) ? node36087 : node36026;
											assign node36026 = (inp[2]) ? node36056 : node36027;
												assign node36027 = (inp[1]) ? node36039 : node36028;
													assign node36028 = (inp[5]) ? node36034 : node36029;
														assign node36029 = (inp[11]) ? 4'b0111 : node36030;
															assign node36030 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node36034 = (inp[10]) ? node36036 : 4'b0010;
															assign node36036 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node36039 = (inp[11]) ? node36045 : node36040;
														assign node36040 = (inp[10]) ? 4'b0011 : node36041;
															assign node36041 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node36045 = (inp[10]) ? node36051 : node36046;
															assign node36046 = (inp[5]) ? node36048 : 4'b0011;
																assign node36048 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node36051 = (inp[5]) ? node36053 : 4'b0010;
																assign node36053 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node36056 = (inp[5]) ? node36076 : node36057;
													assign node36057 = (inp[1]) ? node36067 : node36058;
														assign node36058 = (inp[11]) ? 4'b0011 : node36059;
															assign node36059 = (inp[0]) ? node36063 : node36060;
																assign node36060 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node36063 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node36067 = (inp[0]) ? node36069 : 4'b0111;
															assign node36069 = (inp[10]) ? node36073 : node36070;
																assign node36070 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node36073 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node36076 = (inp[10]) ? node36082 : node36077;
														assign node36077 = (inp[0]) ? 4'b0110 : node36078;
															assign node36078 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node36082 = (inp[11]) ? 4'b0111 : node36083;
															assign node36083 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node36087 = (inp[2]) ? node36117 : node36088;
												assign node36088 = (inp[10]) ? node36100 : node36089;
													assign node36089 = (inp[0]) ? node36095 : node36090;
														assign node36090 = (inp[11]) ? 4'b0111 : node36091;
															assign node36091 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node36095 = (inp[5]) ? 4'b0111 : node36096;
															assign node36096 = (inp[11]) ? 4'b0011 : 4'b0111;
													assign node36100 = (inp[1]) ? node36106 : node36101;
														assign node36101 = (inp[5]) ? node36103 : 4'b0010;
															assign node36103 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node36106 = (inp[0]) ? node36112 : node36107;
															assign node36107 = (inp[5]) ? node36109 : 4'b0110;
																assign node36109 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node36112 = (inp[11]) ? node36114 : 4'b0110;
																assign node36114 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node36117 = (inp[1]) ? node36135 : node36118;
													assign node36118 = (inp[5]) ? node36128 : node36119;
														assign node36119 = (inp[10]) ? node36123 : node36120;
															assign node36120 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node36123 = (inp[11]) ? node36125 : 4'b0111;
																assign node36125 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node36128 = (inp[11]) ? node36132 : node36129;
															assign node36129 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node36132 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node36135 = (inp[10]) ? node36145 : node36136;
														assign node36136 = (inp[0]) ? node36140 : node36137;
															assign node36137 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node36140 = (inp[5]) ? 4'b0010 : node36141;
																assign node36141 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node36145 = (inp[0]) ? node36147 : 4'b0011;
															assign node36147 = (inp[11]) ? 4'b0010 : 4'b0011;
										assign node36150 = (inp[10]) ? node36220 : node36151;
											assign node36151 = (inp[2]) ? node36183 : node36152;
												assign node36152 = (inp[13]) ? node36162 : node36153;
													assign node36153 = (inp[5]) ? 4'b0011 : node36154;
														assign node36154 = (inp[1]) ? node36156 : 4'b0110;
															assign node36156 = (inp[11]) ? 4'b0010 : node36157;
																assign node36157 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node36162 = (inp[1]) ? node36174 : node36163;
														assign node36163 = (inp[5]) ? node36169 : node36164;
															assign node36164 = (inp[11]) ? 4'b0010 : node36165;
																assign node36165 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node36169 = (inp[11]) ? 4'b0110 : node36170;
																assign node36170 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node36174 = (inp[11]) ? node36178 : node36175;
															assign node36175 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node36178 = (inp[0]) ? node36180 : 4'b0110;
																assign node36180 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node36183 = (inp[13]) ? node36201 : node36184;
													assign node36184 = (inp[1]) ? node36192 : node36185;
														assign node36185 = (inp[5]) ? 4'b0111 : node36186;
															assign node36186 = (inp[0]) ? 4'b0011 : node36187;
																assign node36187 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node36192 = (inp[5]) ? node36196 : node36193;
															assign node36193 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node36196 = (inp[11]) ? 4'b0111 : node36197;
																assign node36197 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node36201 = (inp[1]) ? node36209 : node36202;
														assign node36202 = (inp[5]) ? 4'b0011 : node36203;
															assign node36203 = (inp[11]) ? node36205 : 4'b0111;
																assign node36205 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node36209 = (inp[0]) ? node36215 : node36210;
															assign node36210 = (inp[5]) ? node36212 : 4'b0011;
																assign node36212 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node36215 = (inp[5]) ? 4'b0011 : node36216;
																assign node36216 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node36220 = (inp[2]) ? node36254 : node36221;
												assign node36221 = (inp[13]) ? node36241 : node36222;
													assign node36222 = (inp[1]) ? node36230 : node36223;
														assign node36223 = (inp[5]) ? 4'b0010 : node36224;
															assign node36224 = (inp[11]) ? 4'b0111 : node36225;
																assign node36225 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node36230 = (inp[11]) ? node36236 : node36231;
															assign node36231 = (inp[0]) ? node36233 : 4'b0010;
																assign node36233 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node36236 = (inp[0]) ? 4'b0011 : node36237;
																assign node36237 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node36241 = (inp[1]) ? 4'b0111 : node36242;
														assign node36242 = (inp[5]) ? node36248 : node36243;
															assign node36243 = (inp[11]) ? 4'b0011 : node36244;
																assign node36244 = (inp[0]) ? 4'b0011 : 4'b0010;
															assign node36248 = (inp[0]) ? 4'b0111 : node36249;
																assign node36249 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node36254 = (inp[13]) ? node36270 : node36255;
													assign node36255 = (inp[1]) ? node36265 : node36256;
														assign node36256 = (inp[5]) ? node36262 : node36257;
															assign node36257 = (inp[11]) ? 4'b0010 : node36258;
																assign node36258 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node36262 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node36265 = (inp[11]) ? node36267 : 4'b0110;
															assign node36267 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node36270 = (inp[5]) ? node36278 : node36271;
														assign node36271 = (inp[1]) ? 4'b0010 : node36272;
															assign node36272 = (inp[11]) ? node36274 : 4'b0110;
																assign node36274 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node36278 = (inp[0]) ? 4'b0010 : node36279;
															assign node36279 = (inp[11]) ? 4'b0010 : 4'b0011;
								assign node36283 = (inp[9]) ? node36629 : node36284;
									assign node36284 = (inp[5]) ? node36476 : node36285;
										assign node36285 = (inp[11]) ? node36377 : node36286;
											assign node36286 = (inp[10]) ? node36330 : node36287;
												assign node36287 = (inp[15]) ? node36313 : node36288;
													assign node36288 = (inp[0]) ? node36302 : node36289;
														assign node36289 = (inp[1]) ? node36295 : node36290;
															assign node36290 = (inp[13]) ? node36292 : 4'b0110;
																assign node36292 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node36295 = (inp[13]) ? node36299 : node36296;
																assign node36296 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node36299 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node36302 = (inp[1]) ? node36308 : node36303;
															assign node36303 = (inp[13]) ? node36305 : 4'b0010;
																assign node36305 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node36308 = (inp[2]) ? 4'b0111 : node36309;
																assign node36309 = (inp[13]) ? 4'b0010 : 4'b0111;
													assign node36313 = (inp[0]) ? node36321 : node36314;
														assign node36314 = (inp[13]) ? 4'b0110 : node36315;
															assign node36315 = (inp[1]) ? node36317 : 4'b0010;
																assign node36317 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node36321 = (inp[2]) ? 4'b0111 : node36322;
															assign node36322 = (inp[13]) ? node36326 : node36323;
																assign node36323 = (inp[1]) ? 4'b0010 : 4'b0110;
																assign node36326 = (inp[1]) ? 4'b0111 : 4'b0010;
												assign node36330 = (inp[0]) ? node36354 : node36331;
													assign node36331 = (inp[15]) ? node36341 : node36332;
														assign node36332 = (inp[13]) ? node36338 : node36333;
															assign node36333 = (inp[1]) ? 4'b0010 : node36334;
																assign node36334 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node36338 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node36341 = (inp[2]) ? node36347 : node36342;
															assign node36342 = (inp[13]) ? 4'b0011 : node36343;
																assign node36343 = (inp[1]) ? 4'b0011 : 4'b0111;
															assign node36347 = (inp[1]) ? node36351 : node36348;
																assign node36348 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node36351 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node36354 = (inp[2]) ? node36364 : node36355;
														assign node36355 = (inp[1]) ? node36357 : 4'b0011;
															assign node36357 = (inp[15]) ? node36361 : node36358;
																assign node36358 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node36361 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node36364 = (inp[1]) ? node36370 : node36365;
															assign node36365 = (inp[13]) ? node36367 : 4'b0110;
																assign node36367 = (inp[15]) ? 4'b0110 : 4'b0011;
															assign node36370 = (inp[15]) ? node36374 : node36371;
																assign node36371 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node36374 = (inp[13]) ? 4'b0010 : 4'b0110;
											assign node36377 = (inp[10]) ? node36431 : node36378;
												assign node36378 = (inp[0]) ? node36406 : node36379;
													assign node36379 = (inp[1]) ? node36391 : node36380;
														assign node36380 = (inp[13]) ? node36386 : node36381;
															assign node36381 = (inp[15]) ? node36383 : 4'b0111;
																assign node36383 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node36386 = (inp[2]) ? 4'b0010 : node36387;
																assign node36387 = (inp[15]) ? 4'b0010 : 4'b0110;
														assign node36391 = (inp[2]) ? node36399 : node36392;
															assign node36392 = (inp[13]) ? node36396 : node36393;
																assign node36393 = (inp[15]) ? 4'b0010 : 4'b0111;
																assign node36396 = (inp[15]) ? 4'b0111 : 4'b0010;
															assign node36399 = (inp[13]) ? node36403 : node36400;
																assign node36400 = (inp[15]) ? 4'b0111 : 4'b0011;
																assign node36403 = (inp[15]) ? 4'b0011 : 4'b0111;
													assign node36406 = (inp[15]) ? node36418 : node36407;
														assign node36407 = (inp[1]) ? node36411 : node36408;
															assign node36408 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node36411 = (inp[13]) ? node36415 : node36412;
																assign node36412 = (inp[2]) ? 4'b0010 : 4'b0110;
																assign node36415 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node36418 = (inp[13]) ? node36426 : node36419;
															assign node36419 = (inp[1]) ? node36423 : node36420;
																assign node36420 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node36423 = (inp[2]) ? 4'b0111 : 4'b0011;
															assign node36426 = (inp[1]) ? 4'b0011 : node36427;
																assign node36427 = (inp[2]) ? 4'b0111 : 4'b0011;
												assign node36431 = (inp[15]) ? node36455 : node36432;
													assign node36432 = (inp[1]) ? node36440 : node36433;
														assign node36433 = (inp[0]) ? node36435 : 4'b0011;
															assign node36435 = (inp[13]) ? node36437 : 4'b0110;
																assign node36437 = (inp[2]) ? 4'b0011 : 4'b0111;
														assign node36440 = (inp[0]) ? node36448 : node36441;
															assign node36441 = (inp[13]) ? node36445 : node36442;
																assign node36442 = (inp[2]) ? 4'b0010 : 4'b0110;
																assign node36445 = (inp[2]) ? 4'b0110 : 4'b0011;
															assign node36448 = (inp[13]) ? node36452 : node36449;
																assign node36449 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node36452 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node36455 = (inp[0]) ? node36467 : node36456;
														assign node36456 = (inp[1]) ? node36462 : node36457;
															assign node36457 = (inp[13]) ? 4'b0110 : node36458;
																assign node36458 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node36462 = (inp[13]) ? node36464 : 4'b0110;
																assign node36464 = (inp[2]) ? 4'b0010 : 4'b0110;
														assign node36467 = (inp[13]) ? 4'b0010 : node36468;
															assign node36468 = (inp[2]) ? node36472 : node36469;
																assign node36469 = (inp[1]) ? 4'b0010 : 4'b0110;
																assign node36472 = (inp[1]) ? 4'b0110 : 4'b0010;
										assign node36476 = (inp[10]) ? node36554 : node36477;
											assign node36477 = (inp[0]) ? node36519 : node36478;
												assign node36478 = (inp[11]) ? node36498 : node36479;
													assign node36479 = (inp[15]) ? node36491 : node36480;
														assign node36480 = (inp[2]) ? node36488 : node36481;
															assign node36481 = (inp[13]) ? node36485 : node36482;
																assign node36482 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node36485 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node36488 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node36491 = (inp[2]) ? node36495 : node36492;
															assign node36492 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node36495 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node36498 = (inp[2]) ? node36510 : node36499;
														assign node36499 = (inp[1]) ? node36505 : node36500;
															assign node36500 = (inp[15]) ? node36502 : 4'b0011;
																assign node36502 = (inp[13]) ? 4'b0110 : 4'b0011;
															assign node36505 = (inp[15]) ? 4'b0110 : node36506;
																assign node36506 = (inp[13]) ? 4'b0011 : 4'b0110;
														assign node36510 = (inp[13]) ? node36514 : node36511;
															assign node36511 = (inp[15]) ? 4'b0110 : 4'b0010;
															assign node36514 = (inp[15]) ? 4'b0010 : node36515;
																assign node36515 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node36519 = (inp[2]) ? node36543 : node36520;
													assign node36520 = (inp[11]) ? node36534 : node36521;
														assign node36521 = (inp[1]) ? node36529 : node36522;
															assign node36522 = (inp[13]) ? node36526 : node36523;
																assign node36523 = (inp[15]) ? 4'b0011 : 4'b0110;
																assign node36526 = (inp[15]) ? 4'b0110 : 4'b0011;
															assign node36529 = (inp[15]) ? 4'b0110 : node36530;
																assign node36530 = (inp[13]) ? 4'b0011 : 4'b0110;
														assign node36534 = (inp[13]) ? node36538 : node36535;
															assign node36535 = (inp[15]) ? 4'b0010 : 4'b0110;
															assign node36538 = (inp[1]) ? node36540 : 4'b0011;
																assign node36540 = (inp[15]) ? 4'b0110 : 4'b0010;
													assign node36543 = (inp[13]) ? node36551 : node36544;
														assign node36544 = (inp[15]) ? 4'b0110 : node36545;
															assign node36545 = (inp[11]) ? node36547 : 4'b0010;
																assign node36547 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node36551 = (inp[15]) ? 4'b0010 : 4'b0110;
											assign node36554 = (inp[2]) ? node36592 : node36555;
												assign node36555 = (inp[1]) ? node36573 : node36556;
													assign node36556 = (inp[0]) ? node36566 : node36557;
														assign node36557 = (inp[11]) ? 4'b0010 : node36558;
															assign node36558 = (inp[15]) ? node36562 : node36559;
																assign node36559 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node36562 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node36566 = (inp[15]) ? node36570 : node36567;
															assign node36567 = (inp[13]) ? 4'b0010 : 4'b0111;
															assign node36570 = (inp[13]) ? 4'b0111 : 4'b0010;
													assign node36573 = (inp[13]) ? node36585 : node36574;
														assign node36574 = (inp[15]) ? node36580 : node36575;
															assign node36575 = (inp[0]) ? node36577 : 4'b0111;
																assign node36577 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node36580 = (inp[11]) ? node36582 : 4'b0010;
																assign node36582 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node36585 = (inp[15]) ? node36587 : 4'b0010;
															assign node36587 = (inp[0]) ? 4'b0111 : node36588;
																assign node36588 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node36592 = (inp[0]) ? node36616 : node36593;
													assign node36593 = (inp[11]) ? node36607 : node36594;
														assign node36594 = (inp[1]) ? node36602 : node36595;
															assign node36595 = (inp[15]) ? node36599 : node36596;
																assign node36596 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node36599 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node36602 = (inp[13]) ? 4'b0110 : node36603;
																assign node36603 = (inp[15]) ? 4'b0110 : 4'b0011;
														assign node36607 = (inp[15]) ? node36613 : node36608;
															assign node36608 = (inp[13]) ? node36610 : 4'b0011;
																assign node36610 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node36613 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node36616 = (inp[15]) ? node36626 : node36617;
														assign node36617 = (inp[13]) ? node36621 : node36618;
															assign node36618 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node36621 = (inp[11]) ? 4'b0111 : node36622;
																assign node36622 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node36626 = (inp[13]) ? 4'b0011 : 4'b0111;
									assign node36629 = (inp[10]) ? node36787 : node36630;
										assign node36630 = (inp[1]) ? node36712 : node36631;
											assign node36631 = (inp[2]) ? node36677 : node36632;
												assign node36632 = (inp[0]) ? node36652 : node36633;
													assign node36633 = (inp[11]) ? node36643 : node36634;
														assign node36634 = (inp[5]) ? 4'b0011 : node36635;
															assign node36635 = (inp[15]) ? node36639 : node36636;
																assign node36636 = (inp[13]) ? 4'b0110 : 4'b0011;
																assign node36639 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node36643 = (inp[5]) ? 4'b0111 : node36644;
															assign node36644 = (inp[15]) ? node36648 : node36645;
																assign node36645 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node36648 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node36652 = (inp[15]) ? node36666 : node36653;
														assign node36653 = (inp[11]) ? node36659 : node36654;
															assign node36654 = (inp[13]) ? node36656 : 4'b0111;
																assign node36656 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node36659 = (inp[5]) ? node36663 : node36660;
																assign node36660 = (inp[13]) ? 4'b0111 : 4'b0010;
																assign node36663 = (inp[13]) ? 4'b0010 : 4'b0111;
														assign node36666 = (inp[13]) ? node36672 : node36667;
															assign node36667 = (inp[5]) ? node36669 : 4'b0111;
																assign node36669 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node36672 = (inp[5]) ? 4'b0111 : node36673;
																assign node36673 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node36677 = (inp[0]) ? node36695 : node36678;
													assign node36678 = (inp[11]) ? node36686 : node36679;
														assign node36679 = (inp[5]) ? node36683 : node36680;
															assign node36680 = (inp[15]) ? 4'b0011 : 4'b0010;
															assign node36683 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node36686 = (inp[5]) ? 4'b0011 : node36687;
															assign node36687 = (inp[15]) ? node36691 : node36688;
																assign node36688 = (inp[13]) ? 4'b0011 : 4'b0110;
																assign node36691 = (inp[13]) ? 4'b0110 : 4'b0011;
													assign node36695 = (inp[11]) ? node36701 : node36696;
														assign node36696 = (inp[15]) ? node36698 : 4'b0011;
															assign node36698 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node36701 = (inp[5]) ? node36707 : node36702;
															assign node36702 = (inp[13]) ? node36704 : 4'b0110;
																assign node36704 = (inp[15]) ? 4'b0110 : 4'b0011;
															assign node36707 = (inp[13]) ? 4'b0111 : node36708;
																assign node36708 = (inp[15]) ? 4'b0111 : 4'b0011;
											assign node36712 = (inp[5]) ? node36754 : node36713;
												assign node36713 = (inp[2]) ? node36733 : node36714;
													assign node36714 = (inp[11]) ? node36722 : node36715;
														assign node36715 = (inp[15]) ? node36719 : node36716;
															assign node36716 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node36719 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node36722 = (inp[15]) ? node36728 : node36723;
															assign node36723 = (inp[13]) ? 4'b0011 : node36724;
																assign node36724 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node36728 = (inp[13]) ? 4'b0110 : node36729;
																assign node36729 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node36733 = (inp[0]) ? node36745 : node36734;
														assign node36734 = (inp[11]) ? node36742 : node36735;
															assign node36735 = (inp[15]) ? node36739 : node36736;
																assign node36736 = (inp[13]) ? 4'b0111 : 4'b0010;
																assign node36739 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node36742 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node36745 = (inp[15]) ? node36751 : node36746;
															assign node36746 = (inp[13]) ? 4'b0110 : node36747;
																assign node36747 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node36751 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node36754 = (inp[0]) ? node36770 : node36755;
													assign node36755 = (inp[15]) ? node36763 : node36756;
														assign node36756 = (inp[2]) ? node36760 : node36757;
															assign node36757 = (inp[13]) ? 4'b0010 : 4'b0111;
															assign node36760 = (inp[13]) ? 4'b0111 : 4'b0011;
														assign node36763 = (inp[13]) ? node36767 : node36764;
															assign node36764 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node36767 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node36770 = (inp[15]) ? node36778 : node36771;
														assign node36771 = (inp[13]) ? node36775 : node36772;
															assign node36772 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node36775 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node36778 = (inp[11]) ? node36780 : 4'b0111;
															assign node36780 = (inp[13]) ? node36784 : node36781;
																assign node36781 = (inp[2]) ? 4'b0111 : 4'b0011;
																assign node36784 = (inp[2]) ? 4'b0011 : 4'b0111;
										assign node36787 = (inp[1]) ? node36859 : node36788;
											assign node36788 = (inp[5]) ? node36830 : node36789;
												assign node36789 = (inp[0]) ? node36811 : node36790;
													assign node36790 = (inp[15]) ? node36802 : node36791;
														assign node36791 = (inp[2]) ? node36797 : node36792;
															assign node36792 = (inp[13]) ? node36794 : 4'b0010;
																assign node36794 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node36797 = (inp[13]) ? node36799 : 4'b0111;
																assign node36799 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node36802 = (inp[11]) ? 4'b0010 : node36803;
															assign node36803 = (inp[2]) ? node36807 : node36804;
																assign node36804 = (inp[13]) ? 4'b0010 : 4'b0110;
																assign node36807 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node36811 = (inp[11]) ? node36823 : node36812;
														assign node36812 = (inp[15]) ? node36818 : node36813;
															assign node36813 = (inp[13]) ? node36815 : 4'b0010;
																assign node36815 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node36818 = (inp[2]) ? 4'b0111 : node36819;
																assign node36819 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node36823 = (inp[2]) ? 4'b0111 : node36824;
															assign node36824 = (inp[15]) ? node36826 : 4'b0011;
																assign node36826 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node36830 = (inp[0]) ? node36850 : node36831;
													assign node36831 = (inp[11]) ? node36841 : node36832;
														assign node36832 = (inp[13]) ? 4'b0111 : node36833;
															assign node36833 = (inp[15]) ? node36837 : node36834;
																assign node36834 = (inp[2]) ? 4'b0011 : 4'b0111;
																assign node36837 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node36841 = (inp[13]) ? node36845 : node36842;
															assign node36842 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node36845 = (inp[15]) ? 4'b0110 : node36846;
																assign node36846 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node36850 = (inp[2]) ? node36852 : 4'b0110;
														assign node36852 = (inp[13]) ? node36856 : node36853;
															assign node36853 = (inp[15]) ? 4'b0110 : 4'b0010;
															assign node36856 = (inp[15]) ? 4'b0010 : 4'b0111;
											assign node36859 = (inp[5]) ? node36897 : node36860;
												assign node36860 = (inp[0]) ? node36880 : node36861;
													assign node36861 = (inp[15]) ? node36871 : node36862;
														assign node36862 = (inp[13]) ? node36866 : node36863;
															assign node36863 = (inp[2]) ? 4'b0011 : 4'b0111;
															assign node36866 = (inp[2]) ? node36868 : 4'b0010;
																assign node36868 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node36871 = (inp[11]) ? 4'b0010 : node36872;
															assign node36872 = (inp[13]) ? node36876 : node36873;
																assign node36873 = (inp[2]) ? 4'b0110 : 4'b0010;
																assign node36876 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node36880 = (inp[2]) ? node36890 : node36881;
														assign node36881 = (inp[11]) ? 4'b0011 : node36882;
															assign node36882 = (inp[13]) ? node36886 : node36883;
																assign node36883 = (inp[15]) ? 4'b0010 : 4'b0111;
																assign node36886 = (inp[15]) ? 4'b0111 : 4'b0010;
														assign node36890 = (inp[13]) ? node36894 : node36891;
															assign node36891 = (inp[15]) ? 4'b0111 : 4'b0011;
															assign node36894 = (inp[15]) ? 4'b0011 : 4'b0111;
												assign node36897 = (inp[0]) ? node36913 : node36898;
													assign node36898 = (inp[15]) ? node36908 : node36899;
														assign node36899 = (inp[13]) ? node36903 : node36900;
															assign node36900 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node36903 = (inp[2]) ? node36905 : 4'b0011;
																assign node36905 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node36908 = (inp[2]) ? node36910 : 4'b0011;
															assign node36910 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node36913 = (inp[15]) ? node36925 : node36914;
														assign node36914 = (inp[13]) ? node36920 : node36915;
															assign node36915 = (inp[11]) ? 4'b0011 : node36916;
																assign node36916 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node36920 = (inp[11]) ? node36922 : 4'b0011;
																assign node36922 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node36925 = (inp[13]) ? node36929 : node36926;
															assign node36926 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node36929 = (inp[2]) ? 4'b0010 : 4'b0110;
						assign node36932 = (inp[2]) ? node37350 : node36933;
							assign node36933 = (inp[9]) ? node37145 : node36934;
								assign node36934 = (inp[4]) ? node37026 : node36935;
									assign node36935 = (inp[5]) ? node36991 : node36936;
										assign node36936 = (inp[0]) ? node36964 : node36937;
											assign node36937 = (inp[1]) ? node36949 : node36938;
												assign node36938 = (inp[13]) ? node36942 : node36939;
													assign node36939 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node36942 = (inp[12]) ? node36946 : node36943;
														assign node36943 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node36946 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node36949 = (inp[15]) ? node36957 : node36950;
													assign node36950 = (inp[12]) ? node36954 : node36951;
														assign node36951 = (inp[13]) ? 4'b0011 : 4'b0110;
														assign node36954 = (inp[13]) ? 4'b0110 : 4'b0011;
													assign node36957 = (inp[13]) ? node36961 : node36958;
														assign node36958 = (inp[12]) ? 4'b0110 : 4'b0011;
														assign node36961 = (inp[12]) ? 4'b0010 : 4'b0110;
											assign node36964 = (inp[12]) ? node36980 : node36965;
												assign node36965 = (inp[13]) ? node36973 : node36966;
													assign node36966 = (inp[15]) ? node36970 : node36967;
														assign node36967 = (inp[1]) ? 4'b0111 : 4'b0011;
														assign node36970 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node36973 = (inp[1]) ? node36977 : node36974;
														assign node36974 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node36977 = (inp[15]) ? 4'b0110 : 4'b0010;
												assign node36980 = (inp[13]) ? node36986 : node36981;
													assign node36981 = (inp[1]) ? node36983 : 4'b0111;
														assign node36983 = (inp[15]) ? 4'b0111 : 4'b0011;
													assign node36986 = (inp[15]) ? 4'b0011 : node36987;
														assign node36987 = (inp[1]) ? 4'b0111 : 4'b0010;
										assign node36991 = (inp[12]) ? node37013 : node36992;
											assign node36992 = (inp[13]) ? node37000 : node36993;
												assign node36993 = (inp[15]) ? node36997 : node36994;
													assign node36994 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node36997 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node37000 = (inp[1]) ? node37008 : node37001;
													assign node37001 = (inp[0]) ? node37005 : node37002;
														assign node37002 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node37005 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node37008 = (inp[15]) ? node37010 : 4'b0011;
														assign node37010 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node37013 = (inp[13]) ? node37021 : node37014;
												assign node37014 = (inp[1]) ? node37016 : 4'b0110;
													assign node37016 = (inp[15]) ? 4'b0110 : node37017;
														assign node37017 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node37021 = (inp[15]) ? 4'b0010 : node37022;
													assign node37022 = (inp[1]) ? 4'b0110 : 4'b0011;
									assign node37026 = (inp[5]) ? node37084 : node37027;
										assign node37027 = (inp[12]) ? node37069 : node37028;
											assign node37028 = (inp[15]) ? node37040 : node37029;
												assign node37029 = (inp[13]) ? node37035 : node37030;
													assign node37030 = (inp[0]) ? node37032 : 4'b0010;
														assign node37032 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node37035 = (inp[11]) ? node37037 : 4'b0110;
														assign node37037 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node37040 = (inp[13]) ? node37056 : node37041;
													assign node37041 = (inp[11]) ? node37049 : node37042;
														assign node37042 = (inp[0]) ? node37046 : node37043;
															assign node37043 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node37046 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node37049 = (inp[0]) ? node37053 : node37050;
															assign node37050 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node37053 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node37056 = (inp[11]) ? node37064 : node37057;
														assign node37057 = (inp[0]) ? node37061 : node37058;
															assign node37058 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node37061 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node37064 = (inp[1]) ? node37066 : 4'b0010;
															assign node37066 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node37069 = (inp[15]) ? node37081 : node37070;
												assign node37070 = (inp[13]) ? node37076 : node37071;
													assign node37071 = (inp[0]) ? node37073 : 4'b0010;
														assign node37073 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node37076 = (inp[0]) ? 4'b0110 : node37077;
														assign node37077 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node37081 = (inp[13]) ? 4'b0010 : 4'b0110;
										assign node37084 = (inp[12]) ? node37130 : node37085;
											assign node37085 = (inp[15]) ? node37097 : node37086;
												assign node37086 = (inp[13]) ? node37092 : node37087;
													assign node37087 = (inp[0]) ? node37089 : 4'b0011;
														assign node37089 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node37092 = (inp[1]) ? node37094 : 4'b0111;
														assign node37094 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node37097 = (inp[13]) ? node37117 : node37098;
													assign node37098 = (inp[10]) ? node37112 : node37099;
														assign node37099 = (inp[11]) ? node37105 : node37100;
															assign node37100 = (inp[1]) ? 4'b0111 : node37101;
																assign node37101 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node37105 = (inp[1]) ? node37109 : node37106;
																assign node37106 = (inp[0]) ? 4'b0110 : 4'b0111;
																assign node37109 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node37112 = (inp[1]) ? node37114 : 4'b0110;
															assign node37114 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node37117 = (inp[11]) ? node37125 : node37118;
														assign node37118 = (inp[0]) ? node37122 : node37119;
															assign node37119 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node37122 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node37125 = (inp[1]) ? node37127 : 4'b0010;
															assign node37127 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node37130 = (inp[15]) ? node37142 : node37131;
												assign node37131 = (inp[13]) ? node37137 : node37132;
													assign node37132 = (inp[1]) ? node37134 : 4'b0011;
														assign node37134 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node37137 = (inp[0]) ? 4'b0111 : node37138;
														assign node37138 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node37142 = (inp[13]) ? 4'b0011 : 4'b0111;
								assign node37145 = (inp[5]) ? node37261 : node37146;
									assign node37146 = (inp[4]) ? node37198 : node37147;
										assign node37147 = (inp[0]) ? node37173 : node37148;
											assign node37148 = (inp[13]) ? node37158 : node37149;
												assign node37149 = (inp[12]) ? node37153 : node37150;
													assign node37150 = (inp[1]) ? 4'b0111 : 4'b0011;
													assign node37153 = (inp[15]) ? 4'b0111 : node37154;
														assign node37154 = (inp[1]) ? 4'b0010 : 4'b0111;
												assign node37158 = (inp[12]) ? node37166 : node37159;
													assign node37159 = (inp[1]) ? node37163 : node37160;
														assign node37160 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node37163 = (inp[15]) ? 4'b0111 : 4'b0010;
													assign node37166 = (inp[1]) ? node37170 : node37167;
														assign node37167 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node37170 = (inp[15]) ? 4'b0011 : 4'b0111;
											assign node37173 = (inp[13]) ? node37185 : node37174;
												assign node37174 = (inp[12]) ? node37180 : node37175;
													assign node37175 = (inp[1]) ? node37177 : 4'b0010;
														assign node37177 = (inp[15]) ? 4'b0011 : 4'b0110;
													assign node37180 = (inp[15]) ? 4'b0110 : node37181;
														assign node37181 = (inp[1]) ? 4'b0010 : 4'b0110;
												assign node37185 = (inp[12]) ? node37193 : node37186;
													assign node37186 = (inp[15]) ? node37190 : node37187;
														assign node37187 = (inp[1]) ? 4'b0011 : 4'b0111;
														assign node37190 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node37193 = (inp[15]) ? 4'b0010 : node37194;
														assign node37194 = (inp[1]) ? 4'b0110 : 4'b0011;
										assign node37198 = (inp[12]) ? node37246 : node37199;
											assign node37199 = (inp[15]) ? node37211 : node37200;
												assign node37200 = (inp[13]) ? node37206 : node37201;
													assign node37201 = (inp[1]) ? 4'b0011 : node37202;
														assign node37202 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node37206 = (inp[1]) ? node37208 : 4'b0111;
														assign node37208 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node37211 = (inp[13]) ? node37223 : node37212;
													assign node37212 = (inp[10]) ? node37214 : 4'b0110;
														assign node37214 = (inp[11]) ? node37218 : node37215;
															assign node37215 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node37218 = (inp[0]) ? 4'b0111 : node37219;
																assign node37219 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node37223 = (inp[10]) ? node37237 : node37224;
														assign node37224 = (inp[11]) ? node37230 : node37225;
															assign node37225 = (inp[0]) ? 4'b0011 : node37226;
																assign node37226 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node37230 = (inp[0]) ? node37234 : node37231;
																assign node37231 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node37234 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node37237 = (inp[11]) ? 4'b0010 : node37238;
															assign node37238 = (inp[1]) ? node37242 : node37239;
																assign node37239 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node37242 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node37246 = (inp[15]) ? node37258 : node37247;
												assign node37247 = (inp[13]) ? node37253 : node37248;
													assign node37248 = (inp[1]) ? node37250 : 4'b0011;
														assign node37250 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node37253 = (inp[0]) ? 4'b0111 : node37254;
														assign node37254 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node37258 = (inp[13]) ? 4'b0011 : 4'b0111;
									assign node37261 = (inp[4]) ? node37301 : node37262;
										assign node37262 = (inp[13]) ? node37276 : node37263;
											assign node37263 = (inp[12]) ? node37269 : node37264;
												assign node37264 = (inp[1]) ? node37266 : 4'b0011;
													assign node37266 = (inp[15]) ? 4'b0010 : 4'b0111;
												assign node37269 = (inp[15]) ? 4'b0111 : node37270;
													assign node37270 = (inp[1]) ? node37272 : 4'b0111;
														assign node37272 = (inp[0]) ? 4'b0010 : 4'b0011;
											assign node37276 = (inp[12]) ? node37296 : node37277;
												assign node37277 = (inp[15]) ? node37283 : node37278;
													assign node37278 = (inp[1]) ? 4'b0010 : node37279;
														assign node37279 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node37283 = (inp[10]) ? node37289 : node37284;
														assign node37284 = (inp[0]) ? 4'b0110 : node37285;
															assign node37285 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node37289 = (inp[0]) ? node37293 : node37290;
															assign node37290 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node37293 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node37296 = (inp[15]) ? 4'b0011 : node37297;
													assign node37297 = (inp[1]) ? 4'b0111 : 4'b0010;
										assign node37301 = (inp[12]) ? node37335 : node37302;
											assign node37302 = (inp[15]) ? node37314 : node37303;
												assign node37303 = (inp[13]) ? node37309 : node37304;
													assign node37304 = (inp[1]) ? 4'b0010 : node37305;
														assign node37305 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node37309 = (inp[0]) ? 4'b0110 : node37310;
														assign node37310 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node37314 = (inp[13]) ? node37328 : node37315;
													assign node37315 = (inp[11]) ? node37317 : 4'b0111;
														assign node37317 = (inp[10]) ? node37323 : node37318;
															assign node37318 = (inp[1]) ? node37320 : 4'b0111;
																assign node37320 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node37323 = (inp[1]) ? node37325 : 4'b0110;
																assign node37325 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node37328 = (inp[0]) ? node37332 : node37329;
														assign node37329 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node37332 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node37335 = (inp[15]) ? node37347 : node37336;
												assign node37336 = (inp[13]) ? node37342 : node37337;
													assign node37337 = (inp[1]) ? node37339 : 4'b0010;
														assign node37339 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node37342 = (inp[1]) ? 4'b0110 : node37343;
														assign node37343 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node37347 = (inp[13]) ? 4'b0010 : 4'b0110;
							assign node37350 = (inp[9]) ? node37544 : node37351;
								assign node37351 = (inp[5]) ? node37465 : node37352;
									assign node37352 = (inp[4]) ? node37410 : node37353;
										assign node37353 = (inp[0]) ? node37381 : node37354;
											assign node37354 = (inp[13]) ? node37366 : node37355;
												assign node37355 = (inp[1]) ? node37359 : node37356;
													assign node37356 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node37359 = (inp[12]) ? node37363 : node37360;
														assign node37360 = (inp[15]) ? 4'b0010 : 4'b0111;
														assign node37363 = (inp[15]) ? 4'b0111 : 4'b0010;
												assign node37366 = (inp[12]) ? node37374 : node37367;
													assign node37367 = (inp[1]) ? node37371 : node37368;
														assign node37368 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node37371 = (inp[15]) ? 4'b0111 : 4'b0010;
													assign node37374 = (inp[1]) ? node37378 : node37375;
														assign node37375 = (inp[15]) ? 4'b0011 : 4'b0010;
														assign node37378 = (inp[15]) ? 4'b0011 : 4'b0111;
											assign node37381 = (inp[12]) ? node37397 : node37382;
												assign node37382 = (inp[13]) ? node37390 : node37383;
													assign node37383 = (inp[15]) ? node37387 : node37384;
														assign node37384 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node37387 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node37390 = (inp[1]) ? node37394 : node37391;
														assign node37391 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node37394 = (inp[15]) ? 4'b0111 : 4'b0011;
												assign node37397 = (inp[13]) ? node37403 : node37398;
													assign node37398 = (inp[1]) ? node37400 : 4'b0110;
														assign node37400 = (inp[15]) ? 4'b0110 : 4'b0010;
													assign node37403 = (inp[1]) ? node37407 : node37404;
														assign node37404 = (inp[15]) ? 4'b0010 : 4'b0011;
														assign node37407 = (inp[15]) ? 4'b0010 : 4'b0110;
										assign node37410 = (inp[12]) ? node37450 : node37411;
											assign node37411 = (inp[15]) ? node37423 : node37412;
												assign node37412 = (inp[13]) ? node37418 : node37413;
													assign node37413 = (inp[0]) ? node37415 : 4'b0010;
														assign node37415 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node37418 = (inp[0]) ? 4'b0110 : node37419;
														assign node37419 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node37423 = (inp[13]) ? node37437 : node37424;
													assign node37424 = (inp[10]) ? node37430 : node37425;
														assign node37425 = (inp[1]) ? node37427 : 4'b0110;
															assign node37427 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node37430 = (inp[0]) ? node37434 : node37431;
															assign node37431 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node37434 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node37437 = (inp[11]) ? node37443 : node37438;
														assign node37438 = (inp[0]) ? 4'b0011 : node37439;
															assign node37439 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node37443 = (inp[0]) ? node37447 : node37444;
															assign node37444 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node37447 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node37450 = (inp[15]) ? node37462 : node37451;
												assign node37451 = (inp[13]) ? node37457 : node37452;
													assign node37452 = (inp[0]) ? node37454 : 4'b0010;
														assign node37454 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node37457 = (inp[0]) ? 4'b0110 : node37458;
														assign node37458 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node37462 = (inp[13]) ? 4'b0010 : 4'b0110;
									assign node37465 = (inp[12]) ? node37525 : node37466;
										assign node37466 = (inp[13]) ? node37488 : node37467;
											assign node37467 = (inp[15]) ? node37477 : node37468;
												assign node37468 = (inp[1]) ? node37474 : node37469;
													assign node37469 = (inp[0]) ? node37471 : 4'b0011;
														assign node37471 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node37474 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node37477 = (inp[4]) ? node37481 : node37478;
													assign node37478 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node37481 = (inp[1]) ? node37485 : node37482;
														assign node37482 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node37485 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node37488 = (inp[1]) ? node37502 : node37489;
												assign node37489 = (inp[15]) ? node37495 : node37490;
													assign node37490 = (inp[0]) ? 4'b0111 : node37491;
														assign node37491 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node37495 = (inp[0]) ? node37499 : node37496;
														assign node37496 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node37499 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node37502 = (inp[0]) ? node37518 : node37503;
													assign node37503 = (inp[11]) ? node37511 : node37504;
														assign node37504 = (inp[15]) ? node37508 : node37505;
															assign node37505 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node37508 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node37511 = (inp[10]) ? 4'b0010 : node37512;
															assign node37512 = (inp[15]) ? node37514 : 4'b0010;
																assign node37514 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node37518 = (inp[15]) ? node37522 : node37519;
														assign node37519 = (inp[4]) ? 4'b0111 : 4'b0010;
														assign node37522 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node37525 = (inp[15]) ? node37541 : node37526;
											assign node37526 = (inp[13]) ? node37534 : node37527;
												assign node37527 = (inp[1]) ? node37531 : node37528;
													assign node37528 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node37531 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node37534 = (inp[1]) ? 4'b0111 : node37535;
													assign node37535 = (inp[4]) ? node37537 : 4'b0010;
														assign node37537 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node37541 = (inp[13]) ? 4'b0011 : 4'b0111;
								assign node37544 = (inp[5]) ? node37672 : node37545;
									assign node37545 = (inp[4]) ? node37613 : node37546;
										assign node37546 = (inp[0]) ? node37588 : node37547;
											assign node37547 = (inp[1]) ? node37559 : node37548;
												assign node37548 = (inp[13]) ? node37552 : node37549;
													assign node37549 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node37552 = (inp[12]) ? node37556 : node37553;
														assign node37553 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node37556 = (inp[15]) ? 4'b0010 : 4'b0011;
												assign node37559 = (inp[10]) ? node37573 : node37560;
													assign node37560 = (inp[15]) ? node37568 : node37561;
														assign node37561 = (inp[13]) ? node37565 : node37562;
															assign node37562 = (inp[12]) ? 4'b0011 : 4'b0110;
															assign node37565 = (inp[12]) ? 4'b0110 : 4'b0011;
														assign node37568 = (inp[13]) ? 4'b0110 : node37569;
															assign node37569 = (inp[12]) ? 4'b0110 : 4'b0011;
													assign node37573 = (inp[15]) ? node37581 : node37574;
														assign node37574 = (inp[12]) ? node37578 : node37575;
															assign node37575 = (inp[13]) ? 4'b0011 : 4'b0110;
															assign node37578 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node37581 = (inp[12]) ? node37585 : node37582;
															assign node37582 = (inp[13]) ? 4'b0110 : 4'b0011;
															assign node37585 = (inp[13]) ? 4'b0010 : 4'b0110;
											assign node37588 = (inp[12]) ? node37602 : node37589;
												assign node37589 = (inp[13]) ? node37595 : node37590;
													assign node37590 = (inp[1]) ? node37592 : 4'b0011;
														assign node37592 = (inp[15]) ? 4'b0010 : 4'b0111;
													assign node37595 = (inp[1]) ? node37599 : node37596;
														assign node37596 = (inp[15]) ? 4'b0111 : 4'b0110;
														assign node37599 = (inp[15]) ? 4'b0110 : 4'b0010;
												assign node37602 = (inp[13]) ? node37608 : node37603;
													assign node37603 = (inp[15]) ? 4'b0111 : node37604;
														assign node37604 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node37608 = (inp[15]) ? 4'b0011 : node37609;
														assign node37609 = (inp[1]) ? 4'b0111 : 4'b0010;
										assign node37613 = (inp[12]) ? node37657 : node37614;
											assign node37614 = (inp[15]) ? node37626 : node37615;
												assign node37615 = (inp[13]) ? node37621 : node37616;
													assign node37616 = (inp[1]) ? 4'b0011 : node37617;
														assign node37617 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node37621 = (inp[1]) ? node37623 : 4'b0111;
														assign node37623 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node37626 = (inp[13]) ? node37642 : node37627;
													assign node37627 = (inp[10]) ? node37635 : node37628;
														assign node37628 = (inp[1]) ? node37632 : node37629;
															assign node37629 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node37632 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node37635 = (inp[1]) ? node37639 : node37636;
															assign node37636 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node37639 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node37642 = (inp[11]) ? node37648 : node37643;
														assign node37643 = (inp[0]) ? node37645 : 4'b0010;
															assign node37645 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node37648 = (inp[10]) ? 4'b0011 : node37649;
															assign node37649 = (inp[1]) ? node37653 : node37650;
																assign node37650 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node37653 = (inp[0]) ? 4'b0011 : 4'b0010;
											assign node37657 = (inp[15]) ? node37669 : node37658;
												assign node37658 = (inp[13]) ? node37664 : node37659;
													assign node37659 = (inp[1]) ? node37661 : 4'b0011;
														assign node37661 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node37664 = (inp[1]) ? 4'b0111 : node37665;
														assign node37665 = (inp[0]) ? 4'b0111 : 4'b0110;
												assign node37669 = (inp[13]) ? 4'b0011 : 4'b0111;
									assign node37672 = (inp[12]) ? node37732 : node37673;
										assign node37673 = (inp[13]) ? node37699 : node37674;
											assign node37674 = (inp[15]) ? node37684 : node37675;
												assign node37675 = (inp[4]) ? node37679 : node37676;
													assign node37676 = (inp[1]) ? 4'b0110 : 4'b0010;
													assign node37679 = (inp[1]) ? 4'b0010 : node37680;
														assign node37680 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node37684 = (inp[4]) ? node37688 : node37685;
													assign node37685 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node37688 = (inp[11]) ? node37694 : node37689;
														assign node37689 = (inp[1]) ? node37691 : 4'b0111;
															assign node37691 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node37694 = (inp[1]) ? 4'b0111 : node37695;
															assign node37695 = (inp[0]) ? 4'b0111 : 4'b0110;
											assign node37699 = (inp[4]) ? node37719 : node37700;
												assign node37700 = (inp[1]) ? node37714 : node37701;
													assign node37701 = (inp[11]) ? node37707 : node37702;
														assign node37702 = (inp[10]) ? node37704 : 4'b0110;
															assign node37704 = (inp[15]) ? 4'b0110 : 4'b0111;
														assign node37707 = (inp[0]) ? node37711 : node37708;
															assign node37708 = (inp[15]) ? 4'b0110 : 4'b0111;
															assign node37711 = (inp[15]) ? 4'b0111 : 4'b0110;
													assign node37714 = (inp[15]) ? node37716 : 4'b0011;
														assign node37716 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node37719 = (inp[15]) ? node37725 : node37720;
													assign node37720 = (inp[0]) ? 4'b0110 : node37721;
														assign node37721 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node37725 = (inp[1]) ? node37729 : node37726;
														assign node37726 = (inp[0]) ? 4'b0011 : 4'b0010;
														assign node37729 = (inp[0]) ? 4'b0010 : 4'b0011;
										assign node37732 = (inp[15]) ? node37748 : node37733;
											assign node37733 = (inp[13]) ? node37741 : node37734;
												assign node37734 = (inp[1]) ? node37738 : node37735;
													assign node37735 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node37738 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node37741 = (inp[1]) ? 4'b0110 : node37742;
													assign node37742 = (inp[4]) ? node37744 : 4'b0011;
														assign node37744 = (inp[0]) ? 4'b0110 : 4'b0111;
											assign node37748 = (inp[13]) ? 4'b0010 : 4'b0110;
					assign node37751 = (inp[6]) ? node39973 : node37752;
						assign node37752 = (inp[12]) ? node38876 : node37753;
							assign node37753 = (inp[15]) ? node38261 : node37754;
								assign node37754 = (inp[4]) ? node38024 : node37755;
									assign node37755 = (inp[10]) ? node37909 : node37756;
										assign node37756 = (inp[11]) ? node37836 : node37757;
											assign node37757 = (inp[2]) ? node37803 : node37758;
												assign node37758 = (inp[13]) ? node37780 : node37759;
													assign node37759 = (inp[5]) ? node37769 : node37760;
														assign node37760 = (inp[1]) ? node37766 : node37761;
															assign node37761 = (inp[0]) ? node37763 : 4'b0101;
																assign node37763 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node37766 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node37769 = (inp[9]) ? node37775 : node37770;
															assign node37770 = (inp[0]) ? 4'b0001 : node37771;
																assign node37771 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node37775 = (inp[1]) ? node37777 : 4'b0000;
																assign node37777 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node37780 = (inp[5]) ? node37792 : node37781;
														assign node37781 = (inp[1]) ? node37789 : node37782;
															assign node37782 = (inp[9]) ? node37786 : node37783;
																assign node37783 = (inp[0]) ? 4'b0000 : 4'b0001;
																assign node37786 = (inp[0]) ? 4'b0001 : 4'b0000;
															assign node37789 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node37792 = (inp[9]) ? node37798 : node37793;
															assign node37793 = (inp[1]) ? 4'b0100 : node37794;
																assign node37794 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node37798 = (inp[1]) ? 4'b0101 : node37799;
																assign node37799 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node37803 = (inp[13]) ? node37821 : node37804;
													assign node37804 = (inp[1]) ? node37812 : node37805;
														assign node37805 = (inp[5]) ? node37807 : 4'b0000;
															assign node37807 = (inp[9]) ? node37809 : 4'b0100;
																assign node37809 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node37812 = (inp[9]) ? node37816 : node37813;
															assign node37813 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node37816 = (inp[0]) ? 4'b0101 : node37817;
																assign node37817 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node37821 = (inp[1]) ? node37827 : node37822;
														assign node37822 = (inp[5]) ? 4'b0001 : node37823;
															assign node37823 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node37827 = (inp[9]) ? node37831 : node37828;
															assign node37828 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node37831 = (inp[0]) ? 4'b0000 : node37832;
																assign node37832 = (inp[5]) ? 4'b0000 : 4'b0001;
											assign node37836 = (inp[5]) ? node37872 : node37837;
												assign node37837 = (inp[9]) ? node37853 : node37838;
													assign node37838 = (inp[2]) ? node37846 : node37839;
														assign node37839 = (inp[13]) ? node37843 : node37840;
															assign node37840 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node37843 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node37846 = (inp[13]) ? node37850 : node37847;
															assign node37847 = (inp[1]) ? 4'b0100 : 4'b0000;
															assign node37850 = (inp[1]) ? 4'b0001 : 4'b0100;
													assign node37853 = (inp[2]) ? node37863 : node37854;
														assign node37854 = (inp[13]) ? node37860 : node37855;
															assign node37855 = (inp[1]) ? node37857 : 4'b0100;
																assign node37857 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node37860 = (inp[1]) ? 4'b0101 : 4'b0001;
														assign node37863 = (inp[13]) ? node37867 : node37864;
															assign node37864 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node37867 = (inp[1]) ? 4'b0000 : node37868;
																assign node37868 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node37872 = (inp[9]) ? node37890 : node37873;
													assign node37873 = (inp[13]) ? node37881 : node37874;
														assign node37874 = (inp[2]) ? node37878 : node37875;
															assign node37875 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node37878 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node37881 = (inp[2]) ? node37885 : node37882;
															assign node37882 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node37885 = (inp[0]) ? 4'b0000 : node37886;
																assign node37886 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node37890 = (inp[13]) ? node37902 : node37891;
														assign node37891 = (inp[2]) ? node37897 : node37892;
															assign node37892 = (inp[0]) ? node37894 : 4'b0000;
																assign node37894 = (inp[1]) ? 4'b0000 : 4'b0001;
															assign node37897 = (inp[0]) ? 4'b0100 : node37898;
																assign node37898 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node37902 = (inp[2]) ? 4'b0001 : node37903;
															assign node37903 = (inp[1]) ? node37905 : 4'b0100;
																assign node37905 = (inp[0]) ? 4'b0100 : 4'b0101;
										assign node37909 = (inp[2]) ? node37963 : node37910;
											assign node37910 = (inp[13]) ? node37934 : node37911;
												assign node37911 = (inp[5]) ? node37919 : node37912;
													assign node37912 = (inp[1]) ? node37914 : 4'b0100;
														assign node37914 = (inp[0]) ? node37916 : 4'b0000;
															assign node37916 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node37919 = (inp[9]) ? node37925 : node37920;
														assign node37920 = (inp[0]) ? node37922 : 4'b0000;
															assign node37922 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node37925 = (inp[1]) ? node37929 : node37926;
															assign node37926 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node37929 = (inp[11]) ? 4'b0001 : node37930;
																assign node37930 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node37934 = (inp[5]) ? node37948 : node37935;
													assign node37935 = (inp[1]) ? node37945 : node37936;
														assign node37936 = (inp[9]) ? node37942 : node37937;
															assign node37937 = (inp[0]) ? 4'b0001 : node37938;
																assign node37938 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node37942 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node37945 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node37948 = (inp[1]) ? node37958 : node37949;
														assign node37949 = (inp[9]) ? node37955 : node37950;
															assign node37950 = (inp[0]) ? 4'b0100 : node37951;
																assign node37951 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node37955 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node37958 = (inp[0]) ? node37960 : 4'b0101;
															assign node37960 = (inp[9]) ? 4'b0101 : 4'b0100;
											assign node37963 = (inp[13]) ? node37995 : node37964;
												assign node37964 = (inp[1]) ? node37978 : node37965;
													assign node37965 = (inp[5]) ? node37973 : node37966;
														assign node37966 = (inp[9]) ? node37968 : 4'b0001;
															assign node37968 = (inp[0]) ? 4'b0000 : node37969;
																assign node37969 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node37973 = (inp[9]) ? node37975 : 4'b0100;
															assign node37975 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node37978 = (inp[9]) ? node37990 : node37979;
														assign node37979 = (inp[5]) ? node37985 : node37980;
															assign node37980 = (inp[11]) ? 4'b0101 : node37981;
																assign node37981 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node37985 = (inp[0]) ? node37987 : 4'b0101;
																assign node37987 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node37990 = (inp[5]) ? node37992 : 4'b0100;
															assign node37992 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node37995 = (inp[5]) ? node38007 : node37996;
													assign node37996 = (inp[1]) ? node38004 : node37997;
														assign node37997 = (inp[9]) ? node37999 : 4'b0100;
															assign node37999 = (inp[11]) ? node38001 : 4'b0101;
																assign node38001 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node38004 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node38007 = (inp[9]) ? node38019 : node38008;
														assign node38008 = (inp[0]) ? node38014 : node38009;
															assign node38009 = (inp[1]) ? 4'b0000 : node38010;
																assign node38010 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node38014 = (inp[1]) ? node38016 : 4'b0001;
																assign node38016 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node38019 = (inp[0]) ? 4'b0000 : node38020;
															assign node38020 = (inp[1]) ? 4'b0001 : 4'b0000;
									assign node38024 = (inp[2]) ? node38148 : node38025;
										assign node38025 = (inp[13]) ? node38089 : node38026;
											assign node38026 = (inp[1]) ? node38060 : node38027;
												assign node38027 = (inp[5]) ? node38045 : node38028;
													assign node38028 = (inp[10]) ? node38034 : node38029;
														assign node38029 = (inp[0]) ? node38031 : 4'b0110;
															assign node38031 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node38034 = (inp[9]) ? node38040 : node38035;
															assign node38035 = (inp[11]) ? 4'b0110 : node38036;
																assign node38036 = (inp[0]) ? 4'b0110 : 4'b0111;
															assign node38040 = (inp[11]) ? 4'b0111 : node38041;
																assign node38041 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node38045 = (inp[9]) ? node38053 : node38046;
														assign node38046 = (inp[10]) ? node38050 : node38047;
															assign node38047 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node38050 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node38053 = (inp[10]) ? node38055 : 4'b0010;
															assign node38055 = (inp[0]) ? 4'b0011 : node38056;
																assign node38056 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node38060 = (inp[10]) ? node38078 : node38061;
													assign node38061 = (inp[5]) ? node38071 : node38062;
														assign node38062 = (inp[9]) ? node38068 : node38063;
															assign node38063 = (inp[0]) ? node38065 : 4'b0010;
																assign node38065 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node38068 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node38071 = (inp[0]) ? node38073 : 4'b0011;
															assign node38073 = (inp[9]) ? node38075 : 4'b0011;
																assign node38075 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node38078 = (inp[9]) ? node38084 : node38079;
														assign node38079 = (inp[11]) ? node38081 : 4'b0011;
															assign node38081 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node38084 = (inp[0]) ? node38086 : 4'b0010;
															assign node38086 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node38089 = (inp[1]) ? node38125 : node38090;
												assign node38090 = (inp[5]) ? node38108 : node38091;
													assign node38091 = (inp[10]) ? node38097 : node38092;
														assign node38092 = (inp[9]) ? node38094 : 4'b0010;
															assign node38094 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node38097 = (inp[9]) ? node38103 : node38098;
															assign node38098 = (inp[0]) ? 4'b0011 : node38099;
																assign node38099 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node38103 = (inp[11]) ? 4'b0010 : node38104;
																assign node38104 = (inp[0]) ? 4'b0010 : 4'b0011;
													assign node38108 = (inp[9]) ? node38120 : node38109;
														assign node38109 = (inp[10]) ? node38115 : node38110;
															assign node38110 = (inp[11]) ? node38112 : 4'b0110;
																assign node38112 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node38115 = (inp[0]) ? node38117 : 4'b0111;
																assign node38117 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node38120 = (inp[10]) ? node38122 : 4'b0111;
															assign node38122 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node38125 = (inp[10]) ? node38137 : node38126;
													assign node38126 = (inp[9]) ? node38132 : node38127;
														assign node38127 = (inp[0]) ? 4'b0110 : node38128;
															assign node38128 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node38132 = (inp[11]) ? 4'b0111 : node38133;
															assign node38133 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node38137 = (inp[9]) ? node38143 : node38138;
														assign node38138 = (inp[11]) ? 4'b0111 : node38139;
															assign node38139 = (inp[0]) ? 4'b0111 : 4'b0110;
														assign node38143 = (inp[11]) ? 4'b0110 : node38144;
															assign node38144 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node38148 = (inp[13]) ? node38208 : node38149;
											assign node38149 = (inp[1]) ? node38187 : node38150;
												assign node38150 = (inp[5]) ? node38172 : node38151;
													assign node38151 = (inp[10]) ? node38161 : node38152;
														assign node38152 = (inp[11]) ? 4'b0010 : node38153;
															assign node38153 = (inp[0]) ? node38157 : node38154;
																assign node38154 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node38157 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node38161 = (inp[9]) ? node38167 : node38162;
															assign node38162 = (inp[11]) ? 4'b0010 : node38163;
																assign node38163 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node38167 = (inp[0]) ? 4'b0011 : node38168;
																assign node38168 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node38172 = (inp[9]) ? node38182 : node38173;
														assign node38173 = (inp[11]) ? node38177 : node38174;
															assign node38174 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node38177 = (inp[10]) ? 4'b0111 : node38178;
																assign node38178 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node38182 = (inp[11]) ? 4'b0110 : node38183;
															assign node38183 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node38187 = (inp[10]) ? node38199 : node38188;
													assign node38188 = (inp[9]) ? node38194 : node38189;
														assign node38189 = (inp[0]) ? 4'b0111 : node38190;
															assign node38190 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node38194 = (inp[0]) ? 4'b0110 : node38195;
															assign node38195 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node38199 = (inp[9]) ? node38205 : node38200;
														assign node38200 = (inp[11]) ? 4'b0110 : node38201;
															assign node38201 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node38205 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node38208 = (inp[1]) ? node38240 : node38209;
												assign node38209 = (inp[5]) ? node38225 : node38210;
													assign node38210 = (inp[10]) ? node38216 : node38211;
														assign node38211 = (inp[0]) ? node38213 : 4'b0111;
															assign node38213 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node38216 = (inp[9]) ? node38220 : node38217;
															assign node38217 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node38220 = (inp[0]) ? node38222 : 4'b0110;
																assign node38222 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node38225 = (inp[10]) ? node38233 : node38226;
														assign node38226 = (inp[0]) ? node38230 : node38227;
															assign node38227 = (inp[9]) ? 4'b0011 : 4'b0010;
															assign node38230 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node38233 = (inp[9]) ? 4'b0010 : node38234;
															assign node38234 = (inp[11]) ? node38236 : 4'b0011;
																assign node38236 = (inp[0]) ? 4'b0010 : 4'b0011;
												assign node38240 = (inp[10]) ? node38250 : node38241;
													assign node38241 = (inp[9]) ? node38247 : node38242;
														assign node38242 = (inp[0]) ? 4'b0010 : node38243;
															assign node38243 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node38247 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node38250 = (inp[9]) ? node38256 : node38251;
														assign node38251 = (inp[0]) ? 4'b0011 : node38252;
															assign node38252 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node38256 = (inp[0]) ? 4'b0010 : node38257;
															assign node38257 = (inp[11]) ? 4'b0010 : 4'b0011;
								assign node38261 = (inp[2]) ? node38565 : node38262;
									assign node38262 = (inp[1]) ? node38418 : node38263;
										assign node38263 = (inp[11]) ? node38335 : node38264;
											assign node38264 = (inp[5]) ? node38300 : node38265;
												assign node38265 = (inp[4]) ? node38281 : node38266;
													assign node38266 = (inp[13]) ? node38274 : node38267;
														assign node38267 = (inp[9]) ? node38271 : node38268;
															assign node38268 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node38271 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node38274 = (inp[0]) ? node38276 : 4'b0110;
															assign node38276 = (inp[10]) ? 4'b0110 : node38277;
																assign node38277 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node38281 = (inp[13]) ? node38293 : node38282;
														assign node38282 = (inp[0]) ? node38288 : node38283;
															assign node38283 = (inp[9]) ? node38285 : 4'b0111;
																assign node38285 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node38288 = (inp[10]) ? 4'b0110 : node38289;
																assign node38289 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node38293 = (inp[9]) ? node38297 : node38294;
															assign node38294 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node38297 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node38300 = (inp[9]) ? node38318 : node38301;
													assign node38301 = (inp[10]) ? node38309 : node38302;
														assign node38302 = (inp[4]) ? node38306 : node38303;
															assign node38303 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node38306 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node38309 = (inp[4]) ? node38313 : node38310;
															assign node38310 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node38313 = (inp[13]) ? node38315 : 4'b0011;
																assign node38315 = (inp[0]) ? 4'b0110 : 4'b0111;
													assign node38318 = (inp[10]) ? node38328 : node38319;
														assign node38319 = (inp[4]) ? node38323 : node38320;
															assign node38320 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node38323 = (inp[13]) ? node38325 : 4'b0011;
																assign node38325 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node38328 = (inp[4]) ? node38332 : node38329;
															assign node38329 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node38332 = (inp[13]) ? 4'b0110 : 4'b0010;
											assign node38335 = (inp[4]) ? node38375 : node38336;
												assign node38336 = (inp[10]) ? node38362 : node38337;
													assign node38337 = (inp[0]) ? node38351 : node38338;
														assign node38338 = (inp[9]) ? node38346 : node38339;
															assign node38339 = (inp[13]) ? node38343 : node38340;
																assign node38340 = (inp[5]) ? 4'b0111 : 4'b0010;
																assign node38343 = (inp[5]) ? 4'b0011 : 4'b0111;
															assign node38346 = (inp[5]) ? node38348 : 4'b0011;
																assign node38348 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node38351 = (inp[5]) ? node38357 : node38352;
															assign node38352 = (inp[9]) ? 4'b0110 : node38353;
																assign node38353 = (inp[13]) ? 4'b0111 : 4'b0011;
															assign node38357 = (inp[9]) ? node38359 : 4'b0110;
																assign node38359 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node38362 = (inp[9]) ? node38370 : node38363;
														assign node38363 = (inp[0]) ? 4'b0111 : node38364;
															assign node38364 = (inp[5]) ? 4'b0110 : node38365;
																assign node38365 = (inp[13]) ? 4'b0110 : 4'b0011;
														assign node38370 = (inp[5]) ? node38372 : 4'b0111;
															assign node38372 = (inp[13]) ? 4'b0011 : 4'b0111;
												assign node38375 = (inp[13]) ? node38403 : node38376;
													assign node38376 = (inp[5]) ? node38388 : node38377;
														assign node38377 = (inp[0]) ? node38383 : node38378;
															assign node38378 = (inp[10]) ? node38380 : 4'b0110;
																assign node38380 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node38383 = (inp[10]) ? node38385 : 4'b0111;
																assign node38385 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node38388 = (inp[10]) ? node38396 : node38389;
															assign node38389 = (inp[0]) ? node38393 : node38390;
																assign node38390 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node38393 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node38396 = (inp[9]) ? node38400 : node38397;
																assign node38397 = (inp[0]) ? 4'b0010 : 4'b0011;
																assign node38400 = (inp[0]) ? 4'b0011 : 4'b0010;
													assign node38403 = (inp[5]) ? node38411 : node38404;
														assign node38404 = (inp[10]) ? node38406 : 4'b0010;
															assign node38406 = (inp[9]) ? 4'b0011 : node38407;
																assign node38407 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node38411 = (inp[9]) ? node38415 : node38412;
															assign node38412 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node38415 = (inp[10]) ? 4'b0111 : 4'b0110;
										assign node38418 = (inp[0]) ? node38496 : node38419;
											assign node38419 = (inp[5]) ? node38465 : node38420;
												assign node38420 = (inp[4]) ? node38446 : node38421;
													assign node38421 = (inp[13]) ? node38437 : node38422;
														assign node38422 = (inp[10]) ? node38430 : node38423;
															assign node38423 = (inp[9]) ? node38427 : node38424;
																assign node38424 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node38427 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node38430 = (inp[11]) ? node38434 : node38431;
																assign node38431 = (inp[9]) ? 4'b0111 : 4'b0110;
																assign node38434 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node38437 = (inp[11]) ? 4'b0011 : node38438;
															assign node38438 = (inp[9]) ? node38442 : node38439;
																assign node38439 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node38442 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node38446 = (inp[13]) ? node38454 : node38447;
														assign node38447 = (inp[9]) ? node38451 : node38448;
															assign node38448 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node38451 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node38454 = (inp[9]) ? node38460 : node38455;
															assign node38455 = (inp[10]) ? node38457 : 4'b0110;
																assign node38457 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node38460 = (inp[10]) ? node38462 : 4'b0111;
																assign node38462 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node38465 = (inp[10]) ? node38479 : node38466;
													assign node38466 = (inp[9]) ? node38474 : node38467;
														assign node38467 = (inp[4]) ? node38471 : node38468;
															assign node38468 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node38471 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node38474 = (inp[4]) ? node38476 : 4'b0111;
															assign node38476 = (inp[13]) ? 4'b0110 : 4'b0010;
													assign node38479 = (inp[9]) ? node38487 : node38480;
														assign node38480 = (inp[4]) ? node38484 : node38481;
															assign node38481 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node38484 = (inp[13]) ? 4'b0111 : 4'b0010;
														assign node38487 = (inp[4]) ? node38491 : node38488;
															assign node38488 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node38491 = (inp[13]) ? node38493 : 4'b0011;
																assign node38493 = (inp[11]) ? 4'b0110 : 4'b0111;
											assign node38496 = (inp[9]) ? node38528 : node38497;
												assign node38497 = (inp[10]) ? node38517 : node38498;
													assign node38498 = (inp[5]) ? node38506 : node38499;
														assign node38499 = (inp[13]) ? node38503 : node38500;
															assign node38500 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node38503 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node38506 = (inp[4]) ? node38512 : node38507;
															assign node38507 = (inp[13]) ? node38509 : 4'b0111;
																assign node38509 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node38512 = (inp[13]) ? 4'b0110 : node38513;
																assign node38513 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node38517 = (inp[13]) ? node38525 : node38518;
														assign node38518 = (inp[4]) ? node38522 : node38519;
															assign node38519 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node38522 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node38525 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node38528 = (inp[10]) ? node38542 : node38529;
													assign node38529 = (inp[13]) ? node38537 : node38530;
														assign node38530 = (inp[4]) ? node38534 : node38531;
															assign node38531 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node38534 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node38537 = (inp[4]) ? 4'b0111 : node38538;
															assign node38538 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node38542 = (inp[5]) ? node38552 : node38543;
														assign node38543 = (inp[13]) ? node38549 : node38544;
															assign node38544 = (inp[4]) ? node38546 : 4'b0110;
																assign node38546 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node38549 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node38552 = (inp[11]) ? node38560 : node38553;
															assign node38553 = (inp[13]) ? node38557 : node38554;
																assign node38554 = (inp[4]) ? 4'b0011 : 4'b0110;
																assign node38557 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node38560 = (inp[4]) ? 4'b0010 : node38561;
																assign node38561 = (inp[13]) ? 4'b0011 : 4'b0111;
									assign node38565 = (inp[0]) ? node38719 : node38566;
										assign node38566 = (inp[10]) ? node38642 : node38567;
											assign node38567 = (inp[11]) ? node38605 : node38568;
												assign node38568 = (inp[9]) ? node38582 : node38569;
													assign node38569 = (inp[4]) ? node38579 : node38570;
														assign node38570 = (inp[13]) ? node38574 : node38571;
															assign node38571 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node38574 = (inp[1]) ? 4'b0111 : node38575;
																assign node38575 = (inp[5]) ? 4'b0110 : 4'b0011;
														assign node38579 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node38582 = (inp[1]) ? node38596 : node38583;
														assign node38583 = (inp[4]) ? node38589 : node38584;
															assign node38584 = (inp[5]) ? 4'b0011 : node38585;
																assign node38585 = (inp[13]) ? 4'b0010 : 4'b0110;
															assign node38589 = (inp[13]) ? node38593 : node38590;
																assign node38590 = (inp[5]) ? 4'b0111 : 4'b0011;
																assign node38593 = (inp[5]) ? 4'b0011 : 4'b0111;
														assign node38596 = (inp[4]) ? node38602 : node38597;
															assign node38597 = (inp[13]) ? 4'b0110 : node38598;
																assign node38598 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node38602 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node38605 = (inp[9]) ? node38627 : node38606;
													assign node38606 = (inp[13]) ? node38616 : node38607;
														assign node38607 = (inp[4]) ? node38613 : node38608;
															assign node38608 = (inp[1]) ? 4'b0011 : node38609;
																assign node38609 = (inp[5]) ? 4'b0010 : 4'b0110;
															assign node38613 = (inp[1]) ? 4'b0110 : 4'b0010;
														assign node38616 = (inp[4]) ? node38624 : node38617;
															assign node38617 = (inp[5]) ? node38621 : node38618;
																assign node38618 = (inp[1]) ? 4'b0111 : 4'b0010;
																assign node38621 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node38624 = (inp[1]) ? 4'b0010 : 4'b0111;
													assign node38627 = (inp[1]) ? node38637 : node38628;
														assign node38628 = (inp[4]) ? node38630 : 4'b0011;
															assign node38630 = (inp[5]) ? node38634 : node38631;
																assign node38631 = (inp[13]) ? 4'b0110 : 4'b0011;
																assign node38634 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node38637 = (inp[4]) ? node38639 : 4'b0110;
															assign node38639 = (inp[13]) ? 4'b0011 : 4'b0111;
											assign node38642 = (inp[1]) ? node38684 : node38643;
												assign node38643 = (inp[9]) ? node38663 : node38644;
													assign node38644 = (inp[5]) ? node38656 : node38645;
														assign node38645 = (inp[13]) ? node38651 : node38646;
															assign node38646 = (inp[4]) ? 4'b0011 : node38647;
																assign node38647 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node38651 = (inp[4]) ? 4'b0110 : node38652;
																assign node38652 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node38656 = (inp[11]) ? node38658 : 4'b0111;
															assign node38658 = (inp[4]) ? 4'b0110 : node38659;
																assign node38659 = (inp[13]) ? 4'b0110 : 4'b0011;
													assign node38663 = (inp[11]) ? node38671 : node38664;
														assign node38664 = (inp[5]) ? 4'b0010 : node38665;
															assign node38665 = (inp[4]) ? node38667 : 4'b0111;
																assign node38667 = (inp[13]) ? 4'b0110 : 4'b0010;
														assign node38671 = (inp[13]) ? node38677 : node38672;
															assign node38672 = (inp[4]) ? node38674 : 4'b0010;
																assign node38674 = (inp[5]) ? 4'b0111 : 4'b0010;
															assign node38677 = (inp[4]) ? node38681 : node38678;
																assign node38678 = (inp[5]) ? 4'b0111 : 4'b0010;
																assign node38681 = (inp[5]) ? 4'b0011 : 4'b0111;
												assign node38684 = (inp[9]) ? node38700 : node38685;
													assign node38685 = (inp[11]) ? node38695 : node38686;
														assign node38686 = (inp[4]) ? node38692 : node38687;
															assign node38687 = (inp[13]) ? 4'b0110 : node38688;
																assign node38688 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node38692 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node38695 = (inp[4]) ? node38697 : 4'b0010;
															assign node38697 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node38700 = (inp[11]) ? node38710 : node38701;
														assign node38701 = (inp[5]) ? node38705 : node38702;
															assign node38702 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node38705 = (inp[4]) ? node38707 : 4'b0111;
																assign node38707 = (inp[13]) ? 4'b0011 : 4'b0111;
														assign node38710 = (inp[4]) ? node38716 : node38711;
															assign node38711 = (inp[13]) ? node38713 : 4'b0011;
																assign node38713 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node38716 = (inp[13]) ? 4'b0010 : 4'b0110;
										assign node38719 = (inp[1]) ? node38793 : node38720;
											assign node38720 = (inp[5]) ? node38758 : node38721;
												assign node38721 = (inp[13]) ? node38743 : node38722;
													assign node38722 = (inp[4]) ? node38730 : node38723;
														assign node38723 = (inp[11]) ? node38725 : 4'b0110;
															assign node38725 = (inp[9]) ? 4'b0111 : node38726;
																assign node38726 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node38730 = (inp[9]) ? node38738 : node38731;
															assign node38731 = (inp[10]) ? node38735 : node38732;
																assign node38732 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node38735 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node38738 = (inp[10]) ? 4'b0010 : node38739;
																assign node38739 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node38743 = (inp[4]) ? node38751 : node38744;
														assign node38744 = (inp[9]) ? node38748 : node38745;
															assign node38745 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node38748 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node38751 = (inp[10]) ? node38755 : node38752;
															assign node38752 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node38755 = (inp[9]) ? 4'b0111 : 4'b0110;
												assign node38758 = (inp[13]) ? node38778 : node38759;
													assign node38759 = (inp[4]) ? node38773 : node38760;
														assign node38760 = (inp[9]) ? node38768 : node38761;
															assign node38761 = (inp[10]) ? node38765 : node38762;
																assign node38762 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node38765 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node38768 = (inp[11]) ? node38770 : 4'b0011;
																assign node38770 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node38773 = (inp[10]) ? node38775 : 4'b0111;
															assign node38775 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node38778 = (inp[4]) ? node38786 : node38779;
														assign node38779 = (inp[10]) ? node38783 : node38780;
															assign node38780 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node38783 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node38786 = (inp[10]) ? node38790 : node38787;
															assign node38787 = (inp[9]) ? 4'b0010 : 4'b0011;
															assign node38790 = (inp[9]) ? 4'b0011 : 4'b0010;
											assign node38793 = (inp[5]) ? node38833 : node38794;
												assign node38794 = (inp[9]) ? node38812 : node38795;
													assign node38795 = (inp[4]) ? node38807 : node38796;
														assign node38796 = (inp[13]) ? node38800 : node38797;
															assign node38797 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node38800 = (inp[11]) ? node38804 : node38801;
																assign node38801 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node38804 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node38807 = (inp[13]) ? 4'b0011 : node38808;
															assign node38808 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node38812 = (inp[11]) ? node38828 : node38813;
														assign node38813 = (inp[10]) ? node38821 : node38814;
															assign node38814 = (inp[4]) ? node38818 : node38815;
																assign node38815 = (inp[13]) ? 4'b0110 : 4'b0010;
																assign node38818 = (inp[13]) ? 4'b0011 : 4'b0111;
															assign node38821 = (inp[4]) ? node38825 : node38822;
																assign node38822 = (inp[13]) ? 4'b0111 : 4'b0011;
																assign node38825 = (inp[13]) ? 4'b0010 : 4'b0110;
														assign node38828 = (inp[10]) ? node38830 : 4'b0011;
															assign node38830 = (inp[4]) ? 4'b0110 : 4'b0011;
												assign node38833 = (inp[4]) ? node38855 : node38834;
													assign node38834 = (inp[13]) ? node38848 : node38835;
														assign node38835 = (inp[9]) ? node38843 : node38836;
															assign node38836 = (inp[10]) ? node38840 : node38837;
																assign node38837 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node38840 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node38843 = (inp[10]) ? node38845 : 4'b0011;
																assign node38845 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node38848 = (inp[10]) ? node38852 : node38849;
															assign node38849 = (inp[9]) ? 4'b0111 : 4'b0110;
															assign node38852 = (inp[9]) ? 4'b0110 : 4'b0111;
													assign node38855 = (inp[13]) ? node38869 : node38856;
														assign node38856 = (inp[11]) ? node38864 : node38857;
															assign node38857 = (inp[9]) ? node38861 : node38858;
																assign node38858 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node38861 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node38864 = (inp[10]) ? node38866 : 4'b0110;
																assign node38866 = (inp[9]) ? 4'b0110 : 4'b0111;
														assign node38869 = (inp[9]) ? node38873 : node38870;
															assign node38870 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node38873 = (inp[10]) ? 4'b0010 : 4'b0011;
							assign node38876 = (inp[4]) ? node39398 : node38877;
								assign node38877 = (inp[15]) ? node39167 : node38878;
									assign node38878 = (inp[2]) ? node39026 : node38879;
										assign node38879 = (inp[13]) ? node38951 : node38880;
											assign node38880 = (inp[1]) ? node38916 : node38881;
												assign node38881 = (inp[9]) ? node38899 : node38882;
													assign node38882 = (inp[5]) ? node38890 : node38883;
														assign node38883 = (inp[10]) ? node38885 : 4'b0110;
															assign node38885 = (inp[11]) ? node38887 : 4'b0111;
																assign node38887 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node38890 = (inp[0]) ? 4'b0111 : node38891;
															assign node38891 = (inp[10]) ? node38895 : node38892;
																assign node38892 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node38895 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node38899 = (inp[5]) ? node38911 : node38900;
														assign node38900 = (inp[10]) ? node38906 : node38901;
															assign node38901 = (inp[0]) ? node38903 : 4'b0111;
																assign node38903 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node38906 = (inp[0]) ? node38908 : 4'b0110;
																assign node38908 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node38911 = (inp[10]) ? node38913 : 4'b0110;
															assign node38913 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node38916 = (inp[5]) ? node38932 : node38917;
													assign node38917 = (inp[11]) ? node38925 : node38918;
														assign node38918 = (inp[10]) ? node38920 : 4'b0111;
															assign node38920 = (inp[0]) ? node38922 : 4'b0110;
																assign node38922 = (inp[9]) ? 4'b0111 : 4'b0110;
														assign node38925 = (inp[10]) ? node38929 : node38926;
															assign node38926 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node38929 = (inp[9]) ? 4'b0111 : 4'b0110;
													assign node38932 = (inp[9]) ? node38942 : node38933;
														assign node38933 = (inp[10]) ? node38937 : node38934;
															assign node38934 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node38937 = (inp[0]) ? node38939 : 4'b0010;
																assign node38939 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node38942 = (inp[0]) ? node38944 : 4'b0011;
															assign node38944 = (inp[11]) ? node38948 : node38945;
																assign node38945 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node38948 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node38951 = (inp[1]) ? node38991 : node38952;
												assign node38952 = (inp[10]) ? node38976 : node38953;
													assign node38953 = (inp[9]) ? node38965 : node38954;
														assign node38954 = (inp[11]) ? node38960 : node38955;
															assign node38955 = (inp[0]) ? node38957 : 4'b0011;
																assign node38957 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node38960 = (inp[5]) ? 4'b0010 : node38961;
																assign node38961 = (inp[0]) ? 4'b0010 : 4'b0011;
														assign node38965 = (inp[0]) ? node38971 : node38966;
															assign node38966 = (inp[5]) ? node38968 : 4'b0010;
																assign node38968 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node38971 = (inp[5]) ? 4'b0011 : node38972;
																assign node38972 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node38976 = (inp[5]) ? node38986 : node38977;
														assign node38977 = (inp[11]) ? node38979 : 4'b0010;
															assign node38979 = (inp[0]) ? node38983 : node38980;
																assign node38980 = (inp[9]) ? 4'b0011 : 4'b0010;
																assign node38983 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node38986 = (inp[9]) ? 4'b0010 : node38987;
															assign node38987 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node38991 = (inp[5]) ? node39007 : node38992;
													assign node38992 = (inp[0]) ? node39000 : node38993;
														assign node38993 = (inp[10]) ? 4'b0010 : node38994;
															assign node38994 = (inp[9]) ? 4'b0010 : node38995;
																assign node38995 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node39000 = (inp[9]) ? node39004 : node39001;
															assign node39001 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node39004 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node39007 = (inp[10]) ? node39019 : node39008;
														assign node39008 = (inp[9]) ? node39014 : node39009;
															assign node39009 = (inp[0]) ? 4'b0111 : node39010;
																assign node39010 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node39014 = (inp[11]) ? 4'b0110 : node39015;
																assign node39015 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node39019 = (inp[11]) ? 4'b0110 : node39020;
															assign node39020 = (inp[9]) ? 4'b0110 : node39021;
																assign node39021 = (inp[0]) ? 4'b0110 : 4'b0111;
										assign node39026 = (inp[13]) ? node39096 : node39027;
											assign node39027 = (inp[5]) ? node39059 : node39028;
												assign node39028 = (inp[10]) ? node39044 : node39029;
													assign node39029 = (inp[11]) ? node39035 : node39030;
														assign node39030 = (inp[9]) ? 4'b0010 : node39031;
															assign node39031 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node39035 = (inp[0]) ? 4'b0011 : node39036;
															assign node39036 = (inp[1]) ? node39040 : node39037;
																assign node39037 = (inp[9]) ? 4'b0010 : 4'b0011;
																assign node39040 = (inp[9]) ? 4'b0011 : 4'b0010;
													assign node39044 = (inp[1]) ? node39048 : node39045;
														assign node39045 = (inp[9]) ? 4'b0011 : 4'b0010;
														assign node39048 = (inp[9]) ? node39054 : node39049;
															assign node39049 = (inp[0]) ? 4'b0011 : node39050;
																assign node39050 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node39054 = (inp[0]) ? 4'b0010 : node39055;
																assign node39055 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node39059 = (inp[1]) ? node39081 : node39060;
													assign node39060 = (inp[0]) ? node39076 : node39061;
														assign node39061 = (inp[9]) ? node39069 : node39062;
															assign node39062 = (inp[11]) ? node39066 : node39063;
																assign node39063 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node39066 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node39069 = (inp[11]) ? node39073 : node39070;
																assign node39070 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node39073 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node39076 = (inp[10]) ? node39078 : 4'b0011;
															assign node39078 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node39081 = (inp[0]) ? node39089 : node39082;
														assign node39082 = (inp[9]) ? node39084 : 4'b0110;
															assign node39084 = (inp[11]) ? node39086 : 4'b0110;
																assign node39086 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node39089 = (inp[10]) ? node39093 : node39090;
															assign node39090 = (inp[9]) ? 4'b0110 : 4'b0111;
															assign node39093 = (inp[9]) ? 4'b0111 : 4'b0110;
											assign node39096 = (inp[1]) ? node39132 : node39097;
												assign node39097 = (inp[5]) ? node39113 : node39098;
													assign node39098 = (inp[11]) ? node39108 : node39099;
														assign node39099 = (inp[0]) ? 4'b0110 : node39100;
															assign node39100 = (inp[9]) ? node39104 : node39101;
																assign node39101 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node39104 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node39108 = (inp[9]) ? node39110 : 4'b0111;
															assign node39110 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node39113 = (inp[9]) ? node39121 : node39114;
														assign node39114 = (inp[10]) ? 4'b0110 : node39115;
															assign node39115 = (inp[11]) ? node39117 : 4'b0111;
																assign node39117 = (inp[0]) ? 4'b0110 : 4'b0111;
														assign node39121 = (inp[10]) ? node39127 : node39122;
															assign node39122 = (inp[11]) ? node39124 : 4'b0110;
																assign node39124 = (inp[0]) ? 4'b0111 : 4'b0110;
															assign node39127 = (inp[11]) ? node39129 : 4'b0111;
																assign node39129 = (inp[0]) ? 4'b0110 : 4'b0111;
												assign node39132 = (inp[5]) ? node39146 : node39133;
													assign node39133 = (inp[9]) ? node39139 : node39134;
														assign node39134 = (inp[0]) ? 4'b0110 : node39135;
															assign node39135 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node39139 = (inp[10]) ? 4'b0111 : node39140;
															assign node39140 = (inp[11]) ? node39142 : 4'b0110;
																assign node39142 = (inp[0]) ? 4'b0111 : 4'b0110;
													assign node39146 = (inp[9]) ? node39156 : node39147;
														assign node39147 = (inp[10]) ? node39151 : node39148;
															assign node39148 = (inp[0]) ? 4'b0010 : 4'b0011;
															assign node39151 = (inp[0]) ? 4'b0011 : node39152;
																assign node39152 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node39156 = (inp[10]) ? node39162 : node39157;
															assign node39157 = (inp[0]) ? 4'b0011 : node39158;
																assign node39158 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node39162 = (inp[11]) ? 4'b0010 : node39163;
																assign node39163 = (inp[0]) ? 4'b0010 : 4'b0011;
									assign node39167 = (inp[10]) ? node39291 : node39168;
										assign node39168 = (inp[9]) ? node39228 : node39169;
											assign node39169 = (inp[0]) ? node39203 : node39170;
												assign node39170 = (inp[5]) ? node39192 : node39171;
													assign node39171 = (inp[2]) ? node39181 : node39172;
														assign node39172 = (inp[11]) ? 4'b0000 : node39173;
															assign node39173 = (inp[1]) ? node39177 : node39174;
																assign node39174 = (inp[13]) ? 4'b0001 : 4'b0101;
																assign node39177 = (inp[13]) ? 4'b0100 : 4'b0001;
														assign node39181 = (inp[11]) ? node39187 : node39182;
															assign node39182 = (inp[1]) ? node39184 : 4'b0000;
																assign node39184 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node39187 = (inp[1]) ? 4'b0101 : node39188;
																assign node39188 = (inp[13]) ? 4'b0101 : 4'b0001;
													assign node39192 = (inp[13]) ? node39196 : node39193;
														assign node39193 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node39196 = (inp[2]) ? node39200 : node39197;
															assign node39197 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node39200 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node39203 = (inp[2]) ? node39219 : node39204;
													assign node39204 = (inp[13]) ? node39212 : node39205;
														assign node39205 = (inp[5]) ? node39209 : node39206;
															assign node39206 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node39209 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node39212 = (inp[5]) ? 4'b0101 : node39213;
															assign node39213 = (inp[1]) ? node39215 : 4'b0000;
																assign node39215 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node39219 = (inp[13]) ? node39225 : node39220;
														assign node39220 = (inp[1]) ? 4'b0100 : node39221;
															assign node39221 = (inp[5]) ? 4'b0100 : 4'b0001;
														assign node39225 = (inp[5]) ? 4'b0000 : 4'b0100;
											assign node39228 = (inp[11]) ? node39262 : node39229;
												assign node39229 = (inp[2]) ? node39245 : node39230;
													assign node39230 = (inp[13]) ? node39236 : node39231;
														assign node39231 = (inp[1]) ? 4'b0001 : node39232;
															assign node39232 = (inp[5]) ? 4'b0001 : 4'b0100;
														assign node39236 = (inp[1]) ? node39240 : node39237;
															assign node39237 = (inp[0]) ? 4'b0100 : 4'b0000;
															assign node39240 = (inp[5]) ? node39242 : 4'b0101;
																assign node39242 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node39245 = (inp[13]) ? node39255 : node39246;
														assign node39246 = (inp[5]) ? node39252 : node39247;
															assign node39247 = (inp[1]) ? 4'b0100 : node39248;
																assign node39248 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node39252 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node39255 = (inp[5]) ? node39259 : node39256;
															assign node39256 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node39259 = (inp[0]) ? 4'b0001 : 4'b0000;
												assign node39262 = (inp[13]) ? node39278 : node39263;
													assign node39263 = (inp[2]) ? node39271 : node39264;
														assign node39264 = (inp[5]) ? node39268 : node39265;
															assign node39265 = (inp[1]) ? 4'b0001 : 4'b0101;
															assign node39268 = (inp[0]) ? 4'b0000 : 4'b0001;
														assign node39271 = (inp[5]) ? 4'b0101 : node39272;
															assign node39272 = (inp[1]) ? node39274 : 4'b0000;
																assign node39274 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node39278 = (inp[2]) ? node39284 : node39279;
														assign node39279 = (inp[1]) ? node39281 : 4'b0001;
															assign node39281 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node39284 = (inp[5]) ? 4'b0001 : node39285;
															assign node39285 = (inp[1]) ? node39287 : 4'b0100;
																assign node39287 = (inp[0]) ? 4'b0001 : 4'b0000;
										assign node39291 = (inp[9]) ? node39341 : node39292;
											assign node39292 = (inp[13]) ? node39324 : node39293;
												assign node39293 = (inp[2]) ? node39309 : node39294;
													assign node39294 = (inp[1]) ? node39302 : node39295;
														assign node39295 = (inp[5]) ? 4'b0001 : node39296;
															assign node39296 = (inp[0]) ? 4'b0101 : node39297;
																assign node39297 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node39302 = (inp[5]) ? 4'b0001 : node39303;
															assign node39303 = (inp[0]) ? 4'b0001 : node39304;
																assign node39304 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node39309 = (inp[5]) ? node39319 : node39310;
														assign node39310 = (inp[1]) ? node39316 : node39311;
															assign node39311 = (inp[0]) ? 4'b0000 : node39312;
																assign node39312 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node39316 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node39319 = (inp[11]) ? 4'b0101 : node39320;
															assign node39320 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node39324 = (inp[2]) ? node39332 : node39325;
													assign node39325 = (inp[11]) ? 4'b0100 : node39326;
														assign node39326 = (inp[5]) ? node39328 : 4'b0001;
															assign node39328 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node39332 = (inp[5]) ? node39338 : node39333;
														assign node39333 = (inp[1]) ? 4'b0000 : node39334;
															assign node39334 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node39338 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node39341 = (inp[2]) ? node39371 : node39342;
												assign node39342 = (inp[13]) ? node39358 : node39343;
													assign node39343 = (inp[1]) ? node39351 : node39344;
														assign node39344 = (inp[5]) ? 4'b0000 : node39345;
															assign node39345 = (inp[11]) ? 4'b0100 : node39346;
																assign node39346 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node39351 = (inp[11]) ? node39353 : 4'b0000;
															assign node39353 = (inp[5]) ? node39355 : 4'b0000;
																assign node39355 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node39358 = (inp[0]) ? node39366 : node39359;
														assign node39359 = (inp[1]) ? 4'b0100 : node39360;
															assign node39360 = (inp[5]) ? node39362 : 4'b0000;
																assign node39362 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node39366 = (inp[5]) ? 4'b0101 : node39367;
															assign node39367 = (inp[1]) ? 4'b0101 : 4'b0000;
												assign node39371 = (inp[11]) ? node39385 : node39372;
													assign node39372 = (inp[1]) ? node39382 : node39373;
														assign node39373 = (inp[13]) ? 4'b0101 : node39374;
															assign node39374 = (inp[5]) ? node39378 : node39375;
																assign node39375 = (inp[0]) ? 4'b0001 : 4'b0000;
																assign node39378 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node39382 = (inp[13]) ? 4'b0001 : 4'b0101;
													assign node39385 = (inp[13]) ? node39391 : node39386;
														assign node39386 = (inp[5]) ? 4'b0100 : node39387;
															assign node39387 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node39391 = (inp[5]) ? 4'b0000 : node39392;
															assign node39392 = (inp[1]) ? node39394 : 4'b0101;
																assign node39394 = (inp[0]) ? 4'b0000 : 4'b0001;
								assign node39398 = (inp[10]) ? node39668 : node39399;
									assign node39399 = (inp[9]) ? node39545 : node39400;
										assign node39400 = (inp[11]) ? node39476 : node39401;
											assign node39401 = (inp[0]) ? node39439 : node39402;
												assign node39402 = (inp[15]) ? node39422 : node39403;
													assign node39403 = (inp[13]) ? node39415 : node39404;
														assign node39404 = (inp[1]) ? node39412 : node39405;
															assign node39405 = (inp[5]) ? node39409 : node39406;
																assign node39406 = (inp[2]) ? 4'b0001 : 4'b0101;
																assign node39409 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node39412 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node39415 = (inp[2]) ? node39417 : 4'b0101;
															assign node39417 = (inp[1]) ? 4'b0001 : node39418;
																assign node39418 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node39422 = (inp[2]) ? node39430 : node39423;
														assign node39423 = (inp[13]) ? 4'b0101 : node39424;
															assign node39424 = (inp[1]) ? 4'b0001 : node39425;
																assign node39425 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node39430 = (inp[1]) ? 4'b0101 : node39431;
															assign node39431 = (inp[13]) ? node39435 : node39432;
																assign node39432 = (inp[5]) ? 4'b0101 : 4'b0001;
																assign node39435 = (inp[5]) ? 4'b0001 : 4'b0101;
												assign node39439 = (inp[5]) ? node39457 : node39440;
													assign node39440 = (inp[1]) ? node39448 : node39441;
														assign node39441 = (inp[2]) ? node39445 : node39442;
															assign node39442 = (inp[13]) ? 4'b0001 : 4'b0101;
															assign node39445 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node39448 = (inp[13]) ? node39454 : node39449;
															assign node39449 = (inp[2]) ? 4'b0101 : node39450;
																assign node39450 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node39454 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node39457 = (inp[15]) ? node39469 : node39458;
														assign node39458 = (inp[2]) ? node39464 : node39459;
															assign node39459 = (inp[1]) ? node39461 : 4'b0101;
																assign node39461 = (inp[13]) ? 4'b0100 : 4'b0000;
															assign node39464 = (inp[13]) ? 4'b0001 : node39465;
																assign node39465 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node39469 = (inp[1]) ? 4'b0001 : node39470;
															assign node39470 = (inp[2]) ? node39472 : 4'b0100;
																assign node39472 = (inp[13]) ? 4'b0000 : 4'b0100;
											assign node39476 = (inp[0]) ? node39512 : node39477;
												assign node39477 = (inp[1]) ? node39501 : node39478;
													assign node39478 = (inp[13]) ? node39492 : node39479;
														assign node39479 = (inp[15]) ? node39485 : node39480;
															assign node39480 = (inp[2]) ? node39482 : 4'b0100;
																assign node39482 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node39485 = (inp[2]) ? node39489 : node39486;
																assign node39486 = (inp[5]) ? 4'b0001 : 4'b0101;
																assign node39489 = (inp[5]) ? 4'b0100 : 4'b0001;
														assign node39492 = (inp[15]) ? 4'b0001 : node39493;
															assign node39493 = (inp[5]) ? node39497 : node39494;
																assign node39494 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node39497 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node39501 = (inp[13]) ? node39509 : node39502;
														assign node39502 = (inp[2]) ? node39506 : node39503;
															assign node39503 = (inp[15]) ? 4'b0001 : 4'b0000;
															assign node39506 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node39509 = (inp[2]) ? 4'b0000 : 4'b0100;
												assign node39512 = (inp[15]) ? node39526 : node39513;
													assign node39513 = (inp[13]) ? node39521 : node39514;
														assign node39514 = (inp[1]) ? 4'b0101 : node39515;
															assign node39515 = (inp[2]) ? node39517 : 4'b0000;
																assign node39517 = (inp[5]) ? 4'b0101 : 4'b0000;
														assign node39521 = (inp[2]) ? node39523 : 4'b0100;
															assign node39523 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node39526 = (inp[13]) ? node39538 : node39527;
														assign node39527 = (inp[2]) ? node39533 : node39528;
															assign node39528 = (inp[5]) ? 4'b0000 : node39529;
																assign node39529 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node39533 = (inp[5]) ? 4'b0100 : node39534;
																assign node39534 = (inp[1]) ? 4'b0100 : 4'b0000;
														assign node39538 = (inp[2]) ? 4'b0000 : node39539;
															assign node39539 = (inp[5]) ? 4'b0100 : node39540;
																assign node39540 = (inp[1]) ? 4'b0100 : 4'b0000;
										assign node39545 = (inp[0]) ? node39611 : node39546;
											assign node39546 = (inp[11]) ? node39582 : node39547;
												assign node39547 = (inp[15]) ? node39567 : node39548;
													assign node39548 = (inp[13]) ? node39558 : node39549;
														assign node39549 = (inp[5]) ? 4'b0101 : node39550;
															assign node39550 = (inp[1]) ? node39554 : node39551;
																assign node39551 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node39554 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node39558 = (inp[5]) ? node39564 : node39559;
															assign node39559 = (inp[2]) ? node39561 : 4'b0001;
																assign node39561 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node39564 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node39567 = (inp[2]) ? node39575 : node39568;
														assign node39568 = (inp[13]) ? node39570 : 4'b0000;
															assign node39570 = (inp[1]) ? 4'b0100 : node39571;
																assign node39571 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node39575 = (inp[13]) ? node39577 : 4'b0100;
															assign node39577 = (inp[1]) ? 4'b0000 : node39578;
																assign node39578 = (inp[5]) ? 4'b0000 : 4'b0100;
												assign node39582 = (inp[2]) ? node39594 : node39583;
													assign node39583 = (inp[13]) ? node39587 : node39584;
														assign node39584 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node39587 = (inp[1]) ? 4'b0101 : node39588;
															assign node39588 = (inp[5]) ? node39590 : 4'b0000;
																assign node39590 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node39594 = (inp[13]) ? node39604 : node39595;
														assign node39595 = (inp[5]) ? node39599 : node39596;
															assign node39596 = (inp[1]) ? 4'b0101 : 4'b0001;
															assign node39599 = (inp[15]) ? 4'b0101 : node39600;
																assign node39600 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node39604 = (inp[1]) ? 4'b0001 : node39605;
															assign node39605 = (inp[5]) ? 4'b0000 : node39606;
																assign node39606 = (inp[15]) ? 4'b0101 : 4'b0100;
											assign node39611 = (inp[13]) ? node39649 : node39612;
												assign node39612 = (inp[2]) ? node39634 : node39613;
													assign node39613 = (inp[1]) ? node39625 : node39614;
														assign node39614 = (inp[5]) ? node39620 : node39615;
															assign node39615 = (inp[11]) ? 4'b0101 : node39616;
																assign node39616 = (inp[15]) ? 4'b0100 : 4'b0101;
															assign node39620 = (inp[11]) ? 4'b0001 : node39621;
																assign node39621 = (inp[15]) ? 4'b0000 : 4'b0001;
														assign node39625 = (inp[5]) ? 4'b0000 : node39626;
															assign node39626 = (inp[11]) ? node39630 : node39627;
																assign node39627 = (inp[15]) ? 4'b0000 : 4'b0001;
																assign node39630 = (inp[15]) ? 4'b0001 : 4'b0000;
													assign node39634 = (inp[1]) ? node39646 : node39635;
														assign node39635 = (inp[5]) ? node39641 : node39636;
															assign node39636 = (inp[11]) ? 4'b0001 : node39637;
																assign node39637 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node39641 = (inp[11]) ? node39643 : 4'b0101;
																assign node39643 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node39646 = (inp[15]) ? 4'b0101 : 4'b0100;
												assign node39649 = (inp[2]) ? node39659 : node39650;
													assign node39650 = (inp[1]) ? 4'b0101 : node39651;
														assign node39651 = (inp[5]) ? node39655 : node39652;
															assign node39652 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node39655 = (inp[15]) ? 4'b0101 : 4'b0100;
													assign node39659 = (inp[1]) ? 4'b0001 : node39660;
														assign node39660 = (inp[5]) ? 4'b0001 : node39661;
															assign node39661 = (inp[11]) ? 4'b0101 : node39662;
																assign node39662 = (inp[15]) ? 4'b0101 : 4'b0100;
									assign node39668 = (inp[9]) ? node39824 : node39669;
										assign node39669 = (inp[11]) ? node39753 : node39670;
											assign node39670 = (inp[0]) ? node39714 : node39671;
												assign node39671 = (inp[15]) ? node39693 : node39672;
													assign node39672 = (inp[13]) ? node39684 : node39673;
														assign node39673 = (inp[1]) ? node39681 : node39674;
															assign node39674 = (inp[5]) ? node39678 : node39675;
																assign node39675 = (inp[2]) ? 4'b0000 : 4'b0100;
																assign node39678 = (inp[2]) ? 4'b0101 : 4'b0000;
															assign node39681 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node39684 = (inp[1]) ? node39690 : node39685;
															assign node39685 = (inp[5]) ? 4'b0100 : node39686;
																assign node39686 = (inp[2]) ? 4'b0100 : 4'b0001;
															assign node39690 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node39693 = (inp[2]) ? node39705 : node39694;
														assign node39694 = (inp[13]) ? node39700 : node39695;
															assign node39695 = (inp[5]) ? 4'b0000 : node39696;
																assign node39696 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node39700 = (inp[1]) ? 4'b0100 : node39701;
																assign node39701 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node39705 = (inp[13]) ? node39709 : node39706;
															assign node39706 = (inp[5]) ? 4'b0100 : 4'b0000;
															assign node39709 = (inp[1]) ? 4'b0000 : node39710;
																assign node39710 = (inp[5]) ? 4'b0000 : 4'b0100;
												assign node39714 = (inp[1]) ? node39742 : node39715;
													assign node39715 = (inp[2]) ? node39729 : node39716;
														assign node39716 = (inp[5]) ? node39722 : node39717;
															assign node39717 = (inp[13]) ? 4'b0000 : node39718;
																assign node39718 = (inp[15]) ? 4'b0100 : 4'b0101;
															assign node39722 = (inp[13]) ? node39726 : node39723;
																assign node39723 = (inp[15]) ? 4'b0000 : 4'b0001;
																assign node39726 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node39729 = (inp[15]) ? node39735 : node39730;
															assign node39730 = (inp[13]) ? node39732 : 4'b0001;
																assign node39732 = (inp[5]) ? 4'b0000 : 4'b0100;
															assign node39735 = (inp[13]) ? node39739 : node39736;
																assign node39736 = (inp[5]) ? 4'b0101 : 4'b0000;
																assign node39739 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node39742 = (inp[13]) ? node39750 : node39743;
														assign node39743 = (inp[2]) ? node39747 : node39744;
															assign node39744 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node39747 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node39750 = (inp[2]) ? 4'b0001 : 4'b0101;
											assign node39753 = (inp[0]) ? node39789 : node39754;
												assign node39754 = (inp[1]) ? node39778 : node39755;
													assign node39755 = (inp[13]) ? node39769 : node39756;
														assign node39756 = (inp[15]) ? node39764 : node39757;
															assign node39757 = (inp[2]) ? node39761 : node39758;
																assign node39758 = (inp[5]) ? 4'b0001 : 4'b0101;
																assign node39761 = (inp[5]) ? 4'b0101 : 4'b0001;
															assign node39764 = (inp[5]) ? 4'b0000 : node39765;
																assign node39765 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node39769 = (inp[15]) ? 4'b0101 : node39770;
															assign node39770 = (inp[2]) ? node39774 : node39771;
																assign node39771 = (inp[5]) ? 4'b0100 : 4'b0000;
																assign node39774 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node39778 = (inp[13]) ? node39786 : node39779;
														assign node39779 = (inp[2]) ? node39783 : node39780;
															assign node39780 = (inp[15]) ? 4'b0000 : 4'b0001;
															assign node39783 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node39786 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node39789 = (inp[15]) ? node39807 : node39790;
													assign node39790 = (inp[13]) ? node39798 : node39791;
														assign node39791 = (inp[2]) ? 4'b0100 : node39792;
															assign node39792 = (inp[1]) ? 4'b0000 : node39793;
																assign node39793 = (inp[5]) ? 4'b0001 : 4'b0101;
														assign node39798 = (inp[2]) ? node39804 : node39799;
															assign node39799 = (inp[1]) ? 4'b0101 : node39800;
																assign node39800 = (inp[5]) ? 4'b0101 : 4'b0000;
															assign node39804 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node39807 = (inp[1]) ? node39819 : node39808;
														assign node39808 = (inp[5]) ? node39814 : node39809;
															assign node39809 = (inp[13]) ? 4'b0001 : node39810;
																assign node39810 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node39814 = (inp[13]) ? 4'b0101 : node39815;
																assign node39815 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node39819 = (inp[13]) ? 4'b0001 : node39820;
															assign node39820 = (inp[2]) ? 4'b0101 : 4'b0001;
										assign node39824 = (inp[0]) ? node39894 : node39825;
											assign node39825 = (inp[11]) ? node39859 : node39826;
												assign node39826 = (inp[15]) ? node39848 : node39827;
													assign node39827 = (inp[13]) ? node39837 : node39828;
														assign node39828 = (inp[1]) ? node39834 : node39829;
															assign node39829 = (inp[5]) ? 4'b0100 : node39830;
																assign node39830 = (inp[2]) ? 4'b0001 : 4'b0101;
															assign node39834 = (inp[2]) ? 4'b0100 : 4'b0000;
														assign node39837 = (inp[2]) ? node39843 : node39838;
															assign node39838 = (inp[1]) ? 4'b0101 : node39839;
																assign node39839 = (inp[5]) ? 4'b0101 : 4'b0000;
															assign node39843 = (inp[1]) ? 4'b0001 : node39844;
																assign node39844 = (inp[5]) ? 4'b0001 : 4'b0101;
													assign node39848 = (inp[1]) ? node39850 : 4'b0001;
														assign node39850 = (inp[5]) ? node39852 : 4'b0001;
															assign node39852 = (inp[13]) ? node39856 : node39853;
																assign node39853 = (inp[2]) ? 4'b0101 : 4'b0001;
																assign node39856 = (inp[2]) ? 4'b0001 : 4'b0101;
												assign node39859 = (inp[1]) ? node39883 : node39860;
													assign node39860 = (inp[2]) ? node39872 : node39861;
														assign node39861 = (inp[13]) ? node39867 : node39862;
															assign node39862 = (inp[5]) ? 4'b0001 : node39863;
																assign node39863 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node39867 = (inp[5]) ? node39869 : 4'b0001;
																assign node39869 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node39872 = (inp[5]) ? node39880 : node39873;
															assign node39873 = (inp[13]) ? node39877 : node39874;
																assign node39874 = (inp[15]) ? 4'b0001 : 4'b0000;
																assign node39877 = (inp[15]) ? 4'b0100 : 4'b0101;
															assign node39880 = (inp[13]) ? 4'b0000 : 4'b0100;
													assign node39883 = (inp[13]) ? node39891 : node39884;
														assign node39884 = (inp[2]) ? node39888 : node39885;
															assign node39885 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node39888 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node39891 = (inp[2]) ? 4'b0000 : 4'b0100;
											assign node39894 = (inp[15]) ? node39936 : node39895;
												assign node39895 = (inp[11]) ? node39913 : node39896;
													assign node39896 = (inp[13]) ? node39908 : node39897;
														assign node39897 = (inp[2]) ? node39903 : node39898;
															assign node39898 = (inp[5]) ? 4'b0000 : node39899;
																assign node39899 = (inp[1]) ? 4'b0000 : 4'b0100;
															assign node39903 = (inp[1]) ? 4'b0101 : node39904;
																assign node39904 = (inp[5]) ? 4'b0100 : 4'b0000;
														assign node39908 = (inp[1]) ? node39910 : 4'b0001;
															assign node39910 = (inp[2]) ? 4'b0000 : 4'b0100;
													assign node39913 = (inp[13]) ? node39925 : node39914;
														assign node39914 = (inp[1]) ? node39922 : node39915;
															assign node39915 = (inp[2]) ? node39919 : node39916;
																assign node39916 = (inp[5]) ? 4'b0000 : 4'b0100;
																assign node39919 = (inp[5]) ? 4'b0101 : 4'b0000;
															assign node39922 = (inp[2]) ? 4'b0101 : 4'b0001;
														assign node39925 = (inp[2]) ? node39931 : node39926;
															assign node39926 = (inp[1]) ? 4'b0100 : node39927;
																assign node39927 = (inp[5]) ? 4'b0100 : 4'b0001;
															assign node39931 = (inp[5]) ? 4'b0000 : node39932;
																assign node39932 = (inp[1]) ? 4'b0000 : 4'b0100;
												assign node39936 = (inp[11]) ? node39956 : node39937;
													assign node39937 = (inp[13]) ? node39945 : node39938;
														assign node39938 = (inp[2]) ? node39940 : 4'b0001;
															assign node39940 = (inp[1]) ? 4'b0100 : node39941;
																assign node39941 = (inp[5]) ? 4'b0100 : 4'b0001;
														assign node39945 = (inp[2]) ? node39951 : node39946;
															assign node39946 = (inp[5]) ? 4'b0100 : node39947;
																assign node39947 = (inp[1]) ? 4'b0100 : 4'b0001;
															assign node39951 = (inp[1]) ? 4'b0000 : node39952;
																assign node39952 = (inp[5]) ? 4'b0000 : 4'b0100;
													assign node39956 = (inp[5]) ? node39966 : node39957;
														assign node39957 = (inp[1]) ? node39959 : 4'b0100;
															assign node39959 = (inp[13]) ? node39963 : node39960;
																assign node39960 = (inp[2]) ? 4'b0100 : 4'b0000;
																assign node39963 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node39966 = (inp[13]) ? node39970 : node39967;
															assign node39967 = (inp[2]) ? 4'b0100 : 4'b0000;
															assign node39970 = (inp[2]) ? 4'b0000 : 4'b0100;
						assign node39973 = (inp[13]) ? node40589 : node39974;
							assign node39974 = (inp[4]) ? node40390 : node39975;
								assign node39975 = (inp[12]) ? node40153 : node39976;
									assign node39976 = (inp[1]) ? node40048 : node39977;
										assign node39977 = (inp[15]) ? node40025 : node39978;
											assign node39978 = (inp[0]) ? node40010 : node39979;
												assign node39979 = (inp[5]) ? node40003 : node39980;
													assign node39980 = (inp[10]) ? node39988 : node39981;
														assign node39981 = (inp[2]) ? node39985 : node39982;
															assign node39982 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node39985 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node39988 = (inp[11]) ? node39996 : node39989;
															assign node39989 = (inp[9]) ? node39993 : node39990;
																assign node39990 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node39993 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node39996 = (inp[2]) ? node40000 : node39997;
																assign node39997 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node40000 = (inp[9]) ? 4'b0100 : 4'b0101;
													assign node40003 = (inp[2]) ? node40007 : node40004;
														assign node40004 = (inp[9]) ? 4'b0100 : 4'b0101;
														assign node40007 = (inp[9]) ? 4'b0101 : 4'b0100;
												assign node40010 = (inp[5]) ? node40018 : node40011;
													assign node40011 = (inp[9]) ? node40015 : node40012;
														assign node40012 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node40015 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node40018 = (inp[9]) ? node40022 : node40019;
														assign node40019 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node40022 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node40025 = (inp[2]) ? node40037 : node40026;
												assign node40026 = (inp[9]) ? node40032 : node40027;
													assign node40027 = (inp[5]) ? node40029 : 4'b0000;
														assign node40029 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node40032 = (inp[0]) ? node40034 : 4'b0001;
														assign node40034 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node40037 = (inp[9]) ? node40043 : node40038;
													assign node40038 = (inp[0]) ? node40040 : 4'b0001;
														assign node40040 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node40043 = (inp[0]) ? node40045 : 4'b0000;
														assign node40045 = (inp[5]) ? 4'b0001 : 4'b0000;
										assign node40048 = (inp[0]) ? node40078 : node40049;
											assign node40049 = (inp[9]) ? node40071 : node40050;
												assign node40050 = (inp[11]) ? node40058 : node40051;
													assign node40051 = (inp[2]) ? node40055 : node40052;
														assign node40052 = (inp[15]) ? 4'b0001 : 4'b0000;
														assign node40055 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node40058 = (inp[10]) ? node40064 : node40059;
														assign node40059 = (inp[15]) ? 4'b0000 : node40060;
															assign node40060 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node40064 = (inp[15]) ? node40068 : node40065;
															assign node40065 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node40068 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node40071 = (inp[2]) ? node40075 : node40072;
													assign node40072 = (inp[15]) ? 4'b0000 : 4'b0001;
													assign node40075 = (inp[15]) ? 4'b0001 : 4'b0000;
											assign node40078 = (inp[11]) ? node40114 : node40079;
												assign node40079 = (inp[9]) ? node40099 : node40080;
													assign node40080 = (inp[15]) ? node40092 : node40081;
														assign node40081 = (inp[10]) ? node40087 : node40082;
															assign node40082 = (inp[5]) ? 4'b0000 : node40083;
																assign node40083 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node40087 = (inp[2]) ? node40089 : 4'b0001;
																assign node40089 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node40092 = (inp[2]) ? node40096 : node40093;
															assign node40093 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node40096 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node40099 = (inp[15]) ? node40107 : node40100;
														assign node40100 = (inp[2]) ? node40104 : node40101;
															assign node40101 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node40104 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node40107 = (inp[2]) ? node40111 : node40108;
															assign node40108 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node40111 = (inp[5]) ? 4'b0000 : 4'b0001;
												assign node40114 = (inp[10]) ? node40140 : node40115;
													assign node40115 = (inp[2]) ? node40131 : node40116;
														assign node40116 = (inp[15]) ? node40124 : node40117;
															assign node40117 = (inp[9]) ? node40121 : node40118;
																assign node40118 = (inp[5]) ? 4'b0001 : 4'b0000;
																assign node40121 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node40124 = (inp[9]) ? node40128 : node40125;
																assign node40125 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node40128 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node40131 = (inp[5]) ? 4'b0001 : node40132;
															assign node40132 = (inp[15]) ? node40136 : node40133;
																assign node40133 = (inp[9]) ? 4'b0000 : 4'b0001;
																assign node40136 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node40140 = (inp[15]) ? node40142 : 4'b0000;
														assign node40142 = (inp[2]) ? node40148 : node40143;
															assign node40143 = (inp[9]) ? node40145 : 4'b0000;
																assign node40145 = (inp[5]) ? 4'b0001 : 4'b0000;
															assign node40148 = (inp[9]) ? node40150 : 4'b0001;
																assign node40150 = (inp[5]) ? 4'b0000 : 4'b0001;
									assign node40153 = (inp[1]) ? node40241 : node40154;
										assign node40154 = (inp[15]) ? node40178 : node40155;
											assign node40155 = (inp[9]) ? node40167 : node40156;
												assign node40156 = (inp[2]) ? node40162 : node40157;
													assign node40157 = (inp[0]) ? 4'b0000 : node40158;
														assign node40158 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node40162 = (inp[0]) ? 4'b0001 : node40163;
														assign node40163 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node40167 = (inp[2]) ? node40173 : node40168;
													assign node40168 = (inp[5]) ? 4'b0001 : node40169;
														assign node40169 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node40173 = (inp[5]) ? 4'b0000 : node40174;
														assign node40174 = (inp[0]) ? 4'b0000 : 4'b0001;
											assign node40178 = (inp[10]) ? node40220 : node40179;
												assign node40179 = (inp[11]) ? node40197 : node40180;
													assign node40180 = (inp[2]) ? node40188 : node40181;
														assign node40181 = (inp[9]) ? node40183 : 4'b0100;
															assign node40183 = (inp[5]) ? 4'b0101 : node40184;
																assign node40184 = (inp[0]) ? 4'b0101 : 4'b0100;
														assign node40188 = (inp[9]) ? node40194 : node40189;
															assign node40189 = (inp[0]) ? 4'b0101 : node40190;
																assign node40190 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node40194 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node40197 = (inp[0]) ? node40211 : node40198;
														assign node40198 = (inp[5]) ? node40204 : node40199;
															assign node40199 = (inp[2]) ? 4'b0100 : node40200;
																assign node40200 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node40204 = (inp[9]) ? node40208 : node40205;
																assign node40205 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node40208 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node40211 = (inp[5]) ? node40213 : 4'b0101;
															assign node40213 = (inp[2]) ? node40217 : node40214;
																assign node40214 = (inp[9]) ? 4'b0101 : 4'b0100;
																assign node40217 = (inp[9]) ? 4'b0100 : 4'b0101;
												assign node40220 = (inp[2]) ? node40230 : node40221;
													assign node40221 = (inp[9]) ? node40225 : node40222;
														assign node40222 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node40225 = (inp[5]) ? 4'b0101 : node40226;
															assign node40226 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node40230 = (inp[9]) ? node40236 : node40231;
														assign node40231 = (inp[0]) ? 4'b0101 : node40232;
															assign node40232 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node40236 = (inp[0]) ? 4'b0100 : node40237;
															assign node40237 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node40241 = (inp[11]) ? node40315 : node40242;
											assign node40242 = (inp[10]) ? node40274 : node40243;
												assign node40243 = (inp[0]) ? node40261 : node40244;
													assign node40244 = (inp[15]) ? node40252 : node40245;
														assign node40245 = (inp[9]) ? node40247 : 4'b0101;
															assign node40247 = (inp[2]) ? node40249 : 4'b0101;
																assign node40249 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node40252 = (inp[9]) ? 4'b0101 : node40253;
															assign node40253 = (inp[5]) ? node40257 : node40254;
																assign node40254 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node40257 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node40261 = (inp[9]) ? node40267 : node40262;
														assign node40262 = (inp[5]) ? 4'b0101 : node40263;
															assign node40263 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node40267 = (inp[2]) ? node40271 : node40268;
															assign node40268 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node40271 = (inp[15]) ? 4'b0100 : 4'b0101;
												assign node40274 = (inp[9]) ? node40298 : node40275;
													assign node40275 = (inp[2]) ? node40287 : node40276;
														assign node40276 = (inp[15]) ? node40282 : node40277;
															assign node40277 = (inp[5]) ? 4'b0101 : node40278;
																assign node40278 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node40282 = (inp[5]) ? 4'b0100 : node40283;
																assign node40283 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node40287 = (inp[15]) ? node40293 : node40288;
															assign node40288 = (inp[0]) ? 4'b0100 : node40289;
																assign node40289 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node40293 = (inp[0]) ? 4'b0101 : node40294;
																assign node40294 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node40298 = (inp[0]) ? node40308 : node40299;
														assign node40299 = (inp[5]) ? 4'b0100 : node40300;
															assign node40300 = (inp[15]) ? node40304 : node40301;
																assign node40301 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node40304 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node40308 = (inp[2]) ? node40312 : node40309;
															assign node40309 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node40312 = (inp[15]) ? 4'b0100 : 4'b0101;
											assign node40315 = (inp[10]) ? node40351 : node40316;
												assign node40316 = (inp[2]) ? node40336 : node40317;
													assign node40317 = (inp[15]) ? node40329 : node40318;
														assign node40318 = (inp[9]) ? node40324 : node40319;
															assign node40319 = (inp[0]) ? 4'b0101 : node40320;
																assign node40320 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node40324 = (inp[5]) ? 4'b0100 : node40325;
																assign node40325 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node40329 = (inp[9]) ? node40331 : 4'b0100;
															assign node40331 = (inp[0]) ? 4'b0101 : node40332;
																assign node40332 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node40336 = (inp[0]) ? 4'b0100 : node40337;
														assign node40337 = (inp[15]) ? node40343 : node40338;
															assign node40338 = (inp[9]) ? node40340 : 4'b0100;
																assign node40340 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node40343 = (inp[9]) ? node40347 : node40344;
																assign node40344 = (inp[5]) ? 4'b0101 : 4'b0100;
																assign node40347 = (inp[5]) ? 4'b0100 : 4'b0101;
												assign node40351 = (inp[9]) ? node40373 : node40352;
													assign node40352 = (inp[2]) ? node40364 : node40353;
														assign node40353 = (inp[15]) ? node40359 : node40354;
															assign node40354 = (inp[5]) ? 4'b0101 : node40355;
																assign node40355 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node40359 = (inp[0]) ? 4'b0100 : node40360;
																assign node40360 = (inp[5]) ? 4'b0100 : 4'b0101;
														assign node40364 = (inp[15]) ? node40370 : node40365;
															assign node40365 = (inp[5]) ? 4'b0100 : node40366;
																assign node40366 = (inp[0]) ? 4'b0100 : 4'b0101;
															assign node40370 = (inp[5]) ? 4'b0101 : 4'b0100;
													assign node40373 = (inp[5]) ? node40383 : node40374;
														assign node40374 = (inp[15]) ? node40376 : 4'b0101;
															assign node40376 = (inp[0]) ? node40380 : node40377;
																assign node40377 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node40380 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node40383 = (inp[2]) ? node40387 : node40384;
															assign node40384 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node40387 = (inp[15]) ? 4'b0100 : 4'b0101;
								assign node40390 = (inp[5]) ? node40554 : node40391;
									assign node40391 = (inp[2]) ? node40513 : node40392;
										assign node40392 = (inp[0]) ? node40438 : node40393;
											assign node40393 = (inp[10]) ? node40409 : node40394;
												assign node40394 = (inp[9]) ? node40402 : node40395;
													assign node40395 = (inp[15]) ? node40397 : 4'b0100;
														assign node40397 = (inp[12]) ? 4'b0101 : node40398;
															assign node40398 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node40402 = (inp[15]) ? node40404 : 4'b0101;
														assign node40404 = (inp[1]) ? 4'b0100 : node40405;
															assign node40405 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node40409 = (inp[11]) ? node40421 : node40410;
													assign node40410 = (inp[15]) ? node40416 : node40411;
														assign node40411 = (inp[9]) ? 4'b0101 : node40412;
															assign node40412 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node40416 = (inp[9]) ? node40418 : 4'b0101;
															assign node40418 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node40421 = (inp[12]) ? node40431 : node40422;
														assign node40422 = (inp[1]) ? node40424 : 4'b0100;
															assign node40424 = (inp[9]) ? node40428 : node40425;
																assign node40425 = (inp[15]) ? 4'b0101 : 4'b0100;
																assign node40428 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node40431 = (inp[9]) ? node40433 : 4'b0101;
															assign node40433 = (inp[15]) ? 4'b0100 : node40434;
																assign node40434 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node40438 = (inp[11]) ? node40472 : node40439;
												assign node40439 = (inp[10]) ? node40461 : node40440;
													assign node40440 = (inp[9]) ? node40452 : node40441;
														assign node40441 = (inp[15]) ? node40447 : node40442;
															assign node40442 = (inp[1]) ? 4'b0100 : node40443;
																assign node40443 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node40447 = (inp[12]) ? 4'b0101 : node40448;
																assign node40448 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node40452 = (inp[1]) ? 4'b0101 : node40453;
															assign node40453 = (inp[15]) ? node40457 : node40454;
																assign node40454 = (inp[12]) ? 4'b0101 : 4'b0100;
																assign node40457 = (inp[12]) ? 4'b0100 : 4'b0101;
													assign node40461 = (inp[9]) ? 4'b0100 : node40462;
														assign node40462 = (inp[15]) ? node40468 : node40463;
															assign node40463 = (inp[12]) ? 4'b0100 : node40464;
																assign node40464 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node40468 = (inp[12]) ? 4'b0101 : 4'b0100;
												assign node40472 = (inp[1]) ? node40490 : node40473;
													assign node40473 = (inp[12]) ? node40483 : node40474;
														assign node40474 = (inp[10]) ? node40476 : 4'b0101;
															assign node40476 = (inp[9]) ? node40480 : node40477;
																assign node40477 = (inp[15]) ? 4'b0100 : 4'b0101;
																assign node40480 = (inp[15]) ? 4'b0101 : 4'b0100;
														assign node40483 = (inp[9]) ? node40487 : node40484;
															assign node40484 = (inp[15]) ? 4'b0101 : 4'b0100;
															assign node40487 = (inp[15]) ? 4'b0100 : 4'b0101;
													assign node40490 = (inp[10]) ? node40500 : node40491;
														assign node40491 = (inp[12]) ? node40493 : 4'b0100;
															assign node40493 = (inp[9]) ? node40497 : node40494;
																assign node40494 = (inp[15]) ? 4'b0101 : 4'b0100;
																assign node40497 = (inp[15]) ? 4'b0100 : 4'b0101;
														assign node40500 = (inp[12]) ? node40506 : node40501;
															assign node40501 = (inp[15]) ? 4'b0101 : node40502;
																assign node40502 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node40506 = (inp[9]) ? node40510 : node40507;
																assign node40507 = (inp[15]) ? 4'b0101 : 4'b0100;
																assign node40510 = (inp[15]) ? 4'b0100 : 4'b0101;
										assign node40513 = (inp[9]) ? node40539 : node40514;
											assign node40514 = (inp[15]) ? node40534 : node40515;
												assign node40515 = (inp[1]) ? 4'b0100 : node40516;
													assign node40516 = (inp[10]) ? node40522 : node40517;
														assign node40517 = (inp[0]) ? 4'b0101 : node40518;
															assign node40518 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node40522 = (inp[11]) ? node40528 : node40523;
															assign node40523 = (inp[0]) ? node40525 : 4'b0100;
																assign node40525 = (inp[12]) ? 4'b0100 : 4'b0101;
															assign node40528 = (inp[0]) ? node40530 : 4'b0101;
																assign node40530 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node40534 = (inp[1]) ? 4'b0101 : node40535;
													assign node40535 = (inp[12]) ? 4'b0101 : 4'b0100;
											assign node40539 = (inp[15]) ? node40549 : node40540;
												assign node40540 = (inp[1]) ? 4'b0101 : node40541;
													assign node40541 = (inp[12]) ? node40545 : node40542;
														assign node40542 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node40545 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node40549 = (inp[12]) ? 4'b0100 : node40550;
													assign node40550 = (inp[1]) ? 4'b0100 : 4'b0101;
									assign node40554 = (inp[12]) ? node40574 : node40555;
										assign node40555 = (inp[9]) ? node40565 : node40556;
											assign node40556 = (inp[15]) ? node40562 : node40557;
												assign node40557 = (inp[0]) ? node40559 : 4'b0100;
													assign node40559 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node40562 = (inp[1]) ? 4'b0101 : 4'b0100;
											assign node40565 = (inp[1]) ? node40571 : node40566;
												assign node40566 = (inp[15]) ? 4'b0101 : node40567;
													assign node40567 = (inp[0]) ? 4'b0100 : 4'b0101;
												assign node40571 = (inp[15]) ? 4'b0100 : 4'b0101;
										assign node40574 = (inp[9]) ? node40582 : node40575;
											assign node40575 = (inp[15]) ? 4'b0101 : node40576;
												assign node40576 = (inp[1]) ? 4'b0100 : node40577;
													assign node40577 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node40582 = (inp[15]) ? 4'b0100 : node40583;
												assign node40583 = (inp[1]) ? 4'b0101 : node40584;
													assign node40584 = (inp[0]) ? 4'b0101 : 4'b0100;
							assign node40589 = (inp[4]) ? node40911 : node40590;
								assign node40590 = (inp[12]) ? node40792 : node40591;
									assign node40591 = (inp[1]) ? node40693 : node40592;
										assign node40592 = (inp[15]) ? node40650 : node40593;
											assign node40593 = (inp[5]) ? node40619 : node40594;
												assign node40594 = (inp[2]) ? node40610 : node40595;
													assign node40595 = (inp[11]) ? node40603 : node40596;
														assign node40596 = (inp[9]) ? node40600 : node40597;
															assign node40597 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node40600 = (inp[0]) ? 4'b0001 : 4'b0000;
														assign node40603 = (inp[9]) ? node40607 : node40604;
															assign node40604 = (inp[0]) ? 4'b0000 : 4'b0001;
															assign node40607 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node40610 = (inp[10]) ? 4'b0000 : node40611;
														assign node40611 = (inp[0]) ? node40615 : node40612;
															assign node40612 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node40615 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node40619 = (inp[0]) ? node40635 : node40620;
													assign node40620 = (inp[11]) ? node40628 : node40621;
														assign node40621 = (inp[9]) ? node40625 : node40622;
															assign node40622 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node40625 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node40628 = (inp[9]) ? node40632 : node40629;
															assign node40629 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node40632 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node40635 = (inp[10]) ? node40643 : node40636;
														assign node40636 = (inp[9]) ? node40640 : node40637;
															assign node40637 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node40640 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node40643 = (inp[11]) ? node40645 : 4'b0001;
															assign node40645 = (inp[2]) ? 4'b0001 : node40646;
																assign node40646 = (inp[9]) ? 4'b0001 : 4'b0000;
											assign node40650 = (inp[5]) ? node40678 : node40651;
												assign node40651 = (inp[0]) ? node40657 : node40652;
													assign node40652 = (inp[2]) ? 4'b0101 : node40653;
														assign node40653 = (inp[9]) ? 4'b0101 : 4'b0100;
													assign node40657 = (inp[11]) ? node40665 : node40658;
														assign node40658 = (inp[9]) ? node40662 : node40659;
															assign node40659 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node40662 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node40665 = (inp[10]) ? node40671 : node40666;
															assign node40666 = (inp[2]) ? 4'b0100 : node40667;
																assign node40667 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node40671 = (inp[9]) ? node40675 : node40672;
																assign node40672 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node40675 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node40678 = (inp[11]) ? node40686 : node40679;
													assign node40679 = (inp[9]) ? node40683 : node40680;
														assign node40680 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node40683 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node40686 = (inp[9]) ? node40690 : node40687;
														assign node40687 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node40690 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node40693 = (inp[11]) ? node40743 : node40694;
											assign node40694 = (inp[15]) ? node40726 : node40695;
												assign node40695 = (inp[0]) ? node40711 : node40696;
													assign node40696 = (inp[2]) ? node40704 : node40697;
														assign node40697 = (inp[9]) ? node40701 : node40698;
															assign node40698 = (inp[5]) ? 4'b0100 : 4'b0101;
															assign node40701 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node40704 = (inp[9]) ? node40708 : node40705;
															assign node40705 = (inp[5]) ? 4'b0101 : 4'b0100;
															assign node40708 = (inp[5]) ? 4'b0100 : 4'b0101;
													assign node40711 = (inp[10]) ? node40717 : node40712;
														assign node40712 = (inp[2]) ? 4'b0101 : node40713;
															assign node40713 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node40717 = (inp[5]) ? node40721 : node40718;
															assign node40718 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node40721 = (inp[9]) ? 4'b0100 : node40722;
																assign node40722 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node40726 = (inp[9]) ? node40732 : node40727;
													assign node40727 = (inp[2]) ? 4'b0101 : node40728;
														assign node40728 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node40732 = (inp[2]) ? node40738 : node40733;
														assign node40733 = (inp[0]) ? 4'b0101 : node40734;
															assign node40734 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node40738 = (inp[5]) ? 4'b0100 : node40739;
															assign node40739 = (inp[0]) ? 4'b0100 : 4'b0101;
											assign node40743 = (inp[10]) ? node40769 : node40744;
												assign node40744 = (inp[15]) ? node40760 : node40745;
													assign node40745 = (inp[2]) ? node40749 : node40746;
														assign node40746 = (inp[9]) ? 4'b0101 : 4'b0100;
														assign node40749 = (inp[9]) ? node40755 : node40750;
															assign node40750 = (inp[5]) ? 4'b0101 : node40751;
																assign node40751 = (inp[0]) ? 4'b0101 : 4'b0100;
															assign node40755 = (inp[5]) ? 4'b0100 : node40756;
																assign node40756 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node40760 = (inp[5]) ? node40762 : 4'b0100;
														assign node40762 = (inp[9]) ? node40766 : node40763;
															assign node40763 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node40766 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node40769 = (inp[2]) ? node40781 : node40770;
													assign node40770 = (inp[9]) ? node40776 : node40771;
														assign node40771 = (inp[5]) ? 4'b0100 : node40772;
															assign node40772 = (inp[0]) ? 4'b0100 : 4'b0101;
														assign node40776 = (inp[5]) ? 4'b0101 : node40777;
															assign node40777 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node40781 = (inp[9]) ? node40787 : node40782;
														assign node40782 = (inp[0]) ? 4'b0101 : node40783;
															assign node40783 = (inp[5]) ? 4'b0101 : 4'b0100;
														assign node40787 = (inp[0]) ? 4'b0100 : node40788;
															assign node40788 = (inp[5]) ? 4'b0100 : 4'b0101;
									assign node40792 = (inp[1]) ? node40840 : node40793;
										assign node40793 = (inp[15]) ? node40817 : node40794;
											assign node40794 = (inp[2]) ? node40806 : node40795;
												assign node40795 = (inp[9]) ? node40801 : node40796;
													assign node40796 = (inp[5]) ? node40798 : 4'b0101;
														assign node40798 = (inp[0]) ? 4'b0100 : 4'b0101;
													assign node40801 = (inp[5]) ? node40803 : 4'b0100;
														assign node40803 = (inp[0]) ? 4'b0101 : 4'b0100;
												assign node40806 = (inp[9]) ? node40812 : node40807;
													assign node40807 = (inp[5]) ? node40809 : 4'b0100;
														assign node40809 = (inp[0]) ? 4'b0101 : 4'b0100;
													assign node40812 = (inp[0]) ? node40814 : 4'b0101;
														assign node40814 = (inp[5]) ? 4'b0100 : 4'b0101;
											assign node40817 = (inp[2]) ? node40829 : node40818;
												assign node40818 = (inp[9]) ? node40824 : node40819;
													assign node40819 = (inp[5]) ? 4'b0000 : node40820;
														assign node40820 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node40824 = (inp[0]) ? 4'b0001 : node40825;
														assign node40825 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node40829 = (inp[9]) ? node40835 : node40830;
													assign node40830 = (inp[5]) ? 4'b0001 : node40831;
														assign node40831 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node40835 = (inp[0]) ? 4'b0000 : node40836;
														assign node40836 = (inp[5]) ? 4'b0000 : 4'b0001;
										assign node40840 = (inp[11]) ? node40888 : node40841;
											assign node40841 = (inp[0]) ? node40881 : node40842;
												assign node40842 = (inp[10]) ? node40858 : node40843;
													assign node40843 = (inp[5]) ? node40851 : node40844;
														assign node40844 = (inp[2]) ? node40848 : node40845;
															assign node40845 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node40848 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node40851 = (inp[2]) ? node40855 : node40852;
															assign node40852 = (inp[9]) ? 4'b0001 : 4'b0000;
															assign node40855 = (inp[9]) ? 4'b0000 : 4'b0001;
													assign node40858 = (inp[5]) ? node40866 : node40859;
														assign node40859 = (inp[2]) ? node40863 : node40860;
															assign node40860 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node40863 = (inp[9]) ? 4'b0001 : 4'b0000;
														assign node40866 = (inp[15]) ? node40874 : node40867;
															assign node40867 = (inp[2]) ? node40871 : node40868;
																assign node40868 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node40871 = (inp[9]) ? 4'b0000 : 4'b0001;
															assign node40874 = (inp[2]) ? node40878 : node40875;
																assign node40875 = (inp[9]) ? 4'b0001 : 4'b0000;
																assign node40878 = (inp[9]) ? 4'b0000 : 4'b0001;
												assign node40881 = (inp[2]) ? node40885 : node40882;
													assign node40882 = (inp[9]) ? 4'b0001 : 4'b0000;
													assign node40885 = (inp[9]) ? 4'b0000 : 4'b0001;
											assign node40888 = (inp[2]) ? node40900 : node40889;
												assign node40889 = (inp[9]) ? node40895 : node40890;
													assign node40890 = (inp[5]) ? 4'b0000 : node40891;
														assign node40891 = (inp[0]) ? 4'b0000 : 4'b0001;
													assign node40895 = (inp[0]) ? 4'b0001 : node40896;
														assign node40896 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node40900 = (inp[9]) ? node40906 : node40901;
													assign node40901 = (inp[5]) ? 4'b0001 : node40902;
														assign node40902 = (inp[0]) ? 4'b0001 : 4'b0000;
													assign node40906 = (inp[5]) ? 4'b0000 : node40907;
														assign node40907 = (inp[0]) ? 4'b0000 : 4'b0001;
								assign node40911 = (inp[9]) ? node40925 : node40912;
									assign node40912 = (inp[1]) ? 4'b0001 : node40913;
										assign node40913 = (inp[12]) ? node40919 : node40914;
											assign node40914 = (inp[0]) ? 4'b0000 : node40915;
												assign node40915 = (inp[15]) ? 4'b0000 : 4'b0001;
											assign node40919 = (inp[0]) ? 4'b0001 : node40920;
												assign node40920 = (inp[15]) ? 4'b0001 : 4'b0000;
									assign node40925 = (inp[1]) ? 4'b0000 : node40926;
										assign node40926 = (inp[12]) ? node40932 : node40927;
											assign node40927 = (inp[15]) ? 4'b0001 : node40928;
												assign node40928 = (inp[0]) ? 4'b0001 : 4'b0000;
											assign node40932 = (inp[0]) ? 4'b0000 : node40933;
												assign node40933 = (inp[15]) ? 4'b0000 : 4'b0001;
			assign node40938 = (inp[12]) ? node45034 : node40939;
				assign node40939 = (inp[6]) ? node43689 : node40940;
					assign node40940 = (inp[15]) ? node42280 : node40941;
						assign node40941 = (inp[14]) ? node41751 : node40942;
							assign node40942 = (inp[2]) ? node41316 : node40943;
								assign node40943 = (inp[7]) ? node41157 : node40944;
									assign node40944 = (inp[5]) ? node41040 : node40945;
										assign node40945 = (inp[4]) ? node41017 : node40946;
											assign node40946 = (inp[9]) ? node40986 : node40947;
												assign node40947 = (inp[11]) ? node40961 : node40948;
													assign node40948 = (inp[1]) ? node40954 : node40949;
														assign node40949 = (inp[13]) ? 4'b0001 : node40950;
															assign node40950 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node40954 = (inp[13]) ? node40958 : node40955;
															assign node40955 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node40958 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node40961 = (inp[13]) ? node40977 : node40962;
														assign node40962 = (inp[0]) ? node40970 : node40963;
															assign node40963 = (inp[1]) ? node40967 : node40964;
																assign node40964 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node40967 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node40970 = (inp[1]) ? node40974 : node40971;
																assign node40971 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node40974 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node40977 = (inp[0]) ? node40979 : 4'b0000;
															assign node40979 = (inp[1]) ? node40983 : node40980;
																assign node40980 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node40983 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node40986 = (inp[11]) ? node40994 : node40987;
													assign node40987 = (inp[10]) ? node40991 : node40988;
														assign node40988 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node40991 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node40994 = (inp[0]) ? node41004 : node40995;
														assign node40995 = (inp[1]) ? 4'b0001 : node40996;
															assign node40996 = (inp[10]) ? node41000 : node40997;
																assign node40997 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node41000 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node41004 = (inp[1]) ? node41010 : node41005;
															assign node41005 = (inp[13]) ? 4'b0001 : node41006;
																assign node41006 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node41010 = (inp[13]) ? node41014 : node41011;
																assign node41011 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node41014 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node41017 = (inp[10]) ? node41029 : node41018;
												assign node41018 = (inp[13]) ? node41024 : node41019;
													assign node41019 = (inp[11]) ? node41021 : 4'b0000;
														assign node41021 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node41024 = (inp[11]) ? node41026 : 4'b0001;
														assign node41026 = (inp[1]) ? 4'b0000 : 4'b0001;
												assign node41029 = (inp[13]) ? node41035 : node41030;
													assign node41030 = (inp[1]) ? node41032 : 4'b0001;
														assign node41032 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node41035 = (inp[1]) ? node41037 : 4'b0000;
														assign node41037 = (inp[11]) ? 4'b0001 : 4'b0000;
										assign node41040 = (inp[4]) ? node41094 : node41041;
											assign node41041 = (inp[11]) ? node41077 : node41042;
												assign node41042 = (inp[9]) ? node41064 : node41043;
													assign node41043 = (inp[1]) ? node41057 : node41044;
														assign node41044 = (inp[0]) ? node41052 : node41045;
															assign node41045 = (inp[13]) ? node41049 : node41046;
																assign node41046 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node41049 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node41052 = (inp[10]) ? node41054 : 4'b0001;
																assign node41054 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node41057 = (inp[13]) ? node41061 : node41058;
															assign node41058 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node41061 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node41064 = (inp[1]) ? node41070 : node41065;
														assign node41065 = (inp[10]) ? 4'b0000 : node41066;
															assign node41066 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node41070 = (inp[10]) ? node41074 : node41071;
															assign node41071 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node41074 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node41077 = (inp[13]) ? node41085 : node41078;
													assign node41078 = (inp[1]) ? node41082 : node41079;
														assign node41079 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node41082 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node41085 = (inp[9]) ? node41087 : 4'b0001;
														assign node41087 = (inp[1]) ? node41091 : node41088;
															assign node41088 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node41091 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node41094 = (inp[0]) ? node41134 : node41095;
												assign node41095 = (inp[9]) ? node41111 : node41096;
													assign node41096 = (inp[10]) ? node41100 : node41097;
														assign node41097 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node41100 = (inp[13]) ? node41106 : node41101;
															assign node41101 = (inp[11]) ? 4'b0100 : node41102;
																assign node41102 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node41106 = (inp[1]) ? 4'b0101 : node41107;
																assign node41107 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node41111 = (inp[11]) ? node41127 : node41112;
														assign node41112 = (inp[13]) ? node41120 : node41113;
															assign node41113 = (inp[10]) ? node41117 : node41114;
																assign node41114 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node41117 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node41120 = (inp[10]) ? node41124 : node41121;
																assign node41121 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node41124 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node41127 = (inp[13]) ? node41131 : node41128;
															assign node41128 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node41131 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node41134 = (inp[11]) ? node41150 : node41135;
													assign node41135 = (inp[10]) ? node41143 : node41136;
														assign node41136 = (inp[1]) ? node41140 : node41137;
															assign node41137 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node41140 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node41143 = (inp[13]) ? node41147 : node41144;
															assign node41144 = (inp[9]) ? 4'b0100 : 4'b0101;
															assign node41147 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node41150 = (inp[13]) ? node41154 : node41151;
														assign node41151 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41154 = (inp[10]) ? 4'b0101 : 4'b0100;
									assign node41157 = (inp[5]) ? node41251 : node41158;
										assign node41158 = (inp[4]) ? node41198 : node41159;
											assign node41159 = (inp[1]) ? node41175 : node41160;
												assign node41160 = (inp[11]) ? node41168 : node41161;
													assign node41161 = (inp[10]) ? node41165 : node41162;
														assign node41162 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node41165 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node41168 = (inp[10]) ? node41172 : node41169;
														assign node41169 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node41172 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node41175 = (inp[11]) ? node41191 : node41176;
													assign node41176 = (inp[0]) ? node41184 : node41177;
														assign node41177 = (inp[13]) ? node41181 : node41178;
															assign node41178 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node41181 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41184 = (inp[10]) ? node41188 : node41185;
															assign node41185 = (inp[9]) ? 4'b0101 : 4'b0100;
															assign node41188 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node41191 = (inp[13]) ? node41195 : node41192;
														assign node41192 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41195 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node41198 = (inp[9]) ? node41220 : node41199;
												assign node41199 = (inp[10]) ? node41209 : node41200;
													assign node41200 = (inp[13]) ? node41204 : node41201;
														assign node41201 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node41204 = (inp[11]) ? node41206 : 4'b0101;
															assign node41206 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node41209 = (inp[13]) ? node41215 : node41210;
														assign node41210 = (inp[11]) ? node41212 : 4'b0101;
															assign node41212 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node41215 = (inp[1]) ? node41217 : 4'b0100;
															assign node41217 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node41220 = (inp[1]) ? node41228 : node41221;
													assign node41221 = (inp[10]) ? node41225 : node41222;
														assign node41222 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node41225 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node41228 = (inp[11]) ? node41238 : node41229;
														assign node41229 = (inp[0]) ? node41235 : node41230;
															assign node41230 = (inp[10]) ? node41232 : 4'b0101;
																assign node41232 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node41235 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node41238 = (inp[0]) ? node41246 : node41239;
															assign node41239 = (inp[13]) ? node41243 : node41240;
																assign node41240 = (inp[10]) ? 4'b0100 : 4'b0101;
																assign node41243 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node41246 = (inp[10]) ? node41248 : 4'b0101;
																assign node41248 = (inp[13]) ? 4'b0101 : 4'b0100;
										assign node41251 = (inp[4]) ? node41293 : node41252;
											assign node41252 = (inp[11]) ? node41260 : node41253;
												assign node41253 = (inp[10]) ? node41257 : node41254;
													assign node41254 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node41257 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node41260 = (inp[0]) ? node41270 : node41261;
													assign node41261 = (inp[1]) ? 4'b0101 : node41262;
														assign node41262 = (inp[9]) ? node41264 : 4'b0101;
															assign node41264 = (inp[13]) ? 4'b0100 : node41265;
																assign node41265 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node41270 = (inp[9]) ? node41280 : node41271;
														assign node41271 = (inp[10]) ? node41273 : 4'b0100;
															assign node41273 = (inp[13]) ? node41277 : node41274;
																assign node41274 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node41277 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node41280 = (inp[10]) ? node41288 : node41281;
															assign node41281 = (inp[13]) ? node41285 : node41282;
																assign node41282 = (inp[1]) ? 4'b0100 : 4'b0101;
																assign node41285 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node41288 = (inp[1]) ? node41290 : 4'b0101;
																assign node41290 = (inp[13]) ? 4'b0100 : 4'b0101;
											assign node41293 = (inp[13]) ? node41305 : node41294;
												assign node41294 = (inp[10]) ? node41300 : node41295;
													assign node41295 = (inp[11]) ? node41297 : 4'b0000;
														assign node41297 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node41300 = (inp[1]) ? node41302 : 4'b0001;
														assign node41302 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node41305 = (inp[10]) ? node41311 : node41306;
													assign node41306 = (inp[1]) ? node41308 : 4'b0001;
														assign node41308 = (inp[11]) ? 4'b0000 : 4'b0001;
													assign node41311 = (inp[1]) ? node41313 : 4'b0000;
														assign node41313 = (inp[11]) ? 4'b0001 : 4'b0000;
								assign node41316 = (inp[7]) ? node41558 : node41317;
									assign node41317 = (inp[4]) ? node41471 : node41318;
										assign node41318 = (inp[11]) ? node41382 : node41319;
											assign node41319 = (inp[0]) ? node41355 : node41320;
												assign node41320 = (inp[5]) ? node41340 : node41321;
													assign node41321 = (inp[1]) ? node41333 : node41322;
														assign node41322 = (inp[9]) ? node41328 : node41323;
															assign node41323 = (inp[10]) ? 4'b0101 : node41324;
																assign node41324 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node41328 = (inp[10]) ? node41330 : 4'b0101;
																assign node41330 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node41333 = (inp[13]) ? node41337 : node41334;
															assign node41334 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node41337 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node41340 = (inp[9]) ? node41348 : node41341;
														assign node41341 = (inp[13]) ? node41345 : node41342;
															assign node41342 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node41345 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41348 = (inp[10]) ? node41352 : node41349;
															assign node41349 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node41352 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node41355 = (inp[9]) ? node41369 : node41356;
													assign node41356 = (inp[1]) ? node41364 : node41357;
														assign node41357 = (inp[13]) ? node41361 : node41358;
															assign node41358 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node41361 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41364 = (inp[13]) ? node41366 : 4'b0100;
															assign node41366 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node41369 = (inp[5]) ? node41377 : node41370;
														assign node41370 = (inp[10]) ? node41374 : node41371;
															assign node41371 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node41374 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node41377 = (inp[13]) ? 4'b0100 : node41378;
															assign node41378 = (inp[10]) ? 4'b0101 : 4'b0100;
											assign node41382 = (inp[5]) ? node41428 : node41383;
												assign node41383 = (inp[0]) ? node41407 : node41384;
													assign node41384 = (inp[13]) ? node41396 : node41385;
														assign node41385 = (inp[9]) ? node41391 : node41386;
															assign node41386 = (inp[10]) ? node41388 : 4'b0100;
																assign node41388 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node41391 = (inp[1]) ? node41393 : 4'b0100;
																assign node41393 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41396 = (inp[9]) ? node41402 : node41397;
															assign node41397 = (inp[10]) ? node41399 : 4'b0100;
																assign node41399 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node41402 = (inp[1]) ? 4'b0100 : node41403;
																assign node41403 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node41407 = (inp[1]) ? node41423 : node41408;
														assign node41408 = (inp[9]) ? node41416 : node41409;
															assign node41409 = (inp[10]) ? node41413 : node41410;
																assign node41410 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node41413 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node41416 = (inp[13]) ? node41420 : node41417;
																assign node41417 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node41420 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41423 = (inp[10]) ? node41425 : 4'b0101;
															assign node41425 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node41428 = (inp[0]) ? node41450 : node41429;
													assign node41429 = (inp[9]) ? node41443 : node41430;
														assign node41430 = (inp[1]) ? node41438 : node41431;
															assign node41431 = (inp[10]) ? node41435 : node41432;
																assign node41432 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node41435 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node41438 = (inp[10]) ? 4'b0101 : node41439;
																assign node41439 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node41443 = (inp[13]) ? 4'b0101 : node41444;
															assign node41444 = (inp[10]) ? node41446 : 4'b0101;
																assign node41446 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node41450 = (inp[13]) ? node41464 : node41451;
														assign node41451 = (inp[9]) ? node41457 : node41452;
															assign node41452 = (inp[10]) ? node41454 : 4'b0101;
																assign node41454 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node41457 = (inp[10]) ? node41461 : node41458;
																assign node41458 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node41461 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node41464 = (inp[1]) ? node41468 : node41465;
															assign node41465 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node41468 = (inp[10]) ? 4'b0101 : 4'b0100;
										assign node41471 = (inp[5]) ? node41511 : node41472;
											assign node41472 = (inp[11]) ? node41480 : node41473;
												assign node41473 = (inp[13]) ? node41477 : node41474;
													assign node41474 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node41477 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node41480 = (inp[1]) ? node41488 : node41481;
													assign node41481 = (inp[13]) ? node41485 : node41482;
														assign node41482 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41485 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node41488 = (inp[0]) ? node41498 : node41489;
														assign node41489 = (inp[9]) ? 4'b0101 : node41490;
															assign node41490 = (inp[10]) ? node41494 : node41491;
																assign node41491 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node41494 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node41498 = (inp[9]) ? node41506 : node41499;
															assign node41499 = (inp[10]) ? node41503 : node41500;
																assign node41500 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node41503 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node41506 = (inp[10]) ? 4'b0100 : node41507;
																assign node41507 = (inp[13]) ? 4'b0101 : 4'b0100;
											assign node41511 = (inp[1]) ? node41535 : node41512;
												assign node41512 = (inp[11]) ? node41520 : node41513;
													assign node41513 = (inp[10]) ? node41517 : node41514;
														assign node41514 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node41517 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node41520 = (inp[9]) ? node41528 : node41521;
														assign node41521 = (inp[0]) ? node41523 : 4'b0001;
															assign node41523 = (inp[10]) ? 4'b0001 : node41524;
																assign node41524 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node41528 = (inp[10]) ? node41532 : node41529;
															assign node41529 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node41532 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node41535 = (inp[10]) ? node41551 : node41536;
													assign node41536 = (inp[0]) ? node41544 : node41537;
														assign node41537 = (inp[11]) ? node41541 : node41538;
															assign node41538 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node41541 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node41544 = (inp[11]) ? node41548 : node41545;
															assign node41545 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node41548 = (inp[13]) ? 4'b0000 : 4'b0001;
													assign node41551 = (inp[13]) ? node41555 : node41552;
														assign node41552 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node41555 = (inp[11]) ? 4'b0001 : 4'b0000;
									assign node41558 = (inp[5]) ? node41652 : node41559;
										assign node41559 = (inp[1]) ? node41607 : node41560;
											assign node41560 = (inp[11]) ? node41592 : node41561;
												assign node41561 = (inp[4]) ? node41569 : node41562;
													assign node41562 = (inp[13]) ? node41566 : node41563;
														assign node41563 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node41566 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node41569 = (inp[9]) ? node41585 : node41570;
														assign node41570 = (inp[0]) ? node41578 : node41571;
															assign node41571 = (inp[13]) ? node41575 : node41572;
																assign node41572 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node41575 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node41578 = (inp[13]) ? node41582 : node41579;
																assign node41579 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node41582 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node41585 = (inp[10]) ? node41589 : node41586;
															assign node41586 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node41589 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node41592 = (inp[4]) ? node41600 : node41593;
													assign node41593 = (inp[9]) ? 4'b0000 : node41594;
														assign node41594 = (inp[10]) ? node41596 : 4'b0000;
															assign node41596 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node41600 = (inp[13]) ? node41604 : node41601;
														assign node41601 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node41604 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node41607 = (inp[13]) ? node41615 : node41608;
												assign node41608 = (inp[4]) ? node41612 : node41609;
													assign node41609 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node41612 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node41615 = (inp[0]) ? node41637 : node41616;
													assign node41616 = (inp[11]) ? node41624 : node41617;
														assign node41617 = (inp[4]) ? node41621 : node41618;
															assign node41618 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node41621 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node41624 = (inp[9]) ? node41632 : node41625;
															assign node41625 = (inp[4]) ? node41629 : node41626;
																assign node41626 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node41629 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node41632 = (inp[10]) ? 4'b0001 : node41633;
																assign node41633 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node41637 = (inp[9]) ? node41645 : node41638;
														assign node41638 = (inp[10]) ? node41642 : node41639;
															assign node41639 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node41642 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node41645 = (inp[4]) ? node41649 : node41646;
															assign node41646 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node41649 = (inp[10]) ? 4'b0000 : 4'b0001;
										assign node41652 = (inp[4]) ? node41676 : node41653;
											assign node41653 = (inp[10]) ? node41665 : node41654;
												assign node41654 = (inp[13]) ? node41660 : node41655;
													assign node41655 = (inp[11]) ? 4'b0000 : node41656;
														assign node41656 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node41660 = (inp[1]) ? 4'b0001 : node41661;
														assign node41661 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node41665 = (inp[13]) ? node41671 : node41666;
													assign node41666 = (inp[1]) ? 4'b0001 : node41667;
														assign node41667 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node41671 = (inp[11]) ? 4'b0000 : node41672;
														assign node41672 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node41676 = (inp[9]) ? node41724 : node41677;
												assign node41677 = (inp[1]) ? node41697 : node41678;
													assign node41678 = (inp[0]) ? node41684 : node41679;
														assign node41679 = (inp[13]) ? node41681 : 4'b0101;
															assign node41681 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node41684 = (inp[11]) ? node41692 : node41685;
															assign node41685 = (inp[10]) ? node41689 : node41686;
																assign node41686 = (inp[13]) ? 4'b0100 : 4'b0101;
																assign node41689 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node41692 = (inp[13]) ? node41694 : 4'b0100;
																assign node41694 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node41697 = (inp[0]) ? node41711 : node41698;
														assign node41698 = (inp[11]) ? node41704 : node41699;
															assign node41699 = (inp[10]) ? node41701 : 4'b0100;
																assign node41701 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node41704 = (inp[13]) ? node41708 : node41705;
																assign node41705 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node41708 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41711 = (inp[10]) ? node41717 : node41712;
															assign node41712 = (inp[11]) ? node41714 : 4'b0101;
																assign node41714 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node41717 = (inp[11]) ? node41721 : node41718;
																assign node41718 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node41721 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node41724 = (inp[1]) ? node41732 : node41725;
													assign node41725 = (inp[13]) ? node41729 : node41726;
														assign node41726 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node41729 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node41732 = (inp[10]) ? node41740 : node41733;
														assign node41733 = (inp[0]) ? 4'b0100 : node41734;
															assign node41734 = (inp[13]) ? node41736 : 4'b0100;
																assign node41736 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node41740 = (inp[0]) ? node41746 : node41741;
															assign node41741 = (inp[13]) ? 4'b0100 : node41742;
																assign node41742 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node41746 = (inp[11]) ? 4'b0100 : node41747;
																assign node41747 = (inp[13]) ? 4'b0101 : 4'b0100;
							assign node41751 = (inp[5]) ? node41925 : node41752;
								assign node41752 = (inp[13]) ? node41828 : node41753;
									assign node41753 = (inp[10]) ? node41789 : node41754;
										assign node41754 = (inp[2]) ? node41766 : node41755;
											assign node41755 = (inp[7]) ? node41761 : node41756;
												assign node41756 = (inp[1]) ? 4'b0010 : node41757;
													assign node41757 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node41761 = (inp[1]) ? 4'b0110 : node41762;
													assign node41762 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node41766 = (inp[7]) ? node41778 : node41767;
												assign node41767 = (inp[4]) ? node41773 : node41768;
													assign node41768 = (inp[1]) ? node41770 : 4'b0110;
														assign node41770 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node41773 = (inp[1]) ? node41775 : 4'b0111;
														assign node41775 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node41778 = (inp[4]) ? node41784 : node41779;
													assign node41779 = (inp[11]) ? node41781 : 4'b0011;
														assign node41781 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node41784 = (inp[11]) ? node41786 : 4'b0010;
														assign node41786 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node41789 = (inp[11]) ? node41805 : node41790;
											assign node41790 = (inp[2]) ? node41794 : node41791;
												assign node41791 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node41794 = (inp[7]) ? node41802 : node41795;
													assign node41795 = (inp[4]) ? node41799 : node41796;
														assign node41796 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node41799 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node41802 = (inp[4]) ? 4'b0011 : 4'b0010;
											assign node41805 = (inp[1]) ? node41817 : node41806;
												assign node41806 = (inp[2]) ? node41810 : node41807;
													assign node41807 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node41810 = (inp[7]) ? node41814 : node41811;
														assign node41811 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node41814 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node41817 = (inp[2]) ? node41821 : node41818;
													assign node41818 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node41821 = (inp[7]) ? node41825 : node41822;
														assign node41822 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node41825 = (inp[4]) ? 4'b0011 : 4'b0010;
									assign node41828 = (inp[10]) ? node41878 : node41829;
										assign node41829 = (inp[1]) ? node41851 : node41830;
											assign node41830 = (inp[11]) ? node41842 : node41831;
												assign node41831 = (inp[2]) ? node41835 : node41832;
													assign node41832 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node41835 = (inp[7]) ? node41839 : node41836;
														assign node41836 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node41839 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node41842 = (inp[2]) ? node41846 : node41843;
													assign node41843 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node41846 = (inp[4]) ? 4'b0110 : node41847;
														assign node41847 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node41851 = (inp[2]) ? node41855 : node41852;
												assign node41852 = (inp[7]) ? 4'b0111 : 4'b0011;
												assign node41855 = (inp[7]) ? node41875 : node41856;
													assign node41856 = (inp[0]) ? node41862 : node41857;
														assign node41857 = (inp[4]) ? 4'b0110 : node41858;
															assign node41858 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node41862 = (inp[9]) ? node41870 : node41863;
															assign node41863 = (inp[4]) ? node41867 : node41864;
																assign node41864 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node41867 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node41870 = (inp[4]) ? 4'b0111 : node41871;
																assign node41871 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node41875 = (inp[4]) ? 4'b0011 : 4'b0010;
										assign node41878 = (inp[11]) ? node41902 : node41879;
											assign node41879 = (inp[7]) ? node41897 : node41880;
												assign node41880 = (inp[2]) ? node41882 : 4'b0010;
													assign node41882 = (inp[0]) ? node41890 : node41883;
														assign node41883 = (inp[9]) ? 4'b0110 : node41884;
															assign node41884 = (inp[4]) ? node41886 : 4'b0110;
																assign node41886 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node41890 = (inp[9]) ? node41892 : 4'b0110;
															assign node41892 = (inp[1]) ? node41894 : 4'b0111;
																assign node41894 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node41897 = (inp[2]) ? node41899 : 4'b0110;
													assign node41899 = (inp[4]) ? 4'b0010 : 4'b0011;
											assign node41902 = (inp[1]) ? node41914 : node41903;
												assign node41903 = (inp[2]) ? node41907 : node41904;
													assign node41904 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node41907 = (inp[4]) ? node41911 : node41908;
														assign node41908 = (inp[7]) ? 4'b0010 : 4'b0110;
														assign node41911 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node41914 = (inp[2]) ? node41918 : node41915;
													assign node41915 = (inp[7]) ? 4'b0110 : 4'b0010;
													assign node41918 = (inp[7]) ? node41922 : node41919;
														assign node41919 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node41922 = (inp[4]) ? 4'b0010 : 4'b0011;
								assign node41925 = (inp[7]) ? node42173 : node41926;
									assign node41926 = (inp[9]) ? node42038 : node41927;
										assign node41927 = (inp[4]) ? node41985 : node41928;
											assign node41928 = (inp[2]) ? node41952 : node41929;
												assign node41929 = (inp[0]) ? node41937 : node41930;
													assign node41930 = (inp[13]) ? 4'b0111 : node41931;
														assign node41931 = (inp[10]) ? 4'b0111 : node41932;
															assign node41932 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node41937 = (inp[10]) ? node41945 : node41938;
														assign node41938 = (inp[13]) ? 4'b0111 : node41939;
															assign node41939 = (inp[1]) ? 4'b0110 : node41940;
																assign node41940 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node41945 = (inp[13]) ? 4'b0110 : node41946;
															assign node41946 = (inp[11]) ? node41948 : 4'b0111;
																assign node41948 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node41952 = (inp[0]) ? node41972 : node41953;
													assign node41953 = (inp[10]) ? node41963 : node41954;
														assign node41954 = (inp[1]) ? node41960 : node41955;
															assign node41955 = (inp[11]) ? node41957 : 4'b0010;
																assign node41957 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node41960 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node41963 = (inp[1]) ? 4'b0010 : node41964;
															assign node41964 = (inp[13]) ? node41968 : node41965;
																assign node41965 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node41968 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node41972 = (inp[13]) ? node41978 : node41973;
														assign node41973 = (inp[10]) ? node41975 : 4'b0011;
															assign node41975 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node41978 = (inp[10]) ? node41980 : 4'b0010;
															assign node41980 = (inp[11]) ? node41982 : 4'b0011;
																assign node41982 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node41985 = (inp[2]) ? node42005 : node41986;
												assign node41986 = (inp[13]) ? node41994 : node41987;
													assign node41987 = (inp[10]) ? 4'b0010 : node41988;
														assign node41988 = (inp[11]) ? node41990 : 4'b0011;
															assign node41990 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node41994 = (inp[10]) ? node42000 : node41995;
														assign node41995 = (inp[1]) ? 4'b0010 : node41996;
															assign node41996 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node42000 = (inp[1]) ? 4'b0011 : node42001;
															assign node42001 = (inp[0]) ? 4'b0011 : 4'b0010;
												assign node42005 = (inp[11]) ? node42031 : node42006;
													assign node42006 = (inp[13]) ? node42016 : node42007;
														assign node42007 = (inp[0]) ? 4'b0111 : node42008;
															assign node42008 = (inp[10]) ? node42012 : node42009;
																assign node42009 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node42012 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node42016 = (inp[0]) ? node42024 : node42017;
															assign node42017 = (inp[10]) ? node42021 : node42018;
																assign node42018 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node42021 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node42024 = (inp[1]) ? node42028 : node42025;
																assign node42025 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node42028 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node42031 = (inp[13]) ? node42035 : node42032;
														assign node42032 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node42035 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node42038 = (inp[0]) ? node42096 : node42039;
											assign node42039 = (inp[4]) ? node42067 : node42040;
												assign node42040 = (inp[2]) ? node42052 : node42041;
													assign node42041 = (inp[13]) ? node42049 : node42042;
														assign node42042 = (inp[10]) ? 4'b0111 : node42043;
															assign node42043 = (inp[11]) ? node42045 : 4'b0110;
																assign node42045 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node42049 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node42052 = (inp[1]) ? node42060 : node42053;
														assign node42053 = (inp[13]) ? 4'b0011 : node42054;
															assign node42054 = (inp[10]) ? 4'b0011 : node42055;
																assign node42055 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node42060 = (inp[13]) ? node42064 : node42061;
															assign node42061 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node42064 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node42067 = (inp[2]) ? node42085 : node42068;
													assign node42068 = (inp[10]) ? node42080 : node42069;
														assign node42069 = (inp[13]) ? node42075 : node42070;
															assign node42070 = (inp[1]) ? 4'b0011 : node42071;
																assign node42071 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node42075 = (inp[1]) ? 4'b0010 : node42076;
																assign node42076 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node42080 = (inp[11]) ? node42082 : 4'b0010;
															assign node42082 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node42085 = (inp[10]) ? node42091 : node42086;
														assign node42086 = (inp[13]) ? node42088 : 4'b0110;
															assign node42088 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42091 = (inp[13]) ? node42093 : 4'b0111;
															assign node42093 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node42096 = (inp[4]) ? node42142 : node42097;
												assign node42097 = (inp[2]) ? node42113 : node42098;
													assign node42098 = (inp[11]) ? node42104 : node42099;
														assign node42099 = (inp[13]) ? node42101 : 4'b0110;
															assign node42101 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node42104 = (inp[13]) ? node42106 : 4'b0111;
															assign node42106 = (inp[1]) ? node42110 : node42107;
																assign node42107 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node42110 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node42113 = (inp[1]) ? node42127 : node42114;
														assign node42114 = (inp[11]) ? node42122 : node42115;
															assign node42115 = (inp[13]) ? node42119 : node42116;
																assign node42116 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node42119 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node42122 = (inp[10]) ? 4'b0010 : node42123;
																assign node42123 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node42127 = (inp[11]) ? node42135 : node42128;
															assign node42128 = (inp[13]) ? node42132 : node42129;
																assign node42129 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node42132 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node42135 = (inp[10]) ? node42139 : node42136;
																assign node42136 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node42139 = (inp[13]) ? 4'b0011 : 4'b0010;
												assign node42142 = (inp[2]) ? node42158 : node42143;
													assign node42143 = (inp[10]) ? node42151 : node42144;
														assign node42144 = (inp[13]) ? node42146 : 4'b0011;
															assign node42146 = (inp[1]) ? 4'b0010 : node42147;
																assign node42147 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node42151 = (inp[13]) ? 4'b0011 : node42152;
															assign node42152 = (inp[1]) ? 4'b0010 : node42153;
																assign node42153 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node42158 = (inp[11]) ? node42166 : node42159;
														assign node42159 = (inp[1]) ? 4'b0111 : node42160;
															assign node42160 = (inp[10]) ? node42162 : 4'b0111;
																assign node42162 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node42166 = (inp[10]) ? node42170 : node42167;
															assign node42167 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node42170 = (inp[13]) ? 4'b0110 : 4'b0111;
									assign node42173 = (inp[1]) ? node42241 : node42174;
										assign node42174 = (inp[10]) ? node42208 : node42175;
											assign node42175 = (inp[13]) ? node42191 : node42176;
												assign node42176 = (inp[11]) ? node42184 : node42177;
													assign node42177 = (inp[4]) ? node42181 : node42178;
														assign node42178 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node42181 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node42184 = (inp[2]) ? node42188 : node42185;
														assign node42185 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node42188 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node42191 = (inp[11]) ? node42199 : node42192;
													assign node42192 = (inp[4]) ? node42196 : node42193;
														assign node42193 = (inp[2]) ? 4'b0111 : 4'b0010;
														assign node42196 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node42199 = (inp[0]) ? 4'b0010 : node42200;
														assign node42200 = (inp[4]) ? node42204 : node42201;
															assign node42201 = (inp[2]) ? 4'b0110 : 4'b0010;
															assign node42204 = (inp[2]) ? 4'b0010 : 4'b0110;
											assign node42208 = (inp[13]) ? node42224 : node42209;
												assign node42209 = (inp[11]) ? node42217 : node42210;
													assign node42210 = (inp[2]) ? node42214 : node42211;
														assign node42211 = (inp[4]) ? 4'b0111 : 4'b0010;
														assign node42214 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node42217 = (inp[4]) ? node42221 : node42218;
														assign node42218 = (inp[2]) ? 4'b0110 : 4'b0010;
														assign node42221 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node42224 = (inp[11]) ? node42234 : node42225;
													assign node42225 = (inp[0]) ? node42227 : 4'b0110;
														assign node42227 = (inp[4]) ? node42231 : node42228;
															assign node42228 = (inp[2]) ? 4'b0110 : 4'b0011;
															assign node42231 = (inp[2]) ? 4'b0010 : 4'b0110;
													assign node42234 = (inp[2]) ? node42238 : node42235;
														assign node42235 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node42238 = (inp[4]) ? 4'b0011 : 4'b0111;
										assign node42241 = (inp[10]) ? node42261 : node42242;
											assign node42242 = (inp[13]) ? node42252 : node42243;
												assign node42243 = (inp[4]) ? node42249 : node42244;
													assign node42244 = (inp[2]) ? 4'b0110 : node42245;
														assign node42245 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node42249 = (inp[2]) ? 4'b0010 : 4'b0110;
												assign node42252 = (inp[2]) ? node42258 : node42253;
													assign node42253 = (inp[4]) ? 4'b0111 : node42254;
														assign node42254 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node42258 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node42261 = (inp[13]) ? node42271 : node42262;
												assign node42262 = (inp[4]) ? node42268 : node42263;
													assign node42263 = (inp[2]) ? 4'b0111 : node42264;
														assign node42264 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node42268 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node42271 = (inp[4]) ? node42277 : node42272;
													assign node42272 = (inp[2]) ? 4'b0110 : node42273;
														assign node42273 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node42277 = (inp[2]) ? 4'b0010 : 4'b0110;
						assign node42280 = (inp[13]) ? node43022 : node42281;
							assign node42281 = (inp[2]) ? node42749 : node42282;
								assign node42282 = (inp[4]) ? node42540 : node42283;
									assign node42283 = (inp[0]) ? node42445 : node42284;
										assign node42284 = (inp[9]) ? node42362 : node42285;
											assign node42285 = (inp[14]) ? node42311 : node42286;
												assign node42286 = (inp[10]) ? node42298 : node42287;
													assign node42287 = (inp[1]) ? 4'b0011 : node42288;
														assign node42288 = (inp[7]) ? node42290 : 4'b0010;
															assign node42290 = (inp[11]) ? node42294 : node42291;
																assign node42291 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node42294 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node42298 = (inp[1]) ? node42304 : node42299;
														assign node42299 = (inp[11]) ? node42301 : 4'b0011;
															assign node42301 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node42304 = (inp[5]) ? 4'b0010 : node42305;
															assign node42305 = (inp[7]) ? node42307 : 4'b0010;
																assign node42307 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node42311 = (inp[11]) ? node42333 : node42312;
													assign node42312 = (inp[7]) ? node42320 : node42313;
														assign node42313 = (inp[10]) ? node42317 : node42314;
															assign node42314 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node42317 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node42320 = (inp[5]) ? node42328 : node42321;
															assign node42321 = (inp[1]) ? node42325 : node42322;
																assign node42322 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node42325 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node42328 = (inp[1]) ? node42330 : 4'b0010;
																assign node42330 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node42333 = (inp[10]) ? node42347 : node42334;
														assign node42334 = (inp[5]) ? node42340 : node42335;
															assign node42335 = (inp[1]) ? node42337 : 4'b0011;
																assign node42337 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node42340 = (inp[7]) ? node42344 : node42341;
																assign node42341 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node42344 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node42347 = (inp[7]) ? node42355 : node42348;
															assign node42348 = (inp[1]) ? node42352 : node42349;
																assign node42349 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node42352 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node42355 = (inp[5]) ? node42359 : node42356;
																assign node42356 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node42359 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node42362 = (inp[14]) ? node42412 : node42363;
												assign node42363 = (inp[5]) ? node42381 : node42364;
													assign node42364 = (inp[7]) ? node42372 : node42365;
														assign node42365 = (inp[1]) ? node42369 : node42366;
															assign node42366 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node42369 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node42372 = (inp[10]) ? node42374 : 4'b0011;
															assign node42374 = (inp[11]) ? node42378 : node42375;
																assign node42375 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node42378 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node42381 = (inp[11]) ? node42397 : node42382;
														assign node42382 = (inp[10]) ? node42390 : node42383;
															assign node42383 = (inp[1]) ? node42387 : node42384;
																assign node42384 = (inp[7]) ? 4'b0011 : 4'b0010;
																assign node42387 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node42390 = (inp[7]) ? node42394 : node42391;
																assign node42391 = (inp[1]) ? 4'b0010 : 4'b0011;
																assign node42394 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node42397 = (inp[7]) ? node42405 : node42398;
															assign node42398 = (inp[10]) ? node42402 : node42399;
																assign node42399 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node42402 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node42405 = (inp[1]) ? node42409 : node42406;
																assign node42406 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node42409 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node42412 = (inp[10]) ? node42430 : node42413;
													assign node42413 = (inp[1]) ? node42421 : node42414;
														assign node42414 = (inp[11]) ? node42416 : 4'b0010;
															assign node42416 = (inp[5]) ? 4'b0011 : node42417;
																assign node42417 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node42421 = (inp[11]) ? node42423 : 4'b0011;
															assign node42423 = (inp[7]) ? node42427 : node42424;
																assign node42424 = (inp[5]) ? 4'b0011 : 4'b0010;
																assign node42427 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node42430 = (inp[1]) ? node42438 : node42431;
														assign node42431 = (inp[11]) ? node42433 : 4'b0011;
															assign node42433 = (inp[5]) ? node42435 : 4'b0011;
																assign node42435 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node42438 = (inp[11]) ? node42440 : 4'b0010;
															assign node42440 = (inp[7]) ? node42442 : 4'b0011;
																assign node42442 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node42445 = (inp[10]) ? node42497 : node42446;
											assign node42446 = (inp[1]) ? node42474 : node42447;
												assign node42447 = (inp[11]) ? node42455 : node42448;
													assign node42448 = (inp[7]) ? node42450 : 4'b0010;
														assign node42450 = (inp[14]) ? 4'b0010 : node42451;
															assign node42451 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node42455 = (inp[5]) ? node42469 : node42456;
														assign node42456 = (inp[9]) ? node42464 : node42457;
															assign node42457 = (inp[7]) ? node42461 : node42458;
																assign node42458 = (inp[14]) ? 4'b0011 : 4'b0010;
																assign node42461 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node42464 = (inp[7]) ? 4'b0011 : node42465;
																assign node42465 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node42469 = (inp[7]) ? node42471 : 4'b0010;
															assign node42471 = (inp[14]) ? 4'b0011 : 4'b0010;
												assign node42474 = (inp[11]) ? node42484 : node42475;
													assign node42475 = (inp[9]) ? node42477 : 4'b0011;
														assign node42477 = (inp[5]) ? node42479 : 4'b0011;
															assign node42479 = (inp[7]) ? node42481 : 4'b0011;
																assign node42481 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node42484 = (inp[5]) ? node42492 : node42485;
														assign node42485 = (inp[14]) ? node42489 : node42486;
															assign node42486 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node42489 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node42492 = (inp[7]) ? node42494 : 4'b0011;
															assign node42494 = (inp[14]) ? 4'b0010 : 4'b0011;
											assign node42497 = (inp[1]) ? node42519 : node42498;
												assign node42498 = (inp[11]) ? node42508 : node42499;
													assign node42499 = (inp[9]) ? node42501 : 4'b0011;
														assign node42501 = (inp[7]) ? node42503 : 4'b0011;
															assign node42503 = (inp[5]) ? node42505 : 4'b0011;
																assign node42505 = (inp[14]) ? 4'b0011 : 4'b0010;
													assign node42508 = (inp[5]) ? node42516 : node42509;
														assign node42509 = (inp[14]) ? node42513 : node42510;
															assign node42510 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node42513 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node42516 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node42519 = (inp[11]) ? node42527 : node42520;
													assign node42520 = (inp[14]) ? 4'b0010 : node42521;
														assign node42521 = (inp[5]) ? node42523 : 4'b0010;
															assign node42523 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node42527 = (inp[5]) ? node42535 : node42528;
														assign node42528 = (inp[14]) ? node42532 : node42529;
															assign node42529 = (inp[7]) ? 4'b0011 : 4'b0010;
															assign node42532 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node42535 = (inp[14]) ? node42537 : 4'b0010;
															assign node42537 = (inp[7]) ? 4'b0011 : 4'b0010;
									assign node42540 = (inp[14]) ? node42612 : node42541;
										assign node42541 = (inp[10]) ? node42571 : node42542;
											assign node42542 = (inp[1]) ? node42562 : node42543;
												assign node42543 = (inp[11]) ? node42545 : 4'b0110;
													assign node42545 = (inp[0]) ? node42555 : node42546;
														assign node42546 = (inp[9]) ? node42548 : 4'b0110;
															assign node42548 = (inp[5]) ? node42552 : node42549;
																assign node42549 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node42552 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node42555 = (inp[7]) ? node42559 : node42556;
															assign node42556 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node42559 = (inp[9]) ? 4'b0110 : 4'b0111;
												assign node42562 = (inp[11]) ? node42564 : 4'b0111;
													assign node42564 = (inp[7]) ? node42568 : node42565;
														assign node42565 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node42568 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node42571 = (inp[1]) ? node42589 : node42572;
												assign node42572 = (inp[11]) ? node42574 : 4'b0111;
													assign node42574 = (inp[0]) ? node42582 : node42575;
														assign node42575 = (inp[7]) ? node42579 : node42576;
															assign node42576 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node42579 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node42582 = (inp[7]) ? node42586 : node42583;
															assign node42583 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node42586 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node42589 = (inp[11]) ? node42591 : 4'b0110;
													assign node42591 = (inp[0]) ? node42603 : node42592;
														assign node42592 = (inp[9]) ? node42598 : node42593;
															assign node42593 = (inp[7]) ? node42595 : 4'b0111;
																assign node42595 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node42598 = (inp[5]) ? 4'b0111 : node42599;
																assign node42599 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node42603 = (inp[9]) ? node42609 : node42604;
															assign node42604 = (inp[7]) ? 4'b0110 : node42605;
																assign node42605 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node42609 = (inp[5]) ? 4'b0110 : 4'b0111;
										assign node42612 = (inp[11]) ? node42672 : node42613;
											assign node42613 = (inp[7]) ? node42643 : node42614;
												assign node42614 = (inp[5]) ? node42630 : node42615;
													assign node42615 = (inp[9]) ? node42623 : node42616;
														assign node42616 = (inp[1]) ? node42620 : node42617;
															assign node42617 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node42620 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node42623 = (inp[10]) ? node42627 : node42624;
															assign node42624 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node42627 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node42630 = (inp[0]) ? node42638 : node42631;
														assign node42631 = (inp[1]) ? node42635 : node42632;
															assign node42632 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node42635 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node42638 = (inp[10]) ? 4'b0110 : node42639;
															assign node42639 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node42643 = (inp[5]) ? node42661 : node42644;
													assign node42644 = (inp[0]) ? node42654 : node42645;
														assign node42645 = (inp[9]) ? node42647 : 4'b0110;
															assign node42647 = (inp[10]) ? node42651 : node42648;
																assign node42648 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node42651 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node42654 = (inp[10]) ? node42658 : node42655;
															assign node42655 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node42658 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node42661 = (inp[9]) ? node42667 : node42662;
														assign node42662 = (inp[1]) ? node42664 : 4'b0111;
															assign node42664 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node42667 = (inp[10]) ? 4'b0111 : node42668;
															assign node42668 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node42672 = (inp[9]) ? node42712 : node42673;
												assign node42673 = (inp[0]) ? node42695 : node42674;
													assign node42674 = (inp[1]) ? node42686 : node42675;
														assign node42675 = (inp[10]) ? node42681 : node42676;
															assign node42676 = (inp[5]) ? 4'b0110 : node42677;
																assign node42677 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node42681 = (inp[7]) ? 4'b0111 : node42682;
																assign node42682 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node42686 = (inp[10]) ? node42690 : node42687;
															assign node42687 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node42690 = (inp[5]) ? 4'b0110 : node42691;
																assign node42691 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node42695 = (inp[1]) ? node42703 : node42696;
														assign node42696 = (inp[10]) ? node42700 : node42697;
															assign node42697 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node42700 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node42703 = (inp[10]) ? node42709 : node42704;
															assign node42704 = (inp[7]) ? 4'b0111 : node42705;
																assign node42705 = (inp[5]) ? 4'b0111 : 4'b0110;
															assign node42709 = (inp[5]) ? 4'b0110 : 4'b0111;
												assign node42712 = (inp[7]) ? node42732 : node42713;
													assign node42713 = (inp[0]) ? node42719 : node42714;
														assign node42714 = (inp[5]) ? node42716 : 4'b0111;
															assign node42716 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node42719 = (inp[5]) ? node42727 : node42720;
															assign node42720 = (inp[10]) ? node42724 : node42721;
																assign node42721 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node42724 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node42727 = (inp[10]) ? node42729 : 4'b0111;
																assign node42729 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node42732 = (inp[5]) ? node42740 : node42733;
														assign node42733 = (inp[1]) ? node42737 : node42734;
															assign node42734 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node42737 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node42740 = (inp[0]) ? node42744 : node42741;
															assign node42741 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node42744 = (inp[1]) ? node42746 : 4'b0111;
																assign node42746 = (inp[10]) ? 4'b0110 : 4'b0111;
								assign node42749 = (inp[4]) ? node42863 : node42750;
									assign node42750 = (inp[7]) ? node42782 : node42751;
										assign node42751 = (inp[11]) ? node42775 : node42752;
											assign node42752 = (inp[10]) ? node42764 : node42753;
												assign node42753 = (inp[1]) ? node42759 : node42754;
													assign node42754 = (inp[14]) ? node42756 : 4'b0110;
														assign node42756 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node42759 = (inp[5]) ? node42761 : 4'b0111;
														assign node42761 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node42764 = (inp[1]) ? node42770 : node42765;
													assign node42765 = (inp[14]) ? node42767 : 4'b0111;
														assign node42767 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node42770 = (inp[14]) ? node42772 : 4'b0110;
														assign node42772 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node42775 = (inp[10]) ? node42779 : node42776;
												assign node42776 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node42779 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node42782 = (inp[1]) ? node42824 : node42783;
											assign node42783 = (inp[10]) ? node42797 : node42784;
												assign node42784 = (inp[5]) ? node42792 : node42785;
													assign node42785 = (inp[11]) ? node42789 : node42786;
														assign node42786 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node42789 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node42792 = (inp[11]) ? 4'b0110 : node42793;
														assign node42793 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node42797 = (inp[14]) ? node42819 : node42798;
													assign node42798 = (inp[0]) ? node42806 : node42799;
														assign node42799 = (inp[5]) ? node42803 : node42800;
															assign node42800 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node42803 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node42806 = (inp[9]) ? node42812 : node42807;
															assign node42807 = (inp[11]) ? 4'b0110 : node42808;
																assign node42808 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node42812 = (inp[11]) ? node42816 : node42813;
																assign node42813 = (inp[5]) ? 4'b0110 : 4'b0111;
																assign node42816 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node42819 = (inp[5]) ? 4'b0111 : node42820;
														assign node42820 = (inp[11]) ? 4'b0111 : 4'b0110;
											assign node42824 = (inp[10]) ? node42850 : node42825;
												assign node42825 = (inp[11]) ? node42845 : node42826;
													assign node42826 = (inp[9]) ? node42838 : node42827;
														assign node42827 = (inp[0]) ? node42833 : node42828;
															assign node42828 = (inp[5]) ? 4'b0111 : node42829;
																assign node42829 = (inp[14]) ? 4'b0110 : 4'b0111;
															assign node42833 = (inp[5]) ? 4'b0110 : node42834;
																assign node42834 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node42838 = (inp[14]) ? node42842 : node42839;
															assign node42839 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node42842 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node42845 = (inp[14]) ? 4'b0111 : node42846;
														assign node42846 = (inp[5]) ? 4'b0111 : 4'b0110;
												assign node42850 = (inp[14]) ? node42858 : node42851;
													assign node42851 = (inp[11]) ? node42855 : node42852;
														assign node42852 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node42855 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node42858 = (inp[11]) ? 4'b0110 : node42859;
														assign node42859 = (inp[5]) ? 4'b0110 : 4'b0111;
									assign node42863 = (inp[7]) ? node42991 : node42864;
										assign node42864 = (inp[14]) ? node42918 : node42865;
											assign node42865 = (inp[5]) ? node42901 : node42866;
												assign node42866 = (inp[9]) ? node42878 : node42867;
													assign node42867 = (inp[11]) ? node42873 : node42868;
														assign node42868 = (inp[10]) ? 4'b0010 : node42869;
															assign node42869 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node42873 = (inp[1]) ? 4'b0011 : node42874;
															assign node42874 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node42878 = (inp[1]) ? node42886 : node42879;
														assign node42879 = (inp[11]) ? node42883 : node42880;
															assign node42880 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node42883 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node42886 = (inp[0]) ? node42894 : node42887;
															assign node42887 = (inp[11]) ? node42891 : node42888;
																assign node42888 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node42891 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node42894 = (inp[11]) ? node42898 : node42895;
																assign node42895 = (inp[10]) ? 4'b0011 : 4'b0010;
																assign node42898 = (inp[10]) ? 4'b0010 : 4'b0011;
												assign node42901 = (inp[11]) ? node42911 : node42902;
													assign node42902 = (inp[0]) ? node42904 : 4'b0011;
														assign node42904 = (inp[1]) ? node42908 : node42905;
															assign node42905 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node42908 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node42911 = (inp[1]) ? node42915 : node42912;
														assign node42912 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node42915 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node42918 = (inp[10]) ? node42962 : node42919;
												assign node42919 = (inp[0]) ? node42935 : node42920;
													assign node42920 = (inp[1]) ? node42928 : node42921;
														assign node42921 = (inp[11]) ? node42925 : node42922;
															assign node42922 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node42925 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node42928 = (inp[5]) ? node42932 : node42929;
															assign node42929 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node42932 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node42935 = (inp[9]) ? node42949 : node42936;
														assign node42936 = (inp[5]) ? node42942 : node42937;
															assign node42937 = (inp[11]) ? 4'b0011 : node42938;
																assign node42938 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node42942 = (inp[1]) ? node42946 : node42943;
																assign node42943 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node42946 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node42949 = (inp[5]) ? node42955 : node42950;
															assign node42950 = (inp[11]) ? 4'b0010 : node42951;
																assign node42951 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node42955 = (inp[1]) ? node42959 : node42956;
																assign node42956 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node42959 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node42962 = (inp[0]) ? node42974 : node42963;
													assign node42963 = (inp[1]) ? node42969 : node42964;
														assign node42964 = (inp[11]) ? 4'b0011 : node42965;
															assign node42965 = (inp[5]) ? 4'b0010 : 4'b0011;
														assign node42969 = (inp[11]) ? 4'b0010 : node42970;
															assign node42970 = (inp[9]) ? 4'b0010 : 4'b0011;
													assign node42974 = (inp[1]) ? node42984 : node42975;
														assign node42975 = (inp[9]) ? node42977 : 4'b0010;
															assign node42977 = (inp[11]) ? node42981 : node42978;
																assign node42978 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node42981 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node42984 = (inp[11]) ? node42988 : node42985;
															assign node42985 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node42988 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node42991 = (inp[10]) ? node43007 : node42992;
											assign node42992 = (inp[1]) ? node43000 : node42993;
												assign node42993 = (inp[5]) ? node42995 : 4'b0010;
													assign node42995 = (inp[11]) ? 4'b0010 : node42996;
														assign node42996 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node43000 = (inp[5]) ? node43002 : 4'b0011;
													assign node43002 = (inp[11]) ? 4'b0011 : node43003;
														assign node43003 = (inp[14]) ? 4'b0011 : 4'b0010;
											assign node43007 = (inp[1]) ? node43015 : node43008;
												assign node43008 = (inp[11]) ? 4'b0011 : node43009;
													assign node43009 = (inp[14]) ? 4'b0011 : node43010;
														assign node43010 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node43015 = (inp[14]) ? 4'b0010 : node43016;
													assign node43016 = (inp[5]) ? node43018 : 4'b0010;
														assign node43018 = (inp[11]) ? 4'b0010 : 4'b0011;
							assign node43022 = (inp[4]) ? node43366 : node43023;
								assign node43023 = (inp[2]) ? node43151 : node43024;
									assign node43024 = (inp[10]) ? node43088 : node43025;
										assign node43025 = (inp[1]) ? node43055 : node43026;
											assign node43026 = (inp[11]) ? node43034 : node43027;
												assign node43027 = (inp[5]) ? node43029 : 4'b0010;
													assign node43029 = (inp[7]) ? node43031 : 4'b0010;
														assign node43031 = (inp[14]) ? 4'b0010 : 4'b0011;
												assign node43034 = (inp[14]) ? node43040 : node43035;
													assign node43035 = (inp[7]) ? node43037 : 4'b0010;
														assign node43037 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node43040 = (inp[0]) ? node43048 : node43041;
														assign node43041 = (inp[9]) ? 4'b0011 : node43042;
															assign node43042 = (inp[5]) ? node43044 : 4'b0010;
																assign node43044 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node43048 = (inp[5]) ? node43052 : node43049;
															assign node43049 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node43052 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node43055 = (inp[7]) ? node43063 : node43056;
												assign node43056 = (inp[14]) ? node43058 : 4'b0011;
													assign node43058 = (inp[5]) ? 4'b0011 : node43059;
														assign node43059 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node43063 = (inp[5]) ? node43069 : node43064;
													assign node43064 = (inp[14]) ? 4'b0011 : node43065;
														assign node43065 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node43069 = (inp[9]) ? node43083 : node43070;
														assign node43070 = (inp[0]) ? node43078 : node43071;
															assign node43071 = (inp[11]) ? node43075 : node43072;
																assign node43072 = (inp[14]) ? 4'b0011 : 4'b0010;
																assign node43075 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node43078 = (inp[11]) ? 4'b0011 : node43079;
																assign node43079 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node43083 = (inp[11]) ? node43085 : 4'b0010;
															assign node43085 = (inp[14]) ? 4'b0010 : 4'b0011;
										assign node43088 = (inp[1]) ? node43118 : node43089;
											assign node43089 = (inp[7]) ? node43097 : node43090;
												assign node43090 = (inp[11]) ? node43092 : 4'b0011;
													assign node43092 = (inp[14]) ? node43094 : 4'b0011;
														assign node43094 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node43097 = (inp[14]) ? node43113 : node43098;
													assign node43098 = (inp[0]) ? node43106 : node43099;
														assign node43099 = (inp[5]) ? node43103 : node43100;
															assign node43100 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node43103 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node43106 = (inp[11]) ? node43110 : node43107;
															assign node43107 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node43110 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node43113 = (inp[5]) ? node43115 : 4'b0011;
														assign node43115 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node43118 = (inp[7]) ? node43126 : node43119;
												assign node43119 = (inp[14]) ? node43121 : 4'b0010;
													assign node43121 = (inp[11]) ? node43123 : 4'b0010;
														assign node43123 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node43126 = (inp[5]) ? node43132 : node43127;
													assign node43127 = (inp[11]) ? node43129 : 4'b0010;
														assign node43129 = (inp[14]) ? 4'b0010 : 4'b0011;
													assign node43132 = (inp[0]) ? node43146 : node43133;
														assign node43133 = (inp[9]) ? node43141 : node43134;
															assign node43134 = (inp[14]) ? node43138 : node43135;
																assign node43135 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node43138 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node43141 = (inp[14]) ? 4'b0010 : node43142;
																assign node43142 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node43146 = (inp[11]) ? node43148 : 4'b0011;
															assign node43148 = (inp[9]) ? 4'b0011 : 4'b0010;
									assign node43151 = (inp[0]) ? node43257 : node43152;
										assign node43152 = (inp[14]) ? node43190 : node43153;
											assign node43153 = (inp[1]) ? node43173 : node43154;
												assign node43154 = (inp[10]) ? node43166 : node43155;
													assign node43155 = (inp[7]) ? node43157 : 4'b0110;
														assign node43157 = (inp[9]) ? node43161 : node43158;
															assign node43158 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node43161 = (inp[5]) ? node43163 : 4'b0110;
																assign node43163 = (inp[11]) ? 4'b0110 : 4'b0111;
													assign node43166 = (inp[7]) ? node43168 : 4'b0111;
														assign node43168 = (inp[5]) ? node43170 : 4'b0110;
															assign node43170 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node43173 = (inp[10]) ? node43183 : node43174;
													assign node43174 = (inp[7]) ? node43176 : 4'b0111;
														assign node43176 = (inp[11]) ? node43180 : node43177;
															assign node43177 = (inp[5]) ? 4'b0110 : 4'b0111;
															assign node43180 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node43183 = (inp[7]) ? node43185 : 4'b0110;
														assign node43185 = (inp[11]) ? 4'b0110 : node43186;
															assign node43186 = (inp[5]) ? 4'b0111 : 4'b0110;
											assign node43190 = (inp[5]) ? node43230 : node43191;
												assign node43191 = (inp[9]) ? node43213 : node43192;
													assign node43192 = (inp[11]) ? node43206 : node43193;
														assign node43193 = (inp[10]) ? node43201 : node43194;
															assign node43194 = (inp[1]) ? node43198 : node43195;
																assign node43195 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node43198 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node43201 = (inp[1]) ? 4'b0111 : node43202;
																assign node43202 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node43206 = (inp[10]) ? node43210 : node43207;
															assign node43207 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node43210 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node43213 = (inp[10]) ? node43223 : node43214;
														assign node43214 = (inp[1]) ? node43220 : node43215;
															assign node43215 = (inp[7]) ? node43217 : 4'b0110;
																assign node43217 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node43220 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node43223 = (inp[1]) ? node43227 : node43224;
															assign node43224 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node43227 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node43230 = (inp[11]) ? node43240 : node43231;
													assign node43231 = (inp[7]) ? node43233 : 4'b0110;
														assign node43233 = (inp[10]) ? node43237 : node43234;
															assign node43234 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node43237 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node43240 = (inp[7]) ? node43248 : node43241;
														assign node43241 = (inp[10]) ? node43245 : node43242;
															assign node43242 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node43245 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node43248 = (inp[9]) ? node43254 : node43249;
															assign node43249 = (inp[10]) ? node43251 : 4'b0110;
																assign node43251 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node43254 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node43257 = (inp[5]) ? node43329 : node43258;
											assign node43258 = (inp[11]) ? node43298 : node43259;
												assign node43259 = (inp[14]) ? node43279 : node43260;
													assign node43260 = (inp[7]) ? node43266 : node43261;
														assign node43261 = (inp[10]) ? 4'b0110 : node43262;
															assign node43262 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node43266 = (inp[9]) ? node43272 : node43267;
															assign node43267 = (inp[1]) ? node43269 : 4'b0111;
																assign node43269 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node43272 = (inp[1]) ? node43276 : node43273;
																assign node43273 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node43276 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node43279 = (inp[7]) ? node43287 : node43280;
														assign node43280 = (inp[10]) ? node43284 : node43281;
															assign node43281 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node43284 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node43287 = (inp[9]) ? node43293 : node43288;
															assign node43288 = (inp[10]) ? node43290 : 4'b0110;
																assign node43290 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node43293 = (inp[10]) ? 4'b0111 : node43294;
																assign node43294 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node43298 = (inp[14]) ? node43314 : node43299;
													assign node43299 = (inp[1]) ? node43307 : node43300;
														assign node43300 = (inp[7]) ? node43304 : node43301;
															assign node43301 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node43304 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node43307 = (inp[7]) ? node43311 : node43308;
															assign node43308 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node43311 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node43314 = (inp[9]) ? node43322 : node43315;
														assign node43315 = (inp[1]) ? node43319 : node43316;
															assign node43316 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node43319 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node43322 = (inp[1]) ? node43326 : node43323;
															assign node43323 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node43326 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node43329 = (inp[11]) ? node43359 : node43330;
												assign node43330 = (inp[1]) ? node43344 : node43331;
													assign node43331 = (inp[9]) ? node43333 : 4'b0111;
														assign node43333 = (inp[14]) ? node43339 : node43334;
															assign node43334 = (inp[10]) ? node43336 : 4'b0111;
																assign node43336 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node43339 = (inp[10]) ? node43341 : 4'b0110;
																assign node43341 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node43344 = (inp[14]) ? node43352 : node43345;
														assign node43345 = (inp[7]) ? node43349 : node43346;
															assign node43346 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node43349 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node43352 = (inp[10]) ? node43356 : node43353;
															assign node43353 = (inp[7]) ? 4'b0111 : 4'b0110;
															assign node43356 = (inp[7]) ? 4'b0110 : 4'b0111;
												assign node43359 = (inp[10]) ? node43363 : node43360;
													assign node43360 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node43363 = (inp[1]) ? 4'b0110 : 4'b0111;
								assign node43366 = (inp[2]) ? node43566 : node43367;
									assign node43367 = (inp[11]) ? node43445 : node43368;
										assign node43368 = (inp[5]) ? node43376 : node43369;
											assign node43369 = (inp[1]) ? node43373 : node43370;
												assign node43370 = (inp[10]) ? 4'b0111 : 4'b0110;
												assign node43373 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node43376 = (inp[14]) ? node43400 : node43377;
												assign node43377 = (inp[7]) ? node43387 : node43378;
													assign node43378 = (inp[9]) ? 4'b0110 : node43379;
														assign node43379 = (inp[0]) ? node43381 : 4'b0111;
															assign node43381 = (inp[10]) ? 4'b0110 : node43382;
																assign node43382 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node43387 = (inp[9]) ? node43393 : node43388;
														assign node43388 = (inp[10]) ? node43390 : 4'b0110;
															assign node43390 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node43393 = (inp[10]) ? node43397 : node43394;
															assign node43394 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node43397 = (inp[1]) ? 4'b0110 : 4'b0111;
												assign node43400 = (inp[9]) ? node43424 : node43401;
													assign node43401 = (inp[0]) ? node43417 : node43402;
														assign node43402 = (inp[7]) ? node43410 : node43403;
															assign node43403 = (inp[10]) ? node43407 : node43404;
																assign node43404 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node43407 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node43410 = (inp[1]) ? node43414 : node43411;
																assign node43411 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node43414 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node43417 = (inp[7]) ? node43419 : 4'b0110;
															assign node43419 = (inp[1]) ? 4'b0110 : node43420;
																assign node43420 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node43424 = (inp[7]) ? node43432 : node43425;
														assign node43425 = (inp[10]) ? node43429 : node43426;
															assign node43426 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node43429 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node43432 = (inp[0]) ? node43438 : node43433;
															assign node43433 = (inp[10]) ? node43435 : 4'b0110;
																assign node43435 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node43438 = (inp[10]) ? node43442 : node43439;
																assign node43439 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node43442 = (inp[1]) ? 4'b0110 : 4'b0111;
										assign node43445 = (inp[0]) ? node43505 : node43446;
											assign node43446 = (inp[5]) ? node43486 : node43447;
												assign node43447 = (inp[9]) ? node43463 : node43448;
													assign node43448 = (inp[10]) ? 4'b0111 : node43449;
														assign node43449 = (inp[1]) ? node43457 : node43450;
															assign node43450 = (inp[14]) ? node43454 : node43451;
																assign node43451 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node43454 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node43457 = (inp[14]) ? node43459 : 4'b0111;
																assign node43459 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node43463 = (inp[1]) ? node43473 : node43464;
														assign node43464 = (inp[7]) ? 4'b0110 : node43465;
															assign node43465 = (inp[10]) ? node43469 : node43466;
																assign node43466 = (inp[14]) ? 4'b0111 : 4'b0110;
																assign node43469 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node43473 = (inp[7]) ? node43481 : node43474;
															assign node43474 = (inp[10]) ? node43478 : node43475;
																assign node43475 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node43478 = (inp[14]) ? 4'b0111 : 4'b0110;
															assign node43481 = (inp[10]) ? node43483 : 4'b0111;
																assign node43483 = (inp[14]) ? 4'b0110 : 4'b0111;
												assign node43486 = (inp[1]) ? node43494 : node43487;
													assign node43487 = (inp[10]) ? 4'b0111 : node43488;
														assign node43488 = (inp[7]) ? 4'b0110 : node43489;
															assign node43489 = (inp[14]) ? 4'b0110 : 4'b0111;
													assign node43494 = (inp[10]) ? node43500 : node43495;
														assign node43495 = (inp[14]) ? 4'b0111 : node43496;
															assign node43496 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node43500 = (inp[14]) ? 4'b0110 : node43501;
															assign node43501 = (inp[9]) ? 4'b0110 : 4'b0111;
											assign node43505 = (inp[7]) ? node43543 : node43506;
												assign node43506 = (inp[9]) ? node43524 : node43507;
													assign node43507 = (inp[10]) ? node43517 : node43508;
														assign node43508 = (inp[5]) ? 4'b0110 : node43509;
															assign node43509 = (inp[1]) ? node43513 : node43510;
																assign node43510 = (inp[14]) ? 4'b0111 : 4'b0110;
																assign node43513 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node43517 = (inp[5]) ? node43519 : 4'b0110;
															assign node43519 = (inp[14]) ? node43521 : 4'b0111;
																assign node43521 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node43524 = (inp[5]) ? node43534 : node43525;
														assign node43525 = (inp[10]) ? 4'b0110 : node43526;
															assign node43526 = (inp[1]) ? node43530 : node43527;
																assign node43527 = (inp[14]) ? 4'b0111 : 4'b0110;
																assign node43530 = (inp[14]) ? 4'b0110 : 4'b0111;
														assign node43534 = (inp[1]) ? 4'b0111 : node43535;
															assign node43535 = (inp[10]) ? node43539 : node43536;
																assign node43536 = (inp[14]) ? 4'b0110 : 4'b0111;
																assign node43539 = (inp[14]) ? 4'b0111 : 4'b0110;
												assign node43543 = (inp[1]) ? node43555 : node43544;
													assign node43544 = (inp[10]) ? node43550 : node43545;
														assign node43545 = (inp[14]) ? 4'b0110 : node43546;
															assign node43546 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node43550 = (inp[14]) ? 4'b0111 : node43551;
															assign node43551 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node43555 = (inp[10]) ? node43561 : node43556;
														assign node43556 = (inp[5]) ? 4'b0111 : node43557;
															assign node43557 = (inp[14]) ? 4'b0111 : 4'b0110;
														assign node43561 = (inp[14]) ? 4'b0110 : node43562;
															assign node43562 = (inp[5]) ? 4'b0110 : 4'b0111;
									assign node43566 = (inp[10]) ? node43620 : node43567;
										assign node43567 = (inp[1]) ? node43599 : node43568;
											assign node43568 = (inp[7]) ? node43592 : node43569;
												assign node43569 = (inp[14]) ? node43577 : node43570;
													assign node43570 = (inp[9]) ? 4'b0010 : node43571;
														assign node43571 = (inp[11]) ? 4'b0010 : node43572;
															assign node43572 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node43577 = (inp[9]) ? node43585 : node43578;
														assign node43578 = (inp[5]) ? node43582 : node43579;
															assign node43579 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node43582 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node43585 = (inp[11]) ? node43589 : node43586;
															assign node43586 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node43589 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node43592 = (inp[5]) ? node43594 : 4'b0010;
													assign node43594 = (inp[14]) ? 4'b0010 : node43595;
														assign node43595 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node43599 = (inp[11]) ? node43613 : node43600;
												assign node43600 = (inp[14]) ? node43608 : node43601;
													assign node43601 = (inp[7]) ? node43605 : node43602;
														assign node43602 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node43605 = (inp[5]) ? 4'b0010 : 4'b0011;
													assign node43608 = (inp[5]) ? node43610 : 4'b0011;
														assign node43610 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node43613 = (inp[14]) ? node43615 : 4'b0011;
													assign node43615 = (inp[7]) ? 4'b0011 : node43616;
														assign node43616 = (inp[5]) ? 4'b0011 : 4'b0010;
										assign node43620 = (inp[1]) ? node43658 : node43621;
											assign node43621 = (inp[7]) ? node43651 : node43622;
												assign node43622 = (inp[14]) ? node43628 : node43623;
													assign node43623 = (inp[11]) ? 4'b0011 : node43624;
														assign node43624 = (inp[5]) ? 4'b0011 : 4'b0010;
													assign node43628 = (inp[9]) ? node43644 : node43629;
														assign node43629 = (inp[0]) ? node43637 : node43630;
															assign node43630 = (inp[11]) ? node43634 : node43631;
																assign node43631 = (inp[5]) ? 4'b0010 : 4'b0011;
																assign node43634 = (inp[5]) ? 4'b0011 : 4'b0010;
															assign node43637 = (inp[5]) ? node43641 : node43638;
																assign node43638 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node43641 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node43644 = (inp[11]) ? node43648 : node43645;
															assign node43645 = (inp[5]) ? 4'b0010 : 4'b0011;
															assign node43648 = (inp[5]) ? 4'b0011 : 4'b0010;
												assign node43651 = (inp[11]) ? 4'b0011 : node43652;
													assign node43652 = (inp[14]) ? 4'b0011 : node43653;
														assign node43653 = (inp[5]) ? 4'b0010 : 4'b0011;
											assign node43658 = (inp[7]) ? node43682 : node43659;
												assign node43659 = (inp[5]) ? node43677 : node43660;
													assign node43660 = (inp[9]) ? node43668 : node43661;
														assign node43661 = (inp[11]) ? node43665 : node43662;
															assign node43662 = (inp[14]) ? 4'b0010 : 4'b0011;
															assign node43665 = (inp[14]) ? 4'b0011 : 4'b0010;
														assign node43668 = (inp[0]) ? node43670 : 4'b0011;
															assign node43670 = (inp[14]) ? node43674 : node43671;
																assign node43671 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node43674 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node43677 = (inp[14]) ? node43679 : 4'b0010;
														assign node43679 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node43682 = (inp[11]) ? 4'b0010 : node43683;
													assign node43683 = (inp[14]) ? 4'b0010 : node43684;
														assign node43684 = (inp[5]) ? 4'b0011 : 4'b0010;
					assign node43689 = (inp[15]) ? node44523 : node43690;
						assign node43690 = (inp[14]) ? node44280 : node43691;
							assign node43691 = (inp[4]) ? node43861 : node43692;
								assign node43692 = (inp[5]) ? node43740 : node43693;
									assign node43693 = (inp[7]) ? node43717 : node43694;
										assign node43694 = (inp[1]) ? node43702 : node43695;
											assign node43695 = (inp[13]) ? node43699 : node43696;
												assign node43696 = (inp[11]) ? 4'b0011 : 4'b0010;
												assign node43699 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node43702 = (inp[11]) ? node43710 : node43703;
												assign node43703 = (inp[13]) ? node43707 : node43704;
													assign node43704 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node43707 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node43710 = (inp[13]) ? node43714 : node43711;
													assign node43711 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node43714 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node43717 = (inp[13]) ? node43729 : node43718;
											assign node43718 = (inp[11]) ? node43724 : node43719;
												assign node43719 = (inp[2]) ? node43721 : 4'b0110;
													assign node43721 = (inp[1]) ? 4'b0111 : 4'b0110;
												assign node43724 = (inp[2]) ? node43726 : 4'b0111;
													assign node43726 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node43729 = (inp[11]) ? node43735 : node43730;
												assign node43730 = (inp[1]) ? node43732 : 4'b0111;
													assign node43732 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node43735 = (inp[2]) ? node43737 : 4'b0110;
													assign node43737 = (inp[1]) ? 4'b0111 : 4'b0110;
									assign node43740 = (inp[7]) ? node43838 : node43741;
										assign node43741 = (inp[10]) ? node43795 : node43742;
											assign node43742 = (inp[2]) ? node43780 : node43743;
												assign node43743 = (inp[9]) ? node43761 : node43744;
													assign node43744 = (inp[1]) ? node43754 : node43745;
														assign node43745 = (inp[0]) ? node43751 : node43746;
															assign node43746 = (inp[11]) ? node43748 : 4'b0110;
																assign node43748 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node43751 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node43754 = (inp[11]) ? node43758 : node43755;
															assign node43755 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node43758 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node43761 = (inp[1]) ? node43767 : node43762;
														assign node43762 = (inp[0]) ? node43764 : 4'b0111;
															assign node43764 = (inp[11]) ? 4'b0111 : 4'b0110;
														assign node43767 = (inp[0]) ? node43773 : node43768;
															assign node43768 = (inp[11]) ? 4'b0110 : node43769;
																assign node43769 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node43773 = (inp[11]) ? node43777 : node43774;
																assign node43774 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node43777 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node43780 = (inp[11]) ? node43788 : node43781;
													assign node43781 = (inp[1]) ? node43785 : node43782;
														assign node43782 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node43785 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node43788 = (inp[13]) ? node43792 : node43789;
														assign node43789 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node43792 = (inp[1]) ? 4'b0111 : 4'b0110;
											assign node43795 = (inp[1]) ? node43803 : node43796;
												assign node43796 = (inp[11]) ? node43800 : node43797;
													assign node43797 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node43800 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node43803 = (inp[9]) ? node43829 : node43804;
													assign node43804 = (inp[0]) ? node43820 : node43805;
														assign node43805 = (inp[2]) ? node43813 : node43806;
															assign node43806 = (inp[11]) ? node43810 : node43807;
																assign node43807 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node43810 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node43813 = (inp[11]) ? node43817 : node43814;
																assign node43814 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node43817 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node43820 = (inp[13]) ? node43822 : 4'b0111;
															assign node43822 = (inp[2]) ? node43826 : node43823;
																assign node43823 = (inp[11]) ? 4'b0110 : 4'b0111;
																assign node43826 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node43829 = (inp[13]) ? 4'b0111 : node43830;
														assign node43830 = (inp[11]) ? node43834 : node43831;
															assign node43831 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node43834 = (inp[2]) ? 4'b0110 : 4'b0111;
										assign node43838 = (inp[13]) ? node43850 : node43839;
											assign node43839 = (inp[11]) ? node43845 : node43840;
												assign node43840 = (inp[2]) ? 4'b0010 : node43841;
													assign node43841 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node43845 = (inp[2]) ? 4'b0011 : node43846;
													assign node43846 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node43850 = (inp[11]) ? node43856 : node43851;
												assign node43851 = (inp[1]) ? 4'b0011 : node43852;
													assign node43852 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node43856 = (inp[2]) ? 4'b0010 : node43857;
													assign node43857 = (inp[1]) ? 4'b0010 : 4'b0011;
								assign node43861 = (inp[1]) ? node44103 : node43862;
									assign node43862 = (inp[7]) ? node43966 : node43863;
										assign node43863 = (inp[5]) ? node43925 : node43864;
											assign node43864 = (inp[13]) ? node43888 : node43865;
												assign node43865 = (inp[9]) ? node43881 : node43866;
													assign node43866 = (inp[10]) ? node43874 : node43867;
														assign node43867 = (inp[11]) ? node43871 : node43868;
															assign node43868 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node43871 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node43874 = (inp[2]) ? node43878 : node43875;
															assign node43875 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node43878 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node43881 = (inp[11]) ? node43885 : node43882;
														assign node43882 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node43885 = (inp[2]) ? 4'b0010 : 4'b0011;
												assign node43888 = (inp[9]) ? node43912 : node43889;
													assign node43889 = (inp[0]) ? node43899 : node43890;
														assign node43890 = (inp[10]) ? 4'b0010 : node43891;
															assign node43891 = (inp[2]) ? node43895 : node43892;
																assign node43892 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node43895 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node43899 = (inp[10]) ? node43905 : node43900;
															assign node43900 = (inp[2]) ? node43902 : 4'b0011;
																assign node43902 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node43905 = (inp[11]) ? node43909 : node43906;
																assign node43906 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node43909 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node43912 = (inp[0]) ? node43918 : node43913;
														assign node43913 = (inp[11]) ? 4'b0011 : node43914;
															assign node43914 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node43918 = (inp[11]) ? node43922 : node43919;
															assign node43919 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node43922 = (inp[2]) ? 4'b0011 : 4'b0010;
											assign node43925 = (inp[9]) ? node43959 : node43926;
												assign node43926 = (inp[2]) ? node43942 : node43927;
													assign node43927 = (inp[0]) ? node43935 : node43928;
														assign node43928 = (inp[11]) ? node43932 : node43929;
															assign node43929 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node43932 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node43935 = (inp[11]) ? node43939 : node43936;
															assign node43936 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node43939 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node43942 = (inp[0]) ? node43948 : node43943;
														assign node43943 = (inp[10]) ? 4'b0111 : node43944;
															assign node43944 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node43948 = (inp[10]) ? node43954 : node43949;
															assign node43949 = (inp[13]) ? 4'b0111 : node43950;
																assign node43950 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node43954 = (inp[11]) ? node43956 : 4'b0110;
																assign node43956 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node43959 = (inp[13]) ? node43963 : node43960;
													assign node43960 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node43963 = (inp[11]) ? 4'b0110 : 4'b0111;
										assign node43966 = (inp[5]) ? node44024 : node43967;
											assign node43967 = (inp[0]) ? node43983 : node43968;
												assign node43968 = (inp[13]) ? node43976 : node43969;
													assign node43969 = (inp[11]) ? node43973 : node43970;
														assign node43970 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node43973 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node43976 = (inp[2]) ? node43980 : node43977;
														assign node43977 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node43980 = (inp[11]) ? 4'b0111 : 4'b0110;
												assign node43983 = (inp[11]) ? node44009 : node43984;
													assign node43984 = (inp[10]) ? node43994 : node43985;
														assign node43985 = (inp[9]) ? node43991 : node43986;
															assign node43986 = (inp[2]) ? 4'b0110 : node43987;
																assign node43987 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node43991 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node43994 = (inp[9]) ? node44002 : node43995;
															assign node43995 = (inp[13]) ? node43999 : node43996;
																assign node43996 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node43999 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node44002 = (inp[2]) ? node44006 : node44003;
																assign node44003 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node44006 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node44009 = (inp[10]) ? node44017 : node44010;
														assign node44010 = (inp[2]) ? node44014 : node44011;
															assign node44011 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node44014 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node44017 = (inp[2]) ? node44021 : node44018;
															assign node44018 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node44021 = (inp[13]) ? 4'b0111 : 4'b0110;
											assign node44024 = (inp[10]) ? node44060 : node44025;
												assign node44025 = (inp[0]) ? node44047 : node44026;
													assign node44026 = (inp[9]) ? node44032 : node44027;
														assign node44027 = (inp[13]) ? 4'b0010 : node44028;
															assign node44028 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node44032 = (inp[2]) ? node44040 : node44033;
															assign node44033 = (inp[11]) ? node44037 : node44034;
																assign node44034 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node44037 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node44040 = (inp[11]) ? node44044 : node44041;
																assign node44041 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node44044 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node44047 = (inp[11]) ? node44055 : node44048;
														assign node44048 = (inp[13]) ? node44052 : node44049;
															assign node44049 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node44052 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node44055 = (inp[2]) ? 4'b0011 : node44056;
															assign node44056 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node44060 = (inp[9]) ? node44078 : node44061;
													assign node44061 = (inp[0]) ? 4'b0010 : node44062;
														assign node44062 = (inp[11]) ? node44070 : node44063;
															assign node44063 = (inp[13]) ? node44067 : node44064;
																assign node44064 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node44067 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node44070 = (inp[13]) ? node44074 : node44071;
																assign node44071 = (inp[2]) ? 4'b0010 : 4'b0011;
																assign node44074 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node44078 = (inp[0]) ? node44088 : node44079;
														assign node44079 = (inp[13]) ? node44081 : 4'b0010;
															assign node44081 = (inp[2]) ? node44085 : node44082;
																assign node44082 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node44085 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node44088 = (inp[2]) ? node44096 : node44089;
															assign node44089 = (inp[13]) ? node44093 : node44090;
																assign node44090 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node44093 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node44096 = (inp[11]) ? node44100 : node44097;
																assign node44097 = (inp[13]) ? 4'b0010 : 4'b0011;
																assign node44100 = (inp[13]) ? 4'b0011 : 4'b0010;
									assign node44103 = (inp[0]) ? node44189 : node44104;
										assign node44104 = (inp[7]) ? node44148 : node44105;
											assign node44105 = (inp[5]) ? node44113 : node44106;
												assign node44106 = (inp[11]) ? node44110 : node44107;
													assign node44107 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node44110 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node44113 = (inp[2]) ? node44129 : node44114;
													assign node44114 = (inp[9]) ? node44122 : node44115;
														assign node44115 = (inp[11]) ? node44119 : node44116;
															assign node44116 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node44119 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node44122 = (inp[11]) ? node44126 : node44123;
															assign node44123 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node44126 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node44129 = (inp[10]) ? node44135 : node44130;
														assign node44130 = (inp[11]) ? node44132 : 4'b0110;
															assign node44132 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node44135 = (inp[9]) ? node44141 : node44136;
															assign node44136 = (inp[13]) ? node44138 : 4'b0110;
																assign node44138 = (inp[11]) ? 4'b0110 : 4'b0111;
															assign node44141 = (inp[11]) ? node44145 : node44142;
																assign node44142 = (inp[13]) ? 4'b0111 : 4'b0110;
																assign node44145 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node44148 = (inp[5]) ? node44174 : node44149;
												assign node44149 = (inp[2]) ? node44157 : node44150;
													assign node44150 = (inp[11]) ? node44154 : node44151;
														assign node44151 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node44154 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node44157 = (inp[9]) ? node44165 : node44158;
														assign node44158 = (inp[11]) ? node44162 : node44159;
															assign node44159 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node44162 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node44165 = (inp[10]) ? node44167 : 4'b0111;
															assign node44167 = (inp[13]) ? node44171 : node44168;
																assign node44168 = (inp[11]) ? 4'b0111 : 4'b0110;
																assign node44171 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node44174 = (inp[9]) ? node44182 : node44175;
													assign node44175 = (inp[11]) ? node44179 : node44176;
														assign node44176 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node44179 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node44182 = (inp[13]) ? node44186 : node44183;
														assign node44183 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node44186 = (inp[11]) ? 4'b0010 : 4'b0011;
										assign node44189 = (inp[2]) ? node44229 : node44190;
											assign node44190 = (inp[5]) ? node44216 : node44191;
												assign node44191 = (inp[7]) ? node44199 : node44192;
													assign node44192 = (inp[11]) ? node44196 : node44193;
														assign node44193 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node44196 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node44199 = (inp[9]) ? node44207 : node44200;
														assign node44200 = (inp[13]) ? node44204 : node44201;
															assign node44201 = (inp[11]) ? 4'b0111 : 4'b0110;
															assign node44204 = (inp[11]) ? 4'b0110 : 4'b0111;
														assign node44207 = (inp[10]) ? node44211 : node44208;
															assign node44208 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node44211 = (inp[13]) ? node44213 : 4'b0111;
																assign node44213 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node44216 = (inp[7]) ? node44222 : node44217;
													assign node44217 = (inp[13]) ? node44219 : 4'b0110;
														assign node44219 = (inp[11]) ? 4'b0111 : 4'b0110;
													assign node44222 = (inp[11]) ? node44226 : node44223;
														assign node44223 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node44226 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node44229 = (inp[5]) ? node44251 : node44230;
												assign node44230 = (inp[7]) ? node44238 : node44231;
													assign node44231 = (inp[11]) ? node44235 : node44232;
														assign node44232 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node44235 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node44238 = (inp[10]) ? node44246 : node44239;
														assign node44239 = (inp[11]) ? node44243 : node44240;
															assign node44240 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node44243 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node44246 = (inp[13]) ? node44248 : 4'b0110;
															assign node44248 = (inp[11]) ? 4'b0110 : 4'b0111;
												assign node44251 = (inp[7]) ? node44259 : node44252;
													assign node44252 = (inp[11]) ? node44256 : node44253;
														assign node44253 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node44256 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node44259 = (inp[10]) ? node44273 : node44260;
														assign node44260 = (inp[9]) ? node44266 : node44261;
															assign node44261 = (inp[13]) ? node44263 : 4'b0011;
																assign node44263 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node44266 = (inp[13]) ? node44270 : node44267;
																assign node44267 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node44270 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node44273 = (inp[13]) ? node44277 : node44274;
															assign node44274 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node44277 = (inp[11]) ? 4'b0010 : 4'b0011;
							assign node44280 = (inp[11]) ? node44406 : node44281;
								assign node44281 = (inp[1]) ? node44333 : node44282;
									assign node44282 = (inp[13]) ? node44306 : node44283;
										assign node44283 = (inp[5]) ? node44295 : node44284;
											assign node44284 = (inp[4]) ? node44292 : node44285;
												assign node44285 = (inp[2]) ? node44289 : node44286;
													assign node44286 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node44289 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node44292 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node44295 = (inp[7]) ? node44301 : node44296;
												assign node44296 = (inp[4]) ? 4'b0101 : node44297;
													assign node44297 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node44301 = (inp[4]) ? 4'b0000 : node44302;
													assign node44302 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node44306 = (inp[5]) ? node44322 : node44307;
											assign node44307 = (inp[2]) ? node44315 : node44308;
												assign node44308 = (inp[4]) ? node44312 : node44309;
													assign node44309 = (inp[7]) ? 4'b0101 : 4'b0001;
													assign node44312 = (inp[7]) ? 4'b0001 : 4'b0101;
												assign node44315 = (inp[4]) ? node44319 : node44316;
													assign node44316 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node44319 = (inp[7]) ? 4'b0001 : 4'b0101;
											assign node44322 = (inp[7]) ? node44328 : node44323;
												assign node44323 = (inp[4]) ? 4'b0100 : node44324;
													assign node44324 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node44328 = (inp[4]) ? 4'b0001 : node44329;
													assign node44329 = (inp[2]) ? 4'b0101 : 4'b0100;
									assign node44333 = (inp[13]) ? node44357 : node44334;
										assign node44334 = (inp[5]) ? node44346 : node44335;
											assign node44335 = (inp[7]) ? node44341 : node44336;
												assign node44336 = (inp[4]) ? 4'b0100 : node44337;
													assign node44337 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node44341 = (inp[4]) ? 4'b0001 : node44342;
													assign node44342 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node44346 = (inp[4]) ? node44354 : node44347;
												assign node44347 = (inp[7]) ? node44351 : node44348;
													assign node44348 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node44351 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node44354 = (inp[7]) ? 4'b0001 : 4'b0101;
										assign node44357 = (inp[4]) ? node44401 : node44358;
											assign node44358 = (inp[7]) ? node44398 : node44359;
												assign node44359 = (inp[0]) ? node44367 : node44360;
													assign node44360 = (inp[5]) ? node44364 : node44361;
														assign node44361 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node44364 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node44367 = (inp[10]) ? node44383 : node44368;
														assign node44368 = (inp[9]) ? node44376 : node44369;
															assign node44369 = (inp[5]) ? node44373 : node44370;
																assign node44370 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node44373 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node44376 = (inp[2]) ? node44380 : node44377;
																assign node44377 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node44380 = (inp[5]) ? 4'b0001 : 4'b0000;
														assign node44383 = (inp[9]) ? node44391 : node44384;
															assign node44384 = (inp[5]) ? node44388 : node44385;
																assign node44385 = (inp[2]) ? 4'b0000 : 4'b0001;
																assign node44388 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node44391 = (inp[2]) ? node44395 : node44392;
																assign node44392 = (inp[5]) ? 4'b0000 : 4'b0001;
																assign node44395 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node44398 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node44401 = (inp[7]) ? 4'b0000 : node44402;
												assign node44402 = (inp[5]) ? 4'b0100 : 4'b0101;
								assign node44406 = (inp[1]) ? node44468 : node44407;
									assign node44407 = (inp[13]) ? node44431 : node44408;
										assign node44408 = (inp[5]) ? node44420 : node44409;
											assign node44409 = (inp[4]) ? node44417 : node44410;
												assign node44410 = (inp[2]) ? node44414 : node44411;
													assign node44411 = (inp[7]) ? 4'b0100 : 4'b0000;
													assign node44414 = (inp[7]) ? 4'b0101 : 4'b0001;
												assign node44417 = (inp[7]) ? 4'b0000 : 4'b0100;
											assign node44420 = (inp[7]) ? node44426 : node44421;
												assign node44421 = (inp[4]) ? 4'b0101 : node44422;
													assign node44422 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node44426 = (inp[4]) ? 4'b0000 : node44427;
													assign node44427 = (inp[2]) ? 4'b0100 : 4'b0101;
										assign node44431 = (inp[4]) ? node44463 : node44432;
											assign node44432 = (inp[7]) ? node44436 : node44433;
												assign node44433 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node44436 = (inp[0]) ? node44444 : node44437;
													assign node44437 = (inp[5]) ? node44441 : node44438;
														assign node44438 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node44441 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node44444 = (inp[10]) ? node44458 : node44445;
														assign node44445 = (inp[9]) ? node44451 : node44446;
															assign node44446 = (inp[5]) ? node44448 : 4'b0100;
																assign node44448 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node44451 = (inp[5]) ? node44455 : node44452;
																assign node44452 = (inp[2]) ? 4'b0100 : 4'b0101;
																assign node44455 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node44458 = (inp[2]) ? node44460 : 4'b0100;
															assign node44460 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node44463 = (inp[7]) ? 4'b0001 : node44464;
												assign node44464 = (inp[5]) ? 4'b0100 : 4'b0101;
									assign node44468 = (inp[13]) ? node44492 : node44469;
										assign node44469 = (inp[2]) ? node44481 : node44470;
											assign node44470 = (inp[4]) ? node44476 : node44471;
												assign node44471 = (inp[7]) ? 4'b0100 : node44472;
													assign node44472 = (inp[5]) ? 4'b0001 : 4'b0000;
												assign node44476 = (inp[7]) ? 4'b0001 : node44477;
													assign node44477 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node44481 = (inp[7]) ? node44489 : node44482;
												assign node44482 = (inp[4]) ? node44486 : node44483;
													assign node44483 = (inp[5]) ? 4'b0000 : 4'b0001;
													assign node44486 = (inp[5]) ? 4'b0101 : 4'b0100;
												assign node44489 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node44492 = (inp[4]) ? node44518 : node44493;
											assign node44493 = (inp[7]) ? node44515 : node44494;
												assign node44494 = (inp[9]) ? node44502 : node44495;
													assign node44495 = (inp[2]) ? node44499 : node44496;
														assign node44496 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node44499 = (inp[5]) ? 4'b0001 : 4'b0000;
													assign node44502 = (inp[10]) ? node44508 : node44503;
														assign node44503 = (inp[2]) ? 4'b0001 : node44504;
															assign node44504 = (inp[5]) ? 4'b0000 : 4'b0001;
														assign node44508 = (inp[5]) ? node44512 : node44509;
															assign node44509 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node44512 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node44515 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node44518 = (inp[7]) ? 4'b0000 : node44519;
												assign node44519 = (inp[5]) ? 4'b0100 : 4'b0101;
						assign node44523 = (inp[4]) ? node44839 : node44524;
							assign node44524 = (inp[5]) ? node44708 : node44525;
								assign node44525 = (inp[14]) ? node44549 : node44526;
									assign node44526 = (inp[11]) ? node44538 : node44527;
										assign node44527 = (inp[1]) ? node44533 : node44528;
											assign node44528 = (inp[2]) ? node44530 : 4'b0000;
												assign node44530 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node44533 = (inp[2]) ? node44535 : 4'b0001;
												assign node44535 = (inp[7]) ? 4'b0000 : 4'b0001;
										assign node44538 = (inp[1]) ? node44544 : node44539;
											assign node44539 = (inp[7]) ? node44541 : 4'b0001;
												assign node44541 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node44544 = (inp[7]) ? node44546 : 4'b0000;
												assign node44546 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node44549 = (inp[0]) ? node44645 : node44550;
										assign node44550 = (inp[13]) ? node44576 : node44551;
											assign node44551 = (inp[11]) ? node44569 : node44552;
												assign node44552 = (inp[10]) ? node44560 : node44553;
													assign node44553 = (inp[1]) ? node44557 : node44554;
														assign node44554 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node44557 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node44560 = (inp[7]) ? 4'b0101 : node44561;
														assign node44561 = (inp[2]) ? node44565 : node44562;
															assign node44562 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node44565 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node44569 = (inp[1]) ? node44573 : node44570;
													assign node44570 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node44573 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node44576 = (inp[7]) ? node44606 : node44577;
												assign node44577 = (inp[9]) ? node44593 : node44578;
													assign node44578 = (inp[11]) ? node44586 : node44579;
														assign node44579 = (inp[2]) ? node44583 : node44580;
															assign node44580 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node44583 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node44586 = (inp[1]) ? node44590 : node44587;
															assign node44587 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node44590 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node44593 = (inp[10]) ? node44599 : node44594;
														assign node44594 = (inp[2]) ? node44596 : 4'b0101;
															assign node44596 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node44599 = (inp[1]) ? node44603 : node44600;
															assign node44600 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node44603 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node44606 = (inp[10]) ? node44628 : node44607;
													assign node44607 = (inp[11]) ? node44621 : node44608;
														assign node44608 = (inp[9]) ? node44614 : node44609;
															assign node44609 = (inp[2]) ? 4'b0101 : node44610;
																assign node44610 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node44614 = (inp[1]) ? node44618 : node44615;
																assign node44615 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node44618 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node44621 = (inp[1]) ? node44625 : node44622;
															assign node44622 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node44625 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node44628 = (inp[9]) ? node44638 : node44629;
														assign node44629 = (inp[11]) ? node44631 : 4'b0100;
															assign node44631 = (inp[1]) ? node44635 : node44632;
																assign node44632 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node44635 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node44638 = (inp[2]) ? node44642 : node44639;
															assign node44639 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node44642 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node44645 = (inp[11]) ? node44681 : node44646;
											assign node44646 = (inp[7]) ? node44660 : node44647;
												assign node44647 = (inp[10]) ? node44653 : node44648;
													assign node44648 = (inp[2]) ? 4'b0100 : node44649;
														assign node44649 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node44653 = (inp[2]) ? node44657 : node44654;
														assign node44654 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node44657 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node44660 = (inp[10]) ? node44674 : node44661;
													assign node44661 = (inp[9]) ? node44669 : node44662;
														assign node44662 = (inp[1]) ? node44666 : node44663;
															assign node44663 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node44666 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node44669 = (inp[2]) ? 4'b0101 : node44670;
															assign node44670 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node44674 = (inp[2]) ? node44678 : node44675;
														assign node44675 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node44678 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node44681 = (inp[9]) ? node44701 : node44682;
												assign node44682 = (inp[7]) ? node44690 : node44683;
													assign node44683 = (inp[2]) ? node44687 : node44684;
														assign node44684 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node44687 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node44690 = (inp[10]) ? node44694 : node44691;
														assign node44691 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node44694 = (inp[2]) ? node44698 : node44695;
															assign node44695 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node44698 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node44701 = (inp[1]) ? node44705 : node44702;
													assign node44702 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node44705 = (inp[2]) ? 4'b0100 : 4'b0101;
								assign node44708 = (inp[9]) ? node44780 : node44709;
									assign node44709 = (inp[13]) ? node44749 : node44710;
										assign node44710 = (inp[2]) ? node44738 : node44711;
											assign node44711 = (inp[1]) ? node44721 : node44712;
												assign node44712 = (inp[14]) ? 4'b0100 : node44713;
													assign node44713 = (inp[7]) ? node44717 : node44714;
														assign node44714 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node44717 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node44721 = (inp[14]) ? 4'b0101 : node44722;
													assign node44722 = (inp[0]) ? node44728 : node44723;
														assign node44723 = (inp[11]) ? node44725 : 4'b0100;
															assign node44725 = (inp[7]) ? 4'b0101 : 4'b0100;
														assign node44728 = (inp[10]) ? 4'b0101 : node44729;
															assign node44729 = (inp[11]) ? node44733 : node44730;
																assign node44730 = (inp[7]) ? 4'b0100 : 4'b0101;
																assign node44733 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node44738 = (inp[1]) ? node44744 : node44739;
												assign node44739 = (inp[11]) ? 4'b0101 : node44740;
													assign node44740 = (inp[14]) ? 4'b0101 : 4'b0100;
												assign node44744 = (inp[14]) ? 4'b0100 : node44745;
													assign node44745 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node44749 = (inp[14]) ? node44773 : node44750;
											assign node44750 = (inp[11]) ? node44762 : node44751;
												assign node44751 = (inp[1]) ? node44757 : node44752;
													assign node44752 = (inp[7]) ? node44754 : 4'b0100;
														assign node44754 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node44757 = (inp[2]) ? 4'b0101 : node44758;
														assign node44758 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node44762 = (inp[1]) ? node44768 : node44763;
													assign node44763 = (inp[7]) ? node44765 : 4'b0101;
														assign node44765 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node44768 = (inp[2]) ? 4'b0100 : node44769;
														assign node44769 = (inp[7]) ? 4'b0101 : 4'b0100;
											assign node44773 = (inp[1]) ? node44777 : node44774;
												assign node44774 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node44777 = (inp[2]) ? 4'b0100 : 4'b0101;
									assign node44780 = (inp[11]) ? node44824 : node44781;
										assign node44781 = (inp[1]) ? node44791 : node44782;
											assign node44782 = (inp[14]) ? node44788 : node44783;
												assign node44783 = (inp[7]) ? node44785 : 4'b0100;
													assign node44785 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node44788 = (inp[2]) ? 4'b0101 : 4'b0100;
											assign node44791 = (inp[7]) ? node44797 : node44792;
												assign node44792 = (inp[14]) ? node44794 : 4'b0101;
													assign node44794 = (inp[2]) ? 4'b0100 : 4'b0101;
												assign node44797 = (inp[13]) ? node44811 : node44798;
													assign node44798 = (inp[0]) ? node44804 : node44799;
														assign node44799 = (inp[2]) ? node44801 : 4'b0101;
															assign node44801 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node44804 = (inp[2]) ? node44808 : node44805;
															assign node44805 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node44808 = (inp[14]) ? 4'b0100 : 4'b0101;
													assign node44811 = (inp[0]) ? node44819 : node44812;
														assign node44812 = (inp[2]) ? node44816 : node44813;
															assign node44813 = (inp[14]) ? 4'b0101 : 4'b0100;
															assign node44816 = (inp[14]) ? 4'b0100 : 4'b0101;
														assign node44819 = (inp[14]) ? 4'b0101 : node44820;
															assign node44820 = (inp[2]) ? 4'b0101 : 4'b0100;
										assign node44824 = (inp[1]) ? node44832 : node44825;
											assign node44825 = (inp[2]) ? 4'b0101 : node44826;
												assign node44826 = (inp[7]) ? 4'b0100 : node44827;
													assign node44827 = (inp[14]) ? 4'b0100 : 4'b0101;
											assign node44832 = (inp[2]) ? 4'b0100 : node44833;
												assign node44833 = (inp[7]) ? 4'b0101 : node44834;
													assign node44834 = (inp[14]) ? 4'b0101 : 4'b0100;
							assign node44839 = (inp[5]) ? node45007 : node44840;
								assign node44840 = (inp[14]) ? node45000 : node44841;
									assign node44841 = (inp[2]) ? node44953 : node44842;
										assign node44842 = (inp[13]) ? node44910 : node44843;
											assign node44843 = (inp[7]) ? node44885 : node44844;
												assign node44844 = (inp[10]) ? node44864 : node44845;
													assign node44845 = (inp[9]) ? node44859 : node44846;
														assign node44846 = (inp[0]) ? node44854 : node44847;
															assign node44847 = (inp[11]) ? node44851 : node44848;
																assign node44848 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node44851 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node44854 = (inp[11]) ? node44856 : 4'b0100;
																assign node44856 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node44859 = (inp[11]) ? node44861 : 4'b0100;
															assign node44861 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node44864 = (inp[0]) ? node44872 : node44865;
														assign node44865 = (inp[1]) ? node44869 : node44866;
															assign node44866 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node44869 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node44872 = (inp[9]) ? node44880 : node44873;
															assign node44873 = (inp[11]) ? node44877 : node44874;
																assign node44874 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node44877 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node44880 = (inp[1]) ? 4'b0101 : node44881;
																assign node44881 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node44885 = (inp[0]) ? node44893 : node44886;
													assign node44886 = (inp[11]) ? node44890 : node44887;
														assign node44887 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node44890 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node44893 = (inp[9]) ? node44899 : node44894;
														assign node44894 = (inp[1]) ? 4'b0101 : node44895;
															assign node44895 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node44899 = (inp[10]) ? node44905 : node44900;
															assign node44900 = (inp[11]) ? node44902 : 4'b0101;
																assign node44902 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node44905 = (inp[11]) ? node44907 : 4'b0100;
																assign node44907 = (inp[1]) ? 4'b0100 : 4'b0101;
											assign node44910 = (inp[9]) ? node44938 : node44911;
												assign node44911 = (inp[0]) ? node44919 : node44912;
													assign node44912 = (inp[1]) ? node44916 : node44913;
														assign node44913 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node44916 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node44919 = (inp[7]) ? node44925 : node44920;
														assign node44920 = (inp[11]) ? node44922 : 4'b0100;
															assign node44922 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node44925 = (inp[10]) ? node44933 : node44926;
															assign node44926 = (inp[11]) ? node44930 : node44927;
																assign node44927 = (inp[1]) ? 4'b0101 : 4'b0100;
																assign node44930 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node44933 = (inp[11]) ? 4'b0100 : node44934;
																assign node44934 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node44938 = (inp[7]) ? node44946 : node44939;
													assign node44939 = (inp[11]) ? node44943 : node44940;
														assign node44940 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node44943 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node44946 = (inp[11]) ? node44950 : node44947;
														assign node44947 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node44950 = (inp[1]) ? 4'b0100 : 4'b0101;
										assign node44953 = (inp[1]) ? node44961 : node44954;
											assign node44954 = (inp[7]) ? node44958 : node44955;
												assign node44955 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node44958 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node44961 = (inp[10]) ? node44993 : node44962;
												assign node44962 = (inp[13]) ? node44986 : node44963;
													assign node44963 = (inp[9]) ? node44979 : node44964;
														assign node44964 = (inp[0]) ? node44972 : node44965;
															assign node44965 = (inp[11]) ? node44969 : node44966;
																assign node44966 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node44969 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node44972 = (inp[7]) ? node44976 : node44973;
																assign node44973 = (inp[11]) ? 4'b0101 : 4'b0100;
																assign node44976 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node44979 = (inp[7]) ? node44983 : node44980;
															assign node44980 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node44983 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node44986 = (inp[7]) ? node44990 : node44987;
														assign node44987 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node44990 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node44993 = (inp[11]) ? node44997 : node44994;
													assign node44994 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node44997 = (inp[7]) ? 4'b0100 : 4'b0101;
									assign node45000 = (inp[1]) ? node45004 : node45001;
										assign node45001 = (inp[7]) ? 4'b0001 : 4'b0000;
										assign node45004 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node45007 = (inp[1]) ? node45021 : node45008;
									assign node45008 = (inp[14]) ? 4'b0001 : node45009;
										assign node45009 = (inp[11]) ? node45015 : node45010;
											assign node45010 = (inp[7]) ? 4'b0000 : node45011;
												assign node45011 = (inp[2]) ? 4'b0000 : 4'b0001;
											assign node45015 = (inp[7]) ? 4'b0001 : node45016;
												assign node45016 = (inp[2]) ? 4'b0001 : 4'b0000;
									assign node45021 = (inp[14]) ? 4'b0000 : node45022;
										assign node45022 = (inp[11]) ? node45028 : node45023;
											assign node45023 = (inp[2]) ? 4'b0001 : node45024;
												assign node45024 = (inp[7]) ? 4'b0001 : 4'b0000;
											assign node45028 = (inp[2]) ? 4'b0000 : node45029;
												assign node45029 = (inp[7]) ? 4'b0000 : 4'b0001;
				assign node45034 = (inp[14]) ? node46782 : node45035;
					assign node45035 = (inp[15]) ? node46277 : node45036;
						assign node45036 = (inp[6]) ? node45716 : node45037;
							assign node45037 = (inp[11]) ? node45397 : node45038;
								assign node45038 = (inp[13]) ? node45280 : node45039;
									assign node45039 = (inp[4]) ? node45135 : node45040;
										assign node45040 = (inp[7]) ? node45104 : node45041;
											assign node45041 = (inp[2]) ? node45073 : node45042;
												assign node45042 = (inp[5]) ? node45058 : node45043;
													assign node45043 = (inp[0]) ? node45051 : node45044;
														assign node45044 = (inp[1]) ? node45048 : node45045;
															assign node45045 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node45048 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node45051 = (inp[1]) ? node45055 : node45052;
															assign node45052 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node45055 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node45058 = (inp[0]) ? node45064 : node45059;
														assign node45059 = (inp[1]) ? 4'b0010 : node45060;
															assign node45060 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node45064 = (inp[9]) ? node45066 : 4'b0010;
															assign node45066 = (inp[10]) ? node45070 : node45067;
																assign node45067 = (inp[1]) ? 4'b0011 : 4'b0010;
																assign node45070 = (inp[1]) ? 4'b0010 : 4'b0011;
												assign node45073 = (inp[0]) ? node45091 : node45074;
													assign node45074 = (inp[9]) ? node45080 : node45075;
														assign node45075 = (inp[1]) ? node45077 : 4'b0110;
															assign node45077 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node45080 = (inp[5]) ? node45086 : node45081;
															assign node45081 = (inp[10]) ? node45083 : 4'b0111;
																assign node45083 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node45086 = (inp[1]) ? 4'b0110 : node45087;
																assign node45087 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node45091 = (inp[9]) ? node45097 : node45092;
														assign node45092 = (inp[10]) ? 4'b0111 : node45093;
															assign node45093 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node45097 = (inp[10]) ? node45101 : node45098;
															assign node45098 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node45101 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node45104 = (inp[2]) ? node45120 : node45105;
												assign node45105 = (inp[1]) ? node45113 : node45106;
													assign node45106 = (inp[10]) ? node45110 : node45107;
														assign node45107 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node45110 = (inp[5]) ? 4'b0110 : 4'b0111;
													assign node45113 = (inp[5]) ? node45117 : node45114;
														assign node45114 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node45117 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node45120 = (inp[1]) ? node45128 : node45121;
													assign node45121 = (inp[5]) ? node45125 : node45122;
														assign node45122 = (inp[10]) ? 4'b0010 : 4'b0011;
														assign node45125 = (inp[10]) ? 4'b0011 : 4'b0010;
													assign node45128 = (inp[10]) ? node45132 : node45129;
														assign node45129 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node45132 = (inp[5]) ? 4'b0010 : 4'b0011;
										assign node45135 = (inp[0]) ? node45213 : node45136;
											assign node45136 = (inp[5]) ? node45170 : node45137;
												assign node45137 = (inp[10]) ? node45151 : node45138;
													assign node45138 = (inp[1]) ? node45144 : node45139;
														assign node45139 = (inp[2]) ? 4'b0110 : node45140;
															assign node45140 = (inp[7]) ? 4'b0011 : 4'b0110;
														assign node45144 = (inp[2]) ? node45148 : node45145;
															assign node45145 = (inp[7]) ? 4'b0010 : 4'b0111;
															assign node45148 = (inp[7]) ? 4'b0111 : 4'b0011;
													assign node45151 = (inp[1]) ? node45163 : node45152;
														assign node45152 = (inp[9]) ? node45158 : node45153;
															assign node45153 = (inp[2]) ? node45155 : 4'b0111;
																assign node45155 = (inp[7]) ? 4'b0111 : 4'b0010;
															assign node45158 = (inp[7]) ? node45160 : 4'b0111;
																assign node45160 = (inp[2]) ? 4'b0111 : 4'b0010;
														assign node45163 = (inp[7]) ? node45167 : node45164;
															assign node45164 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node45167 = (inp[2]) ? 4'b0110 : 4'b0011;
												assign node45170 = (inp[2]) ? node45188 : node45171;
													assign node45171 = (inp[7]) ? node45185 : node45172;
														assign node45172 = (inp[9]) ? node45178 : node45173;
															assign node45173 = (inp[1]) ? node45175 : 4'b0010;
																assign node45175 = (inp[10]) ? 4'b0011 : 4'b0010;
															assign node45178 = (inp[1]) ? node45182 : node45179;
																assign node45179 = (inp[10]) ? 4'b0010 : 4'b0011;
																assign node45182 = (inp[10]) ? 4'b0011 : 4'b0010;
														assign node45185 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node45188 = (inp[7]) ? node45202 : node45189;
														assign node45189 = (inp[9]) ? node45195 : node45190;
															assign node45190 = (inp[10]) ? node45192 : 4'b0111;
																assign node45192 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node45195 = (inp[1]) ? node45199 : node45196;
																assign node45196 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node45199 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node45202 = (inp[9]) ? node45208 : node45203;
															assign node45203 = (inp[10]) ? node45205 : 4'b0011;
																assign node45205 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node45208 = (inp[10]) ? 4'b0010 : node45209;
																assign node45209 = (inp[1]) ? 4'b0011 : 4'b0010;
											assign node45213 = (inp[1]) ? node45251 : node45214;
												assign node45214 = (inp[2]) ? node45236 : node45215;
													assign node45215 = (inp[9]) ? node45223 : node45216;
														assign node45216 = (inp[10]) ? 4'b0010 : node45217;
															assign node45217 = (inp[5]) ? 4'b0110 : node45218;
																assign node45218 = (inp[7]) ? 4'b0011 : 4'b0110;
														assign node45223 = (inp[5]) ? node45231 : node45224;
															assign node45224 = (inp[7]) ? node45228 : node45225;
																assign node45225 = (inp[10]) ? 4'b0111 : 4'b0110;
																assign node45228 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node45231 = (inp[7]) ? 4'b0111 : node45232;
																assign node45232 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node45236 = (inp[10]) ? node45244 : node45237;
														assign node45237 = (inp[7]) ? node45241 : node45238;
															assign node45238 = (inp[5]) ? 4'b0110 : 4'b0011;
															assign node45241 = (inp[5]) ? 4'b0010 : 4'b0110;
														assign node45244 = (inp[5]) ? node45248 : node45245;
															assign node45245 = (inp[7]) ? 4'b0111 : 4'b0010;
															assign node45248 = (inp[7]) ? 4'b0011 : 4'b0111;
												assign node45251 = (inp[2]) ? node45267 : node45252;
													assign node45252 = (inp[10]) ? node45260 : node45253;
														assign node45253 = (inp[7]) ? node45257 : node45254;
															assign node45254 = (inp[5]) ? 4'b0010 : 4'b0111;
															assign node45257 = (inp[5]) ? 4'b0110 : 4'b0010;
														assign node45260 = (inp[7]) ? node45264 : node45261;
															assign node45261 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node45264 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node45267 = (inp[10]) ? node45273 : node45268;
														assign node45268 = (inp[5]) ? node45270 : 4'b0111;
															assign node45270 = (inp[7]) ? 4'b0011 : 4'b0111;
														assign node45273 = (inp[5]) ? node45277 : node45274;
															assign node45274 = (inp[7]) ? 4'b0110 : 4'b0010;
															assign node45277 = (inp[7]) ? 4'b0010 : 4'b0110;
									assign node45280 = (inp[1]) ? node45344 : node45281;
										assign node45281 = (inp[10]) ? node45311 : node45282;
											assign node45282 = (inp[5]) ? node45300 : node45283;
												assign node45283 = (inp[4]) ? node45291 : node45284;
													assign node45284 = (inp[7]) ? node45288 : node45285;
														assign node45285 = (inp[2]) ? 4'b0111 : 4'b0011;
														assign node45288 = (inp[2]) ? 4'b0010 : 4'b0111;
													assign node45291 = (inp[9]) ? node45293 : 4'b0010;
														assign node45293 = (inp[2]) ? node45297 : node45294;
															assign node45294 = (inp[7]) ? 4'b0010 : 4'b0111;
															assign node45297 = (inp[7]) ? 4'b0111 : 4'b0010;
												assign node45300 = (inp[2]) ? node45308 : node45301;
													assign node45301 = (inp[7]) ? node45305 : node45302;
														assign node45302 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node45305 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node45308 = (inp[7]) ? 4'b0011 : 4'b0111;
											assign node45311 = (inp[4]) ? node45323 : node45312;
												assign node45312 = (inp[7]) ? node45316 : node45313;
													assign node45313 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node45316 = (inp[2]) ? node45320 : node45317;
														assign node45317 = (inp[5]) ? 4'b0111 : 4'b0110;
														assign node45320 = (inp[5]) ? 4'b0010 : 4'b0011;
												assign node45323 = (inp[7]) ? node45337 : node45324;
													assign node45324 = (inp[9]) ? node45330 : node45325;
														assign node45325 = (inp[5]) ? 4'b0011 : node45326;
															assign node45326 = (inp[2]) ? 4'b0011 : 4'b0110;
														assign node45330 = (inp[2]) ? node45334 : node45331;
															assign node45331 = (inp[5]) ? 4'b0011 : 4'b0110;
															assign node45334 = (inp[5]) ? 4'b0110 : 4'b0011;
													assign node45337 = (inp[5]) ? node45341 : node45338;
														assign node45338 = (inp[2]) ? 4'b0110 : 4'b0011;
														assign node45341 = (inp[2]) ? 4'b0010 : 4'b0110;
										assign node45344 = (inp[10]) ? node45370 : node45345;
											assign node45345 = (inp[7]) ? node45357 : node45346;
												assign node45346 = (inp[2]) ? node45352 : node45347;
													assign node45347 = (inp[4]) ? node45349 : 4'b0010;
														assign node45349 = (inp[5]) ? 4'b0011 : 4'b0110;
													assign node45352 = (inp[4]) ? node45354 : 4'b0110;
														assign node45354 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node45357 = (inp[2]) ? node45365 : node45358;
													assign node45358 = (inp[4]) ? node45362 : node45359;
														assign node45359 = (inp[5]) ? 4'b0110 : 4'b0111;
														assign node45362 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node45365 = (inp[5]) ? 4'b0010 : node45366;
														assign node45366 = (inp[4]) ? 4'b0110 : 4'b0011;
											assign node45370 = (inp[2]) ? node45384 : node45371;
												assign node45371 = (inp[4]) ? node45377 : node45372;
													assign node45372 = (inp[7]) ? node45374 : 4'b0011;
														assign node45374 = (inp[5]) ? 4'b0111 : 4'b0110;
													assign node45377 = (inp[7]) ? node45381 : node45378;
														assign node45378 = (inp[5]) ? 4'b0010 : 4'b0111;
														assign node45381 = (inp[5]) ? 4'b0110 : 4'b0010;
												assign node45384 = (inp[7]) ? node45390 : node45385;
													assign node45385 = (inp[4]) ? node45387 : 4'b0111;
														assign node45387 = (inp[5]) ? 4'b0111 : 4'b0011;
													assign node45390 = (inp[4]) ? node45394 : node45391;
														assign node45391 = (inp[5]) ? 4'b0011 : 4'b0010;
														assign node45394 = (inp[5]) ? 4'b0011 : 4'b0111;
								assign node45397 = (inp[2]) ? node45563 : node45398;
									assign node45398 = (inp[7]) ? node45446 : node45399;
										assign node45399 = (inp[4]) ? node45407 : node45400;
											assign node45400 = (inp[13]) ? node45404 : node45401;
												assign node45401 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node45404 = (inp[10]) ? 4'b0010 : 4'b0011;
											assign node45407 = (inp[5]) ? node45439 : node45408;
												assign node45408 = (inp[0]) ? node45424 : node45409;
													assign node45409 = (inp[9]) ? node45417 : node45410;
														assign node45410 = (inp[13]) ? node45414 : node45411;
															assign node45411 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node45414 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node45417 = (inp[10]) ? node45421 : node45418;
															assign node45418 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node45421 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node45424 = (inp[9]) ? node45432 : node45425;
														assign node45425 = (inp[10]) ? node45429 : node45426;
															assign node45426 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node45429 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node45432 = (inp[13]) ? node45436 : node45433;
															assign node45433 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node45436 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node45439 = (inp[10]) ? node45443 : node45440;
													assign node45440 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node45443 = (inp[13]) ? 4'b0011 : 4'b0010;
										assign node45446 = (inp[5]) ? node45494 : node45447;
											assign node45447 = (inp[4]) ? node45487 : node45448;
												assign node45448 = (inp[0]) ? node45470 : node45449;
													assign node45449 = (inp[9]) ? node45459 : node45450;
														assign node45450 = (inp[13]) ? node45452 : 4'b0110;
															assign node45452 = (inp[10]) ? node45456 : node45453;
																assign node45453 = (inp[1]) ? 4'b0111 : 4'b0110;
																assign node45456 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node45459 = (inp[13]) ? node45465 : node45460;
															assign node45460 = (inp[10]) ? node45462 : 4'b0111;
																assign node45462 = (inp[1]) ? 4'b0111 : 4'b0110;
															assign node45465 = (inp[10]) ? node45467 : 4'b0110;
																assign node45467 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node45470 = (inp[1]) ? node45480 : node45471;
														assign node45471 = (inp[9]) ? node45473 : 4'b0111;
															assign node45473 = (inp[13]) ? node45477 : node45474;
																assign node45474 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node45477 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node45480 = (inp[10]) ? node45484 : node45481;
															assign node45481 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node45484 = (inp[13]) ? 4'b0110 : 4'b0111;
												assign node45487 = (inp[13]) ? node45491 : node45488;
													assign node45488 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node45491 = (inp[10]) ? 4'b0011 : 4'b0010;
											assign node45494 = (inp[0]) ? node45532 : node45495;
												assign node45495 = (inp[1]) ? node45517 : node45496;
													assign node45496 = (inp[4]) ? node45502 : node45497;
														assign node45497 = (inp[13]) ? node45499 : 4'b0110;
															assign node45499 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node45502 = (inp[9]) ? node45510 : node45503;
															assign node45503 = (inp[13]) ? node45507 : node45504;
																assign node45504 = (inp[10]) ? 4'b0110 : 4'b0111;
																assign node45507 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node45510 = (inp[10]) ? node45514 : node45511;
																assign node45511 = (inp[13]) ? 4'b0110 : 4'b0111;
																assign node45514 = (inp[13]) ? 4'b0111 : 4'b0110;
													assign node45517 = (inp[13]) ? node45525 : node45518;
														assign node45518 = (inp[4]) ? node45522 : node45519;
															assign node45519 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node45522 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node45525 = (inp[10]) ? node45529 : node45526;
															assign node45526 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node45529 = (inp[4]) ? 4'b0110 : 4'b0111;
												assign node45532 = (inp[1]) ? node45548 : node45533;
													assign node45533 = (inp[4]) ? node45541 : node45534;
														assign node45534 = (inp[9]) ? node45536 : 4'b0111;
															assign node45536 = (inp[13]) ? node45538 : 4'b0111;
																assign node45538 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node45541 = (inp[13]) ? node45545 : node45542;
															assign node45542 = (inp[10]) ? 4'b0110 : 4'b0111;
															assign node45545 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node45548 = (inp[10]) ? node45556 : node45549;
														assign node45549 = (inp[4]) ? node45553 : node45550;
															assign node45550 = (inp[13]) ? 4'b0110 : 4'b0111;
															assign node45553 = (inp[13]) ? 4'b0111 : 4'b0110;
														assign node45556 = (inp[4]) ? node45560 : node45557;
															assign node45557 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node45560 = (inp[13]) ? 4'b0110 : 4'b0111;
									assign node45563 = (inp[7]) ? node45647 : node45564;
										assign node45564 = (inp[4]) ? node45594 : node45565;
											assign node45565 = (inp[5]) ? node45587 : node45566;
												assign node45566 = (inp[9]) ? node45580 : node45567;
													assign node45567 = (inp[1]) ? node45575 : node45568;
														assign node45568 = (inp[10]) ? node45572 : node45569;
															assign node45569 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node45572 = (inp[13]) ? 4'b0110 : 4'b0111;
														assign node45575 = (inp[13]) ? 4'b0110 : node45576;
															assign node45576 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node45580 = (inp[13]) ? node45584 : node45581;
														assign node45581 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node45584 = (inp[10]) ? 4'b0110 : 4'b0111;
												assign node45587 = (inp[13]) ? node45591 : node45588;
													assign node45588 = (inp[10]) ? 4'b0111 : 4'b0110;
													assign node45591 = (inp[10]) ? 4'b0110 : 4'b0111;
											assign node45594 = (inp[5]) ? node45624 : node45595;
												assign node45595 = (inp[0]) ? node45611 : node45596;
													assign node45596 = (inp[10]) ? node45606 : node45597;
														assign node45597 = (inp[9]) ? node45601 : node45598;
															assign node45598 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node45601 = (inp[13]) ? 4'b0010 : node45602;
																assign node45602 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node45606 = (inp[9]) ? node45608 : 4'b0010;
															assign node45608 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node45611 = (inp[13]) ? node45617 : node45612;
														assign node45612 = (inp[10]) ? node45614 : 4'b0011;
															assign node45614 = (inp[1]) ? 4'b0010 : 4'b0011;
														assign node45617 = (inp[1]) ? node45621 : node45618;
															assign node45618 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node45621 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node45624 = (inp[1]) ? node45640 : node45625;
													assign node45625 = (inp[0]) ? node45633 : node45626;
														assign node45626 = (inp[13]) ? node45630 : node45627;
															assign node45627 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node45630 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node45633 = (inp[13]) ? node45637 : node45634;
															assign node45634 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node45637 = (inp[10]) ? 4'b0110 : 4'b0111;
													assign node45640 = (inp[13]) ? node45644 : node45641;
														assign node45641 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node45644 = (inp[10]) ? 4'b0110 : 4'b0111;
										assign node45647 = (inp[5]) ? node45701 : node45648;
											assign node45648 = (inp[4]) ? node45670 : node45649;
												assign node45649 = (inp[1]) ? node45657 : node45650;
													assign node45650 = (inp[10]) ? node45654 : node45651;
														assign node45651 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node45654 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node45657 = (inp[0]) ? node45663 : node45658;
														assign node45658 = (inp[13]) ? node45660 : 4'b0011;
															assign node45660 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node45663 = (inp[13]) ? node45667 : node45664;
															assign node45664 = (inp[10]) ? 4'b0010 : 4'b0011;
															assign node45667 = (inp[10]) ? 4'b0011 : 4'b0010;
												assign node45670 = (inp[0]) ? node45686 : node45671;
													assign node45671 = (inp[9]) ? node45679 : node45672;
														assign node45672 = (inp[1]) ? node45674 : 4'b0111;
															assign node45674 = (inp[13]) ? node45676 : 4'b0111;
																assign node45676 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node45679 = (inp[10]) ? node45683 : node45680;
															assign node45680 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node45683 = (inp[13]) ? 4'b0110 : 4'b0111;
													assign node45686 = (inp[1]) ? node45694 : node45687;
														assign node45687 = (inp[13]) ? node45691 : node45688;
															assign node45688 = (inp[10]) ? 4'b0111 : 4'b0110;
															assign node45691 = (inp[10]) ? 4'b0110 : 4'b0111;
														assign node45694 = (inp[10]) ? node45698 : node45695;
															assign node45695 = (inp[13]) ? 4'b0111 : 4'b0110;
															assign node45698 = (inp[13]) ? 4'b0110 : 4'b0111;
											assign node45701 = (inp[1]) ? node45709 : node45702;
												assign node45702 = (inp[10]) ? node45706 : node45703;
													assign node45703 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node45706 = (inp[13]) ? 4'b0010 : 4'b0011;
												assign node45709 = (inp[10]) ? node45713 : node45710;
													assign node45710 = (inp[13]) ? 4'b0011 : 4'b0010;
													assign node45713 = (inp[13]) ? 4'b0010 : 4'b0011;
							assign node45716 = (inp[7]) ? node46000 : node45717;
								assign node45717 = (inp[5]) ? node45901 : node45718;
									assign node45718 = (inp[2]) ? node45804 : node45719;
										assign node45719 = (inp[10]) ? node45763 : node45720;
											assign node45720 = (inp[9]) ? node45742 : node45721;
												assign node45721 = (inp[1]) ? node45729 : node45722;
													assign node45722 = (inp[11]) ? node45726 : node45723;
														assign node45723 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node45726 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node45729 = (inp[4]) ? node45735 : node45730;
														assign node45730 = (inp[11]) ? 4'b0010 : node45731;
															assign node45731 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node45735 = (inp[13]) ? node45739 : node45736;
															assign node45736 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node45739 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node45742 = (inp[4]) ? node45756 : node45743;
													assign node45743 = (inp[13]) ? node45749 : node45744;
														assign node45744 = (inp[1]) ? node45746 : 4'b0011;
															assign node45746 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node45749 = (inp[1]) ? node45753 : node45750;
															assign node45750 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node45753 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node45756 = (inp[13]) ? node45760 : node45757;
														assign node45757 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node45760 = (inp[11]) ? 4'b0010 : 4'b0011;
											assign node45763 = (inp[1]) ? node45789 : node45764;
												assign node45764 = (inp[0]) ? node45772 : node45765;
													assign node45765 = (inp[13]) ? node45769 : node45766;
														assign node45766 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node45769 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node45772 = (inp[4]) ? node45782 : node45773;
														assign node45773 = (inp[9]) ? node45775 : 4'b0011;
															assign node45775 = (inp[13]) ? node45779 : node45776;
																assign node45776 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node45779 = (inp[11]) ? 4'b0010 : 4'b0011;
														assign node45782 = (inp[13]) ? node45786 : node45783;
															assign node45783 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node45786 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node45789 = (inp[0]) ? node45791 : 4'b0011;
													assign node45791 = (inp[11]) ? node45799 : node45792;
														assign node45792 = (inp[4]) ? node45796 : node45793;
															assign node45793 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node45796 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node45799 = (inp[4]) ? 4'b0011 : node45800;
															assign node45800 = (inp[13]) ? 4'b0011 : 4'b0010;
										assign node45804 = (inp[0]) ? node45858 : node45805;
											assign node45805 = (inp[10]) ? node45831 : node45806;
												assign node45806 = (inp[1]) ? node45822 : node45807;
													assign node45807 = (inp[9]) ? node45813 : node45808;
														assign node45808 = (inp[13]) ? node45810 : 4'b0010;
															assign node45810 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node45813 = (inp[4]) ? node45817 : node45814;
															assign node45814 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node45817 = (inp[13]) ? 4'b0011 : node45818;
																assign node45818 = (inp[11]) ? 4'b0011 : 4'b0010;
													assign node45822 = (inp[11]) ? node45824 : 4'b0010;
														assign node45824 = (inp[13]) ? node45828 : node45825;
															assign node45825 = (inp[4]) ? 4'b0010 : 4'b0011;
															assign node45828 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node45831 = (inp[4]) ? node45839 : node45832;
													assign node45832 = (inp[11]) ? node45836 : node45833;
														assign node45833 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node45836 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node45839 = (inp[11]) ? node45853 : node45840;
														assign node45840 = (inp[9]) ? node45848 : node45841;
															assign node45841 = (inp[1]) ? node45845 : node45842;
																assign node45842 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node45845 = (inp[13]) ? 4'b0010 : 4'b0011;
															assign node45848 = (inp[13]) ? 4'b0010 : node45849;
																assign node45849 = (inp[1]) ? 4'b0011 : 4'b0010;
														assign node45853 = (inp[13]) ? 4'b0011 : node45854;
															assign node45854 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node45858 = (inp[10]) ? node45878 : node45859;
												assign node45859 = (inp[13]) ? node45867 : node45860;
													assign node45860 = (inp[11]) ? 4'b0011 : node45861;
														assign node45861 = (inp[1]) ? node45863 : 4'b0010;
															assign node45863 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node45867 = (inp[11]) ? node45873 : node45868;
														assign node45868 = (inp[1]) ? node45870 : 4'b0011;
															assign node45870 = (inp[9]) ? 4'b0010 : 4'b0011;
														assign node45873 = (inp[1]) ? node45875 : 4'b0010;
															assign node45875 = (inp[4]) ? 4'b0011 : 4'b0010;
												assign node45878 = (inp[1]) ? node45886 : node45879;
													assign node45879 = (inp[11]) ? node45883 : node45880;
														assign node45880 = (inp[13]) ? 4'b0011 : 4'b0010;
														assign node45883 = (inp[13]) ? 4'b0010 : 4'b0011;
													assign node45886 = (inp[4]) ? node45896 : node45887;
														assign node45887 = (inp[9]) ? 4'b0010 : node45888;
															assign node45888 = (inp[11]) ? node45892 : node45889;
																assign node45889 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node45892 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node45896 = (inp[13]) ? node45898 : 4'b0010;
															assign node45898 = (inp[11]) ? 4'b0011 : 4'b0010;
									assign node45901 = (inp[11]) ? node45957 : node45902;
										assign node45902 = (inp[13]) ? node45926 : node45903;
											assign node45903 = (inp[2]) ? 4'b0110 : node45904;
												assign node45904 = (inp[9]) ? node45912 : node45905;
													assign node45905 = (inp[4]) ? node45909 : node45906;
														assign node45906 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node45909 = (inp[1]) ? 4'b0110 : 4'b0111;
													assign node45912 = (inp[10]) ? node45920 : node45913;
														assign node45913 = (inp[1]) ? node45917 : node45914;
															assign node45914 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node45917 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node45920 = (inp[4]) ? node45922 : 4'b0111;
															assign node45922 = (inp[1]) ? 4'b0110 : 4'b0111;
											assign node45926 = (inp[2]) ? 4'b0111 : node45927;
												assign node45927 = (inp[9]) ? node45947 : node45928;
													assign node45928 = (inp[0]) ? node45938 : node45929;
														assign node45929 = (inp[10]) ? 4'b0111 : node45930;
															assign node45930 = (inp[1]) ? node45934 : node45931;
																assign node45931 = (inp[4]) ? 4'b0110 : 4'b0111;
																assign node45934 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node45938 = (inp[10]) ? node45940 : 4'b0111;
															assign node45940 = (inp[4]) ? node45944 : node45941;
																assign node45941 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node45944 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node45947 = (inp[10]) ? node45949 : 4'b0110;
														assign node45949 = (inp[4]) ? node45953 : node45950;
															assign node45950 = (inp[1]) ? 4'b0110 : 4'b0111;
															assign node45953 = (inp[1]) ? 4'b0111 : 4'b0110;
										assign node45957 = (inp[13]) ? node45991 : node45958;
											assign node45958 = (inp[2]) ? 4'b0111 : node45959;
												assign node45959 = (inp[0]) ? node45967 : node45960;
													assign node45960 = (inp[4]) ? node45964 : node45961;
														assign node45961 = (inp[1]) ? 4'b0110 : 4'b0111;
														assign node45964 = (inp[1]) ? 4'b0111 : 4'b0110;
													assign node45967 = (inp[9]) ? node45977 : node45968;
														assign node45968 = (inp[10]) ? 4'b0111 : node45969;
															assign node45969 = (inp[4]) ? node45973 : node45970;
																assign node45970 = (inp[1]) ? 4'b0110 : 4'b0111;
																assign node45973 = (inp[1]) ? 4'b0111 : 4'b0110;
														assign node45977 = (inp[10]) ? node45985 : node45978;
															assign node45978 = (inp[1]) ? node45982 : node45979;
																assign node45979 = (inp[4]) ? 4'b0110 : 4'b0111;
																assign node45982 = (inp[4]) ? 4'b0111 : 4'b0110;
															assign node45985 = (inp[1]) ? 4'b0110 : node45986;
																assign node45986 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node45991 = (inp[2]) ? 4'b0110 : node45992;
												assign node45992 = (inp[1]) ? node45996 : node45993;
													assign node45993 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node45996 = (inp[4]) ? 4'b0110 : 4'b0111;
								assign node46000 = (inp[5]) ? node46060 : node46001;
									assign node46001 = (inp[11]) ? node46041 : node46002;
										assign node46002 = (inp[13]) ? node46018 : node46003;
											assign node46003 = (inp[1]) ? 4'b0110 : node46004;
												assign node46004 = (inp[9]) ? node46010 : node46005;
													assign node46005 = (inp[2]) ? node46007 : 4'b0111;
														assign node46007 = (inp[4]) ? 4'b0110 : 4'b0111;
													assign node46010 = (inp[2]) ? node46014 : node46011;
														assign node46011 = (inp[4]) ? 4'b0111 : 4'b0110;
														assign node46014 = (inp[4]) ? 4'b0110 : 4'b0111;
											assign node46018 = (inp[1]) ? 4'b0111 : node46019;
												assign node46019 = (inp[0]) ? node46031 : node46020;
													assign node46020 = (inp[9]) ? node46026 : node46021;
														assign node46021 = (inp[2]) ? 4'b0110 : node46022;
															assign node46022 = (inp[4]) ? 4'b0110 : 4'b0111;
														assign node46026 = (inp[4]) ? 4'b0111 : node46027;
															assign node46027 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node46031 = (inp[10]) ? 4'b0110 : node46032;
														assign node46032 = (inp[2]) ? node46036 : node46033;
															assign node46033 = (inp[4]) ? 4'b0110 : 4'b0111;
															assign node46036 = (inp[4]) ? 4'b0111 : 4'b0110;
										assign node46041 = (inp[13]) ? node46051 : node46042;
											assign node46042 = (inp[1]) ? 4'b0111 : node46043;
												assign node46043 = (inp[4]) ? node46047 : node46044;
													assign node46044 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node46047 = (inp[2]) ? 4'b0111 : 4'b0110;
											assign node46051 = (inp[1]) ? 4'b0110 : node46052;
												assign node46052 = (inp[2]) ? node46056 : node46053;
													assign node46053 = (inp[4]) ? 4'b0111 : 4'b0110;
													assign node46056 = (inp[4]) ? 4'b0110 : 4'b0111;
									assign node46060 = (inp[10]) ? node46146 : node46061;
										assign node46061 = (inp[0]) ? node46099 : node46062;
											assign node46062 = (inp[13]) ? node46082 : node46063;
												assign node46063 = (inp[11]) ? node46073 : node46064;
													assign node46064 = (inp[2]) ? 4'b0010 : node46065;
														assign node46065 = (inp[4]) ? node46069 : node46066;
															assign node46066 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node46069 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node46073 = (inp[2]) ? 4'b0011 : node46074;
														assign node46074 = (inp[4]) ? node46078 : node46075;
															assign node46075 = (inp[1]) ? 4'b0010 : 4'b0011;
															assign node46078 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node46082 = (inp[11]) ? node46090 : node46083;
													assign node46083 = (inp[2]) ? 4'b0011 : node46084;
														assign node46084 = (inp[1]) ? 4'b0010 : node46085;
															assign node46085 = (inp[4]) ? 4'b0010 : 4'b0011;
													assign node46090 = (inp[2]) ? 4'b0010 : node46091;
														assign node46091 = (inp[4]) ? node46095 : node46092;
															assign node46092 = (inp[1]) ? 4'b0011 : 4'b0010;
															assign node46095 = (inp[1]) ? 4'b0010 : 4'b0011;
											assign node46099 = (inp[4]) ? node46123 : node46100;
												assign node46100 = (inp[11]) ? node46112 : node46101;
													assign node46101 = (inp[13]) ? node46107 : node46102;
														assign node46102 = (inp[1]) ? node46104 : 4'b0010;
															assign node46104 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node46107 = (inp[2]) ? 4'b0011 : node46108;
															assign node46108 = (inp[1]) ? 4'b0010 : 4'b0011;
													assign node46112 = (inp[13]) ? node46118 : node46113;
														assign node46113 = (inp[1]) ? node46115 : 4'b0011;
															assign node46115 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node46118 = (inp[2]) ? 4'b0010 : node46119;
															assign node46119 = (inp[1]) ? 4'b0011 : 4'b0010;
												assign node46123 = (inp[13]) ? node46135 : node46124;
													assign node46124 = (inp[11]) ? node46130 : node46125;
														assign node46125 = (inp[1]) ? 4'b0010 : node46126;
															assign node46126 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node46130 = (inp[2]) ? 4'b0011 : node46131;
															assign node46131 = (inp[1]) ? 4'b0011 : 4'b0010;
													assign node46135 = (inp[11]) ? node46141 : node46136;
														assign node46136 = (inp[1]) ? 4'b0011 : node46137;
															assign node46137 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node46141 = (inp[2]) ? 4'b0010 : node46142;
															assign node46142 = (inp[1]) ? 4'b0010 : 4'b0011;
										assign node46146 = (inp[1]) ? node46230 : node46147;
											assign node46147 = (inp[4]) ? node46185 : node46148;
												assign node46148 = (inp[9]) ? node46156 : node46149;
													assign node46149 = (inp[13]) ? node46153 : node46150;
														assign node46150 = (inp[11]) ? 4'b0011 : 4'b0010;
														assign node46153 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node46156 = (inp[0]) ? node46172 : node46157;
														assign node46157 = (inp[2]) ? node46165 : node46158;
															assign node46158 = (inp[13]) ? node46162 : node46159;
																assign node46159 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node46162 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node46165 = (inp[11]) ? node46169 : node46166;
																assign node46166 = (inp[13]) ? 4'b0011 : 4'b0010;
																assign node46169 = (inp[13]) ? 4'b0010 : 4'b0011;
														assign node46172 = (inp[2]) ? node46178 : node46173;
															assign node46173 = (inp[13]) ? 4'b0010 : node46174;
																assign node46174 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node46178 = (inp[13]) ? node46182 : node46179;
																assign node46179 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node46182 = (inp[11]) ? 4'b0010 : 4'b0011;
												assign node46185 = (inp[0]) ? node46215 : node46186;
													assign node46186 = (inp[9]) ? node46200 : node46187;
														assign node46187 = (inp[13]) ? node46193 : node46188;
															assign node46188 = (inp[2]) ? 4'b0010 : node46189;
																assign node46189 = (inp[11]) ? 4'b0010 : 4'b0011;
															assign node46193 = (inp[11]) ? node46197 : node46194;
																assign node46194 = (inp[2]) ? 4'b0011 : 4'b0010;
																assign node46197 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node46200 = (inp[2]) ? node46208 : node46201;
															assign node46201 = (inp[13]) ? node46205 : node46202;
																assign node46202 = (inp[11]) ? 4'b0010 : 4'b0011;
																assign node46205 = (inp[11]) ? 4'b0011 : 4'b0010;
															assign node46208 = (inp[13]) ? node46212 : node46209;
																assign node46209 = (inp[11]) ? 4'b0011 : 4'b0010;
																assign node46212 = (inp[11]) ? 4'b0010 : 4'b0011;
													assign node46215 = (inp[11]) ? node46223 : node46216;
														assign node46216 = (inp[13]) ? node46220 : node46217;
															assign node46217 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node46220 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node46223 = (inp[2]) ? node46227 : node46224;
															assign node46224 = (inp[13]) ? 4'b0011 : 4'b0010;
															assign node46227 = (inp[13]) ? 4'b0010 : 4'b0011;
											assign node46230 = (inp[9]) ? node46254 : node46231;
												assign node46231 = (inp[13]) ? node46243 : node46232;
													assign node46232 = (inp[11]) ? node46238 : node46233;
														assign node46233 = (inp[2]) ? 4'b0010 : node46234;
															assign node46234 = (inp[4]) ? 4'b0010 : 4'b0011;
														assign node46238 = (inp[2]) ? 4'b0011 : node46239;
															assign node46239 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node46243 = (inp[2]) ? 4'b0010 : node46244;
														assign node46244 = (inp[0]) ? 4'b0010 : node46245;
															assign node46245 = (inp[11]) ? node46249 : node46246;
																assign node46246 = (inp[4]) ? 4'b0011 : 4'b0010;
																assign node46249 = (inp[4]) ? 4'b0010 : 4'b0011;
												assign node46254 = (inp[13]) ? node46266 : node46255;
													assign node46255 = (inp[11]) ? node46261 : node46256;
														assign node46256 = (inp[4]) ? 4'b0010 : node46257;
															assign node46257 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node46261 = (inp[2]) ? 4'b0011 : node46262;
															assign node46262 = (inp[4]) ? 4'b0011 : 4'b0010;
													assign node46266 = (inp[11]) ? node46272 : node46267;
														assign node46267 = (inp[2]) ? 4'b0011 : node46268;
															assign node46268 = (inp[4]) ? 4'b0011 : 4'b0010;
														assign node46272 = (inp[4]) ? 4'b0010 : node46273;
															assign node46273 = (inp[2]) ? 4'b0010 : 4'b0011;
						assign node46277 = (inp[5]) ? node46611 : node46278;
							assign node46278 = (inp[2]) ? node46474 : node46279;
								assign node46279 = (inp[6]) ? node46467 : node46280;
									assign node46280 = (inp[13]) ? node46398 : node46281;
										assign node46281 = (inp[0]) ? node46337 : node46282;
											assign node46282 = (inp[11]) ? node46298 : node46283;
												assign node46283 = (inp[9]) ? node46291 : node46284;
													assign node46284 = (inp[10]) ? node46288 : node46285;
														assign node46285 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node46288 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node46291 = (inp[10]) ? node46295 : node46292;
														assign node46292 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node46295 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node46298 = (inp[9]) ? node46314 : node46299;
													assign node46299 = (inp[10]) ? node46307 : node46300;
														assign node46300 = (inp[4]) ? node46304 : node46301;
															assign node46301 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node46304 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node46307 = (inp[7]) ? node46311 : node46308;
															assign node46308 = (inp[4]) ? 4'b0000 : 4'b0001;
															assign node46311 = (inp[4]) ? 4'b0001 : 4'b0000;
													assign node46314 = (inp[1]) ? node46328 : node46315;
														assign node46315 = (inp[4]) ? node46321 : node46316;
															assign node46316 = (inp[7]) ? node46318 : 4'b0001;
																assign node46318 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node46321 = (inp[10]) ? node46325 : node46322;
																assign node46322 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node46325 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node46328 = (inp[4]) ? 4'b0001 : node46329;
															assign node46329 = (inp[10]) ? node46333 : node46330;
																assign node46330 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node46333 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node46337 = (inp[4]) ? node46367 : node46338;
												assign node46338 = (inp[11]) ? node46346 : node46339;
													assign node46339 = (inp[7]) ? node46343 : node46340;
														assign node46340 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node46343 = (inp[10]) ? 4'b0000 : 4'b0001;
													assign node46346 = (inp[1]) ? node46356 : node46347;
														assign node46347 = (inp[9]) ? 4'b0001 : node46348;
															assign node46348 = (inp[7]) ? node46352 : node46349;
																assign node46349 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node46352 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node46356 = (inp[9]) ? node46362 : node46357;
															assign node46357 = (inp[10]) ? node46359 : 4'b0001;
																assign node46359 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node46362 = (inp[10]) ? 4'b0000 : node46363;
																assign node46363 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node46367 = (inp[1]) ? node46385 : node46368;
													assign node46368 = (inp[11]) ? node46378 : node46369;
														assign node46369 = (inp[9]) ? node46371 : 4'b0001;
															assign node46371 = (inp[10]) ? node46375 : node46372;
																assign node46372 = (inp[7]) ? 4'b0001 : 4'b0000;
																assign node46375 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node46378 = (inp[7]) ? node46382 : node46379;
															assign node46379 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node46382 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node46385 = (inp[11]) ? node46391 : node46386;
														assign node46386 = (inp[10]) ? node46388 : 4'b0000;
															assign node46388 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node46391 = (inp[7]) ? node46395 : node46392;
															assign node46392 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node46395 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node46398 = (inp[4]) ? node46406 : node46399;
											assign node46399 = (inp[7]) ? node46403 : node46400;
												assign node46400 = (inp[10]) ? 4'b0001 : 4'b0000;
												assign node46403 = (inp[10]) ? 4'b0000 : 4'b0001;
											assign node46406 = (inp[9]) ? node46430 : node46407;
												assign node46407 = (inp[11]) ? node46415 : node46408;
													assign node46408 = (inp[10]) ? node46412 : node46409;
														assign node46409 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node46412 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node46415 = (inp[1]) ? node46423 : node46416;
														assign node46416 = (inp[10]) ? node46420 : node46417;
															assign node46417 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node46420 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node46423 = (inp[10]) ? node46427 : node46424;
															assign node46424 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node46427 = (inp[7]) ? 4'b0001 : 4'b0000;
												assign node46430 = (inp[1]) ? node46446 : node46431;
													assign node46431 = (inp[7]) ? node46439 : node46432;
														assign node46432 = (inp[11]) ? node46436 : node46433;
															assign node46433 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node46436 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node46439 = (inp[11]) ? node46443 : node46440;
															assign node46440 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node46443 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node46446 = (inp[11]) ? node46454 : node46447;
														assign node46447 = (inp[10]) ? node46451 : node46448;
															assign node46448 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node46451 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node46454 = (inp[0]) ? node46462 : node46455;
															assign node46455 = (inp[10]) ? node46459 : node46456;
																assign node46456 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node46459 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node46462 = (inp[7]) ? 4'b0001 : node46463;
																assign node46463 = (inp[10]) ? 4'b0000 : 4'b0001;
									assign node46467 = (inp[7]) ? node46471 : node46468;
										assign node46468 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node46471 = (inp[11]) ? 4'b0100 : 4'b0101;
								assign node46474 = (inp[11]) ? node46600 : node46475;
									assign node46475 = (inp[7]) ? node46559 : node46476;
										assign node46476 = (inp[6]) ? 4'b0100 : node46477;
											assign node46477 = (inp[9]) ? node46513 : node46478;
												assign node46478 = (inp[13]) ? node46498 : node46479;
													assign node46479 = (inp[0]) ? node46485 : node46480;
														assign node46480 = (inp[4]) ? 4'b0100 : node46481;
															assign node46481 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node46485 = (inp[1]) ? node46491 : node46486;
															assign node46486 = (inp[10]) ? 4'b0101 : node46487;
																assign node46487 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node46491 = (inp[10]) ? node46495 : node46492;
																assign node46492 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node46495 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node46498 = (inp[0]) ? node46506 : node46499;
														assign node46499 = (inp[4]) ? node46503 : node46500;
															assign node46500 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node46503 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node46506 = (inp[1]) ? 4'b0100 : node46507;
															assign node46507 = (inp[10]) ? 4'b0100 : node46508;
																assign node46508 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node46513 = (inp[0]) ? node46537 : node46514;
													assign node46514 = (inp[13]) ? node46522 : node46515;
														assign node46515 = (inp[10]) ? node46519 : node46516;
															assign node46516 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node46519 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node46522 = (inp[1]) ? node46530 : node46523;
															assign node46523 = (inp[10]) ? node46527 : node46524;
																assign node46524 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node46527 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node46530 = (inp[10]) ? node46534 : node46531;
																assign node46531 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node46534 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node46537 = (inp[13]) ? node46543 : node46538;
														assign node46538 = (inp[10]) ? node46540 : 4'b0101;
															assign node46540 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node46543 = (inp[1]) ? node46551 : node46544;
															assign node46544 = (inp[4]) ? node46548 : node46545;
																assign node46545 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node46548 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node46551 = (inp[4]) ? node46555 : node46552;
																assign node46552 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node46555 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node46559 = (inp[6]) ? 4'b0101 : node46560;
											assign node46560 = (inp[0]) ? node46592 : node46561;
												assign node46561 = (inp[13]) ? node46577 : node46562;
													assign node46562 = (inp[1]) ? node46570 : node46563;
														assign node46563 = (inp[4]) ? node46567 : node46564;
															assign node46564 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node46567 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node46570 = (inp[4]) ? node46574 : node46571;
															assign node46571 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node46574 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node46577 = (inp[9]) ? node46585 : node46578;
														assign node46578 = (inp[4]) ? node46582 : node46579;
															assign node46579 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node46582 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node46585 = (inp[4]) ? node46589 : node46586;
															assign node46586 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node46589 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node46592 = (inp[4]) ? node46596 : node46593;
													assign node46593 = (inp[10]) ? 4'b0100 : 4'b0101;
													assign node46596 = (inp[10]) ? 4'b0101 : 4'b0100;
									assign node46600 = (inp[7]) ? node46606 : node46601;
										assign node46601 = (inp[10]) ? 4'b0101 : node46602;
											assign node46602 = (inp[6]) ? 4'b0101 : 4'b0100;
										assign node46606 = (inp[6]) ? 4'b0100 : node46607;
											assign node46607 = (inp[10]) ? 4'b0100 : 4'b0101;
							assign node46611 = (inp[2]) ? node46771 : node46612;
								assign node46612 = (inp[6]) ? node46704 : node46613;
									assign node46613 = (inp[13]) ? node46629 : node46614;
										assign node46614 = (inp[11]) ? node46622 : node46615;
											assign node46615 = (inp[4]) ? node46619 : node46616;
												assign node46616 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node46619 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node46622 = (inp[4]) ? node46626 : node46623;
												assign node46623 = (inp[10]) ? 4'b0101 : 4'b0100;
												assign node46626 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node46629 = (inp[1]) ? node46653 : node46630;
											assign node46630 = (inp[0]) ? node46638 : node46631;
												assign node46631 = (inp[4]) ? node46635 : node46632;
													assign node46632 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node46635 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node46638 = (inp[7]) ? node46646 : node46639;
													assign node46639 = (inp[10]) ? node46643 : node46640;
														assign node46640 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node46643 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node46646 = (inp[4]) ? node46650 : node46647;
														assign node46647 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node46650 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node46653 = (inp[0]) ? node46677 : node46654;
												assign node46654 = (inp[7]) ? node46670 : node46655;
													assign node46655 = (inp[9]) ? node46663 : node46656;
														assign node46656 = (inp[10]) ? node46660 : node46657;
															assign node46657 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node46660 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node46663 = (inp[10]) ? node46667 : node46664;
															assign node46664 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node46667 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node46670 = (inp[10]) ? node46674 : node46671;
														assign node46671 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node46674 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node46677 = (inp[9]) ? node46699 : node46678;
													assign node46678 = (inp[11]) ? node46686 : node46679;
														assign node46679 = (inp[10]) ? node46683 : node46680;
															assign node46680 = (inp[4]) ? 4'b0101 : 4'b0100;
															assign node46683 = (inp[4]) ? 4'b0100 : 4'b0101;
														assign node46686 = (inp[7]) ? node46692 : node46687;
															assign node46687 = (inp[10]) ? node46689 : 4'b0100;
																assign node46689 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node46692 = (inp[10]) ? node46696 : node46693;
																assign node46693 = (inp[4]) ? 4'b0101 : 4'b0100;
																assign node46696 = (inp[4]) ? 4'b0100 : 4'b0101;
													assign node46699 = (inp[4]) ? node46701 : 4'b0100;
														assign node46701 = (inp[10]) ? 4'b0100 : 4'b0101;
									assign node46704 = (inp[10]) ? node46712 : node46705;
										assign node46705 = (inp[4]) ? node46709 : node46706;
											assign node46706 = (inp[11]) ? 4'b0001 : 4'b0000;
											assign node46709 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node46712 = (inp[1]) ? node46720 : node46713;
											assign node46713 = (inp[11]) ? node46717 : node46714;
												assign node46714 = (inp[4]) ? 4'b0001 : 4'b0000;
												assign node46717 = (inp[4]) ? 4'b0000 : 4'b0001;
											assign node46720 = (inp[13]) ? node46764 : node46721;
												assign node46721 = (inp[0]) ? node46749 : node46722;
													assign node46722 = (inp[7]) ? node46734 : node46723;
														assign node46723 = (inp[9]) ? node46729 : node46724;
															assign node46724 = (inp[11]) ? 4'b0000 : node46725;
																assign node46725 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node46729 = (inp[4]) ? 4'b0000 : node46730;
																assign node46730 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node46734 = (inp[9]) ? node46742 : node46735;
															assign node46735 = (inp[4]) ? node46739 : node46736;
																assign node46736 = (inp[11]) ? 4'b0001 : 4'b0000;
																assign node46739 = (inp[11]) ? 4'b0000 : 4'b0001;
															assign node46742 = (inp[11]) ? node46746 : node46743;
																assign node46743 = (inp[4]) ? 4'b0001 : 4'b0000;
																assign node46746 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node46749 = (inp[9]) ? node46757 : node46750;
														assign node46750 = (inp[11]) ? node46754 : node46751;
															assign node46751 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node46754 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node46757 = (inp[4]) ? node46761 : node46758;
															assign node46758 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node46761 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node46764 = (inp[4]) ? node46768 : node46765;
													assign node46765 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node46768 = (inp[11]) ? 4'b0000 : 4'b0001;
								assign node46771 = (inp[11]) ? node46777 : node46772;
									assign node46772 = (inp[10]) ? 4'b0001 : node46773;
										assign node46773 = (inp[6]) ? 4'b0001 : 4'b0000;
									assign node46777 = (inp[10]) ? 4'b0000 : node46778;
										assign node46778 = (inp[6]) ? 4'b0000 : 4'b0001;
					assign node46782 = (inp[15]) ? node47754 : node46783;
						assign node46783 = (inp[7]) ? node47279 : node46784;
							assign node46784 = (inp[6]) ? node47172 : node46785;
								assign node46785 = (inp[2]) ? node46975 : node46786;
									assign node46786 = (inp[5]) ? node46844 : node46787;
										assign node46787 = (inp[4]) ? node46811 : node46788;
											assign node46788 = (inp[10]) ? node46800 : node46789;
												assign node46789 = (inp[13]) ? node46795 : node46790;
													assign node46790 = (inp[11]) ? 4'b0101 : node46791;
														assign node46791 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node46795 = (inp[1]) ? 4'b0100 : node46796;
														assign node46796 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node46800 = (inp[13]) ? node46806 : node46801;
													assign node46801 = (inp[11]) ? 4'b0100 : node46802;
														assign node46802 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node46806 = (inp[1]) ? 4'b0101 : node46807;
														assign node46807 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node46811 = (inp[11]) ? node46819 : node46812;
												assign node46812 = (inp[13]) ? node46816 : node46813;
													assign node46813 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node46816 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node46819 = (inp[0]) ? node46835 : node46820;
													assign node46820 = (inp[13]) ? node46828 : node46821;
														assign node46821 = (inp[10]) ? node46825 : node46822;
															assign node46822 = (inp[1]) ? 4'b0001 : 4'b0000;
															assign node46825 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node46828 = (inp[1]) ? node46832 : node46829;
															assign node46829 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node46832 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node46835 = (inp[1]) ? node46837 : 4'b0000;
														assign node46837 = (inp[13]) ? node46841 : node46838;
															assign node46838 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node46841 = (inp[10]) ? 4'b0001 : 4'b0000;
										assign node46844 = (inp[9]) ? node46902 : node46845;
											assign node46845 = (inp[11]) ? node46863 : node46846;
												assign node46846 = (inp[10]) ? node46856 : node46847;
													assign node46847 = (inp[1]) ? node46849 : 4'b0001;
														assign node46849 = (inp[13]) ? node46853 : node46850;
															assign node46850 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node46853 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node46856 = (inp[4]) ? node46860 : node46857;
														assign node46857 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node46860 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node46863 = (inp[13]) ? node46879 : node46864;
													assign node46864 = (inp[4]) ? node46872 : node46865;
														assign node46865 = (inp[0]) ? node46867 : 4'b0000;
															assign node46867 = (inp[10]) ? 4'b0000 : node46868;
																assign node46868 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node46872 = (inp[1]) ? node46876 : node46873;
															assign node46873 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node46876 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node46879 = (inp[0]) ? node46893 : node46880;
														assign node46880 = (inp[10]) ? node46886 : node46881;
															assign node46881 = (inp[1]) ? node46883 : 4'b0000;
																assign node46883 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node46886 = (inp[4]) ? node46890 : node46887;
																assign node46887 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node46890 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node46893 = (inp[1]) ? node46895 : 4'b0001;
															assign node46895 = (inp[10]) ? node46899 : node46896;
																assign node46896 = (inp[4]) ? 4'b0001 : 4'b0000;
																assign node46899 = (inp[4]) ? 4'b0000 : 4'b0001;
											assign node46902 = (inp[10]) ? node46952 : node46903;
												assign node46903 = (inp[0]) ? node46931 : node46904;
													assign node46904 = (inp[11]) ? node46918 : node46905;
														assign node46905 = (inp[1]) ? node46913 : node46906;
															assign node46906 = (inp[4]) ? node46910 : node46907;
																assign node46907 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node46910 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node46913 = (inp[13]) ? 4'b0000 : node46914;
																assign node46914 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node46918 = (inp[4]) ? node46926 : node46919;
															assign node46919 = (inp[1]) ? node46923 : node46920;
																assign node46920 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node46923 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node46926 = (inp[13]) ? node46928 : 4'b0000;
																assign node46928 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node46931 = (inp[1]) ? node46939 : node46932;
														assign node46932 = (inp[13]) ? node46936 : node46933;
															assign node46933 = (inp[4]) ? 4'b0001 : 4'b0000;
															assign node46936 = (inp[4]) ? 4'b0000 : 4'b0001;
														assign node46939 = (inp[4]) ? node46945 : node46940;
															assign node46940 = (inp[13]) ? 4'b0000 : node46941;
																assign node46941 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node46945 = (inp[11]) ? node46949 : node46946;
																assign node46946 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node46949 = (inp[13]) ? 4'b0001 : 4'b0000;
												assign node46952 = (inp[1]) ? node46958 : node46953;
													assign node46953 = (inp[13]) ? 4'b0000 : node46954;
														assign node46954 = (inp[4]) ? 4'b0000 : 4'b0001;
													assign node46958 = (inp[13]) ? node46968 : node46959;
														assign node46959 = (inp[0]) ? node46961 : 4'b0000;
															assign node46961 = (inp[11]) ? node46965 : node46962;
																assign node46962 = (inp[4]) ? 4'b0000 : 4'b0001;
																assign node46965 = (inp[4]) ? 4'b0001 : 4'b0000;
														assign node46968 = (inp[4]) ? node46972 : node46969;
															assign node46969 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node46972 = (inp[11]) ? 4'b0000 : 4'b0001;
									assign node46975 = (inp[4]) ? node47085 : node46976;
										assign node46976 = (inp[5]) ? node47036 : node46977;
											assign node46977 = (inp[9]) ? node46999 : node46978;
												assign node46978 = (inp[13]) ? node46988 : node46979;
													assign node46979 = (inp[10]) ? node46985 : node46980;
														assign node46980 = (inp[11]) ? 4'b0000 : node46981;
															assign node46981 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node46985 = (inp[1]) ? 4'b0001 : 4'b0000;
													assign node46988 = (inp[10]) ? node46994 : node46989;
														assign node46989 = (inp[1]) ? 4'b0001 : node46990;
															assign node46990 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node46994 = (inp[1]) ? 4'b0000 : node46995;
															assign node46995 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node46999 = (inp[11]) ? node47021 : node47000;
													assign node47000 = (inp[1]) ? node47016 : node47001;
														assign node47001 = (inp[0]) ? node47009 : node47002;
															assign node47002 = (inp[10]) ? node47006 : node47003;
																assign node47003 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node47006 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node47009 = (inp[10]) ? node47013 : node47010;
																assign node47010 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node47013 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node47016 = (inp[13]) ? 4'b0001 : node47017;
															assign node47017 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node47021 = (inp[0]) ? node47029 : node47022;
														assign node47022 = (inp[13]) ? node47026 : node47023;
															assign node47023 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node47026 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node47029 = (inp[10]) ? node47033 : node47030;
															assign node47030 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node47033 = (inp[13]) ? 4'b0000 : 4'b0001;
											assign node47036 = (inp[9]) ? node47054 : node47037;
												assign node47037 = (inp[13]) ? node47043 : node47038;
													assign node47038 = (inp[10]) ? 4'b0101 : node47039;
														assign node47039 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node47043 = (inp[10]) ? node47049 : node47044;
														assign node47044 = (inp[11]) ? 4'b0101 : node47045;
															assign node47045 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node47049 = (inp[11]) ? 4'b0100 : node47050;
															assign node47050 = (inp[1]) ? 4'b0100 : 4'b0101;
												assign node47054 = (inp[11]) ? node47078 : node47055;
													assign node47055 = (inp[1]) ? node47063 : node47056;
														assign node47056 = (inp[13]) ? node47060 : node47057;
															assign node47057 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node47060 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node47063 = (inp[0]) ? node47071 : node47064;
															assign node47064 = (inp[10]) ? node47068 : node47065;
																assign node47065 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node47068 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node47071 = (inp[10]) ? node47075 : node47072;
																assign node47072 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node47075 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node47078 = (inp[13]) ? node47082 : node47079;
														assign node47079 = (inp[10]) ? 4'b0101 : 4'b0100;
														assign node47082 = (inp[10]) ? 4'b0100 : 4'b0101;
										assign node47085 = (inp[5]) ? node47149 : node47086;
											assign node47086 = (inp[9]) ? node47114 : node47087;
												assign node47087 = (inp[11]) ? node47107 : node47088;
													assign node47088 = (inp[1]) ? node47100 : node47089;
														assign node47089 = (inp[0]) ? node47095 : node47090;
															assign node47090 = (inp[10]) ? node47092 : 4'b0100;
																assign node47092 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node47095 = (inp[10]) ? 4'b0100 : node47096;
																assign node47096 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node47100 = (inp[13]) ? node47104 : node47101;
															assign node47101 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node47104 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node47107 = (inp[10]) ? node47111 : node47108;
														assign node47108 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node47111 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node47114 = (inp[0]) ? node47134 : node47115;
													assign node47115 = (inp[13]) ? node47127 : node47116;
														assign node47116 = (inp[10]) ? node47122 : node47117;
															assign node47117 = (inp[1]) ? 4'b0101 : node47118;
																assign node47118 = (inp[11]) ? 4'b0101 : 4'b0100;
															assign node47122 = (inp[1]) ? 4'b0100 : node47123;
																assign node47123 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node47127 = (inp[10]) ? node47129 : 4'b0100;
															assign node47129 = (inp[1]) ? 4'b0101 : node47130;
																assign node47130 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node47134 = (inp[13]) ? node47142 : node47135;
														assign node47135 = (inp[10]) ? 4'b0100 : node47136;
															assign node47136 = (inp[11]) ? 4'b0101 : node47137;
																assign node47137 = (inp[1]) ? 4'b0101 : 4'b0100;
														assign node47142 = (inp[10]) ? 4'b0101 : node47143;
															assign node47143 = (inp[1]) ? 4'b0100 : node47144;
																assign node47144 = (inp[11]) ? 4'b0100 : 4'b0101;
											assign node47149 = (inp[13]) ? node47161 : node47150;
												assign node47150 = (inp[10]) ? node47156 : node47151;
													assign node47151 = (inp[1]) ? 4'b0100 : node47152;
														assign node47152 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node47156 = (inp[11]) ? 4'b0101 : node47157;
														assign node47157 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node47161 = (inp[10]) ? node47167 : node47162;
													assign node47162 = (inp[1]) ? 4'b0101 : node47163;
														assign node47163 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node47167 = (inp[1]) ? 4'b0100 : node47168;
														assign node47168 = (inp[11]) ? 4'b0100 : 4'b0101;
								assign node47172 = (inp[1]) ? node47196 : node47173;
									assign node47173 = (inp[2]) ? node47185 : node47174;
										assign node47174 = (inp[13]) ? node47180 : node47175;
											assign node47175 = (inp[5]) ? node47177 : 4'b0100;
												assign node47177 = (inp[4]) ? 4'b0101 : 4'b0100;
											assign node47180 = (inp[4]) ? node47182 : 4'b0101;
												assign node47182 = (inp[5]) ? 4'b0100 : 4'b0101;
										assign node47185 = (inp[13]) ? node47191 : node47186;
											assign node47186 = (inp[4]) ? node47188 : 4'b0101;
												assign node47188 = (inp[5]) ? 4'b0101 : 4'b0100;
											assign node47191 = (inp[4]) ? node47193 : 4'b0100;
												assign node47193 = (inp[5]) ? 4'b0100 : 4'b0101;
									assign node47196 = (inp[9]) ? node47256 : node47197;
										assign node47197 = (inp[2]) ? node47249 : node47198;
											assign node47198 = (inp[5]) ? node47234 : node47199;
												assign node47199 = (inp[11]) ? node47221 : node47200;
													assign node47200 = (inp[0]) ? node47210 : node47201;
														assign node47201 = (inp[10]) ? node47205 : node47202;
															assign node47202 = (inp[13]) ? 4'b0100 : 4'b0101;
															assign node47205 = (inp[4]) ? node47207 : 4'b0101;
																assign node47207 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node47210 = (inp[10]) ? node47216 : node47211;
															assign node47211 = (inp[4]) ? node47213 : 4'b0101;
																assign node47213 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node47216 = (inp[13]) ? node47218 : 4'b0101;
																assign node47218 = (inp[4]) ? 4'b0101 : 4'b0100;
													assign node47221 = (inp[10]) ? node47229 : node47222;
														assign node47222 = (inp[13]) ? node47226 : node47223;
															assign node47223 = (inp[4]) ? 4'b0100 : 4'b0101;
															assign node47226 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node47229 = (inp[13]) ? node47231 : 4'b0100;
															assign node47231 = (inp[4]) ? 4'b0101 : 4'b0100;
												assign node47234 = (inp[0]) ? node47242 : node47235;
													assign node47235 = (inp[4]) ? node47239 : node47236;
														assign node47236 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node47239 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node47242 = (inp[13]) ? node47246 : node47243;
														assign node47243 = (inp[4]) ? 4'b0101 : 4'b0100;
														assign node47246 = (inp[4]) ? 4'b0100 : 4'b0101;
											assign node47249 = (inp[5]) ? node47253 : node47250;
												assign node47250 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node47253 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node47256 = (inp[5]) ? node47268 : node47257;
											assign node47257 = (inp[13]) ? node47263 : node47258;
												assign node47258 = (inp[2]) ? 4'b0100 : node47259;
													assign node47259 = (inp[4]) ? 4'b0100 : 4'b0101;
												assign node47263 = (inp[2]) ? 4'b0101 : node47264;
													assign node47264 = (inp[4]) ? 4'b0101 : 4'b0100;
											assign node47268 = (inp[13]) ? node47274 : node47269;
												assign node47269 = (inp[4]) ? 4'b0101 : node47270;
													assign node47270 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node47274 = (inp[2]) ? 4'b0100 : node47275;
													assign node47275 = (inp[4]) ? 4'b0100 : 4'b0101;
							assign node47279 = (inp[6]) ? node47727 : node47280;
								assign node47280 = (inp[2]) ? node47500 : node47281;
									assign node47281 = (inp[5]) ? node47377 : node47282;
										assign node47282 = (inp[4]) ? node47324 : node47283;
											assign node47283 = (inp[9]) ? node47303 : node47284;
												assign node47284 = (inp[13]) ? node47292 : node47285;
													assign node47285 = (inp[10]) ? 4'b0001 : node47286;
														assign node47286 = (inp[11]) ? 4'b0000 : node47287;
															assign node47287 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node47292 = (inp[10]) ? node47298 : node47293;
														assign node47293 = (inp[1]) ? 4'b0001 : node47294;
															assign node47294 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node47298 = (inp[1]) ? 4'b0000 : node47299;
															assign node47299 = (inp[11]) ? 4'b0000 : 4'b0001;
												assign node47303 = (inp[10]) ? node47315 : node47304;
													assign node47304 = (inp[13]) ? node47310 : node47305;
														assign node47305 = (inp[11]) ? 4'b0000 : node47306;
															assign node47306 = (inp[1]) ? 4'b0000 : 4'b0001;
														assign node47310 = (inp[1]) ? 4'b0001 : node47311;
															assign node47311 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node47315 = (inp[13]) ? node47319 : node47316;
														assign node47316 = (inp[11]) ? 4'b0001 : 4'b0000;
														assign node47319 = (inp[1]) ? 4'b0000 : node47320;
															assign node47320 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node47324 = (inp[9]) ? node47344 : node47325;
												assign node47325 = (inp[10]) ? node47337 : node47326;
													assign node47326 = (inp[13]) ? node47332 : node47327;
														assign node47327 = (inp[11]) ? 4'b0100 : node47328;
															assign node47328 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node47332 = (inp[11]) ? 4'b0101 : node47333;
															assign node47333 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node47337 = (inp[13]) ? 4'b0100 : node47338;
														assign node47338 = (inp[1]) ? 4'b0101 : node47339;
															assign node47339 = (inp[11]) ? 4'b0101 : 4'b0100;
												assign node47344 = (inp[0]) ? node47356 : node47345;
													assign node47345 = (inp[10]) ? node47353 : node47346;
														assign node47346 = (inp[13]) ? 4'b0101 : node47347;
															assign node47347 = (inp[11]) ? 4'b0100 : node47348;
																assign node47348 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node47353 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node47356 = (inp[1]) ? node47370 : node47357;
														assign node47357 = (inp[10]) ? node47363 : node47358;
															assign node47358 = (inp[11]) ? node47360 : 4'b0101;
																assign node47360 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node47363 = (inp[11]) ? node47367 : node47364;
																assign node47364 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node47367 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node47370 = (inp[10]) ? node47374 : node47371;
															assign node47371 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node47374 = (inp[13]) ? 4'b0100 : 4'b0101;
										assign node47377 = (inp[4]) ? node47445 : node47378;
											assign node47378 = (inp[0]) ? node47402 : node47379;
												assign node47379 = (inp[13]) ? node47391 : node47380;
													assign node47380 = (inp[10]) ? node47386 : node47381;
														assign node47381 = (inp[1]) ? 4'b0101 : node47382;
															assign node47382 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node47386 = (inp[11]) ? 4'b0100 : node47387;
															assign node47387 = (inp[1]) ? 4'b0100 : 4'b0101;
													assign node47391 = (inp[10]) ? node47397 : node47392;
														assign node47392 = (inp[11]) ? 4'b0100 : node47393;
															assign node47393 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node47397 = (inp[11]) ? 4'b0101 : node47398;
															assign node47398 = (inp[1]) ? 4'b0101 : 4'b0100;
												assign node47402 = (inp[9]) ? node47424 : node47403;
													assign node47403 = (inp[13]) ? node47415 : node47404;
														assign node47404 = (inp[10]) ? node47410 : node47405;
															assign node47405 = (inp[11]) ? 4'b0101 : node47406;
																assign node47406 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node47410 = (inp[1]) ? 4'b0100 : node47411;
																assign node47411 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node47415 = (inp[10]) ? node47419 : node47416;
															assign node47416 = (inp[1]) ? 4'b0100 : 4'b0101;
															assign node47419 = (inp[11]) ? 4'b0101 : node47420;
																assign node47420 = (inp[1]) ? 4'b0101 : 4'b0100;
													assign node47424 = (inp[10]) ? node47436 : node47425;
														assign node47425 = (inp[13]) ? node47431 : node47426;
															assign node47426 = (inp[11]) ? 4'b0101 : node47427;
																assign node47427 = (inp[1]) ? 4'b0101 : 4'b0100;
															assign node47431 = (inp[1]) ? 4'b0100 : node47432;
																assign node47432 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node47436 = (inp[13]) ? node47440 : node47437;
															assign node47437 = (inp[11]) ? 4'b0100 : 4'b0101;
															assign node47440 = (inp[1]) ? 4'b0101 : node47441;
																assign node47441 = (inp[11]) ? 4'b0101 : 4'b0100;
											assign node47445 = (inp[1]) ? node47469 : node47446;
												assign node47446 = (inp[11]) ? node47454 : node47447;
													assign node47447 = (inp[13]) ? node47451 : node47448;
														assign node47448 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node47451 = (inp[10]) ? 4'b0101 : 4'b0100;
													assign node47454 = (inp[0]) ? node47462 : node47455;
														assign node47455 = (inp[13]) ? node47459 : node47456;
															assign node47456 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node47459 = (inp[10]) ? 4'b0100 : 4'b0101;
														assign node47462 = (inp[10]) ? node47466 : node47463;
															assign node47463 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node47466 = (inp[13]) ? 4'b0100 : 4'b0101;
												assign node47469 = (inp[9]) ? node47477 : node47470;
													assign node47470 = (inp[10]) ? node47474 : node47471;
														assign node47471 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node47474 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node47477 = (inp[11]) ? node47485 : node47478;
														assign node47478 = (inp[10]) ? node47482 : node47479;
															assign node47479 = (inp[13]) ? 4'b0101 : 4'b0100;
															assign node47482 = (inp[13]) ? 4'b0100 : 4'b0101;
														assign node47485 = (inp[0]) ? node47493 : node47486;
															assign node47486 = (inp[13]) ? node47490 : node47487;
																assign node47487 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node47490 = (inp[10]) ? 4'b0100 : 4'b0101;
															assign node47493 = (inp[13]) ? node47497 : node47494;
																assign node47494 = (inp[10]) ? 4'b0101 : 4'b0100;
																assign node47497 = (inp[10]) ? 4'b0100 : 4'b0101;
									assign node47500 = (inp[5]) ? node47626 : node47501;
										assign node47501 = (inp[4]) ? node47539 : node47502;
											assign node47502 = (inp[11]) ? node47510 : node47503;
												assign node47503 = (inp[10]) ? node47507 : node47504;
													assign node47504 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node47507 = (inp[13]) ? 4'b0101 : 4'b0100;
												assign node47510 = (inp[9]) ? node47526 : node47511;
													assign node47511 = (inp[10]) ? node47517 : node47512;
														assign node47512 = (inp[1]) ? node47514 : 4'b0101;
															assign node47514 = (inp[13]) ? 4'b0101 : 4'b0100;
														assign node47517 = (inp[0]) ? 4'b0101 : node47518;
															assign node47518 = (inp[1]) ? node47522 : node47519;
																assign node47519 = (inp[13]) ? 4'b0101 : 4'b0100;
																assign node47522 = (inp[13]) ? 4'b0100 : 4'b0101;
													assign node47526 = (inp[13]) ? node47532 : node47527;
														assign node47527 = (inp[10]) ? 4'b0101 : node47528;
															assign node47528 = (inp[1]) ? 4'b0100 : 4'b0101;
														assign node47532 = (inp[1]) ? node47536 : node47533;
															assign node47533 = (inp[10]) ? 4'b0101 : 4'b0100;
															assign node47536 = (inp[10]) ? 4'b0100 : 4'b0101;
											assign node47539 = (inp[0]) ? node47591 : node47540;
												assign node47540 = (inp[11]) ? node47570 : node47541;
													assign node47541 = (inp[9]) ? node47555 : node47542;
														assign node47542 = (inp[13]) ? node47550 : node47543;
															assign node47543 = (inp[1]) ? node47547 : node47544;
																assign node47544 = (inp[10]) ? 4'b0000 : 4'b0001;
																assign node47547 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node47550 = (inp[1]) ? 4'b0001 : node47551;
																assign node47551 = (inp[10]) ? 4'b0001 : 4'b0000;
														assign node47555 = (inp[10]) ? node47563 : node47556;
															assign node47556 = (inp[1]) ? node47560 : node47557;
																assign node47557 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node47560 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node47563 = (inp[13]) ? node47567 : node47564;
																assign node47564 = (inp[1]) ? 4'b0001 : 4'b0000;
																assign node47567 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node47570 = (inp[9]) ? node47584 : node47571;
														assign node47571 = (inp[1]) ? node47577 : node47572;
															assign node47572 = (inp[10]) ? node47574 : 4'b0001;
																assign node47574 = (inp[13]) ? 4'b0000 : 4'b0001;
															assign node47577 = (inp[13]) ? node47581 : node47578;
																assign node47578 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node47581 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node47584 = (inp[13]) ? node47588 : node47585;
															assign node47585 = (inp[10]) ? 4'b0001 : 4'b0000;
															assign node47588 = (inp[10]) ? 4'b0000 : 4'b0001;
												assign node47591 = (inp[9]) ? node47605 : node47592;
													assign node47592 = (inp[13]) ? node47600 : node47593;
														assign node47593 = (inp[10]) ? 4'b0001 : node47594;
															assign node47594 = (inp[1]) ? 4'b0000 : node47595;
																assign node47595 = (inp[11]) ? 4'b0000 : 4'b0001;
														assign node47600 = (inp[10]) ? 4'b0000 : node47601;
															assign node47601 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node47605 = (inp[13]) ? node47615 : node47606;
														assign node47606 = (inp[11]) ? 4'b0000 : node47607;
															assign node47607 = (inp[10]) ? node47611 : node47608;
																assign node47608 = (inp[1]) ? 4'b0000 : 4'b0001;
																assign node47611 = (inp[1]) ? 4'b0001 : 4'b0000;
														assign node47615 = (inp[10]) ? node47621 : node47616;
															assign node47616 = (inp[1]) ? 4'b0001 : node47617;
																assign node47617 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node47621 = (inp[1]) ? 4'b0000 : node47622;
																assign node47622 = (inp[11]) ? 4'b0000 : 4'b0001;
										assign node47626 = (inp[9]) ? node47704 : node47627;
											assign node47627 = (inp[1]) ? node47665 : node47628;
												assign node47628 = (inp[10]) ? node47658 : node47629;
													assign node47629 = (inp[4]) ? node47643 : node47630;
														assign node47630 = (inp[0]) ? node47636 : node47631;
															assign node47631 = (inp[11]) ? node47633 : 4'b0000;
																assign node47633 = (inp[13]) ? 4'b0001 : 4'b0000;
															assign node47636 = (inp[11]) ? node47640 : node47637;
																assign node47637 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node47640 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node47643 = (inp[0]) ? node47651 : node47644;
															assign node47644 = (inp[13]) ? node47648 : node47645;
																assign node47645 = (inp[11]) ? 4'b0000 : 4'b0001;
																assign node47648 = (inp[11]) ? 4'b0001 : 4'b0000;
															assign node47651 = (inp[11]) ? node47655 : node47652;
																assign node47652 = (inp[13]) ? 4'b0000 : 4'b0001;
																assign node47655 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node47658 = (inp[11]) ? node47662 : node47659;
														assign node47659 = (inp[13]) ? 4'b0001 : 4'b0000;
														assign node47662 = (inp[13]) ? 4'b0000 : 4'b0001;
												assign node47665 = (inp[0]) ? node47685 : node47666;
													assign node47666 = (inp[4]) ? node47676 : node47667;
														assign node47667 = (inp[11]) ? node47669 : 4'b0000;
															assign node47669 = (inp[13]) ? node47673 : node47670;
																assign node47670 = (inp[10]) ? 4'b0001 : 4'b0000;
																assign node47673 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node47676 = (inp[11]) ? node47682 : node47677;
															assign node47677 = (inp[13]) ? node47679 : 4'b0001;
																assign node47679 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node47682 = (inp[13]) ? 4'b0001 : 4'b0000;
													assign node47685 = (inp[11]) ? node47699 : node47686;
														assign node47686 = (inp[4]) ? node47692 : node47687;
															assign node47687 = (inp[13]) ? node47689 : 4'b0000;
																assign node47689 = (inp[10]) ? 4'b0000 : 4'b0001;
															assign node47692 = (inp[10]) ? node47696 : node47693;
																assign node47693 = (inp[13]) ? 4'b0001 : 4'b0000;
																assign node47696 = (inp[13]) ? 4'b0000 : 4'b0001;
														assign node47699 = (inp[13]) ? 4'b0000 : node47700;
															assign node47700 = (inp[10]) ? 4'b0001 : 4'b0000;
											assign node47704 = (inp[10]) ? node47716 : node47705;
												assign node47705 = (inp[13]) ? node47711 : node47706;
													assign node47706 = (inp[11]) ? 4'b0000 : node47707;
														assign node47707 = (inp[1]) ? 4'b0000 : 4'b0001;
													assign node47711 = (inp[1]) ? 4'b0001 : node47712;
														assign node47712 = (inp[11]) ? 4'b0001 : 4'b0000;
												assign node47716 = (inp[13]) ? node47722 : node47717;
													assign node47717 = (inp[1]) ? 4'b0001 : node47718;
														assign node47718 = (inp[11]) ? 4'b0001 : 4'b0000;
													assign node47722 = (inp[11]) ? 4'b0000 : node47723;
														assign node47723 = (inp[1]) ? 4'b0000 : 4'b0001;
								assign node47727 = (inp[13]) ? node47741 : node47728;
									assign node47728 = (inp[4]) ? 4'b0001 : node47729;
										assign node47729 = (inp[2]) ? node47735 : node47730;
											assign node47730 = (inp[5]) ? 4'b0000 : node47731;
												assign node47731 = (inp[1]) ? 4'b0000 : 4'b0001;
											assign node47735 = (inp[1]) ? 4'b0001 : node47736;
												assign node47736 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node47741 = (inp[4]) ? 4'b0000 : node47742;
										assign node47742 = (inp[2]) ? node47748 : node47743;
											assign node47743 = (inp[5]) ? 4'b0001 : node47744;
												assign node47744 = (inp[1]) ? 4'b0001 : 4'b0000;
											assign node47748 = (inp[1]) ? 4'b0000 : node47749;
												assign node47749 = (inp[5]) ? 4'b0000 : 4'b0001;
						assign node47754 = (inp[2]) ? node47830 : node47755;
							assign node47755 = (inp[6]) ? node47819 : node47756;
								assign node47756 = (inp[10]) ? node47788 : node47757;
									assign node47757 = (inp[4]) ? node47783 : node47758;
										assign node47758 = (inp[5]) ? 4'b0100 : node47759;
											assign node47759 = (inp[13]) ? node47767 : node47760;
												assign node47760 = (inp[7]) ? node47764 : node47761;
													assign node47761 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node47764 = (inp[11]) ? 4'b0100 : 4'b0101;
												assign node47767 = (inp[1]) ? node47775 : node47768;
													assign node47768 = (inp[7]) ? node47772 : node47769;
														assign node47769 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node47772 = (inp[11]) ? 4'b0100 : 4'b0101;
													assign node47775 = (inp[7]) ? node47779 : node47776;
														assign node47776 = (inp[11]) ? 4'b0101 : 4'b0100;
														assign node47779 = (inp[11]) ? 4'b0100 : 4'b0101;
										assign node47783 = (inp[5]) ? 4'b0101 : node47784;
											assign node47784 = (inp[7]) ? 4'b0101 : 4'b0100;
									assign node47788 = (inp[4]) ? node47814 : node47789;
										assign node47789 = (inp[5]) ? 4'b0101 : node47790;
											assign node47790 = (inp[9]) ? node47798 : node47791;
												assign node47791 = (inp[11]) ? node47795 : node47792;
													assign node47792 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node47795 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node47798 = (inp[13]) ? node47806 : node47799;
													assign node47799 = (inp[7]) ? node47803 : node47800;
														assign node47800 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node47803 = (inp[11]) ? 4'b0101 : 4'b0100;
													assign node47806 = (inp[7]) ? node47810 : node47807;
														assign node47807 = (inp[11]) ? 4'b0100 : 4'b0101;
														assign node47810 = (inp[11]) ? 4'b0101 : 4'b0100;
										assign node47814 = (inp[5]) ? 4'b0100 : node47815;
											assign node47815 = (inp[7]) ? 4'b0100 : 4'b0101;
								assign node47819 = (inp[4]) ? node47825 : node47820;
									assign node47820 = (inp[7]) ? 4'b0001 : node47821;
										assign node47821 = (inp[5]) ? 4'b0001 : 4'b0000;
									assign node47825 = (inp[5]) ? 4'b0000 : node47826;
										assign node47826 = (inp[7]) ? 4'b0000 : 4'b0001;
							assign node47830 = (inp[10]) ? node47850 : node47831;
								assign node47831 = (inp[6]) ? node47845 : node47832;
									assign node47832 = (inp[5]) ? 4'b0001 : node47833;
										assign node47833 = (inp[7]) ? node47839 : node47834;
											assign node47834 = (inp[4]) ? 4'b0000 : node47835;
												assign node47835 = (inp[11]) ? 4'b0000 : 4'b0001;
											assign node47839 = (inp[11]) ? 4'b0001 : node47840;
												assign node47840 = (inp[4]) ? 4'b0001 : 4'b0000;
									assign node47845 = (inp[5]) ? 4'b0000 : node47846;
										assign node47846 = (inp[7]) ? 4'b0000 : 4'b0001;
								assign node47850 = (inp[5]) ? 4'b0000 : node47851;
									assign node47851 = (inp[7]) ? node47859 : node47852;
										assign node47852 = (inp[11]) ? 4'b0001 : node47853;
											assign node47853 = (inp[6]) ? 4'b0001 : node47854;
												assign node47854 = (inp[4]) ? 4'b0001 : 4'b0000;
										assign node47859 = (inp[6]) ? 4'b0000 : node47860;
											assign node47860 = (inp[4]) ? 4'b0000 : node47861;
												assign node47861 = (inp[11]) ? 4'b0000 : 4'b0001;

endmodule