module dtc_split125_bm89 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node42;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node137;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node172;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node364;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node370;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node387;

	assign outp = (inp[3]) ? node222 : node1;
		assign node1 = (inp[6]) ? node97 : node2;
			assign node2 = (inp[7]) ? node36 : node3;
				assign node3 = (inp[9]) ? 3'b111 : node4;
					assign node4 = (inp[4]) ? node12 : node5;
						assign node5 = (inp[10]) ? 3'b111 : node6;
							assign node6 = (inp[5]) ? node8 : 3'b101;
								assign node8 = (inp[11]) ? 3'b101 : 3'b011;
						assign node12 = (inp[10]) ? node20 : node13;
							assign node13 = (inp[5]) ? node15 : 3'b010;
								assign node15 = (inp[11]) ? node17 : 3'b100;
									assign node17 = (inp[0]) ? 3'b110 : 3'b010;
							assign node20 = (inp[0]) ? node24 : node21;
								assign node21 = (inp[1]) ? 3'b110 : 3'b001;
								assign node24 = (inp[11]) ? node30 : node25;
									assign node25 = (inp[5]) ? 3'b001 : node26;
										assign node26 = (inp[8]) ? 3'b001 : 3'b101;
									assign node30 = (inp[1]) ? 3'b101 : node31;
										assign node31 = (inp[5]) ? 3'b001 : 3'b101;
				assign node36 = (inp[10]) ? node76 : node37;
					assign node37 = (inp[1]) ? node59 : node38;
						assign node38 = (inp[0]) ? node56 : node39;
							assign node39 = (inp[11]) ? node45 : node40;
								assign node40 = (inp[2]) ? node42 : 3'b110;
									assign node42 = (inp[8]) ? 3'b111 : 3'b000;
								assign node45 = (inp[8]) ? node53 : node46;
									assign node46 = (inp[4]) ? node50 : node47;
										assign node47 = (inp[2]) ? 3'b111 : 3'b110;
										assign node50 = (inp[9]) ? 3'b011 : 3'b010;
									assign node53 = (inp[9]) ? 3'b111 : 3'b001;
							assign node56 = (inp[9]) ? 3'b001 : 3'b100;
						assign node59 = (inp[5]) ? node67 : node60;
							assign node60 = (inp[8]) ? node64 : node61;
								assign node61 = (inp[4]) ? 3'b100 : 3'b110;
								assign node64 = (inp[9]) ? 3'b000 : 3'b100;
							assign node67 = (inp[8]) ? node69 : 3'b000;
								assign node69 = (inp[4]) ? node71 : 3'b110;
									assign node71 = (inp[11]) ? 3'b001 : node72;
										assign node72 = (inp[9]) ? 3'b110 : 3'b000;
					assign node76 = (inp[4]) ? node84 : node77;
						assign node77 = (inp[9]) ? 3'b100 : node78;
							assign node78 = (inp[11]) ? node80 : 3'b101;
								assign node80 = (inp[1]) ? 3'b011 : 3'b101;
						assign node84 = (inp[2]) ? node90 : node85;
							assign node85 = (inp[9]) ? node87 : 3'b110;
								assign node87 = (inp[0]) ? 3'b011 : 3'b001;
							assign node90 = (inp[1]) ? node94 : node91;
								assign node91 = (inp[0]) ? 3'b001 : 3'b011;
								assign node94 = (inp[11]) ? 3'b001 : 3'b101;
			assign node97 = (inp[9]) ? node133 : node98;
				assign node98 = (inp[4]) ? node126 : node99;
					assign node99 = (inp[10]) ? node111 : node100;
						assign node100 = (inp[7]) ? 3'b000 : node101;
							assign node101 = (inp[11]) ? node105 : node102;
								assign node102 = (inp[5]) ? 3'b000 : 3'b100;
								assign node105 = (inp[8]) ? 3'b100 : node106;
									assign node106 = (inp[5]) ? 3'b010 : 3'b110;
						assign node111 = (inp[11]) ? node115 : node112;
							assign node112 = (inp[7]) ? 3'b100 : 3'b110;
							assign node115 = (inp[5]) ? node119 : node116;
								assign node116 = (inp[1]) ? 3'b101 : 3'b001;
								assign node119 = (inp[0]) ? node123 : node120;
									assign node120 = (inp[2]) ? 3'b011 : 3'b110;
									assign node123 = (inp[1]) ? 3'b100 : 3'b010;
					assign node126 = (inp[2]) ? 3'b000 : node127;
						assign node127 = (inp[10]) ? node129 : 3'b000;
							assign node129 = (inp[7]) ? 3'b000 : 3'b100;
				assign node133 = (inp[4]) ? node177 : node134;
					assign node134 = (inp[7]) ? node150 : node135;
						assign node135 = (inp[10]) ? 3'b011 : node136;
							assign node136 = (inp[1]) ? node144 : node137;
								assign node137 = (inp[11]) ? node139 : 3'b011;
									assign node139 = (inp[5]) ? 3'b001 : node140;
										assign node140 = (inp[0]) ? 3'b001 : 3'b011;
								assign node144 = (inp[11]) ? node146 : 3'b001;
									assign node146 = (inp[8]) ? 3'b001 : 3'b011;
						assign node150 = (inp[8]) ? node164 : node151;
							assign node151 = (inp[5]) ? node157 : node152;
								assign node152 = (inp[11]) ? node154 : 3'b001;
									assign node154 = (inp[2]) ? 3'b111 : 3'b011;
								assign node157 = (inp[10]) ? node161 : node158;
									assign node158 = (inp[1]) ? 3'b110 : 3'b011;
									assign node161 = (inp[11]) ? 3'b101 : 3'b111;
							assign node164 = (inp[10]) ? node170 : node165;
								assign node165 = (inp[5]) ? node167 : 3'b010;
									assign node167 = (inp[1]) ? 3'b100 : 3'b000;
								assign node170 = (inp[2]) ? node172 : 3'b110;
									assign node172 = (inp[5]) ? node174 : 3'b001;
										assign node174 = (inp[11]) ? 3'b001 : 3'b110;
					assign node177 = (inp[10]) ? node195 : node178;
						assign node178 = (inp[7]) ? node188 : node179;
							assign node179 = (inp[11]) ? node181 : 3'b100;
								assign node181 = (inp[1]) ? node185 : node182;
									assign node182 = (inp[2]) ? 3'b110 : 3'b101;
									assign node185 = (inp[8]) ? 3'b010 : 3'b110;
							assign node188 = (inp[5]) ? 3'b000 : node189;
								assign node189 = (inp[8]) ? node191 : 3'b010;
									assign node191 = (inp[0]) ? 3'b100 : 3'b110;
						assign node195 = (inp[11]) ? node213 : node196;
							assign node196 = (inp[7]) ? node204 : node197;
								assign node197 = (inp[8]) ? node199 : 3'b101;
									assign node199 = (inp[5]) ? 3'b001 : node200;
										assign node200 = (inp[0]) ? 3'b001 : 3'b110;
								assign node204 = (inp[2]) ? node210 : node205;
									assign node205 = (inp[8]) ? node207 : 3'b110;
										assign node207 = (inp[0]) ? 3'b100 : 3'b110;
									assign node210 = (inp[5]) ? 3'b010 : 3'b110;
							assign node213 = (inp[5]) ? node215 : 3'b001;
								assign node215 = (inp[8]) ? node219 : node216;
									assign node216 = (inp[0]) ? 3'b110 : 3'b101;
									assign node219 = (inp[0]) ? 3'b001 : 3'b101;
		assign node222 = (inp[6]) ? node344 : node223;
			assign node223 = (inp[9]) ? node275 : node224;
				assign node224 = (inp[7]) ? node264 : node225;
					assign node225 = (inp[5]) ? node241 : node226;
						assign node226 = (inp[10]) ? node232 : node227;
							assign node227 = (inp[1]) ? node229 : 3'b000;
								assign node229 = (inp[0]) ? 3'b100 : 3'b000;
							assign node232 = (inp[4]) ? 3'b100 : node233;
								assign node233 = (inp[1]) ? node235 : 3'b101;
									assign node235 = (inp[0]) ? 3'b001 : node236;
										assign node236 = (inp[2]) ? 3'b101 : 3'b001;
						assign node241 = (inp[8]) ? node259 : node242;
							assign node242 = (inp[4]) ? node254 : node243;
								assign node243 = (inp[10]) ? node249 : node244;
									assign node244 = (inp[11]) ? 3'b010 : node245;
										assign node245 = (inp[1]) ? 3'b000 : 3'b100;
									assign node249 = (inp[11]) ? node251 : 3'b110;
										assign node251 = (inp[1]) ? 3'b100 : 3'b011;
								assign node254 = (inp[0]) ? 3'b000 : node255;
									assign node255 = (inp[1]) ? 3'b000 : 3'b100;
							assign node259 = (inp[11]) ? node261 : 3'b000;
								assign node261 = (inp[4]) ? 3'b000 : 3'b100;
					assign node264 = (inp[10]) ? node266 : 3'b000;
						assign node266 = (inp[4]) ? 3'b000 : node267;
							assign node267 = (inp[8]) ? node271 : node268;
								assign node268 = (inp[1]) ? 3'b010 : 3'b100;
								assign node271 = (inp[0]) ? 3'b100 : 3'b000;
				assign node275 = (inp[4]) ? node309 : node276;
					assign node276 = (inp[7]) ? node290 : node277;
						assign node277 = (inp[10]) ? 3'b111 : node278;
							assign node278 = (inp[1]) ? node284 : node279;
								assign node279 = (inp[11]) ? 3'b011 : node280;
									assign node280 = (inp[0]) ? 3'b101 : 3'b011;
								assign node284 = (inp[11]) ? 3'b101 : node285;
									assign node285 = (inp[5]) ? 3'b011 : 3'b101;
						assign node290 = (inp[10]) ? node300 : node291;
							assign node291 = (inp[2]) ? node297 : node292;
								assign node292 = (inp[11]) ? node294 : 3'b110;
									assign node294 = (inp[0]) ? 3'b011 : 3'b001;
								assign node297 = (inp[8]) ? 3'b110 : 3'b010;
							assign node300 = (inp[1]) ? node304 : node301;
								assign node301 = (inp[11]) ? 3'b101 : 3'b001;
								assign node304 = (inp[5]) ? node306 : 3'b101;
									assign node306 = (inp[0]) ? 3'b001 : 3'b101;
					assign node309 = (inp[10]) ? node323 : node310;
						assign node310 = (inp[8]) ? node318 : node311;
							assign node311 = (inp[11]) ? node315 : node312;
								assign node312 = (inp[7]) ? 3'b000 : 3'b010;
								assign node315 = (inp[0]) ? 3'b110 : 3'b010;
							assign node318 = (inp[0]) ? 3'b110 : node319;
								assign node319 = (inp[2]) ? 3'b000 : 3'b100;
						assign node323 = (inp[7]) ? node333 : node324;
							assign node324 = (inp[5]) ? 3'b001 : node325;
								assign node325 = (inp[1]) ? node329 : node326;
									assign node326 = (inp[11]) ? 3'b011 : 3'b101;
									assign node329 = (inp[11]) ? 3'b101 : 3'b001;
							assign node333 = (inp[11]) ? node341 : node334;
								assign node334 = (inp[5]) ? node336 : 3'b010;
									assign node336 = (inp[0]) ? 3'b100 : node337;
										assign node337 = (inp[8]) ? 3'b010 : 3'b110;
								assign node341 = (inp[8]) ? 3'b110 : 3'b001;
			assign node344 = (inp[9]) ? node346 : 3'b000;
				assign node346 = (inp[10]) ? node354 : node347;
					assign node347 = (inp[7]) ? 3'b000 : node348;
						assign node348 = (inp[4]) ? 3'b000 : node349;
							assign node349 = (inp[11]) ? 3'b110 : 3'b000;
					assign node354 = (inp[7]) ? node380 : node355;
						assign node355 = (inp[8]) ? node367 : node356;
							assign node356 = (inp[11]) ? node364 : node357;
								assign node357 = (inp[4]) ? 3'b100 : node358;
									assign node358 = (inp[0]) ? 3'b110 : node359;
										assign node359 = (inp[5]) ? 3'b110 : 3'b010;
								assign node364 = (inp[4]) ? 3'b010 : 3'b110;
							assign node367 = (inp[0]) ? node373 : node368;
								assign node368 = (inp[4]) ? node370 : 3'b110;
									assign node370 = (inp[5]) ? 3'b100 : 3'b110;
								assign node373 = (inp[2]) ? 3'b000 : node374;
									assign node374 = (inp[4]) ? 3'b000 : node375;
										assign node375 = (inp[11]) ? 3'b000 : 3'b110;
						assign node380 = (inp[4]) ? 3'b000 : node381;
							assign node381 = (inp[11]) ? node385 : node382;
								assign node382 = (inp[5]) ? 3'b000 : 3'b100;
								assign node385 = (inp[8]) ? node387 : 3'b010;
									assign node387 = (inp[1]) ? 3'b100 : 3'b010;

endmodule