module dtc_split875_bm68 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node61;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node124;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node130;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node145;
	wire [3-1:0] node147;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node248;
	wire [3-1:0] node252;
	wire [3-1:0] node254;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node268;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node307;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node351;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node362;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node418;
	wire [3-1:0] node420;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node430;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node447;
	wire [3-1:0] node449;
	wire [3-1:0] node453;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node459;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node477;
	wire [3-1:0] node479;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node488;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node502;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node510;
	wire [3-1:0] node512;
	wire [3-1:0] node514;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node521;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node532;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node542;
	wire [3-1:0] node544;
	wire [3-1:0] node546;
	wire [3-1:0] node549;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node565;
	wire [3-1:0] node567;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node594;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node599;
	wire [3-1:0] node604;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node624;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node633;
	wire [3-1:0] node635;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node640;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node661;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node685;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node690;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node700;
	wire [3-1:0] node701;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node714;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node729;
	wire [3-1:0] node734;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node772;
	wire [3-1:0] node774;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node790;
	wire [3-1:0] node791;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node825;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node838;
	wire [3-1:0] node839;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node851;
	wire [3-1:0] node853;
	wire [3-1:0] node854;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node864;
	wire [3-1:0] node866;
	wire [3-1:0] node868;
	wire [3-1:0] node870;
	wire [3-1:0] node872;
	wire [3-1:0] node875;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node880;
	wire [3-1:0] node882;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node908;
	wire [3-1:0] node909;

	assign outp = (inp[9]) ? node586 : node1;
		assign node1 = (inp[6]) ? node259 : node2;
			assign node2 = (inp[10]) ? node102 : node3;
				assign node3 = (inp[7]) ? node17 : node4;
					assign node4 = (inp[8]) ? node6 : 3'b111;
						assign node6 = (inp[3]) ? node8 : 3'b111;
							assign node8 = (inp[11]) ? node10 : 3'b111;
								assign node10 = (inp[4]) ? 3'b011 : node11;
									assign node11 = (inp[5]) ? node13 : 3'b111;
										assign node13 = (inp[0]) ? 3'b011 : 3'b111;
					assign node17 = (inp[11]) ? node47 : node18;
						assign node18 = (inp[8]) ? node34 : node19;
							assign node19 = (inp[3]) ? node21 : 3'b111;
								assign node21 = (inp[4]) ? node23 : 3'b111;
									assign node23 = (inp[5]) ? node29 : node24;
										assign node24 = (inp[0]) ? node26 : 3'b111;
											assign node26 = (inp[1]) ? 3'b011 : 3'b111;
										assign node29 = (inp[0]) ? 3'b011 : node30;
											assign node30 = (inp[1]) ? 3'b011 : 3'b111;
							assign node34 = (inp[3]) ? 3'b011 : node35;
								assign node35 = (inp[4]) ? node37 : 3'b111;
									assign node37 = (inp[0]) ? 3'b011 : node38;
										assign node38 = (inp[5]) ? node40 : 3'b111;
											assign node40 = (inp[2]) ? 3'b011 : node41;
												assign node41 = (inp[1]) ? 3'b011 : 3'b111;
						assign node47 = (inp[8]) ? node83 : node48;
							assign node48 = (inp[4]) ? node66 : node49;
								assign node49 = (inp[3]) ? 3'b011 : node50;
									assign node50 = (inp[5]) ? node58 : node51;
										assign node51 = (inp[2]) ? node53 : 3'b111;
											assign node53 = (inp[0]) ? node55 : 3'b111;
												assign node55 = (inp[1]) ? 3'b011 : 3'b111;
										assign node58 = (inp[0]) ? 3'b011 : node59;
											assign node59 = (inp[1]) ? node61 : 3'b111;
												assign node61 = (inp[2]) ? 3'b011 : 3'b111;
								assign node66 = (inp[3]) ? node68 : 3'b011;
									assign node68 = (inp[5]) ? node76 : node69;
										assign node69 = (inp[0]) ? node71 : 3'b011;
											assign node71 = (inp[2]) ? 3'b101 : node72;
												assign node72 = (inp[1]) ? 3'b101 : 3'b011;
										assign node76 = (inp[0]) ? 3'b101 : node77;
											assign node77 = (inp[1]) ? 3'b101 : node78;
												assign node78 = (inp[2]) ? 3'b101 : 3'b011;
							assign node83 = (inp[3]) ? node91 : node84;
								assign node84 = (inp[4]) ? node86 : 3'b011;
									assign node86 = (inp[5]) ? 3'b101 : node87;
										assign node87 = (inp[0]) ? 3'b101 : 3'b011;
								assign node91 = (inp[0]) ? node93 : 3'b101;
									assign node93 = (inp[5]) ? node95 : 3'b101;
										assign node95 = (inp[2]) ? node97 : 3'b101;
											assign node97 = (inp[4]) ? node99 : 3'b101;
												assign node99 = (inp[1]) ? 3'b001 : 3'b101;
				assign node102 = (inp[7]) ? node168 : node103;
					assign node103 = (inp[11]) ? node141 : node104;
						assign node104 = (inp[8]) ? node124 : node105;
							assign node105 = (inp[3]) ? node115 : node106;
								assign node106 = (inp[5]) ? node108 : 3'b111;
									assign node108 = (inp[1]) ? node110 : 3'b111;
										assign node110 = (inp[4]) ? node112 : 3'b111;
											assign node112 = (inp[0]) ? 3'b011 : 3'b111;
								assign node115 = (inp[5]) ? 3'b011 : node116;
									assign node116 = (inp[1]) ? 3'b011 : node117;
										assign node117 = (inp[2]) ? 3'b011 : node118;
											assign node118 = (inp[4]) ? 3'b011 : 3'b111;
							assign node124 = (inp[3]) ? node126 : 3'b011;
								assign node126 = (inp[4]) ? 3'b101 : node127;
									assign node127 = (inp[0]) ? node135 : node128;
										assign node128 = (inp[1]) ? node130 : 3'b011;
											assign node130 = (inp[5]) ? node132 : 3'b011;
												assign node132 = (inp[2]) ? 3'b101 : 3'b011;
										assign node135 = (inp[5]) ? 3'b101 : node136;
											assign node136 = (inp[2]) ? 3'b101 : 3'b011;
						assign node141 = (inp[8]) ? node151 : node142;
							assign node142 = (inp[3]) ? 3'b101 : node143;
								assign node143 = (inp[0]) ? node145 : 3'b011;
									assign node145 = (inp[5]) ? node147 : 3'b011;
										assign node147 = (inp[4]) ? 3'b101 : 3'b011;
							assign node151 = (inp[3]) ? node153 : 3'b101;
								assign node153 = (inp[4]) ? 3'b001 : node154;
									assign node154 = (inp[5]) ? node160 : node155;
										assign node155 = (inp[0]) ? node157 : 3'b101;
											assign node157 = (inp[1]) ? 3'b001 : 3'b101;
										assign node160 = (inp[0]) ? 3'b001 : node161;
											assign node161 = (inp[1]) ? 3'b001 : node162;
												assign node162 = (inp[2]) ? 3'b001 : 3'b101;
					assign node168 = (inp[11]) ? node216 : node169;
						assign node169 = (inp[8]) ? node187 : node170;
							assign node170 = (inp[4]) ? node180 : node171;
								assign node171 = (inp[3]) ? 3'b101 : node172;
									assign node172 = (inp[5]) ? 3'b101 : node173;
										assign node173 = (inp[0]) ? node175 : 3'b011;
											assign node175 = (inp[1]) ? 3'b101 : 3'b011;
								assign node180 = (inp[3]) ? node182 : 3'b101;
									assign node182 = (inp[0]) ? 3'b001 : node183;
										assign node183 = (inp[5]) ? 3'b001 : 3'b101;
							assign node187 = (inp[3]) ? node207 : node188;
								assign node188 = (inp[4]) ? node198 : node189;
									assign node189 = (inp[1]) ? node191 : 3'b101;
										assign node191 = (inp[0]) ? node193 : 3'b101;
											assign node193 = (inp[2]) ? node195 : 3'b101;
												assign node195 = (inp[5]) ? 3'b001 : 3'b101;
									assign node198 = (inp[5]) ? 3'b001 : node199;
										assign node199 = (inp[0]) ? 3'b001 : node200;
											assign node200 = (inp[2]) ? node202 : 3'b101;
												assign node202 = (inp[1]) ? 3'b001 : 3'b101;
								assign node207 = (inp[5]) ? node209 : 3'b001;
									assign node209 = (inp[0]) ? node211 : 3'b001;
										assign node211 = (inp[1]) ? node213 : 3'b001;
											assign node213 = (inp[4]) ? 3'b110 : 3'b001;
						assign node216 = (inp[8]) ? node242 : node217;
							assign node217 = (inp[3]) ? node225 : node218;
								assign node218 = (inp[5]) ? 3'b001 : node219;
									assign node219 = (inp[0]) ? 3'b001 : node220;
										assign node220 = (inp[4]) ? 3'b001 : 3'b101;
								assign node225 = (inp[4]) ? node233 : node226;
									assign node226 = (inp[5]) ? node228 : 3'b001;
										assign node228 = (inp[0]) ? node230 : 3'b001;
											assign node230 = (inp[2]) ? 3'b110 : 3'b001;
									assign node233 = (inp[0]) ? 3'b110 : node234;
										assign node234 = (inp[5]) ? 3'b110 : node235;
											assign node235 = (inp[1]) ? node237 : 3'b001;
												assign node237 = (inp[2]) ? 3'b110 : 3'b001;
							assign node242 = (inp[4]) ? node252 : node243;
								assign node243 = (inp[3]) ? 3'b110 : node244;
									assign node244 = (inp[1]) ? node246 : 3'b001;
										assign node246 = (inp[5]) ? node248 : 3'b001;
											assign node248 = (inp[0]) ? 3'b110 : 3'b001;
								assign node252 = (inp[3]) ? node254 : 3'b110;
									assign node254 = (inp[0]) ? node256 : 3'b110;
										assign node256 = (inp[5]) ? 3'b010 : 3'b110;
			assign node259 = (inp[10]) ? node441 : node260;
				assign node260 = (inp[7]) ? node344 : node261;
					assign node261 = (inp[11]) ? node303 : node262;
						assign node262 = (inp[8]) ? node284 : node263;
							assign node263 = (inp[3]) ? node275 : node264;
								assign node264 = (inp[0]) ? node266 : 3'b011;
									assign node266 = (inp[2]) ? node268 : 3'b011;
										assign node268 = (inp[1]) ? node270 : 3'b011;
											assign node270 = (inp[5]) ? node272 : 3'b011;
												assign node272 = (inp[4]) ? 3'b101 : 3'b011;
								assign node275 = (inp[0]) ? 3'b101 : node276;
									assign node276 = (inp[4]) ? 3'b101 : node277;
										assign node277 = (inp[1]) ? 3'b101 : node278;
											assign node278 = (inp[5]) ? 3'b101 : 3'b011;
							assign node284 = (inp[3]) ? node296 : node285;
								assign node285 = (inp[0]) ? 3'b101 : node286;
									assign node286 = (inp[2]) ? 3'b101 : node287;
										assign node287 = (inp[4]) ? 3'b101 : node288;
											assign node288 = (inp[1]) ? 3'b101 : node289;
												assign node289 = (inp[5]) ? 3'b101 : 3'b011;
								assign node296 = (inp[4]) ? 3'b001 : node297;
									assign node297 = (inp[5]) ? node299 : 3'b101;
										assign node299 = (inp[0]) ? 3'b001 : 3'b101;
						assign node303 = (inp[3]) ? node317 : node304;
							assign node304 = (inp[8]) ? 3'b001 : node305;
								assign node305 = (inp[4]) ? node307 : 3'b101;
									assign node307 = (inp[0]) ? node309 : 3'b101;
										assign node309 = (inp[5]) ? node311 : 3'b101;
											assign node311 = (inp[1]) ? 3'b001 : node312;
												assign node312 = (inp[2]) ? 3'b001 : 3'b101;
							assign node317 = (inp[8]) ? node329 : node318;
								assign node318 = (inp[2]) ? 3'b001 : node319;
									assign node319 = (inp[4]) ? 3'b001 : node320;
										assign node320 = (inp[5]) ? 3'b001 : node321;
											assign node321 = (inp[0]) ? 3'b001 : node322;
												assign node322 = (inp[1]) ? 3'b001 : 3'b101;
								assign node329 = (inp[4]) ? 3'b110 : node330;
									assign node330 = (inp[5]) ? node338 : node331;
										assign node331 = (inp[0]) ? node333 : 3'b001;
											assign node333 = (inp[1]) ? node335 : 3'b001;
												assign node335 = (inp[2]) ? 3'b110 : 3'b001;
										assign node338 = (inp[1]) ? 3'b110 : node339;
											assign node339 = (inp[0]) ? 3'b110 : 3'b001;
					assign node344 = (inp[11]) ? node388 : node345;
						assign node345 = (inp[8]) ? node371 : node346;
							assign node346 = (inp[3]) ? node362 : node347;
								assign node347 = (inp[4]) ? 3'b001 : node348;
									assign node348 = (inp[5]) ? node356 : node349;
										assign node349 = (inp[1]) ? node351 : 3'b101;
											assign node351 = (inp[2]) ? node353 : 3'b101;
												assign node353 = (inp[0]) ? 3'b001 : 3'b101;
										assign node356 = (inp[0]) ? 3'b001 : node357;
											assign node357 = (inp[1]) ? 3'b001 : 3'b101;
								assign node362 = (inp[4]) ? node364 : 3'b001;
									assign node364 = (inp[5]) ? 3'b110 : node365;
										assign node365 = (inp[0]) ? node367 : 3'b001;
											assign node367 = (inp[2]) ? 3'b110 : 3'b001;
							assign node371 = (inp[3]) ? node379 : node372;
								assign node372 = (inp[4]) ? node374 : 3'b001;
									assign node374 = (inp[5]) ? 3'b110 : node375;
										assign node375 = (inp[0]) ? 3'b110 : 3'b001;
								assign node379 = (inp[1]) ? node381 : 3'b110;
									assign node381 = (inp[4]) ? node383 : 3'b110;
										assign node383 = (inp[5]) ? node385 : 3'b110;
											assign node385 = (inp[0]) ? 3'b010 : 3'b110;
						assign node388 = (inp[8]) ? node414 : node389;
							assign node389 = (inp[4]) ? node407 : node390;
								assign node390 = (inp[3]) ? 3'b110 : node391;
									assign node391 = (inp[5]) ? node399 : node392;
										assign node392 = (inp[0]) ? node394 : 3'b001;
											assign node394 = (inp[1]) ? 3'b110 : node395;
												assign node395 = (inp[2]) ? 3'b110 : 3'b001;
										assign node399 = (inp[2]) ? 3'b110 : node400;
											assign node400 = (inp[0]) ? 3'b110 : node401;
												assign node401 = (inp[1]) ? 3'b110 : 3'b001;
								assign node407 = (inp[3]) ? node409 : 3'b110;
									assign node409 = (inp[5]) ? 3'b010 : node410;
										assign node410 = (inp[0]) ? 3'b010 : 3'b110;
							assign node414 = (inp[3]) ? node430 : node415;
								assign node415 = (inp[4]) ? node423 : node416;
									assign node416 = (inp[2]) ? node418 : 3'b110;
										assign node418 = (inp[1]) ? node420 : 3'b110;
											assign node420 = (inp[0]) ? 3'b010 : 3'b110;
									assign node423 = (inp[0]) ? 3'b010 : node424;
										assign node424 = (inp[1]) ? 3'b010 : node425;
											assign node425 = (inp[5]) ? 3'b010 : 3'b110;
								assign node430 = (inp[0]) ? node432 : 3'b010;
									assign node432 = (inp[4]) ? node434 : 3'b010;
										assign node434 = (inp[5]) ? node436 : 3'b010;
											assign node436 = (inp[1]) ? 3'b100 : node437;
												assign node437 = (inp[2]) ? 3'b100 : 3'b010;
				assign node441 = (inp[7]) ? node497 : node442;
					assign node442 = (inp[11]) ? node470 : node443;
						assign node443 = (inp[3]) ? node453 : node444;
							assign node444 = (inp[8]) ? 3'b110 : node445;
								assign node445 = (inp[5]) ? node447 : 3'b001;
									assign node447 = (inp[0]) ? node449 : 3'b001;
										assign node449 = (inp[4]) ? 3'b110 : 3'b001;
							assign node453 = (inp[8]) ? node455 : 3'b110;
								assign node455 = (inp[4]) ? 3'b010 : node456;
									assign node456 = (inp[0]) ? node462 : node457;
										assign node457 = (inp[5]) ? node459 : 3'b110;
											assign node459 = (inp[1]) ? 3'b010 : 3'b110;
										assign node462 = (inp[1]) ? 3'b010 : node463;
											assign node463 = (inp[5]) ? 3'b010 : node464;
												assign node464 = (inp[2]) ? 3'b010 : 3'b110;
						assign node470 = (inp[3]) ? node488 : node471;
							assign node471 = (inp[8]) ? 3'b010 : node472;
								assign node472 = (inp[4]) ? node474 : 3'b110;
									assign node474 = (inp[5]) ? node482 : node475;
										assign node475 = (inp[0]) ? node477 : 3'b110;
											assign node477 = (inp[1]) ? node479 : 3'b110;
												assign node479 = (inp[2]) ? 3'b010 : 3'b110;
										assign node482 = (inp[0]) ? 3'b010 : node483;
											assign node483 = (inp[1]) ? 3'b010 : 3'b110;
							assign node488 = (inp[8]) ? node490 : 3'b010;
								assign node490 = (inp[5]) ? 3'b100 : node491;
									assign node491 = (inp[0]) ? 3'b100 : node492;
										assign node492 = (inp[4]) ? 3'b100 : 3'b010;
					assign node497 = (inp[11]) ? node549 : node498;
						assign node498 = (inp[8]) ? node526 : node499;
							assign node499 = (inp[3]) ? node507 : node500;
								assign node500 = (inp[0]) ? 3'b010 : node501;
									assign node501 = (inp[4]) ? 3'b010 : node502;
										assign node502 = (inp[5]) ? 3'b010 : 3'b110;
								assign node507 = (inp[4]) ? node517 : node508;
									assign node508 = (inp[2]) ? node510 : 3'b010;
										assign node510 = (inp[1]) ? node512 : 3'b010;
											assign node512 = (inp[0]) ? node514 : 3'b010;
												assign node514 = (inp[5]) ? 3'b100 : 3'b010;
									assign node517 = (inp[0]) ? 3'b100 : node518;
										assign node518 = (inp[5]) ? 3'b100 : node519;
											assign node519 = (inp[1]) ? node521 : 3'b010;
												assign node521 = (inp[2]) ? 3'b100 : 3'b010;
							assign node526 = (inp[3]) ? node542 : node527;
								assign node527 = (inp[4]) ? node535 : node528;
									assign node528 = (inp[5]) ? node530 : 3'b010;
										assign node530 = (inp[0]) ? node532 : 3'b010;
											assign node532 = (inp[1]) ? 3'b100 : 3'b010;
									assign node535 = (inp[5]) ? 3'b100 : node536;
										assign node536 = (inp[2]) ? 3'b100 : node537;
											assign node537 = (inp[0]) ? 3'b100 : 3'b010;
								assign node542 = (inp[4]) ? node544 : 3'b100;
									assign node544 = (inp[0]) ? node546 : 3'b100;
										assign node546 = (inp[5]) ? 3'b000 : 3'b100;
						assign node549 = (inp[8]) ? node577 : node550;
							assign node550 = (inp[3]) ? node562 : node551;
								assign node551 = (inp[5]) ? 3'b100 : node552;
									assign node552 = (inp[4]) ? 3'b100 : node553;
										assign node553 = (inp[2]) ? node555 : 3'b010;
											assign node555 = (inp[0]) ? 3'b100 : node556;
												assign node556 = (inp[1]) ? 3'b100 : 3'b010;
								assign node562 = (inp[4]) ? node570 : node563;
									assign node563 = (inp[1]) ? node565 : 3'b100;
										assign node565 = (inp[0]) ? node567 : 3'b100;
											assign node567 = (inp[2]) ? 3'b100 : 3'b000;
									assign node570 = (inp[1]) ? 3'b000 : node571;
										assign node571 = (inp[2]) ? 3'b000 : node572;
											assign node572 = (inp[0]) ? 3'b000 : 3'b100;
							assign node577 = (inp[3]) ? 3'b000 : node578;
								assign node578 = (inp[4]) ? 3'b000 : node579;
									assign node579 = (inp[0]) ? node581 : 3'b100;
										assign node581 = (inp[5]) ? 3'b000 : 3'b100;
		assign node586 = (inp[6]) ? node846 : node587;
			assign node587 = (inp[10]) ? node747 : node588;
				assign node588 = (inp[7]) ? node646 : node589;
					assign node589 = (inp[11]) ? node617 : node590;
						assign node590 = (inp[3]) ? node604 : node591;
							assign node591 = (inp[8]) ? 3'b001 : node592;
								assign node592 = (inp[5]) ? node594 : 3'b101;
									assign node594 = (inp[4]) ? node596 : 3'b101;
										assign node596 = (inp[0]) ? 3'b001 : node597;
											assign node597 = (inp[1]) ? node599 : 3'b101;
												assign node599 = (inp[2]) ? 3'b001 : 3'b101;
							assign node604 = (inp[8]) ? node606 : 3'b001;
								assign node606 = (inp[5]) ? 3'b110 : node607;
									assign node607 = (inp[4]) ? 3'b110 : node608;
										assign node608 = (inp[0]) ? node610 : 3'b001;
											assign node610 = (inp[2]) ? 3'b110 : node611;
												assign node611 = (inp[1]) ? 3'b110 : 3'b001;
						assign node617 = (inp[3]) ? node633 : node618;
							assign node618 = (inp[8]) ? 3'b110 : node619;
								assign node619 = (inp[4]) ? node621 : 3'b001;
									assign node621 = (inp[0]) ? node627 : node622;
										assign node622 = (inp[5]) ? node624 : 3'b001;
											assign node624 = (inp[1]) ? 3'b110 : 3'b001;
										assign node627 = (inp[1]) ? 3'b110 : node628;
											assign node628 = (inp[5]) ? 3'b110 : 3'b001;
							assign node633 = (inp[8]) ? node635 : 3'b110;
								assign node635 = (inp[0]) ? 3'b010 : node636;
									assign node636 = (inp[5]) ? 3'b010 : node637;
										assign node637 = (inp[4]) ? 3'b010 : node638;
											assign node638 = (inp[1]) ? node640 : 3'b110;
												assign node640 = (inp[2]) ? 3'b010 : 3'b110;
					assign node646 = (inp[11]) ? node700 : node647;
						assign node647 = (inp[8]) ? node673 : node648;
							assign node648 = (inp[3]) ? node658 : node649;
								assign node649 = (inp[0]) ? 3'b110 : node650;
									assign node650 = (inp[5]) ? 3'b110 : node651;
										assign node651 = (inp[4]) ? 3'b110 : node652;
											assign node652 = (inp[1]) ? 3'b110 : 3'b001;
								assign node658 = (inp[4]) ? node666 : node659;
									assign node659 = (inp[1]) ? node661 : 3'b110;
										assign node661 = (inp[5]) ? node663 : 3'b110;
											assign node663 = (inp[0]) ? 3'b010 : 3'b110;
									assign node666 = (inp[1]) ? 3'b010 : node667;
										assign node667 = (inp[0]) ? 3'b010 : node668;
											assign node668 = (inp[5]) ? 3'b010 : 3'b110;
							assign node673 = (inp[4]) ? node685 : node674;
								assign node674 = (inp[3]) ? 3'b010 : node675;
									assign node675 = (inp[0]) ? node677 : 3'b110;
										assign node677 = (inp[5]) ? node679 : 3'b110;
											assign node679 = (inp[1]) ? 3'b010 : node680;
												assign node680 = (inp[2]) ? 3'b010 : 3'b110;
								assign node685 = (inp[3]) ? node687 : 3'b010;
									assign node687 = (inp[0]) ? node695 : node688;
										assign node688 = (inp[5]) ? node690 : 3'b010;
											assign node690 = (inp[1]) ? node692 : 3'b010;
												assign node692 = (inp[2]) ? 3'b100 : 3'b010;
										assign node695 = (inp[5]) ? 3'b100 : node696;
											assign node696 = (inp[2]) ? 3'b100 : 3'b010;
						assign node700 = (inp[8]) ? node722 : node701;
							assign node701 = (inp[3]) ? node711 : node702;
								assign node702 = (inp[5]) ? 3'b010 : node703;
									assign node703 = (inp[4]) ? 3'b010 : node704;
										assign node704 = (inp[1]) ? 3'b010 : node705;
											assign node705 = (inp[0]) ? 3'b010 : 3'b110;
								assign node711 = (inp[4]) ? 3'b100 : node712;
									assign node712 = (inp[5]) ? node714 : 3'b010;
										assign node714 = (inp[0]) ? node716 : 3'b010;
											assign node716 = (inp[2]) ? 3'b100 : node717;
												assign node717 = (inp[1]) ? 3'b100 : 3'b010;
							assign node722 = (inp[4]) ? node734 : node723;
								assign node723 = (inp[3]) ? 3'b100 : node724;
									assign node724 = (inp[5]) ? node726 : 3'b010;
										assign node726 = (inp[0]) ? 3'b100 : node727;
											assign node727 = (inp[1]) ? node729 : 3'b010;
												assign node729 = (inp[2]) ? 3'b100 : 3'b010;
								assign node734 = (inp[3]) ? node736 : 3'b100;
									assign node736 = (inp[5]) ? node742 : node737;
										assign node737 = (inp[1]) ? node739 : 3'b100;
											assign node739 = (inp[0]) ? 3'b000 : 3'b100;
										assign node742 = (inp[1]) ? 3'b000 : node743;
											assign node743 = (inp[0]) ? 3'b000 : 3'b100;
				assign node747 = (inp[7]) ? node815 : node748;
					assign node748 = (inp[11]) ? node786 : node749;
						assign node749 = (inp[8]) ? node767 : node750;
							assign node750 = (inp[3]) ? 3'b010 : node751;
								assign node751 = (inp[4]) ? node753 : 3'b110;
									assign node753 = (inp[0]) ? node761 : node754;
										assign node754 = (inp[5]) ? node756 : 3'b110;
											assign node756 = (inp[2]) ? 3'b010 : node757;
												assign node757 = (inp[1]) ? 3'b010 : 3'b110;
										assign node761 = (inp[5]) ? 3'b010 : node762;
											assign node762 = (inp[2]) ? 3'b010 : 3'b110;
							assign node767 = (inp[3]) ? node777 : node768;
								assign node768 = (inp[4]) ? node770 : 3'b010;
									assign node770 = (inp[5]) ? node772 : 3'b010;
										assign node772 = (inp[1]) ? node774 : 3'b010;
											assign node774 = (inp[0]) ? 3'b100 : 3'b010;
								assign node777 = (inp[0]) ? 3'b100 : node778;
									assign node778 = (inp[1]) ? 3'b100 : node779;
										assign node779 = (inp[4]) ? 3'b100 : node780;
											assign node780 = (inp[5]) ? 3'b100 : 3'b010;
						assign node786 = (inp[8]) ? node796 : node787;
							assign node787 = (inp[3]) ? 3'b100 : node788;
								assign node788 = (inp[4]) ? node790 : 3'b010;
									assign node790 = (inp[5]) ? 3'b100 : node791;
										assign node791 = (inp[0]) ? 3'b100 : 3'b010;
							assign node796 = (inp[3]) ? node806 : node797;
								assign node797 = (inp[0]) ? node799 : 3'b100;
									assign node799 = (inp[2]) ? node801 : 3'b100;
										assign node801 = (inp[5]) ? node803 : 3'b100;
											assign node803 = (inp[4]) ? 3'b000 : 3'b100;
								assign node806 = (inp[4]) ? 3'b000 : node807;
									assign node807 = (inp[0]) ? 3'b000 : node808;
										assign node808 = (inp[1]) ? 3'b000 : node809;
											assign node809 = (inp[2]) ? 3'b000 : 3'b100;
					assign node815 = (inp[11]) ? 3'b000 : node816;
						assign node816 = (inp[8]) ? node830 : node817;
							assign node817 = (inp[3]) ? node819 : 3'b100;
								assign node819 = (inp[4]) ? 3'b000 : node820;
									assign node820 = (inp[5]) ? node822 : 3'b100;
										assign node822 = (inp[0]) ? 3'b000 : node823;
											assign node823 = (inp[2]) ? node825 : 3'b100;
												assign node825 = (inp[1]) ? 3'b000 : 3'b100;
							assign node830 = (inp[4]) ? 3'b000 : node831;
								assign node831 = (inp[3]) ? 3'b000 : node832;
									assign node832 = (inp[1]) ? node838 : node833;
										assign node833 = (inp[5]) ? node835 : 3'b100;
											assign node835 = (inp[0]) ? 3'b000 : 3'b100;
										assign node838 = (inp[5]) ? 3'b000 : node839;
											assign node839 = (inp[0]) ? 3'b000 : 3'b100;
			assign node846 = (inp[10]) ? 3'b000 : node847;
				assign node847 = (inp[7]) ? node903 : node848;
					assign node848 = (inp[11]) ? node888 : node849;
						assign node849 = (inp[3]) ? node875 : node850;
							assign node850 = (inp[8]) ? node864 : node851;
								assign node851 = (inp[4]) ? node853 : 3'b010;
									assign node853 = (inp[1]) ? node859 : node854;
										assign node854 = (inp[5]) ? node856 : 3'b010;
											assign node856 = (inp[0]) ? 3'b100 : 3'b010;
										assign node859 = (inp[5]) ? 3'b100 : node860;
											assign node860 = (inp[0]) ? 3'b100 : 3'b010;
								assign node864 = (inp[0]) ? node866 : 3'b100;
									assign node866 = (inp[2]) ? node868 : 3'b100;
										assign node868 = (inp[5]) ? node870 : 3'b100;
											assign node870 = (inp[1]) ? node872 : 3'b100;
												assign node872 = (inp[4]) ? 3'b000 : 3'b100;
							assign node875 = (inp[8]) ? node877 : 3'b100;
								assign node877 = (inp[4]) ? 3'b000 : node878;
									assign node878 = (inp[0]) ? 3'b000 : node879;
										assign node879 = (inp[5]) ? 3'b000 : node880;
											assign node880 = (inp[1]) ? node882 : 3'b100;
												assign node882 = (inp[2]) ? 3'b000 : 3'b100;
						assign node888 = (inp[8]) ? 3'b000 : node889;
							assign node889 = (inp[3]) ? 3'b000 : node890;
								assign node890 = (inp[4]) ? node892 : 3'b100;
									assign node892 = (inp[5]) ? 3'b000 : node893;
										assign node893 = (inp[0]) ? node895 : 3'b100;
											assign node895 = (inp[1]) ? 3'b000 : node896;
												assign node896 = (inp[2]) ? 3'b000 : 3'b100;
					assign node903 = (inp[0]) ? 3'b000 : node904;
						assign node904 = (inp[5]) ? 3'b000 : node905;
							assign node905 = (inp[3]) ? 3'b000 : node906;
								assign node906 = (inp[4]) ? 3'b000 : node907;
									assign node907 = (inp[1]) ? 3'b000 : node908;
										assign node908 = (inp[8]) ? 3'b000 : node909;
											assign node909 = (inp[11]) ? 3'b000 : 3'b100;

endmodule