module dtc_split875_bm91 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node129;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node140;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node184;
	wire [3-1:0] node186;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node250;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node319;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node332;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node340;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node347;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node400;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node426;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node450;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node461;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node468;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node483;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node502;
	wire [3-1:0] node504;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node519;
	wire [3-1:0] node523;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node528;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node542;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node553;
	wire [3-1:0] node556;
	wire [3-1:0] node559;
	wire [3-1:0] node560;
	wire [3-1:0] node562;
	wire [3-1:0] node564;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node573;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node581;
	wire [3-1:0] node585;
	wire [3-1:0] node587;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node608;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node621;
	wire [3-1:0] node622;
	wire [3-1:0] node624;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node635;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node646;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node656;
	wire [3-1:0] node657;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node673;
	wire [3-1:0] node674;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node680;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node690;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node696;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node731;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node740;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node753;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node777;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node785;
	wire [3-1:0] node789;
	wire [3-1:0] node790;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node795;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node802;
	wire [3-1:0] node805;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node812;
	wire [3-1:0] node814;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node822;
	wire [3-1:0] node824;
	wire [3-1:0] node825;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node837;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node842;
	wire [3-1:0] node845;
	wire [3-1:0] node848;
	wire [3-1:0] node850;
	wire [3-1:0] node852;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node862;
	wire [3-1:0] node865;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node872;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node886;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node891;
	wire [3-1:0] node895;
	wire [3-1:0] node897;
	wire [3-1:0] node899;
	wire [3-1:0] node902;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node909;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node917;
	wire [3-1:0] node920;
	wire [3-1:0] node922;
	wire [3-1:0] node925;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node938;
	wire [3-1:0] node941;
	wire [3-1:0] node943;
	wire [3-1:0] node946;
	wire [3-1:0] node948;
	wire [3-1:0] node950;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node960;
	wire [3-1:0] node963;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node969;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node977;
	wire [3-1:0] node979;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node984;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node991;
	wire [3-1:0] node993;
	wire [3-1:0] node995;
	wire [3-1:0] node998;
	wire [3-1:0] node1001;
	wire [3-1:0] node1002;
	wire [3-1:0] node1003;
	wire [3-1:0] node1005;
	wire [3-1:0] node1009;
	wire [3-1:0] node1011;
	wire [3-1:0] node1013;
	wire [3-1:0] node1016;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1021;
	wire [3-1:0] node1023;
	wire [3-1:0] node1025;
	wire [3-1:0] node1026;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1034;
	wire [3-1:0] node1035;
	wire [3-1:0] node1037;
	wire [3-1:0] node1039;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1050;
	wire [3-1:0] node1052;
	wire [3-1:0] node1054;
	wire [3-1:0] node1058;
	wire [3-1:0] node1059;
	wire [3-1:0] node1060;
	wire [3-1:0] node1062;
	wire [3-1:0] node1065;
	wire [3-1:0] node1067;
	wire [3-1:0] node1070;
	wire [3-1:0] node1071;
	wire [3-1:0] node1073;
	wire [3-1:0] node1074;
	wire [3-1:0] node1076;
	wire [3-1:0] node1078;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1085;
	wire [3-1:0] node1086;
	wire [3-1:0] node1090;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1096;
	wire [3-1:0] node1097;
	wire [3-1:0] node1101;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1107;
	wire [3-1:0] node1109;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1115;
	wire [3-1:0] node1117;

	assign outp = (inp[3]) ? node808 : node1;
		assign node1 = (inp[9]) ? node351 : node2;
			assign node2 = (inp[1]) ? node108 : node3;
				assign node3 = (inp[5]) ? node49 : node4;
					assign node4 = (inp[6]) ? node24 : node5;
						assign node5 = (inp[4]) ? node15 : node6;
							assign node6 = (inp[0]) ? node8 : 3'b001;
								assign node8 = (inp[2]) ? 3'b000 : node9;
									assign node9 = (inp[7]) ? 3'b000 : node10;
										assign node10 = (inp[8]) ? 3'b000 : 3'b001;
							assign node15 = (inp[0]) ? node17 : 3'b000;
								assign node17 = (inp[2]) ? 3'b001 : node18;
									assign node18 = (inp[8]) ? 3'b001 : node19;
										assign node19 = (inp[7]) ? 3'b001 : 3'b000;
						assign node24 = (inp[10]) ? node34 : node25;
							assign node25 = (inp[0]) ? 3'b000 : node26;
								assign node26 = (inp[4]) ? node28 : 3'b000;
									assign node28 = (inp[8]) ? node30 : 3'b000;
										assign node30 = (inp[7]) ? 3'b000 : 3'b001;
							assign node34 = (inp[7]) ? node42 : node35;
								assign node35 = (inp[0]) ? 3'b000 : node36;
									assign node36 = (inp[8]) ? node38 : 3'b000;
										assign node38 = (inp[4]) ? 3'b001 : 3'b000;
								assign node42 = (inp[0]) ? node46 : node43;
									assign node43 = (inp[4]) ? 3'b001 : 3'b000;
									assign node46 = (inp[4]) ? 3'b000 : 3'b001;
					assign node49 = (inp[4]) ? node75 : node50;
						assign node50 = (inp[6]) ? node62 : node51;
							assign node51 = (inp[7]) ? 3'b001 : node52;
								assign node52 = (inp[0]) ? node54 : 3'b000;
									assign node54 = (inp[8]) ? node56 : 3'b001;
										assign node56 = (inp[2]) ? 3'b001 : node57;
											assign node57 = (inp[11]) ? 3'b001 : 3'b000;
							assign node62 = (inp[0]) ? node68 : node63;
								assign node63 = (inp[8]) ? node65 : 3'b001;
									assign node65 = (inp[7]) ? 3'b000 : 3'b001;
								assign node68 = (inp[7]) ? node70 : 3'b000;
									assign node70 = (inp[10]) ? node72 : 3'b000;
										assign node72 = (inp[2]) ? 3'b001 : 3'b000;
						assign node75 = (inp[6]) ? node87 : node76;
							assign node76 = (inp[8]) ? node78 : 3'b000;
								assign node78 = (inp[7]) ? 3'b000 : node79;
									assign node79 = (inp[11]) ? 3'b000 : node80;
										assign node80 = (inp[2]) ? 3'b000 : node81;
											assign node81 = (inp[0]) ? 3'b001 : 3'b000;
							assign node87 = (inp[0]) ? 3'b001 : node88;
								assign node88 = (inp[8]) ? node96 : node89;
									assign node89 = (inp[10]) ? node91 : 3'b000;
										assign node91 = (inp[2]) ? node93 : 3'b000;
											assign node93 = (inp[7]) ? 3'b001 : 3'b000;
									assign node96 = (inp[10]) ? node102 : node97;
										assign node97 = (inp[11]) ? 3'b000 : node98;
											assign node98 = (inp[7]) ? 3'b000 : 3'b001;
										assign node102 = (inp[7]) ? 3'b001 : node103;
											assign node103 = (inp[11]) ? 3'b000 : 3'b001;
				assign node108 = (inp[8]) ? node226 : node109;
					assign node109 = (inp[6]) ? node175 : node110;
						assign node110 = (inp[5]) ? node144 : node111;
							assign node111 = (inp[4]) ? node133 : node112;
								assign node112 = (inp[0]) ? 3'b000 : node113;
									assign node113 = (inp[7]) ? node119 : node114;
										assign node114 = (inp[10]) ? 3'b001 : node115;
											assign node115 = (inp[2]) ? 3'b001 : 3'b000;
										assign node119 = (inp[11]) ? node125 : node120;
											assign node120 = (inp[2]) ? node122 : 3'b000;
												assign node122 = (inp[10]) ? 3'b000 : 3'b001;
											assign node125 = (inp[2]) ? node129 : node126;
												assign node126 = (inp[10]) ? 3'b001 : 3'b000;
												assign node129 = (inp[10]) ? 3'b000 : 3'b001;
								assign node133 = (inp[0]) ? 3'b001 : node134;
									assign node134 = (inp[2]) ? node138 : node135;
										assign node135 = (inp[10]) ? 3'b000 : 3'b001;
										assign node138 = (inp[7]) ? node140 : 3'b000;
											assign node140 = (inp[10]) ? 3'b001 : 3'b000;
							assign node144 = (inp[4]) ? node156 : node145;
								assign node145 = (inp[7]) ? node147 : 3'b001;
									assign node147 = (inp[0]) ? 3'b000 : node148;
										assign node148 = (inp[10]) ? node150 : 3'b000;
											assign node150 = (inp[11]) ? 3'b001 : node151;
												assign node151 = (inp[2]) ? 3'b000 : 3'b001;
								assign node156 = (inp[7]) ? node162 : node157;
									assign node157 = (inp[11]) ? 3'b000 : node158;
										assign node158 = (inp[0]) ? 3'b001 : 3'b000;
									assign node162 = (inp[0]) ? 3'b001 : node163;
										assign node163 = (inp[10]) ? node169 : node164;
											assign node164 = (inp[2]) ? node166 : 3'b001;
												assign node166 = (inp[11]) ? 3'b001 : 3'b000;
											assign node169 = (inp[2]) ? node171 : 3'b000;
												assign node171 = (inp[11]) ? 3'b000 : 3'b001;
						assign node175 = (inp[5]) ? node193 : node176;
							assign node176 = (inp[4]) ? node190 : node177;
								assign node177 = (inp[0]) ? 3'b001 : node178;
									assign node178 = (inp[7]) ? node184 : node179;
										assign node179 = (inp[10]) ? 3'b000 : node180;
											assign node180 = (inp[2]) ? 3'b000 : 3'b001;
										assign node184 = (inp[2]) ? node186 : 3'b001;
											assign node186 = (inp[10]) ? 3'b000 : 3'b001;
								assign node190 = (inp[0]) ? 3'b000 : 3'b001;
							assign node193 = (inp[4]) ? node205 : node194;
								assign node194 = (inp[0]) ? 3'b000 : node195;
									assign node195 = (inp[7]) ? node197 : 3'b000;
										assign node197 = (inp[10]) ? 3'b000 : node198;
											assign node198 = (inp[2]) ? 3'b001 : node199;
												assign node199 = (inp[11]) ? 3'b000 : 3'b001;
								assign node205 = (inp[11]) ? node213 : node206;
									assign node206 = (inp[0]) ? node210 : node207;
										assign node207 = (inp[7]) ? 3'b001 : 3'b000;
										assign node210 = (inp[7]) ? 3'b000 : 3'b001;
									assign node213 = (inp[2]) ? node221 : node214;
										assign node214 = (inp[7]) ? node218 : node215;
											assign node215 = (inp[0]) ? 3'b001 : 3'b000;
											assign node218 = (inp[0]) ? 3'b000 : 3'b001;
										assign node221 = (inp[0]) ? node223 : 3'b000;
											assign node223 = (inp[7]) ? 3'b000 : 3'b001;
					assign node226 = (inp[4]) ? node314 : node227;
						assign node227 = (inp[0]) ? node283 : node228;
							assign node228 = (inp[6]) ? node254 : node229;
								assign node229 = (inp[5]) ? node239 : node230;
									assign node230 = (inp[10]) ? node236 : node231;
										assign node231 = (inp[7]) ? node233 : 3'b000;
											assign node233 = (inp[2]) ? 3'b000 : 3'b001;
										assign node236 = (inp[7]) ? 3'b000 : 3'b001;
									assign node239 = (inp[11]) ? node247 : node240;
										assign node240 = (inp[7]) ? node244 : node241;
											assign node241 = (inp[10]) ? 3'b001 : 3'b000;
											assign node244 = (inp[10]) ? 3'b000 : 3'b001;
										assign node247 = (inp[2]) ? 3'b001 : node248;
											assign node248 = (inp[7]) ? node250 : 3'b001;
												assign node250 = (inp[10]) ? 3'b001 : 3'b000;
								assign node254 = (inp[5]) ? node270 : node255;
									assign node255 = (inp[11]) ? node263 : node256;
										assign node256 = (inp[7]) ? node260 : node257;
											assign node257 = (inp[10]) ? 3'b000 : 3'b001;
											assign node260 = (inp[10]) ? 3'b001 : 3'b000;
										assign node263 = (inp[7]) ? node267 : node264;
											assign node264 = (inp[10]) ? 3'b000 : 3'b001;
											assign node267 = (inp[10]) ? 3'b001 : 3'b000;
									assign node270 = (inp[10]) ? 3'b000 : node271;
										assign node271 = (inp[7]) ? node277 : node272;
											assign node272 = (inp[2]) ? node274 : 3'b000;
												assign node274 = (inp[11]) ? 3'b000 : 3'b001;
											assign node277 = (inp[2]) ? node279 : 3'b001;
												assign node279 = (inp[11]) ? 3'b001 : 3'b000;
							assign node283 = (inp[6]) ? 3'b001 : node284;
								assign node284 = (inp[11]) ? node290 : node285;
									assign node285 = (inp[7]) ? 3'b001 : node286;
										assign node286 = (inp[5]) ? 3'b001 : 3'b000;
									assign node290 = (inp[2]) ? node304 : node291;
										assign node291 = (inp[10]) ? node299 : node292;
											assign node292 = (inp[7]) ? node296 : node293;
												assign node293 = (inp[5]) ? 3'b001 : 3'b000;
												assign node296 = (inp[5]) ? 3'b000 : 3'b001;
											assign node299 = (inp[5]) ? 3'b000 : node300;
												assign node300 = (inp[7]) ? 3'b001 : 3'b000;
										assign node304 = (inp[10]) ? 3'b001 : node305;
											assign node305 = (inp[7]) ? node309 : node306;
												assign node306 = (inp[5]) ? 3'b001 : 3'b000;
												assign node309 = (inp[5]) ? 3'b000 : 3'b001;
						assign node314 = (inp[7]) ? node326 : node315;
							assign node315 = (inp[5]) ? node323 : node316;
								assign node316 = (inp[0]) ? 3'b000 : node317;
									assign node317 = (inp[10]) ? node319 : 3'b001;
										assign node319 = (inp[6]) ? 3'b001 : 3'b000;
								assign node323 = (inp[0]) ? 3'b001 : 3'b000;
							assign node326 = (inp[6]) ? node344 : node327;
								assign node327 = (inp[0]) ? 3'b001 : node328;
									assign node328 = (inp[10]) ? node338 : node329;
										assign node329 = (inp[2]) ? node335 : node330;
											assign node330 = (inp[5]) ? node332 : 3'b000;
												assign node332 = (inp[11]) ? 3'b001 : 3'b000;
											assign node335 = (inp[5]) ? 3'b000 : 3'b001;
										assign node338 = (inp[11]) ? node340 : 3'b001;
											assign node340 = (inp[5]) ? 3'b000 : 3'b001;
								assign node344 = (inp[0]) ? 3'b000 : node345;
									assign node345 = (inp[2]) ? node347 : 3'b001;
										assign node347 = (inp[5]) ? 3'b001 : 3'b000;
			assign node351 = (inp[4]) ? node617 : node352;
				assign node352 = (inp[6]) ? node478 : node353;
					assign node353 = (inp[0]) ? node421 : node354;
						assign node354 = (inp[1]) ? node362 : node355;
							assign node355 = (inp[7]) ? node359 : node356;
								assign node356 = (inp[5]) ? 3'b100 : 3'b010;
								assign node359 = (inp[5]) ? 3'b010 : 3'b110;
							assign node362 = (inp[7]) ? node378 : node363;
								assign node363 = (inp[5]) ? node371 : node364;
									assign node364 = (inp[10]) ? 3'b110 : node365;
										assign node365 = (inp[8]) ? 3'b101 : node366;
											assign node366 = (inp[2]) ? 3'b110 : 3'b101;
									assign node371 = (inp[10]) ? 3'b010 : node372;
										assign node372 = (inp[8]) ? node374 : 3'b010;
											assign node374 = (inp[11]) ? 3'b010 : 3'b001;
								assign node378 = (inp[5]) ? node400 : node379;
									assign node379 = (inp[10]) ? node393 : node380;
										assign node380 = (inp[11]) ? node388 : node381;
											assign node381 = (inp[8]) ? node385 : node382;
												assign node382 = (inp[2]) ? 3'b010 : 3'b001;
												assign node385 = (inp[2]) ? 3'b001 : 3'b010;
											assign node388 = (inp[8]) ? 3'b010 : node389;
												assign node389 = (inp[2]) ? 3'b010 : 3'b101;
										assign node393 = (inp[8]) ? 3'b001 : node394;
											assign node394 = (inp[2]) ? 3'b001 : node395;
												assign node395 = (inp[11]) ? 3'b110 : 3'b010;
									assign node400 = (inp[2]) ? node412 : node401;
										assign node401 = (inp[8]) ? node405 : node402;
											assign node402 = (inp[10]) ? 3'b010 : 3'b001;
											assign node405 = (inp[11]) ? node409 : node406;
												assign node406 = (inp[10]) ? 3'b101 : 3'b110;
												assign node409 = (inp[10]) ? 3'b110 : 3'b101;
										assign node412 = (inp[11]) ? node416 : node413;
											assign node413 = (inp[10]) ? 3'b101 : 3'b110;
											assign node416 = (inp[8]) ? 3'b110 : node417;
												assign node417 = (inp[10]) ? 3'b110 : 3'b101;
						assign node421 = (inp[5]) ? node447 : node422;
							assign node422 = (inp[8]) ? node438 : node423;
								assign node423 = (inp[1]) ? node433 : node424;
									assign node424 = (inp[7]) ? node430 : node425;
										assign node425 = (inp[2]) ? 3'b001 : node426;
											assign node426 = (inp[11]) ? 3'b110 : 3'b010;
										assign node430 = (inp[2]) ? 3'b101 : 3'b001;
									assign node433 = (inp[11]) ? node435 : 3'b101;
										assign node435 = (inp[7]) ? 3'b101 : 3'b001;
								assign node438 = (inp[7]) ? node444 : node439;
									assign node439 = (inp[1]) ? node441 : 3'b001;
										assign node441 = (inp[11]) ? 3'b000 : 3'b100;
									assign node444 = (inp[1]) ? 3'b011 : 3'b001;
							assign node447 = (inp[1]) ? node465 : node448;
								assign node448 = (inp[7]) ? node458 : node449;
									assign node449 = (inp[8]) ? node453 : node450;
										assign node450 = (inp[2]) ? 3'b110 : 3'b010;
										assign node453 = (inp[11]) ? 3'b110 : node454;
											assign node454 = (inp[2]) ? 3'b110 : 3'b101;
									assign node458 = (inp[11]) ? 3'b110 : node459;
										assign node459 = (inp[2]) ? node461 : 3'b110;
											assign node461 = (inp[8]) ? 3'b010 : 3'b110;
								assign node465 = (inp[7]) ? node471 : node466;
									assign node466 = (inp[11]) ? node468 : 3'b111;
										assign node468 = (inp[8]) ? 3'b111 : 3'b110;
									assign node471 = (inp[11]) ? node475 : node472;
										assign node472 = (inp[8]) ? 3'b111 : 3'b101;
										assign node475 = (inp[8]) ? 3'b101 : 3'b001;
					assign node478 = (inp[1]) ? node536 : node479;
						assign node479 = (inp[5]) ? node507 : node480;
							assign node480 = (inp[7]) ? node486 : node481;
								assign node481 = (inp[10]) ? node483 : 3'b101;
									assign node483 = (inp[0]) ? 3'b101 : 3'b001;
								assign node486 = (inp[10]) ? node494 : node487;
									assign node487 = (inp[0]) ? node489 : 3'b001;
										assign node489 = (inp[8]) ? node491 : 3'b001;
											assign node491 = (inp[2]) ? 3'b101 : 3'b001;
									assign node494 = (inp[0]) ? node502 : node495;
										assign node495 = (inp[2]) ? 3'b101 : node496;
											assign node496 = (inp[8]) ? 3'b101 : node497;
												assign node497 = (inp[11]) ? 3'b001 : 3'b101;
										assign node502 = (inp[8]) ? node504 : 3'b011;
											assign node504 = (inp[2]) ? 3'b111 : 3'b011;
							assign node507 = (inp[0]) ? node523 : node508;
								assign node508 = (inp[7]) ? node516 : node509;
									assign node509 = (inp[2]) ? 3'b110 : node510;
										assign node510 = (inp[8]) ? 3'b110 : node511;
											assign node511 = (inp[10]) ? 3'b010 : 3'b110;
									assign node516 = (inp[8]) ? 3'b001 : node517;
										assign node517 = (inp[10]) ? node519 : 3'b010;
											assign node519 = (inp[2]) ? 3'b010 : 3'b110;
								assign node523 = (inp[7]) ? node525 : 3'b101;
									assign node525 = (inp[2]) ? node527 : 3'b101;
										assign node527 = (inp[10]) ? node533 : node528;
											assign node528 = (inp[8]) ? node530 : 3'b001;
												assign node530 = (inp[11]) ? 3'b001 : 3'b101;
											assign node533 = (inp[11]) ? 3'b011 : 3'b111;
						assign node536 = (inp[5]) ? node568 : node537;
							assign node537 = (inp[0]) ? node559 : node538;
								assign node538 = (inp[7]) ? node550 : node539;
									assign node539 = (inp[10]) ? node545 : node540;
										assign node540 = (inp[2]) ? node542 : 3'b011;
											assign node542 = (inp[8]) ? 3'b011 : 3'b001;
										assign node545 = (inp[8]) ? 3'b101 : node546;
											assign node546 = (inp[2]) ? 3'b101 : 3'b001;
									assign node550 = (inp[8]) ? node556 : node551;
										assign node551 = (inp[2]) ? node553 : 3'b011;
											assign node553 = (inp[10]) ? 3'b001 : 3'b011;
										assign node556 = (inp[10]) ? 3'b011 : 3'b001;
								assign node559 = (inp[7]) ? 3'b111 : node560;
									assign node560 = (inp[2]) ? node562 : 3'b011;
										assign node562 = (inp[10]) ? node564 : 3'b011;
											assign node564 = (inp[8]) ? 3'b111 : 3'b011;
							assign node568 = (inp[8]) ? node590 : node569;
								assign node569 = (inp[10]) ? node577 : node570;
									assign node570 = (inp[0]) ? 3'b001 : node571;
										assign node571 = (inp[7]) ? node573 : 3'b001;
											assign node573 = (inp[2]) ? 3'b011 : 3'b001;
									assign node577 = (inp[2]) ? node579 : 3'b001;
										assign node579 = (inp[11]) ? node585 : node580;
											assign node580 = (inp[0]) ? 3'b001 : node581;
												assign node581 = (inp[7]) ? 3'b101 : 3'b001;
											assign node585 = (inp[7]) ? node587 : 3'b101;
												assign node587 = (inp[0]) ? 3'b001 : 3'b101;
								assign node590 = (inp[0]) ? 3'b011 : node591;
									assign node591 = (inp[10]) ? node603 : node592;
										assign node592 = (inp[7]) ? node598 : node593;
											assign node593 = (inp[11]) ? 3'b001 : node594;
												assign node594 = (inp[2]) ? 3'b011 : 3'b001;
											assign node598 = (inp[11]) ? 3'b011 : node599;
												assign node599 = (inp[2]) ? 3'b001 : 3'b011;
										assign node603 = (inp[11]) ? node611 : node604;
											assign node604 = (inp[7]) ? node608 : node605;
												assign node605 = (inp[2]) ? 3'b001 : 3'b101;
												assign node608 = (inp[2]) ? 3'b111 : 3'b001;
											assign node611 = (inp[7]) ? node613 : 3'b001;
												assign node613 = (inp[2]) ? 3'b101 : 3'b001;
				assign node617 = (inp[0]) ? node753 : node618;
					assign node618 = (inp[6]) ? node702 : node619;
						assign node619 = (inp[5]) ? node661 : node620;
							assign node620 = (inp[1]) ? node632 : node621;
								assign node621 = (inp[7]) ? 3'b100 : node622;
									assign node622 = (inp[10]) ? node624 : 3'b100;
										assign node624 = (inp[2]) ? node626 : 3'b000;
											assign node626 = (inp[8]) ? 3'b100 : node627;
												assign node627 = (inp[11]) ? 3'b000 : 3'b100;
								assign node632 = (inp[7]) ? node640 : node633;
									assign node633 = (inp[10]) ? 3'b100 : node634;
										assign node634 = (inp[8]) ? 3'b110 : node635;
											assign node635 = (inp[2]) ? 3'b100 : 3'b010;
									assign node640 = (inp[2]) ? node656 : node641;
										assign node641 = (inp[11]) ? node649 : node642;
											assign node642 = (inp[10]) ? node646 : node643;
												assign node643 = (inp[8]) ? 3'b000 : 3'b010;
												assign node646 = (inp[8]) ? 3'b010 : 3'b000;
											assign node649 = (inp[8]) ? node653 : node650;
												assign node650 = (inp[10]) ? 3'b100 : 3'b110;
												assign node653 = (inp[10]) ? 3'b010 : 3'b000;
										assign node656 = (inp[10]) ? 3'b010 : node657;
											assign node657 = (inp[8]) ? 3'b010 : 3'b000;
							assign node661 = (inp[1]) ? node673 : node662;
								assign node662 = (inp[8]) ? 3'b000 : node663;
									assign node663 = (inp[11]) ? 3'b000 : node664;
										assign node664 = (inp[2]) ? node666 : 3'b000;
											assign node666 = (inp[7]) ? 3'b000 : node667;
												assign node667 = (inp[10]) ? 3'b100 : 3'b000;
								assign node673 = (inp[7]) ? node683 : node674;
									assign node674 = (inp[8]) ? node676 : 3'b000;
										assign node676 = (inp[2]) ? node680 : node677;
											assign node677 = (inp[11]) ? 3'b000 : 3'b100;
											assign node680 = (inp[10]) ? 3'b000 : 3'b010;
									assign node683 = (inp[8]) ? node693 : node684;
										assign node684 = (inp[2]) ? node688 : node685;
											assign node685 = (inp[10]) ? 3'b000 : 3'b010;
											assign node688 = (inp[11]) ? node690 : 3'b110;
												assign node690 = (inp[10]) ? 3'b100 : 3'b110;
										assign node693 = (inp[10]) ? node699 : node694;
											assign node694 = (inp[11]) ? node696 : 3'b100;
												assign node696 = (inp[2]) ? 3'b100 : 3'b110;
											assign node699 = (inp[11]) ? 3'b100 : 3'b110;
						assign node702 = (inp[1]) ? node736 : node703;
							assign node703 = (inp[8]) ? node721 : node704;
								assign node704 = (inp[7]) ? node706 : 3'b100;
									assign node706 = (inp[10]) ? node712 : node707;
										assign node707 = (inp[11]) ? node709 : 3'b000;
											assign node709 = (inp[5]) ? 3'b100 : 3'b000;
										assign node712 = (inp[5]) ? node714 : 3'b010;
											assign node714 = (inp[2]) ? node718 : node715;
												assign node715 = (inp[11]) ? 3'b100 : 3'b000;
												assign node718 = (inp[11]) ? 3'b110 : 3'b010;
								assign node721 = (inp[10]) ? node731 : node722;
									assign node722 = (inp[7]) ? node728 : node723;
										assign node723 = (inp[11]) ? node725 : 3'b010;
											assign node725 = (inp[5]) ? 3'b100 : 3'b010;
										assign node728 = (inp[5]) ? 3'b000 : 3'b100;
									assign node731 = (inp[7]) ? node733 : 3'b010;
										assign node733 = (inp[5]) ? 3'b010 : 3'b110;
							assign node736 = (inp[7]) ? node740 : node737;
								assign node737 = (inp[5]) ? 3'b100 : 3'b110;
								assign node740 = (inp[2]) ? node744 : node741;
									assign node741 = (inp[5]) ? 3'b010 : 3'b110;
									assign node744 = (inp[8]) ? node750 : node745;
										assign node745 = (inp[5]) ? node747 : 3'b110;
											assign node747 = (inp[11]) ? 3'b101 : 3'b110;
										assign node750 = (inp[5]) ? 3'b110 : 3'b001;
					assign node753 = (inp[6]) ? node789 : node754;
						assign node754 = (inp[5]) ? node772 : node755;
							assign node755 = (inp[1]) ? node765 : node756;
								assign node756 = (inp[7]) ? 3'b010 : node757;
									assign node757 = (inp[8]) ? 3'b010 : node758;
										assign node758 = (inp[2]) ? 3'b010 : node759;
											assign node759 = (inp[11]) ? 3'b100 : 3'b000;
								assign node765 = (inp[8]) ? node769 : node766;
									assign node766 = (inp[7]) ? 3'b110 : 3'b010;
									assign node769 = (inp[7]) ? 3'b110 : 3'b100;
							assign node772 = (inp[1]) ? node782 : node773;
								assign node773 = (inp[7]) ? 3'b100 : node774;
									assign node774 = (inp[2]) ? 3'b100 : node775;
										assign node775 = (inp[8]) ? node777 : 3'b000;
											assign node777 = (inp[11]) ? 3'b100 : 3'b110;
								assign node782 = (inp[8]) ? 3'b010 : node783;
									assign node783 = (inp[11]) ? node785 : 3'b010;
										assign node785 = (inp[7]) ? 3'b010 : 3'b100;
						assign node789 = (inp[5]) ? node799 : node790;
							assign node790 = (inp[7]) ? node792 : 3'b001;
								assign node792 = (inp[1]) ? 3'b101 : node793;
									assign node793 = (inp[2]) ? node795 : 3'b001;
										assign node795 = (inp[10]) ? 3'b101 : 3'b001;
							assign node799 = (inp[1]) ? node805 : node800;
								assign node800 = (inp[10]) ? node802 : 3'b010;
									assign node802 = (inp[7]) ? 3'b110 : 3'b010;
								assign node805 = (inp[7]) ? 3'b001 : 3'b110;
		assign node808 = (inp[6]) ? node830 : node809;
			assign node809 = (inp[4]) ? 3'b000 : node810;
				assign node810 = (inp[9]) ? node812 : 3'b000;
					assign node812 = (inp[0]) ? node814 : 3'b000;
						assign node814 = (inp[1]) ? node816 : 3'b000;
							assign node816 = (inp[5]) ? node822 : node817;
								assign node817 = (inp[7]) ? 3'b100 : node818;
									assign node818 = (inp[8]) ? 3'b100 : 3'b000;
								assign node822 = (inp[8]) ? node824 : 3'b000;
									assign node824 = (inp[11]) ? 3'b000 : node825;
										assign node825 = (inp[7]) ? 3'b000 : 3'b100;
			assign node830 = (inp[9]) ? node1016 : node831;
				assign node831 = (inp[4]) ? node855 : node832;
					assign node832 = (inp[0]) ? node848 : node833;
						assign node833 = (inp[7]) ? node835 : 3'b010;
							assign node835 = (inp[1]) ? node837 : 3'b010;
								assign node837 = (inp[2]) ? node839 : 3'b010;
									assign node839 = (inp[8]) ? node845 : node840;
										assign node840 = (inp[11]) ? node842 : 3'b010;
											assign node842 = (inp[5]) ? 3'b011 : 3'b010;
										assign node845 = (inp[5]) ? 3'b010 : 3'b011;
						assign node848 = (inp[5]) ? node850 : 3'b011;
							assign node850 = (inp[7]) ? node852 : 3'b010;
								assign node852 = (inp[1]) ? 3'b011 : 3'b010;
					assign node855 = (inp[0]) ? node925 : node856;
						assign node856 = (inp[10]) ? node902 : node857;
							assign node857 = (inp[7]) ? node875 : node858;
								assign node858 = (inp[1]) ? node870 : node859;
									assign node859 = (inp[5]) ? node865 : node860;
										assign node860 = (inp[2]) ? node862 : 3'b010;
											assign node862 = (inp[8]) ? 3'b010 : 3'b000;
										assign node865 = (inp[8]) ? node867 : 3'b000;
											assign node867 = (inp[11]) ? 3'b000 : 3'b010;
									assign node870 = (inp[5]) ? node872 : 3'b000;
										assign node872 = (inp[11]) ? 3'b100 : 3'b000;
								assign node875 = (inp[5]) ? node889 : node876;
									assign node876 = (inp[2]) ? node882 : node877;
										assign node877 = (inp[8]) ? 3'b010 : node878;
											assign node878 = (inp[1]) ? 3'b010 : 3'b110;
										assign node882 = (inp[8]) ? node886 : node883;
											assign node883 = (inp[1]) ? 3'b010 : 3'b100;
											assign node886 = (inp[1]) ? 3'b100 : 3'b010;
									assign node889 = (inp[11]) ? node895 : node890;
										assign node890 = (inp[1]) ? 3'b010 : node891;
											assign node891 = (inp[8]) ? 3'b010 : 3'b100;
										assign node895 = (inp[1]) ? node897 : 3'b100;
											assign node897 = (inp[2]) ? node899 : 3'b100;
												assign node899 = (inp[8]) ? 3'b010 : 3'b100;
							assign node902 = (inp[1]) ? node904 : 3'b000;
								assign node904 = (inp[5]) ? node914 : node905;
									assign node905 = (inp[2]) ? 3'b000 : node906;
										assign node906 = (inp[8]) ? 3'b000 : node907;
											assign node907 = (inp[11]) ? node909 : 3'b000;
												assign node909 = (inp[7]) ? 3'b100 : 3'b000;
									assign node914 = (inp[11]) ? node920 : node915;
										assign node915 = (inp[7]) ? node917 : 3'b000;
											assign node917 = (inp[8]) ? 3'b100 : 3'b000;
										assign node920 = (inp[7]) ? node922 : 3'b100;
											assign node922 = (inp[8]) ? 3'b100 : 3'b000;
						assign node925 = (inp[7]) ? node955 : node926;
							assign node926 = (inp[10]) ? node946 : node927;
								assign node927 = (inp[1]) ? node935 : node928;
									assign node928 = (inp[5]) ? 3'b100 : node929;
										assign node929 = (inp[8]) ? 3'b010 : node930;
											assign node930 = (inp[2]) ? 3'b100 : 3'b010;
									assign node935 = (inp[2]) ? node941 : node936;
										assign node936 = (inp[8]) ? node938 : 3'b010;
											assign node938 = (inp[11]) ? 3'b010 : 3'b110;
										assign node941 = (inp[11]) ? node943 : 3'b110;
											assign node943 = (inp[5]) ? 3'b010 : 3'b110;
								assign node946 = (inp[1]) ? node948 : 3'b100;
									assign node948 = (inp[8]) ? node950 : 3'b100;
										assign node950 = (inp[5]) ? node952 : 3'b010;
											assign node952 = (inp[11]) ? 3'b100 : 3'b010;
							assign node955 = (inp[10]) ? node989 : node956;
								assign node956 = (inp[1]) ? node972 : node957;
									assign node957 = (inp[2]) ? node963 : node958;
										assign node958 = (inp[8]) ? node960 : 3'b010;
											assign node960 = (inp[5]) ? 3'b010 : 3'b110;
										assign node963 = (inp[11]) ? node965 : 3'b110;
											assign node965 = (inp[8]) ? node969 : node966;
												assign node966 = (inp[5]) ? 3'b010 : 3'b110;
												assign node969 = (inp[5]) ? 3'b110 : 3'b010;
									assign node972 = (inp[5]) ? node982 : node973;
										assign node973 = (inp[8]) ? node977 : node974;
											assign node974 = (inp[2]) ? 3'b110 : 3'b101;
											assign node977 = (inp[11]) ? node979 : 3'b101;
												assign node979 = (inp[2]) ? 3'b101 : 3'b001;
										assign node982 = (inp[8]) ? 3'b110 : node983;
											assign node983 = (inp[2]) ? 3'b110 : node984;
												assign node984 = (inp[11]) ? 3'b010 : 3'b110;
								assign node989 = (inp[2]) ? node1001 : node990;
									assign node990 = (inp[1]) ? node998 : node991;
										assign node991 = (inp[8]) ? node993 : 3'b100;
											assign node993 = (inp[5]) ? node995 : 3'b010;
												assign node995 = (inp[11]) ? 3'b100 : 3'b010;
										assign node998 = (inp[5]) ? 3'b010 : 3'b110;
									assign node1001 = (inp[8]) ? node1009 : node1002;
										assign node1002 = (inp[1]) ? 3'b010 : node1003;
											assign node1003 = (inp[5]) ? node1005 : 3'b010;
												assign node1005 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1009 = (inp[1]) ? node1011 : 3'b010;
											assign node1011 = (inp[11]) ? node1013 : 3'b110;
												assign node1013 = (inp[5]) ? 3'b010 : 3'b110;
				assign node1016 = (inp[0]) ? node1058 : node1017;
					assign node1017 = (inp[4]) ? 3'b000 : node1018;
						assign node1018 = (inp[10]) ? node1034 : node1019;
							assign node1019 = (inp[1]) ? node1021 : 3'b000;
								assign node1021 = (inp[2]) ? node1023 : 3'b000;
									assign node1023 = (inp[7]) ? node1025 : 3'b000;
										assign node1025 = (inp[5]) ? node1029 : node1026;
											assign node1026 = (inp[8]) ? 3'b010 : 3'b000;
											assign node1029 = (inp[8]) ? 3'b000 : node1030;
												assign node1030 = (inp[11]) ? 3'b010 : 3'b000;
							assign node1034 = (inp[1]) ? node1042 : node1035;
								assign node1035 = (inp[8]) ? node1037 : 3'b000;
									assign node1037 = (inp[7]) ? node1039 : 3'b000;
										assign node1039 = (inp[5]) ? 3'b000 : 3'b100;
								assign node1042 = (inp[2]) ? node1048 : node1043;
									assign node1043 = (inp[7]) ? node1045 : 3'b000;
										assign node1045 = (inp[5]) ? 3'b000 : 3'b100;
									assign node1048 = (inp[7]) ? node1050 : 3'b100;
										assign node1050 = (inp[8]) ? node1052 : 3'b100;
											assign node1052 = (inp[5]) ? node1054 : 3'b010;
												assign node1054 = (inp[11]) ? 3'b100 : 3'b000;
					assign node1058 = (inp[4]) ? node1070 : node1059;
						assign node1059 = (inp[5]) ? node1065 : node1060;
							assign node1060 = (inp[1]) ? node1062 : 3'b010;
								assign node1062 = (inp[7]) ? 3'b110 : 3'b010;
							assign node1065 = (inp[1]) ? node1067 : 3'b100;
								assign node1067 = (inp[7]) ? 3'b010 : 3'b100;
						assign node1070 = (inp[1]) ? node1082 : node1071;
							assign node1071 = (inp[8]) ? node1073 : 3'b000;
								assign node1073 = (inp[10]) ? 3'b000 : node1074;
									assign node1074 = (inp[7]) ? node1076 : 3'b000;
										assign node1076 = (inp[5]) ? node1078 : 3'b100;
											assign node1078 = (inp[11]) ? 3'b000 : 3'b100;
							assign node1082 = (inp[10]) ? node1112 : node1083;
								assign node1083 = (inp[7]) ? node1095 : node1084;
									assign node1084 = (inp[8]) ? node1090 : node1085;
										assign node1085 = (inp[2]) ? 3'b000 : node1086;
											assign node1086 = (inp[5]) ? 3'b000 : 3'b100;
										assign node1090 = (inp[5]) ? node1092 : 3'b100;
											assign node1092 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1095 = (inp[5]) ? node1101 : node1096;
										assign node1096 = (inp[8]) ? 3'b010 : node1097;
											assign node1097 = (inp[2]) ? 3'b100 : 3'b110;
										assign node1101 = (inp[2]) ? node1107 : node1102;
											assign node1102 = (inp[8]) ? 3'b100 : node1103;
												assign node1103 = (inp[11]) ? 3'b000 : 3'b100;
											assign node1107 = (inp[8]) ? node1109 : 3'b100;
												assign node1109 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1112 = (inp[5]) ? 3'b000 : node1113;
									assign node1113 = (inp[7]) ? node1115 : 3'b000;
										assign node1115 = (inp[2]) ? node1117 : 3'b100;
											assign node1117 = (inp[8]) ? 3'b100 : 3'b000;

endmodule