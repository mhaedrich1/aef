module dtc_split66_bm66 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node9;
	wire [4-1:0] node11;
	wire [4-1:0] node13;
	wire [4-1:0] node14;
	wire [4-1:0] node16;
	wire [4-1:0] node18;
	wire [4-1:0] node21;
	wire [4-1:0] node22;
	wire [4-1:0] node24;
	wire [4-1:0] node26;
	wire [4-1:0] node30;
	wire [4-1:0] node31;
	wire [4-1:0] node32;
	wire [4-1:0] node34;
	wire [4-1:0] node35;
	wire [4-1:0] node37;
	wire [4-1:0] node39;
	wire [4-1:0] node41;
	wire [4-1:0] node45;
	wire [4-1:0] node46;
	wire [4-1:0] node47;
	wire [4-1:0] node48;
	wire [4-1:0] node50;
	wire [4-1:0] node52;
	wire [4-1:0] node59;
	wire [4-1:0] node60;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node66;
	wire [4-1:0] node68;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node74;
	wire [4-1:0] node76;
	wire [4-1:0] node78;
	wire [4-1:0] node79;
	wire [4-1:0] node81;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node87;
	wire [4-1:0] node88;
	wire [4-1:0] node90;
	wire [4-1:0] node92;
	wire [4-1:0] node98;
	wire [4-1:0] node99;
	wire [4-1:0] node100;
	wire [4-1:0] node102;
	wire [4-1:0] node104;
	wire [4-1:0] node105;
	wire [4-1:0] node107;
	wire [4-1:0] node108;
	wire [4-1:0] node110;
	wire [4-1:0] node112;
	wire [4-1:0] node114;
	wire [4-1:0] node118;
	wire [4-1:0] node119;
	wire [4-1:0] node120;
	wire [4-1:0] node121;
	wire [4-1:0] node123;
	wire [4-1:0] node125;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node133;
	wire [4-1:0] node134;
	wire [4-1:0] node136;
	wire [4-1:0] node138;
	wire [4-1:0] node140;
	wire [4-1:0] node142;
	wire [4-1:0] node144;
	wire [4-1:0] node147;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node152;
	wire [4-1:0] node154;
	wire [4-1:0] node155;
	wire [4-1:0] node157;
	wire [4-1:0] node159;
	wire [4-1:0] node166;
	wire [4-1:0] node167;
	wire [4-1:0] node169;
	wire [4-1:0] node171;
	wire [4-1:0] node172;
	wire [4-1:0] node173;
	wire [4-1:0] node175;
	wire [4-1:0] node177;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node184;
	wire [4-1:0] node185;
	wire [4-1:0] node187;
	wire [4-1:0] node189;
	wire [4-1:0] node191;
	wire [4-1:0] node196;
	wire [4-1:0] node198;
	wire [4-1:0] node200;
	wire [4-1:0] node201;
	wire [4-1:0] node203;
	wire [4-1:0] node205;
	wire [4-1:0] node207;
	wire [4-1:0] node209;
	wire [4-1:0] node213;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node218;
	wire [4-1:0] node219;
	wire [4-1:0] node221;
	wire [4-1:0] node222;
	wire [4-1:0] node224;
	wire [4-1:0] node226;
	wire [4-1:0] node231;
	wire [4-1:0] node232;
	wire [4-1:0] node233;
	wire [4-1:0] node235;
	wire [4-1:0] node237;
	wire [4-1:0] node242;
	wire [4-1:0] node243;
	wire [4-1:0] node245;
	wire [4-1:0] node247;
	wire [4-1:0] node250;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node254;
	wire [4-1:0] node259;
	wire [4-1:0] node261;
	wire [4-1:0] node262;
	wire [4-1:0] node264;
	wire [4-1:0] node266;
	wire [4-1:0] node268;
	wire [4-1:0] node270;
	wire [4-1:0] node273;
	wire [4-1:0] node276;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node281;
	wire [4-1:0] node283;
	wire [4-1:0] node284;
	wire [4-1:0] node286;
	wire [4-1:0] node288;
	wire [4-1:0] node290;
	wire [4-1:0] node295;
	wire [4-1:0] node296;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node301;
	wire [4-1:0] node303;
	wire [4-1:0] node305;
	wire [4-1:0] node307;
	wire [4-1:0] node312;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node316;
	wire [4-1:0] node318;
	wire [4-1:0] node320;
	wire [4-1:0] node325;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node332;
	wire [4-1:0] node334;
	wire [4-1:0] node340;
	wire [4-1:0] node342;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node346;
	wire [4-1:0] node348;
	wire [4-1:0] node350;
	wire [4-1:0] node352;
	wire [4-1:0] node357;
	wire [4-1:0] node358;
	wire [4-1:0] node359;
	wire [4-1:0] node360;
	wire [4-1:0] node361;
	wire [4-1:0] node362;
	wire [4-1:0] node364;
	wire [4-1:0] node366;
	wire [4-1:0] node368;
	wire [4-1:0] node372;
	wire [4-1:0] node374;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node378;
	wire [4-1:0] node380;
	wire [4-1:0] node382;
	wire [4-1:0] node385;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node392;
	wire [4-1:0] node393;
	wire [4-1:0] node394;
	wire [4-1:0] node396;
	wire [4-1:0] node398;
	wire [4-1:0] node400;
	wire [4-1:0] node405;
	wire [4-1:0] node407;
	wire [4-1:0] node408;
	wire [4-1:0] node410;
	wire [4-1:0] node412;
	wire [4-1:0] node416;
	wire [4-1:0] node417;
	wire [4-1:0] node418;
	wire [4-1:0] node420;
	wire [4-1:0] node422;
	wire [4-1:0] node426;
	wire [4-1:0] node427;
	wire [4-1:0] node429;
	wire [4-1:0] node431;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node435;
	wire [4-1:0] node440;
	wire [4-1:0] node442;
	wire [4-1:0] node444;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node449;
	wire [4-1:0] node450;
	wire [4-1:0] node451;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node456;
	wire [4-1:0] node458;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node469;
	wire [4-1:0] node471;
	wire [4-1:0] node473;
	wire [4-1:0] node478;
	wire [4-1:0] node480;
	wire [4-1:0] node482;
	wire [4-1:0] node483;
	wire [4-1:0] node484;
	wire [4-1:0] node486;
	wire [4-1:0] node488;
	wire [4-1:0] node490;
	wire [4-1:0] node493;
	wire [4-1:0] node496;
	wire [4-1:0] node498;
	wire [4-1:0] node500;
	wire [4-1:0] node502;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node511;
	wire [4-1:0] node513;
	wire [4-1:0] node515;
	wire [4-1:0] node520;
	wire [4-1:0] node523;
	wire [4-1:0] node525;
	wire [4-1:0] node527;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node532;
	wire [4-1:0] node536;
	wire [4-1:0] node537;
	wire [4-1:0] node538;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node541;
	wire [4-1:0] node543;
	wire [4-1:0] node544;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node548;
	wire [4-1:0] node550;
	wire [4-1:0] node556;
	wire [4-1:0] node557;
	wire [4-1:0] node559;
	wire [4-1:0] node561;
	wire [4-1:0] node562;
	wire [4-1:0] node564;
	wire [4-1:0] node568;
	wire [4-1:0] node570;
	wire [4-1:0] node572;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node578;
	wire [4-1:0] node579;
	wire [4-1:0] node580;
	wire [4-1:0] node582;
	wire [4-1:0] node583;
	wire [4-1:0] node585;
	wire [4-1:0] node587;
	wire [4-1:0] node593;
	wire [4-1:0] node595;
	wire [4-1:0] node596;
	wire [4-1:0] node598;
	wire [4-1:0] node600;
	wire [4-1:0] node601;
	wire [4-1:0] node603;
	wire [4-1:0] node605;
	wire [4-1:0] node610;
	wire [4-1:0] node611;
	wire [4-1:0] node612;
	wire [4-1:0] node613;
	wire [4-1:0] node615;
	wire [4-1:0] node617;
	wire [4-1:0] node620;
	wire [4-1:0] node622;
	wire [4-1:0] node624;
	wire [4-1:0] node626;
	wire [4-1:0] node628;
	wire [4-1:0] node632;
	wire [4-1:0] node633;
	wire [4-1:0] node634;
	wire [4-1:0] node636;
	wire [4-1:0] node638;
	wire [4-1:0] node640;
	wire [4-1:0] node642;
	wire [4-1:0] node644;
	wire [4-1:0] node646;
	wire [4-1:0] node649;
	wire [4-1:0] node650;
	wire [4-1:0] node651;
	wire [4-1:0] node652;
	wire [4-1:0] node653;
	wire [4-1:0] node655;
	wire [4-1:0] node663;
	wire [4-1:0] node664;
	wire [4-1:0] node665;
	wire [4-1:0] node666;
	wire [4-1:0] node667;
	wire [4-1:0] node668;
	wire [4-1:0] node669;
	wire [4-1:0] node673;
	wire [4-1:0] node675;
	wire [4-1:0] node677;
	wire [4-1:0] node679;
	wire [4-1:0] node681;
	wire [4-1:0] node683;
	wire [4-1:0] node686;
	wire [4-1:0] node687;
	wire [4-1:0] node688;
	wire [4-1:0] node689;
	wire [4-1:0] node691;
	wire [4-1:0] node696;
	wire [4-1:0] node698;
	wire [4-1:0] node701;
	wire [4-1:0] node703;
	wire [4-1:0] node706;
	wire [4-1:0] node707;
	wire [4-1:0] node709;
	wire [4-1:0] node711;
	wire [4-1:0] node712;
	wire [4-1:0] node714;
	wire [4-1:0] node716;
	wire [4-1:0] node720;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node726;
	wire [4-1:0] node728;
	wire [4-1:0] node730;
	wire [4-1:0] node737;
	wire [4-1:0] node738;
	wire [4-1:0] node739;
	wire [4-1:0] node741;
	wire [4-1:0] node743;
	wire [4-1:0] node745;
	wire [4-1:0] node747;
	wire [4-1:0] node749;
	wire [4-1:0] node752;
	wire [4-1:0] node753;
	wire [4-1:0] node754;
	wire [4-1:0] node756;
	wire [4-1:0] node758;
	wire [4-1:0] node760;
	wire [4-1:0] node762;
	wire [4-1:0] node764;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node772;
	wire [4-1:0] node774;
	wire [4-1:0] node776;
	wire [4-1:0] node777;
	wire [4-1:0] node779;
	wire [4-1:0] node781;
	wire [4-1:0] node786;
	wire [4-1:0] node788;
	wire [4-1:0] node790;
	wire [4-1:0] node793;
	wire [4-1:0] node795;
	wire [4-1:0] node796;
	wire [4-1:0] node798;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node802;
	wire [4-1:0] node804;
	wire [4-1:0] node810;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node813;
	wire [4-1:0] node814;
	wire [4-1:0] node816;
	wire [4-1:0] node818;
	wire [4-1:0] node820;
	wire [4-1:0] node821;
	wire [4-1:0] node823;
	wire [4-1:0] node825;
	wire [4-1:0] node827;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node833;
	wire [4-1:0] node835;
	wire [4-1:0] node839;
	wire [4-1:0] node840;
	wire [4-1:0] node841;
	wire [4-1:0] node843;
	wire [4-1:0] node844;
	wire [4-1:0] node846;
	wire [4-1:0] node848;
	wire [4-1:0] node850;
	wire [4-1:0] node854;
	wire [4-1:0] node855;
	wire [4-1:0] node856;
	wire [4-1:0] node857;
	wire [4-1:0] node859;
	wire [4-1:0] node861;
	wire [4-1:0] node867;
	wire [4-1:0] node869;
	wire [4-1:0] node871;
	wire [4-1:0] node874;
	wire [4-1:0] node875;
	wire [4-1:0] node877;
	wire [4-1:0] node879;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node884;
	wire [4-1:0] node888;
	wire [4-1:0] node889;
	wire [4-1:0] node890;
	wire [4-1:0] node891;
	wire [4-1:0] node893;
	wire [4-1:0] node895;
	wire [4-1:0] node900;
	wire [4-1:0] node902;
	wire [4-1:0] node903;
	wire [4-1:0] node905;
	wire [4-1:0] node906;
	wire [4-1:0] node908;
	wire [4-1:0] node910;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node917;
	wire [4-1:0] node918;
	wire [4-1:0] node920;
	wire [4-1:0] node922;
	wire [4-1:0] node923;
	wire [4-1:0] node924;
	wire [4-1:0] node926;
	wire [4-1:0] node928;
	wire [4-1:0] node933;
	wire [4-1:0] node934;
	wire [4-1:0] node936;
	wire [4-1:0] node938;
	wire [4-1:0] node940;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node946;
	wire [4-1:0] node948;
	wire [4-1:0] node951;
	wire [4-1:0] node952;
	wire [4-1:0] node956;
	wire [4-1:0] node957;
	wire [4-1:0] node958;
	wire [4-1:0] node960;
	wire [4-1:0] node962;
	wire [4-1:0] node964;
	wire [4-1:0] node966;
	wire [4-1:0] node969;
	wire [4-1:0] node971;
	wire [4-1:0] node973;
	wire [4-1:0] node976;
	wire [4-1:0] node978;
	wire [4-1:0] node981;
	wire [4-1:0] node982;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node989;
	wire [4-1:0] node991;
	wire [4-1:0] node993;
	wire [4-1:0] node998;
	wire [4-1:0] node1001;
	wire [4-1:0] node1002;
	wire [4-1:0] node1003;
	wire [4-1:0] node1006;
	wire [4-1:0] node1008;
	wire [4-1:0] node1010;
	wire [4-1:0] node1011;
	wire [4-1:0] node1013;
	wire [4-1:0] node1015;
	wire [4-1:0] node1019;
	wire [4-1:0] node1020;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1025;
	wire [4-1:0] node1028;
	wire [4-1:0] node1031;
	wire [4-1:0] node1032;
	wire [4-1:0] node1035;
	wire [4-1:0] node1038;
	wire [4-1:0] node1039;
	wire [4-1:0] node1040;
	wire [4-1:0] node1041;
	wire [4-1:0] node1044;
	wire [4-1:0] node1047;
	wire [4-1:0] node1048;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1056;
	wire [4-1:0] node1059;
	wire [4-1:0] node1060;
	wire [4-1:0] node1063;
	wire [4-1:0] node1066;
	wire [4-1:0] node1067;
	wire [4-1:0] node1068;
	wire [4-1:0] node1069;
	wire [4-1:0] node1072;
	wire [4-1:0] node1075;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1078;
	wire [4-1:0] node1081;
	wire [4-1:0] node1084;
	wire [4-1:0] node1085;
	wire [4-1:0] node1088;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1093;
	wire [4-1:0] node1097;
	wire [4-1:0] node1098;
	wire [4-1:0] node1101;
	wire [4-1:0] node1104;
	wire [4-1:0] node1105;
	wire [4-1:0] node1106;
	wire [4-1:0] node1108;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1115;
	wire [4-1:0] node1118;
	wire [4-1:0] node1119;
	wire [4-1:0] node1122;
	wire [4-1:0] node1125;
	wire [4-1:0] node1126;
	wire [4-1:0] node1129;
	wire [4-1:0] node1130;
	wire [4-1:0] node1132;
	wire [4-1:0] node1136;
	wire [4-1:0] node1137;
	wire [4-1:0] node1138;
	wire [4-1:0] node1139;
	wire [4-1:0] node1140;
	wire [4-1:0] node1141;
	wire [4-1:0] node1142;
	wire [4-1:0] node1144;
	wire [4-1:0] node1146;
	wire [4-1:0] node1148;
	wire [4-1:0] node1150;
	wire [4-1:0] node1153;
	wire [4-1:0] node1154;
	wire [4-1:0] node1155;
	wire [4-1:0] node1157;
	wire [4-1:0] node1159;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1168;
	wire [4-1:0] node1170;
	wire [4-1:0] node1172;
	wire [4-1:0] node1175;
	wire [4-1:0] node1176;
	wire [4-1:0] node1180;
	wire [4-1:0] node1181;
	wire [4-1:0] node1183;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1186;
	wire [4-1:0] node1188;
	wire [4-1:0] node1194;
	wire [4-1:0] node1195;
	wire [4-1:0] node1197;
	wire [4-1:0] node1198;
	wire [4-1:0] node1199;
	wire [4-1:0] node1201;
	wire [4-1:0] node1203;
	wire [4-1:0] node1205;
	wire [4-1:0] node1210;
	wire [4-1:0] node1212;
	wire [4-1:0] node1215;
	wire [4-1:0] node1216;
	wire [4-1:0] node1217;
	wire [4-1:0] node1218;
	wire [4-1:0] node1219;
	wire [4-1:0] node1221;
	wire [4-1:0] node1223;
	wire [4-1:0] node1228;
	wire [4-1:0] node1230;
	wire [4-1:0] node1232;
	wire [4-1:0] node1233;
	wire [4-1:0] node1234;
	wire [4-1:0] node1236;
	wire [4-1:0] node1238;
	wire [4-1:0] node1242;
	wire [4-1:0] node1244;
	wire [4-1:0] node1246;
	wire [4-1:0] node1248;
	wire [4-1:0] node1251;
	wire [4-1:0] node1252;
	wire [4-1:0] node1253;
	wire [4-1:0] node1255;
	wire [4-1:0] node1256;
	wire [4-1:0] node1258;
	wire [4-1:0] node1260;
	wire [4-1:0] node1262;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1270;
	wire [4-1:0] node1272;
	wire [4-1:0] node1274;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1280;
	wire [4-1:0] node1281;
	wire [4-1:0] node1283;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1288;
	wire [4-1:0] node1290;
	wire [4-1:0] node1292;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1298;
	wire [4-1:0] node1300;
	wire [4-1:0] node1304;
	wire [4-1:0] node1306;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1311;
	wire [4-1:0] node1315;
	wire [4-1:0] node1316;
	wire [4-1:0] node1317;
	wire [4-1:0] node1318;
	wire [4-1:0] node1320;
	wire [4-1:0] node1321;
	wire [4-1:0] node1325;
	wire [4-1:0] node1326;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1331;
	wire [4-1:0] node1335;
	wire [4-1:0] node1336;
	wire [4-1:0] node1340;
	wire [4-1:0] node1342;
	wire [4-1:0] node1345;
	wire [4-1:0] node1346;
	wire [4-1:0] node1348;
	wire [4-1:0] node1349;
	wire [4-1:0] node1350;
	wire [4-1:0] node1352;
	wire [4-1:0] node1354;
	wire [4-1:0] node1358;
	wire [4-1:0] node1360;
	wire [4-1:0] node1362;
	wire [4-1:0] node1364;
	wire [4-1:0] node1367;
	wire [4-1:0] node1369;
	wire [4-1:0] node1371;
	wire [4-1:0] node1373;
	wire [4-1:0] node1376;
	wire [4-1:0] node1377;
	wire [4-1:0] node1378;
	wire [4-1:0] node1379;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1384;
	wire [4-1:0] node1386;
	wire [4-1:0] node1388;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1395;
	wire [4-1:0] node1397;
	wire [4-1:0] node1399;
	wire [4-1:0] node1405;
	wire [4-1:0] node1406;
	wire [4-1:0] node1407;
	wire [4-1:0] node1409;
	wire [4-1:0] node1411;
	wire [4-1:0] node1415;
	wire [4-1:0] node1417;
	wire [4-1:0] node1418;
	wire [4-1:0] node1419;
	wire [4-1:0] node1421;
	wire [4-1:0] node1423;
	wire [4-1:0] node1425;
	wire [4-1:0] node1430;
	wire [4-1:0] node1431;
	wire [4-1:0] node1432;
	wire [4-1:0] node1434;
	wire [4-1:0] node1435;
	wire [4-1:0] node1437;
	wire [4-1:0] node1439;
	wire [4-1:0] node1441;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1447;
	wire [4-1:0] node1449;
	wire [4-1:0] node1453;
	wire [4-1:0] node1455;
	wire [4-1:0] node1456;
	wire [4-1:0] node1458;
	wire [4-1:0] node1462;
	wire [4-1:0] node1463;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1467;
	wire [4-1:0] node1469;
	wire [4-1:0] node1471;
	wire [4-1:0] node1474;
	wire [4-1:0] node1476;
	wire [4-1:0] node1478;
	wire [4-1:0] node1480;
	wire [4-1:0] node1483;
	wire [4-1:0] node1484;
	wire [4-1:0] node1486;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1492;
	wire [4-1:0] node1494;
	wire [4-1:0] node1496;
	wire [4-1:0] node1498;
	wire [4-1:0] node1501;
	wire [4-1:0] node1502;
	wire [4-1:0] node1504;
	wire [4-1:0] node1506;
	wire [4-1:0] node1510;
	wire [4-1:0] node1511;
	wire [4-1:0] node1513;
	wire [4-1:0] node1516;
	wire [4-1:0] node1517;
	wire [4-1:0] node1520;
	wire [4-1:0] node1522;

	assign outp = (inp[10]) ? node536 : node1;
		assign node1 = (inp[5]) ? node213 : node2;
			assign node2 = (inp[4]) ? node98 : node3;
				assign node3 = (inp[14]) ? node59 : node4;
					assign node4 = (inp[13]) ? node6 : 4'b1111;
						assign node6 = (inp[12]) ? node30 : node7;
							assign node7 = (inp[2]) ? node9 : 4'b1111;
								assign node9 = (inp[9]) ? node11 : 4'b1111;
									assign node11 = (inp[8]) ? node13 : 4'b1111;
										assign node13 = (inp[7]) ? node21 : node14;
											assign node14 = (inp[1]) ? node16 : 4'b1111;
												assign node16 = (inp[15]) ? node18 : 4'b1111;
													assign node18 = (inp[6]) ? 4'b1101 : 4'b1111;
											assign node21 = (inp[6]) ? 4'b1101 : node22;
												assign node22 = (inp[1]) ? node24 : 4'b1111;
													assign node24 = (inp[15]) ? node26 : 4'b1111;
														assign node26 = (inp[11]) ? 4'b1101 : 4'b1111;
							assign node30 = (inp[2]) ? 4'b1101 : node31;
								assign node31 = (inp[6]) ? node45 : node32;
									assign node32 = (inp[9]) ? node34 : 4'b1111;
										assign node34 = (inp[8]) ? 4'b1101 : node35;
											assign node35 = (inp[11]) ? node37 : 4'b1111;
												assign node37 = (inp[15]) ? node39 : 4'b1111;
													assign node39 = (inp[1]) ? node41 : 4'b1111;
														assign node41 = (inp[7]) ? 4'b1101 : 4'b1111;
									assign node45 = (inp[8]) ? 4'b1101 : node46;
										assign node46 = (inp[9]) ? 4'b1101 : node47;
											assign node47 = (inp[7]) ? 4'b1101 : node48;
												assign node48 = (inp[11]) ? node50 : 4'b1111;
													assign node50 = (inp[15]) ? node52 : 4'b1111;
														assign node52 = (inp[1]) ? 4'b1101 : 4'b1111;
					assign node59 = (inp[13]) ? node71 : node60;
						assign node60 = (inp[6]) ? node62 : 4'b1101;
							assign node62 = (inp[9]) ? node64 : 4'b1101;
								assign node64 = (inp[12]) ? node66 : 4'b1101;
									assign node66 = (inp[2]) ? node68 : 4'b1101;
										assign node68 = (inp[8]) ? 4'b1011 : 4'b1101;
						assign node71 = (inp[12]) ? node85 : node72;
							assign node72 = (inp[8]) ? node74 : 4'b1101;
								assign node74 = (inp[2]) ? node76 : 4'b1101;
									assign node76 = (inp[9]) ? node78 : 4'b1101;
										assign node78 = (inp[6]) ? 4'b1011 : node79;
											assign node79 = (inp[7]) ? node81 : 4'b1101;
												assign node81 = (inp[15]) ? 4'b1111 : 4'b1101;
							assign node85 = (inp[6]) ? 4'b1011 : node86;
								assign node86 = (inp[9]) ? 4'b1111 : node87;
									assign node87 = (inp[2]) ? 4'b1111 : node88;
										assign node88 = (inp[15]) ? node90 : 4'b1101;
											assign node90 = (inp[8]) ? node92 : 4'b1101;
												assign node92 = (inp[7]) ? 4'b1111 : 4'b1101;
				assign node98 = (inp[14]) ? node166 : node99;
					assign node99 = (inp[12]) ? node131 : node100;
						assign node100 = (inp[2]) ? node102 : 4'b1011;
							assign node102 = (inp[13]) ? node104 : 4'b1011;
								assign node104 = (inp[9]) ? node118 : node105;
									assign node105 = (inp[6]) ? node107 : 4'b1011;
										assign node107 = (inp[8]) ? 4'b1001 : node108;
											assign node108 = (inp[7]) ? node110 : 4'b1011;
												assign node110 = (inp[11]) ? node112 : 4'b1011;
													assign node112 = (inp[15]) ? node114 : 4'b1011;
														assign node114 = (inp[1]) ? 4'b1001 : 4'b1011;
									assign node118 = (inp[7]) ? 4'b1001 : node119;
										assign node119 = (inp[8]) ? 4'b1001 : node120;
											assign node120 = (inp[6]) ? 4'b1001 : node121;
												assign node121 = (inp[11]) ? node123 : 4'b1011;
													assign node123 = (inp[1]) ? node125 : 4'b1011;
														assign node125 = (inp[15]) ? 4'b1001 : 4'b1011;
						assign node131 = (inp[13]) ? 4'b1001 : node132;
							assign node132 = (inp[2]) ? node150 : node133;
								assign node133 = (inp[9]) ? node147 : node134;
									assign node134 = (inp[11]) ? node136 : 4'b1011;
										assign node136 = (inp[1]) ? node138 : 4'b1011;
											assign node138 = (inp[7]) ? node140 : 4'b1011;
												assign node140 = (inp[6]) ? node142 : 4'b1011;
													assign node142 = (inp[15]) ? node144 : 4'b1011;
														assign node144 = (inp[8]) ? 4'b1001 : 4'b1011;
									assign node147 = (inp[6]) ? 4'b1001 : 4'b1011;
								assign node150 = (inp[6]) ? 4'b1001 : node151;
									assign node151 = (inp[9]) ? 4'b1001 : node152;
										assign node152 = (inp[8]) ? node154 : 4'b1011;
											assign node154 = (inp[7]) ? 4'b1001 : node155;
												assign node155 = (inp[11]) ? node157 : 4'b1011;
													assign node157 = (inp[15]) ? node159 : 4'b1011;
														assign node159 = (inp[1]) ? 4'b1001 : 4'b1011;
					assign node166 = (inp[12]) ? node182 : node167;
						assign node167 = (inp[2]) ? node169 : 4'b1001;
							assign node169 = (inp[13]) ? node171 : 4'b1001;
								assign node171 = (inp[6]) ? 4'b1111 : node172;
									assign node172 = (inp[9]) ? 4'b1011 : node173;
										assign node173 = (inp[8]) ? node175 : 4'b1001;
											assign node175 = (inp[15]) ? node177 : 4'b1001;
												assign node177 = (inp[7]) ? 4'b1011 : 4'b1001;
						assign node182 = (inp[6]) ? node196 : node183;
							assign node183 = (inp[2]) ? 4'b1011 : node184;
								assign node184 = (inp[13]) ? 4'b1011 : node185;
									assign node185 = (inp[9]) ? node187 : 4'b1001;
										assign node187 = (inp[7]) ? node189 : 4'b1001;
											assign node189 = (inp[15]) ? node191 : 4'b1001;
												assign node191 = (inp[8]) ? 4'b1011 : 4'b1001;
							assign node196 = (inp[2]) ? node198 : 4'b1110;
								assign node198 = (inp[13]) ? node200 : 4'b1110;
									assign node200 = (inp[9]) ? 4'b1100 : node201;
										assign node201 = (inp[1]) ? node203 : 4'b1110;
											assign node203 = (inp[8]) ? node205 : 4'b1110;
												assign node205 = (inp[15]) ? node207 : 4'b1110;
													assign node207 = (inp[11]) ? node209 : 4'b1110;
														assign node209 = (inp[7]) ? 4'b1100 : 4'b1110;
			assign node213 = (inp[12]) ? node357 : node214;
				assign node214 = (inp[6]) ? node276 : node215;
					assign node215 = (inp[13]) ? node259 : node216;
						assign node216 = (inp[4]) ? node242 : node217;
							assign node217 = (inp[2]) ? node231 : node218;
								assign node218 = (inp[8]) ? 4'b1001 : node219;
									assign node219 = (inp[14]) ? node221 : 4'b1001;
										assign node221 = (inp[9]) ? 4'b1001 : node222;
											assign node222 = (inp[11]) ? node224 : 4'b1011;
												assign node224 = (inp[0]) ? node226 : 4'b1011;
													assign node226 = (inp[1]) ? 4'b1001 : 4'b1011;
								assign node231 = (inp[14]) ? 4'b1001 : node232;
									assign node232 = (inp[9]) ? 4'b1011 : node233;
										assign node233 = (inp[7]) ? node235 : 4'b1001;
											assign node235 = (inp[15]) ? node237 : 4'b1001;
												assign node237 = (inp[8]) ? 4'b1011 : 4'b1001;
							assign node242 = (inp[14]) ? node250 : node243;
								assign node243 = (inp[8]) ? node245 : 4'b1101;
									assign node245 = (inp[2]) ? node247 : 4'b1101;
										assign node247 = (inp[9]) ? 4'b1011 : 4'b1101;
								assign node250 = (inp[9]) ? 4'b1001 : node251;
									assign node251 = (inp[2]) ? 4'b1001 : node252;
										assign node252 = (inp[8]) ? node254 : 4'b1011;
											assign node254 = (inp[7]) ? 4'b1001 : 4'b1011;
						assign node259 = (inp[14]) ? node261 : 4'b1011;
							assign node261 = (inp[2]) ? node273 : node262;
								assign node262 = (inp[15]) ? node264 : 4'b1001;
									assign node264 = (inp[9]) ? node266 : 4'b1001;
										assign node266 = (inp[4]) ? node268 : 4'b1001;
											assign node268 = (inp[8]) ? node270 : 4'b1001;
												assign node270 = (inp[7]) ? 4'b1011 : 4'b1001;
								assign node273 = (inp[4]) ? 4'b1011 : 4'b1111;
					assign node276 = (inp[14]) ? node312 : node277;
						assign node277 = (inp[4]) ? node295 : node278;
							assign node278 = (inp[13]) ? 4'b1101 : node279;
								assign node279 = (inp[2]) ? node281 : 4'b1111;
									assign node281 = (inp[9]) ? node283 : 4'b1111;
										assign node283 = (inp[8]) ? 4'b1101 : node284;
											assign node284 = (inp[7]) ? node286 : 4'b1111;
												assign node286 = (inp[15]) ? node288 : 4'b1111;
													assign node288 = (inp[1]) ? node290 : 4'b1111;
														assign node290 = (inp[11]) ? 4'b1101 : 4'b1111;
							assign node295 = (inp[13]) ? 4'b1001 : node296;
								assign node296 = (inp[2]) ? node298 : 4'b1011;
									assign node298 = (inp[9]) ? 4'b1001 : node299;
										assign node299 = (inp[15]) ? node301 : 4'b1011;
											assign node301 = (inp[1]) ? node303 : 4'b1011;
												assign node303 = (inp[8]) ? node305 : 4'b1011;
													assign node305 = (inp[7]) ? node307 : 4'b1011;
														assign node307 = (inp[11]) ? 4'b1001 : 4'b1011;
						assign node312 = (inp[4]) ? node340 : node313;
							assign node313 = (inp[2]) ? node325 : node314;
								assign node314 = (inp[9]) ? 4'b1111 : node315;
									assign node315 = (inp[13]) ? 4'b1111 : node316;
										assign node316 = (inp[8]) ? node318 : 4'b1101;
											assign node318 = (inp[7]) ? node320 : 4'b1101;
												assign node320 = (inp[15]) ? 4'b1111 : 4'b1101;
								assign node325 = (inp[13]) ? node327 : 4'b1111;
									assign node327 = (inp[8]) ? 4'b1101 : node328;
										assign node328 = (inp[9]) ? 4'b1101 : node329;
											assign node329 = (inp[7]) ? 4'b1101 : node330;
												assign node330 = (inp[15]) ? node332 : 4'b1111;
													assign node332 = (inp[1]) ? node334 : 4'b1111;
														assign node334 = (inp[11]) ? 4'b1101 : 4'b1111;
							assign node340 = (inp[13]) ? node342 : 4'b1110;
								assign node342 = (inp[9]) ? 4'b1100 : node343;
									assign node343 = (inp[2]) ? 4'b1100 : node344;
										assign node344 = (inp[15]) ? node346 : 4'b1110;
											assign node346 = (inp[1]) ? node348 : 4'b1110;
												assign node348 = (inp[7]) ? node350 : 4'b1110;
													assign node350 = (inp[11]) ? node352 : 4'b1110;
														assign node352 = (inp[8]) ? 4'b1100 : 4'b1110;
				assign node357 = (inp[6]) ? node447 : node358;
					assign node358 = (inp[14]) ? node416 : node359;
						assign node359 = (inp[4]) ? node389 : node360;
							assign node360 = (inp[2]) ? node372 : node361;
								assign node361 = (inp[13]) ? 4'b1110 : node362;
									assign node362 = (inp[7]) ? node364 : 4'b1100;
										assign node364 = (inp[8]) ? node366 : 4'b1100;
											assign node366 = (inp[9]) ? node368 : 4'b1100;
												assign node368 = (inp[15]) ? 4'b1110 : 4'b1100;
								assign node372 = (inp[13]) ? node374 : 4'b1110;
									assign node374 = (inp[9]) ? 4'b1100 : node375;
										assign node375 = (inp[7]) ? node385 : node376;
											assign node376 = (inp[1]) ? node378 : 4'b1110;
												assign node378 = (inp[11]) ? node380 : 4'b1110;
													assign node380 = (inp[8]) ? node382 : 4'b1110;
														assign node382 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node385 = (inp[8]) ? 4'b1100 : 4'b1110;
							assign node389 = (inp[13]) ? node405 : node390;
								assign node390 = (inp[2]) ? node392 : 4'b1110;
									assign node392 = (inp[8]) ? 4'b1100 : node393;
										assign node393 = (inp[9]) ? 4'b1100 : node394;
											assign node394 = (inp[7]) ? node396 : 4'b1110;
												assign node396 = (inp[15]) ? node398 : 4'b1110;
													assign node398 = (inp[11]) ? node400 : 4'b1110;
														assign node400 = (inp[1]) ? 4'b1100 : 4'b1110;
								assign node405 = (inp[2]) ? node407 : 4'b1100;
									assign node407 = (inp[9]) ? 4'b1110 : node408;
										assign node408 = (inp[8]) ? node410 : 4'b1100;
											assign node410 = (inp[15]) ? node412 : 4'b1100;
												assign node412 = (inp[7]) ? 4'b1110 : 4'b1100;
						assign node416 = (inp[4]) ? node426 : node417;
							assign node417 = (inp[13]) ? 4'b1010 : node418;
								assign node418 = (inp[9]) ? node420 : 4'b1100;
									assign node420 = (inp[8]) ? node422 : 4'b1100;
										assign node422 = (inp[2]) ? 4'b1010 : 4'b1100;
							assign node426 = (inp[13]) ? node440 : node427;
								assign node427 = (inp[2]) ? node429 : 4'b1110;
									assign node429 = (inp[9]) ? node431 : 4'b1110;
										assign node431 = (inp[8]) ? 4'b1100 : node432;
											assign node432 = (inp[7]) ? 4'b1100 : node433;
												assign node433 = (inp[11]) ? node435 : 4'b1110;
													assign node435 = (inp[1]) ? 4'b1100 : 4'b1110;
								assign node440 = (inp[9]) ? node442 : 4'b1100;
									assign node442 = (inp[8]) ? node444 : 4'b1100;
										assign node444 = (inp[2]) ? 4'b1010 : 4'b1100;
					assign node447 = (inp[13]) ? node507 : node448;
						assign node448 = (inp[4]) ? node478 : node449;
							assign node449 = (inp[2]) ? 4'b1000 : node450;
								assign node450 = (inp[14]) ? node464 : node451;
									assign node451 = (inp[8]) ? 4'b1000 : node452;
										assign node452 = (inp[9]) ? 4'b1000 : node453;
											assign node453 = (inp[7]) ? 4'b1000 : node454;
												assign node454 = (inp[11]) ? node456 : 4'b1010;
													assign node456 = (inp[15]) ? node458 : 4'b1010;
														assign node458 = (inp[1]) ? 4'b1000 : 4'b1010;
									assign node464 = (inp[9]) ? node466 : 4'b1010;
										assign node466 = (inp[8]) ? 4'b1000 : node467;
											assign node467 = (inp[11]) ? node469 : 4'b1010;
												assign node469 = (inp[7]) ? node471 : 4'b1010;
													assign node471 = (inp[15]) ? node473 : 4'b1010;
														assign node473 = (inp[1]) ? 4'b1000 : 4'b1010;
							assign node478 = (inp[9]) ? node480 : 4'b1010;
								assign node480 = (inp[2]) ? node482 : 4'b1010;
									assign node482 = (inp[14]) ? node496 : node483;
										assign node483 = (inp[7]) ? node493 : node484;
											assign node484 = (inp[1]) ? node486 : 4'b1010;
												assign node486 = (inp[8]) ? node488 : 4'b1010;
													assign node488 = (inp[11]) ? node490 : 4'b1010;
														assign node490 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node493 = (inp[8]) ? 4'b1000 : 4'b1010;
										assign node496 = (inp[7]) ? node498 : 4'b1010;
											assign node498 = (inp[1]) ? node500 : 4'b1010;
												assign node500 = (inp[15]) ? node502 : 4'b1010;
													assign node502 = (inp[11]) ? node504 : 4'b1010;
														assign node504 = (inp[8]) ? 4'b1000 : 4'b1010;
						assign node507 = (inp[4]) ? node523 : node508;
							assign node508 = (inp[2]) ? node520 : node509;
								assign node509 = (inp[14]) ? 4'b1000 : node510;
									assign node510 = (inp[9]) ? 4'b1010 : node511;
										assign node511 = (inp[8]) ? node513 : 4'b1000;
											assign node513 = (inp[7]) ? node515 : 4'b1000;
												assign node515 = (inp[15]) ? 4'b1010 : 4'b1000;
								assign node520 = (inp[14]) ? 4'b1110 : 4'b1010;
							assign node523 = (inp[8]) ? node525 : 4'b1000;
								assign node525 = (inp[2]) ? node527 : 4'b1000;
									assign node527 = (inp[7]) ? node529 : 4'b1000;
										assign node529 = (inp[14]) ? 4'b1000 : node530;
											assign node530 = (inp[9]) ? node532 : 4'b1000;
												assign node532 = (inp[15]) ? 4'b1010 : 4'b1000;
		assign node536 = (inp[5]) ? node810 : node537;
			assign node537 = (inp[4]) ? node663 : node538;
				assign node538 = (inp[6]) ? node610 : node539;
					assign node539 = (inp[14]) ? node575 : node540;
						assign node540 = (inp[13]) ? node556 : node541;
							assign node541 = (inp[12]) ? node543 : 4'b1100;
								assign node543 = (inp[2]) ? 4'b1100 : node544;
									assign node544 = (inp[9]) ? node546 : 4'b1110;
										assign node546 = (inp[8]) ? 4'b1100 : node547;
											assign node547 = (inp[7]) ? 4'b1100 : node548;
												assign node548 = (inp[11]) ? node550 : 4'b1110;
													assign node550 = (inp[1]) ? 4'b1100 : 4'b1110;
							assign node556 = (inp[2]) ? node568 : node557;
								assign node557 = (inp[9]) ? node559 : 4'b1100;
									assign node559 = (inp[7]) ? node561 : 4'b1100;
										assign node561 = (inp[12]) ? 4'b1100 : node562;
											assign node562 = (inp[15]) ? node564 : 4'b1100;
												assign node564 = (inp[8]) ? 4'b1110 : 4'b1100;
								assign node568 = (inp[12]) ? node570 : 4'b1110;
									assign node570 = (inp[8]) ? node572 : 4'b1100;
										assign node572 = (inp[9]) ? 4'b1010 : 4'b1100;
						assign node575 = (inp[12]) ? node593 : node576;
							assign node576 = (inp[13]) ? node578 : 4'b1110;
								assign node578 = (inp[2]) ? 4'b1100 : node579;
									assign node579 = (inp[9]) ? 4'b1100 : node580;
										assign node580 = (inp[8]) ? node582 : 4'b1110;
											assign node582 = (inp[7]) ? 4'b1100 : node583;
												assign node583 = (inp[11]) ? node585 : 4'b1110;
													assign node585 = (inp[1]) ? node587 : 4'b1110;
														assign node587 = (inp[15]) ? 4'b1100 : 4'b1110;
							assign node593 = (inp[13]) ? node595 : 4'b1010;
								assign node595 = (inp[2]) ? 4'b1000 : node596;
									assign node596 = (inp[8]) ? node598 : 4'b1010;
										assign node598 = (inp[9]) ? node600 : 4'b1010;
											assign node600 = (inp[7]) ? 4'b1000 : node601;
												assign node601 = (inp[11]) ? node603 : 4'b1010;
													assign node603 = (inp[1]) ? node605 : 4'b1010;
														assign node605 = (inp[15]) ? 4'b1000 : 4'b1010;
					assign node610 = (inp[14]) ? node632 : node611;
						assign node611 = (inp[13]) ? 4'b1010 : node612;
							assign node612 = (inp[12]) ? node620 : node613;
								assign node613 = (inp[9]) ? node615 : 4'b1100;
									assign node615 = (inp[2]) ? node617 : 4'b1100;
										assign node617 = (inp[8]) ? 4'b1010 : 4'b1100;
								assign node620 = (inp[15]) ? node622 : 4'b1000;
									assign node622 = (inp[9]) ? node624 : 4'b1000;
										assign node624 = (inp[8]) ? node626 : 4'b1000;
											assign node626 = (inp[2]) ? node628 : 4'b1000;
												assign node628 = (inp[7]) ? 4'b1010 : 4'b1000;
						assign node632 = (inp[13]) ? 4'b1000 : node633;
							assign node633 = (inp[2]) ? node649 : node634;
								assign node634 = (inp[12]) ? node636 : 4'b1010;
									assign node636 = (inp[15]) ? node638 : 4'b1010;
										assign node638 = (inp[1]) ? node640 : 4'b1010;
											assign node640 = (inp[11]) ? node642 : 4'b1010;
												assign node642 = (inp[9]) ? node644 : 4'b1010;
													assign node644 = (inp[7]) ? node646 : 4'b1010;
														assign node646 = (inp[8]) ? 4'b1000 : 4'b1010;
								assign node649 = (inp[7]) ? 4'b1000 : node650;
									assign node650 = (inp[12]) ? 4'b1000 : node651;
										assign node651 = (inp[8]) ? 4'b1000 : node652;
											assign node652 = (inp[9]) ? 4'b1000 : node653;
												assign node653 = (inp[11]) ? node655 : 4'b1010;
													assign node655 = (inp[1]) ? 4'b1000 : 4'b1010;
				assign node663 = (inp[12]) ? node737 : node664;
					assign node664 = (inp[6]) ? node706 : node665;
						assign node665 = (inp[14]) ? node701 : node666;
							assign node666 = (inp[8]) ? node686 : node667;
								assign node667 = (inp[9]) ? node673 : node668;
									assign node668 = (inp[2]) ? 4'b1010 : node669;
										assign node669 = (inp[13]) ? 4'b1010 : 4'b1000;
									assign node673 = (inp[11]) ? node675 : 4'b1010;
										assign node675 = (inp[15]) ? node677 : 4'b1010;
											assign node677 = (inp[13]) ? node679 : 4'b1010;
												assign node679 = (inp[1]) ? node681 : 4'b1010;
													assign node681 = (inp[7]) ? node683 : 4'b1010;
														assign node683 = (inp[2]) ? 4'b1000 : 4'b1010;
								assign node686 = (inp[9]) ? node696 : node687;
									assign node687 = (inp[13]) ? 4'b1010 : node688;
										assign node688 = (inp[2]) ? 4'b1010 : node689;
											assign node689 = (inp[7]) ? node691 : 4'b1000;
												assign node691 = (inp[15]) ? 4'b1010 : 4'b1000;
									assign node696 = (inp[13]) ? node698 : 4'b1010;
										assign node698 = (inp[2]) ? 4'b1000 : 4'b1010;
							assign node701 = (inp[2]) ? node703 : 4'b1000;
								assign node703 = (inp[13]) ? 4'b1110 : 4'b1000;
						assign node706 = (inp[13]) ? node720 : node707;
							assign node707 = (inp[14]) ? node709 : 4'b1110;
								assign node709 = (inp[2]) ? node711 : 4'b1100;
									assign node711 = (inp[9]) ? 4'b1110 : node712;
										assign node712 = (inp[8]) ? node714 : 4'b1100;
											assign node714 = (inp[15]) ? node716 : 4'b1100;
												assign node716 = (inp[7]) ? 4'b1110 : 4'b1100;
							assign node720 = (inp[14]) ? 4'b1110 : node721;
								assign node721 = (inp[2]) ? 4'b1100 : node722;
									assign node722 = (inp[8]) ? 4'b1100 : node723;
										assign node723 = (inp[9]) ? 4'b1100 : node724;
											assign node724 = (inp[1]) ? node726 : 4'b1110;
												assign node726 = (inp[11]) ? node728 : 4'b1110;
													assign node728 = (inp[7]) ? node730 : 4'b1110;
														assign node730 = (inp[15]) ? 4'b1100 : 4'b1110;
					assign node737 = (inp[6]) ? node769 : node738;
						assign node738 = (inp[13]) ? node752 : node739;
							assign node739 = (inp[14]) ? node741 : 4'b1111;
								assign node741 = (inp[8]) ? node743 : 4'b1101;
									assign node743 = (inp[15]) ? node745 : 4'b1101;
										assign node745 = (inp[2]) ? node747 : 4'b1101;
											assign node747 = (inp[9]) ? node749 : 4'b1101;
												assign node749 = (inp[7]) ? 4'b1111 : 4'b1101;
							assign node752 = (inp[14]) ? 4'b1111 : node753;
								assign node753 = (inp[2]) ? 4'b1101 : node754;
									assign node754 = (inp[1]) ? node756 : 4'b1111;
										assign node756 = (inp[11]) ? node758 : 4'b1111;
											assign node758 = (inp[15]) ? node760 : 4'b1111;
												assign node760 = (inp[9]) ? node762 : 4'b1111;
													assign node762 = (inp[8]) ? node764 : 4'b1111;
														assign node764 = (inp[7]) ? 4'b1101 : 4'b1111;
						assign node769 = (inp[14]) ? node793 : node770;
							assign node770 = (inp[13]) ? node786 : node771;
								assign node771 = (inp[2]) ? 4'b1101 : node772;
									assign node772 = (inp[8]) ? node774 : 4'b1111;
										assign node774 = (inp[9]) ? node776 : 4'b1111;
											assign node776 = (inp[7]) ? 4'b1101 : node777;
												assign node777 = (inp[1]) ? node779 : 4'b1111;
													assign node779 = (inp[15]) ? node781 : 4'b1111;
														assign node781 = (inp[11]) ? 4'b1101 : 4'b1111;
								assign node786 = (inp[9]) ? node788 : 4'b1101;
									assign node788 = (inp[8]) ? node790 : 4'b1101;
										assign node790 = (inp[2]) ? 4'b1011 : 4'b1101;
							assign node793 = (inp[13]) ? node795 : 4'b1011;
								assign node795 = (inp[2]) ? 4'b1001 : node796;
									assign node796 = (inp[9]) ? node798 : 4'b1011;
										assign node798 = (inp[8]) ? 4'b1001 : node799;
											assign node799 = (inp[7]) ? 4'b1001 : node800;
												assign node800 = (inp[15]) ? node802 : 4'b1011;
													assign node802 = (inp[1]) ? node804 : 4'b1011;
														assign node804 = (inp[11]) ? 4'b1001 : 4'b1011;
			assign node810 = (inp[12]) ? node1136 : node811;
				assign node811 = (inp[6]) ? node915 : node812;
					assign node812 = (inp[13]) ? node874 : node813;
						assign node813 = (inp[4]) ? node839 : node814;
							assign node814 = (inp[8]) ? node816 : 4'b0111;
								assign node816 = (inp[9]) ? node818 : 4'b0111;
									assign node818 = (inp[2]) ? node820 : 4'b0111;
										assign node820 = (inp[14]) ? node830 : node821;
											assign node821 = (inp[11]) ? node823 : 4'b0111;
												assign node823 = (inp[15]) ? node825 : 4'b0111;
													assign node825 = (inp[1]) ? node827 : 4'b0111;
														assign node827 = (inp[7]) ? 4'b0101 : 4'b0111;
											assign node830 = (inp[7]) ? 4'b0101 : node831;
												assign node831 = (inp[11]) ? node833 : 4'b0111;
													assign node833 = (inp[15]) ? node835 : 4'b0111;
														assign node835 = (inp[1]) ? 4'b0101 : 4'b0111;
							assign node839 = (inp[2]) ? node867 : node840;
								assign node840 = (inp[14]) ? node854 : node841;
									assign node841 = (inp[9]) ? node843 : 4'b0111;
										assign node843 = (inp[8]) ? 4'b0101 : node844;
											assign node844 = (inp[11]) ? node846 : 4'b0111;
												assign node846 = (inp[15]) ? node848 : 4'b0111;
													assign node848 = (inp[7]) ? node850 : 4'b0111;
														assign node850 = (inp[1]) ? 4'b0101 : 4'b0111;
									assign node854 = (inp[8]) ? 4'b0101 : node855;
										assign node855 = (inp[7]) ? 4'b0101 : node856;
											assign node856 = (inp[9]) ? 4'b0101 : node857;
												assign node857 = (inp[1]) ? node859 : 4'b0111;
													assign node859 = (inp[15]) ? node861 : 4'b0111;
														assign node861 = (inp[11]) ? 4'b0101 : 4'b0111;
								assign node867 = (inp[14]) ? node869 : 4'b0101;
									assign node869 = (inp[8]) ? node871 : 4'b0101;
										assign node871 = (inp[9]) ? 4'b0011 : 4'b0101;
						assign node874 = (inp[4]) ? node888 : node875;
							assign node875 = (inp[9]) ? node877 : 4'b0101;
								assign node877 = (inp[2]) ? node879 : 4'b0101;
									assign node879 = (inp[8]) ? node881 : 4'b0101;
										assign node881 = (inp[14]) ? 4'b0011 : node882;
											assign node882 = (inp[15]) ? node884 : 4'b0101;
												assign node884 = (inp[7]) ? 4'b0111 : 4'b0101;
							assign node888 = (inp[14]) ? node900 : node889;
								assign node889 = (inp[2]) ? 4'b0111 : node890;
									assign node890 = (inp[9]) ? 4'b0111 : node891;
										assign node891 = (inp[15]) ? node893 : 4'b0101;
											assign node893 = (inp[8]) ? node895 : 4'b0101;
												assign node895 = (inp[7]) ? 4'b0111 : 4'b0101;
								assign node900 = (inp[2]) ? node902 : 4'b0011;
									assign node902 = (inp[9]) ? 4'b0001 : node903;
										assign node903 = (inp[8]) ? node905 : 4'b0011;
											assign node905 = (inp[7]) ? 4'b0001 : node906;
												assign node906 = (inp[11]) ? node908 : 4'b0011;
													assign node908 = (inp[1]) ? node910 : 4'b0011;
														assign node910 = (inp[15]) ? 4'b0001 : 4'b0011;
					assign node915 = (inp[14]) ? node981 : node916;
						assign node916 = (inp[13]) ? node944 : node917;
							assign node917 = (inp[4]) ? node933 : node918;
								assign node918 = (inp[2]) ? node920 : 4'b0011;
									assign node920 = (inp[9]) ? node922 : 4'b0011;
										assign node922 = (inp[8]) ? 4'b0001 : node923;
											assign node923 = (inp[7]) ? 4'b0001 : node924;
												assign node924 = (inp[1]) ? node926 : 4'b0011;
													assign node926 = (inp[11]) ? node928 : 4'b0011;
														assign node928 = (inp[15]) ? 4'b0001 : 4'b0011;
								assign node933 = (inp[2]) ? 4'b0011 : node934;
									assign node934 = (inp[8]) ? node936 : 4'b0001;
										assign node936 = (inp[7]) ? node938 : 4'b0001;
											assign node938 = (inp[9]) ? node940 : 4'b0001;
												assign node940 = (inp[15]) ? 4'b0011 : 4'b0001;
							assign node944 = (inp[7]) ? node956 : node945;
								assign node945 = (inp[4]) ? node951 : node946;
									assign node946 = (inp[9]) ? node948 : 4'b0001;
										assign node948 = (inp[2]) ? 4'b0011 : 4'b0001;
									assign node951 = (inp[2]) ? 4'b0001 : node952;
										assign node952 = (inp[9]) ? 4'b0001 : 4'b0011;
								assign node956 = (inp[9]) ? node976 : node957;
									assign node957 = (inp[2]) ? node969 : node958;
										assign node958 = (inp[4]) ? node960 : 4'b0001;
											assign node960 = (inp[1]) ? node962 : 4'b0011;
												assign node962 = (inp[15]) ? node964 : 4'b0011;
													assign node964 = (inp[8]) ? node966 : 4'b0011;
														assign node966 = (inp[11]) ? 4'b0001 : 4'b0011;
										assign node969 = (inp[8]) ? node971 : 4'b0001;
											assign node971 = (inp[15]) ? node973 : 4'b0001;
												assign node973 = (inp[4]) ? 4'b0001 : 4'b0011;
									assign node976 = (inp[2]) ? node978 : 4'b0001;
										assign node978 = (inp[4]) ? 4'b0001 : 4'b0011;
						assign node981 = (inp[4]) ? node1001 : node982;
							assign node982 = (inp[13]) ? node998 : node983;
								assign node983 = (inp[2]) ? node985 : 4'b0011;
									assign node985 = (inp[8]) ? 4'b0001 : node986;
										assign node986 = (inp[9]) ? 4'b0001 : node987;
											assign node987 = (inp[1]) ? node989 : 4'b0011;
												assign node989 = (inp[15]) ? node991 : 4'b0011;
													assign node991 = (inp[11]) ? node993 : 4'b0011;
														assign node993 = (inp[7]) ? 4'b0001 : 4'b0011;
								assign node998 = (inp[2]) ? 4'b0111 : 4'b0001;
							assign node1001 = (inp[9]) ? node1019 : node1002;
								assign node1002 = (inp[2]) ? node1006 : node1003;
									assign node1003 = (inp[13]) ? 4'b0100 : 4'b0110;
									assign node1006 = (inp[7]) ? node1008 : 4'b0110;
										assign node1008 = (inp[1]) ? node1010 : 4'b0110;
											assign node1010 = (inp[13]) ? 4'b0110 : node1011;
												assign node1011 = (inp[8]) ? node1013 : 4'b0110;
													assign node1013 = (inp[11]) ? node1015 : 4'b0110;
														assign node1015 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node1019 = (inp[8]) ? node1125 : node1020;
									assign node1020 = (inp[15]) ? node1066 : node1021;
										assign node1021 = (inp[11]) ? node1059 : node1022;
											assign node1022 = (inp[3]) ? node1038 : node1023;
												assign node1023 = (inp[1]) ? node1031 : node1024;
													assign node1024 = (inp[13]) ? node1028 : node1025;
														assign node1025 = (inp[2]) ? 4'b0100 : 4'b0110;
														assign node1028 = (inp[2]) ? 4'b0110 : 4'b0100;
													assign node1031 = (inp[13]) ? node1035 : node1032;
														assign node1032 = (inp[2]) ? 4'b0100 : 4'b0110;
														assign node1035 = (inp[2]) ? 4'b0110 : 4'b0100;
												assign node1038 = (inp[0]) ? node1052 : node1039;
													assign node1039 = (inp[1]) ? node1047 : node1040;
														assign node1040 = (inp[13]) ? node1044 : node1041;
															assign node1041 = (inp[2]) ? 4'b0100 : 4'b0110;
															assign node1044 = (inp[2]) ? 4'b0110 : 4'b0100;
														assign node1047 = (inp[13]) ? 4'b0100 : node1048;
															assign node1048 = (inp[2]) ? 4'b0100 : 4'b0110;
													assign node1052 = (inp[2]) ? node1056 : node1053;
														assign node1053 = (inp[13]) ? 4'b0100 : 4'b0110;
														assign node1056 = (inp[13]) ? 4'b0110 : 4'b0100;
											assign node1059 = (inp[13]) ? node1063 : node1060;
												assign node1060 = (inp[2]) ? 4'b0100 : 4'b0110;
												assign node1063 = (inp[2]) ? 4'b0110 : 4'b0100;
										assign node1066 = (inp[1]) ? node1104 : node1067;
											assign node1067 = (inp[3]) ? node1075 : node1068;
												assign node1068 = (inp[2]) ? node1072 : node1069;
													assign node1069 = (inp[13]) ? 4'b0100 : 4'b0110;
													assign node1072 = (inp[13]) ? 4'b0110 : 4'b0100;
												assign node1075 = (inp[7]) ? node1091 : node1076;
													assign node1076 = (inp[11]) ? node1084 : node1077;
														assign node1077 = (inp[2]) ? node1081 : node1078;
															assign node1078 = (inp[13]) ? 4'b0100 : 4'b0110;
															assign node1081 = (inp[13]) ? 4'b0110 : 4'b0100;
														assign node1084 = (inp[13]) ? node1088 : node1085;
															assign node1085 = (inp[2]) ? 4'b0100 : 4'b0110;
															assign node1088 = (inp[2]) ? 4'b0110 : 4'b0100;
													assign node1091 = (inp[11]) ? node1097 : node1092;
														assign node1092 = (inp[0]) ? 4'b0110 : node1093;
															assign node1093 = (inp[13]) ? 4'b0100 : 4'b0110;
														assign node1097 = (inp[13]) ? node1101 : node1098;
															assign node1098 = (inp[2]) ? 4'b0100 : 4'b0110;
															assign node1101 = (inp[2]) ? 4'b0110 : 4'b0100;
											assign node1104 = (inp[7]) ? node1118 : node1105;
												assign node1105 = (inp[0]) ? node1111 : node1106;
													assign node1106 = (inp[13]) ? node1108 : 4'b0110;
														assign node1108 = (inp[2]) ? 4'b0110 : 4'b0100;
													assign node1111 = (inp[2]) ? node1115 : node1112;
														assign node1112 = (inp[13]) ? 4'b0100 : 4'b0110;
														assign node1115 = (inp[13]) ? 4'b0110 : 4'b0100;
												assign node1118 = (inp[2]) ? node1122 : node1119;
													assign node1119 = (inp[13]) ? 4'b0100 : 4'b0110;
													assign node1122 = (inp[13]) ? 4'b0110 : 4'b0100;
									assign node1125 = (inp[13]) ? node1129 : node1126;
										assign node1126 = (inp[2]) ? 4'b0100 : 4'b0110;
										assign node1129 = (inp[2]) ? 4'b0110 : node1130;
											assign node1130 = (inp[15]) ? node1132 : 4'b0100;
												assign node1132 = (inp[7]) ? 4'b0110 : 4'b0100;
				assign node1136 = (inp[4]) ? node1278 : node1137;
					assign node1137 = (inp[14]) ? node1215 : node1138;
						assign node1138 = (inp[13]) ? node1180 : node1139;
							assign node1139 = (inp[2]) ? node1165 : node1140;
								assign node1140 = (inp[9]) ? 4'b0100 : node1141;
									assign node1141 = (inp[8]) ? node1153 : node1142;
										assign node1142 = (inp[15]) ? node1144 : 4'b0110;
											assign node1144 = (inp[7]) ? node1146 : 4'b0110;
												assign node1146 = (inp[11]) ? node1148 : 4'b0110;
													assign node1148 = (inp[6]) ? node1150 : 4'b0110;
														assign node1150 = (inp[1]) ? 4'b0100 : 4'b0110;
										assign node1153 = (inp[6]) ? 4'b0100 : node1154;
											assign node1154 = (inp[7]) ? 4'b0100 : node1155;
												assign node1155 = (inp[1]) ? node1157 : 4'b0110;
													assign node1157 = (inp[11]) ? node1159 : 4'b0110;
														assign node1159 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node1165 = (inp[9]) ? node1175 : node1166;
									assign node1166 = (inp[7]) ? node1168 : 4'b0100;
										assign node1168 = (inp[8]) ? node1170 : 4'b0100;
											assign node1170 = (inp[6]) ? node1172 : 4'b0100;
												assign node1172 = (inp[15]) ? 4'b0110 : 4'b0100;
									assign node1175 = (inp[6]) ? 4'b0110 : node1176;
										assign node1176 = (inp[8]) ? 4'b0010 : 4'b0100;
							assign node1180 = (inp[6]) ? node1194 : node1181;
								assign node1181 = (inp[2]) ? node1183 : 4'b0010;
									assign node1183 = (inp[9]) ? 4'b0000 : node1184;
										assign node1184 = (inp[7]) ? 4'b0000 : node1185;
											assign node1185 = (inp[8]) ? 4'b0000 : node1186;
												assign node1186 = (inp[15]) ? node1188 : 4'b0010;
													assign node1188 = (inp[11]) ? 4'b0000 : 4'b0010;
								assign node1194 = (inp[2]) ? node1210 : node1195;
									assign node1195 = (inp[9]) ? node1197 : 4'b0110;
										assign node1197 = (inp[7]) ? 4'b0100 : node1198;
											assign node1198 = (inp[8]) ? 4'b0100 : node1199;
												assign node1199 = (inp[0]) ? node1201 : 4'b0110;
													assign node1201 = (inp[11]) ? node1203 : 4'b0110;
														assign node1203 = (inp[1]) ? node1205 : 4'b0110;
															assign node1205 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node1210 = (inp[8]) ? node1212 : 4'b0100;
										assign node1212 = (inp[9]) ? 4'b0010 : 4'b0100;
						assign node1215 = (inp[2]) ? node1251 : node1216;
							assign node1216 = (inp[6]) ? node1228 : node1217;
								assign node1217 = (inp[13]) ? 4'b0000 : node1218;
									assign node1218 = (inp[9]) ? 4'b0010 : node1219;
										assign node1219 = (inp[7]) ? node1221 : 4'b0000;
											assign node1221 = (inp[8]) ? node1223 : 4'b0000;
												assign node1223 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node1228 = (inp[9]) ? node1230 : 4'b0010;
									assign node1230 = (inp[8]) ? node1232 : 4'b0010;
										assign node1232 = (inp[13]) ? node1242 : node1233;
											assign node1233 = (inp[7]) ? 4'b0000 : node1234;
												assign node1234 = (inp[15]) ? node1236 : 4'b0010;
													assign node1236 = (inp[1]) ? node1238 : 4'b0010;
														assign node1238 = (inp[11]) ? 4'b0000 : 4'b0010;
											assign node1242 = (inp[7]) ? node1244 : 4'b0010;
												assign node1244 = (inp[15]) ? node1246 : 4'b0010;
													assign node1246 = (inp[1]) ? node1248 : 4'b0010;
														assign node1248 = (inp[11]) ? 4'b0000 : 4'b0010;
							assign node1251 = (inp[6]) ? node1267 : node1252;
								assign node1252 = (inp[13]) ? 4'b0110 : node1253;
									assign node1253 = (inp[9]) ? node1255 : 4'b0010;
										assign node1255 = (inp[8]) ? 4'b0000 : node1256;
											assign node1256 = (inp[11]) ? node1258 : 4'b0010;
												assign node1258 = (inp[7]) ? node1260 : 4'b0010;
													assign node1260 = (inp[1]) ? node1262 : 4'b0010;
														assign node1262 = (inp[15]) ? 4'b0000 : 4'b0010;
								assign node1267 = (inp[13]) ? 4'b0000 : node1268;
									assign node1268 = (inp[15]) ? node1270 : 4'b0000;
										assign node1270 = (inp[8]) ? node1272 : 4'b0000;
											assign node1272 = (inp[7]) ? node1274 : 4'b0000;
												assign node1274 = (inp[9]) ? 4'b0010 : 4'b0000;
					assign node1278 = (inp[14]) ? node1376 : node1279;
						assign node1279 = (inp[6]) ? node1315 : node1280;
							assign node1280 = (inp[2]) ? node1304 : node1281;
								assign node1281 = (inp[9]) ? node1283 : 4'b0111;
									assign node1283 = (inp[8]) ? node1285 : 4'b0111;
										assign node1285 = (inp[13]) ? node1295 : node1286;
											assign node1286 = (inp[7]) ? node1288 : 4'b0111;
												assign node1288 = (inp[1]) ? node1290 : 4'b0111;
													assign node1290 = (inp[15]) ? node1292 : 4'b0111;
														assign node1292 = (inp[11]) ? 4'b0101 : 4'b0111;
											assign node1295 = (inp[7]) ? 4'b0101 : node1296;
												assign node1296 = (inp[1]) ? node1298 : 4'b0111;
													assign node1298 = (inp[15]) ? node1300 : 4'b0111;
														assign node1300 = (inp[11]) ? 4'b0101 : 4'b0111;
								assign node1304 = (inp[9]) ? node1306 : 4'b0101;
									assign node1306 = (inp[8]) ? node1308 : 4'b0101;
										assign node1308 = (inp[13]) ? 4'b0011 : node1309;
											assign node1309 = (inp[7]) ? node1311 : 4'b0101;
												assign node1311 = (inp[15]) ? 4'b0111 : 4'b0101;
							assign node1315 = (inp[13]) ? node1345 : node1316;
								assign node1316 = (inp[9]) ? node1340 : node1317;
									assign node1317 = (inp[15]) ? node1325 : node1318;
										assign node1318 = (inp[2]) ? node1320 : 4'b0101;
											assign node1320 = (inp[7]) ? 4'b0101 : node1321;
												assign node1321 = (inp[8]) ? 4'b0101 : 4'b0111;
										assign node1325 = (inp[7]) ? node1335 : node1326;
											assign node1326 = (inp[2]) ? node1328 : 4'b0101;
												assign node1328 = (inp[8]) ? 4'b0101 : node1329;
													assign node1329 = (inp[1]) ? node1331 : 4'b0111;
														assign node1331 = (inp[11]) ? 4'b0101 : 4'b0111;
											assign node1335 = (inp[2]) ? 4'b0101 : node1336;
												assign node1336 = (inp[8]) ? 4'b0111 : 4'b0101;
									assign node1340 = (inp[2]) ? node1342 : 4'b0111;
										assign node1342 = (inp[8]) ? 4'b0011 : 4'b0101;
								assign node1345 = (inp[9]) ? node1367 : node1346;
									assign node1346 = (inp[8]) ? node1348 : 4'b0011;
										assign node1348 = (inp[2]) ? node1358 : node1349;
											assign node1349 = (inp[7]) ? 4'b0001 : node1350;
												assign node1350 = (inp[11]) ? node1352 : 4'b0011;
													assign node1352 = (inp[1]) ? node1354 : 4'b0011;
														assign node1354 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node1358 = (inp[1]) ? node1360 : 4'b0011;
												assign node1360 = (inp[11]) ? node1362 : 4'b0011;
													assign node1362 = (inp[15]) ? node1364 : 4'b0011;
														assign node1364 = (inp[7]) ? 4'b0001 : 4'b0011;
									assign node1367 = (inp[15]) ? node1369 : 4'b0001;
										assign node1369 = (inp[7]) ? node1371 : 4'b0001;
											assign node1371 = (inp[8]) ? node1373 : 4'b0001;
												assign node1373 = (inp[2]) ? 4'b0001 : 4'b0011;
						assign node1376 = (inp[6]) ? node1430 : node1377;
							assign node1377 = (inp[2]) ? node1405 : node1378;
								assign node1378 = (inp[9]) ? node1392 : node1379;
									assign node1379 = (inp[13]) ? node1381 : 4'b0011;
										assign node1381 = (inp[8]) ? 4'b0001 : node1382;
											assign node1382 = (inp[7]) ? node1384 : 4'b0011;
												assign node1384 = (inp[15]) ? node1386 : 4'b0011;
													assign node1386 = (inp[11]) ? node1388 : 4'b0011;
														assign node1388 = (inp[1]) ? 4'b0001 : 4'b0011;
									assign node1392 = (inp[13]) ? 4'b0001 : node1393;
										assign node1393 = (inp[7]) ? 4'b0001 : node1394;
											assign node1394 = (inp[8]) ? 4'b0001 : node1395;
												assign node1395 = (inp[15]) ? node1397 : 4'b0011;
													assign node1397 = (inp[11]) ? node1399 : 4'b0011;
														assign node1399 = (inp[1]) ? 4'b0001 : 4'b0011;
								assign node1405 = (inp[13]) ? node1415 : node1406;
									assign node1406 = (inp[9]) ? 4'b0011 : node1407;
										assign node1407 = (inp[8]) ? node1409 : 4'b0001;
											assign node1409 = (inp[15]) ? node1411 : 4'b0001;
												assign node1411 = (inp[7]) ? 4'b0011 : 4'b0001;
									assign node1415 = (inp[9]) ? node1417 : 4'b0111;
										assign node1417 = (inp[8]) ? 4'b0101 : node1418;
											assign node1418 = (inp[3]) ? 4'b0111 : node1419;
												assign node1419 = (inp[15]) ? node1421 : 4'b0111;
													assign node1421 = (inp[11]) ? node1423 : 4'b0111;
														assign node1423 = (inp[1]) ? node1425 : 4'b0111;
															assign node1425 = (inp[7]) ? 4'b0101 : 4'b0111;
							assign node1430 = (inp[13]) ? node1462 : node1431;
								assign node1431 = (inp[9]) ? node1453 : node1432;
									assign node1432 = (inp[8]) ? node1434 : 4'b0110;
										assign node1434 = (inp[7]) ? node1444 : node1435;
											assign node1435 = (inp[15]) ? node1437 : 4'b0110;
												assign node1437 = (inp[1]) ? node1439 : 4'b0110;
													assign node1439 = (inp[11]) ? node1441 : 4'b0110;
														assign node1441 = (inp[2]) ? 4'b0100 : 4'b0110;
											assign node1444 = (inp[2]) ? 4'b0100 : node1445;
												assign node1445 = (inp[1]) ? node1447 : 4'b0110;
													assign node1447 = (inp[15]) ? node1449 : 4'b0110;
														assign node1449 = (inp[11]) ? 4'b0100 : 4'b0110;
									assign node1453 = (inp[8]) ? node1455 : 4'b0100;
										assign node1455 = (inp[2]) ? 4'b0010 : node1456;
											assign node1456 = (inp[7]) ? node1458 : 4'b0100;
												assign node1458 = (inp[15]) ? 4'b0110 : 4'b0100;
								assign node1462 = (inp[2]) ? node1490 : node1463;
									assign node1463 = (inp[8]) ? node1483 : node1464;
										assign node1464 = (inp[7]) ? node1474 : node1465;
											assign node1465 = (inp[15]) ? node1467 : 4'b0010;
												assign node1467 = (inp[1]) ? node1469 : 4'b0010;
													assign node1469 = (inp[11]) ? node1471 : 4'b0010;
														assign node1471 = (inp[9]) ? 4'b0010 : 4'b0000;
											assign node1474 = (inp[9]) ? node1476 : 4'b0000;
												assign node1476 = (inp[15]) ? node1478 : 4'b0010;
													assign node1478 = (inp[1]) ? node1480 : 4'b0010;
														assign node1480 = (inp[11]) ? 4'b0000 : 4'b0010;
										assign node1483 = (inp[9]) ? 4'b0000 : node1484;
											assign node1484 = (inp[15]) ? node1486 : 4'b0000;
												assign node1486 = (inp[7]) ? 4'b0010 : 4'b0000;
									assign node1490 = (inp[8]) ? node1510 : node1491;
										assign node1491 = (inp[9]) ? node1501 : node1492;
											assign node1492 = (inp[15]) ? node1494 : 4'b0110;
												assign node1494 = (inp[7]) ? node1496 : 4'b0110;
													assign node1496 = (inp[11]) ? node1498 : 4'b0110;
														assign node1498 = (inp[1]) ? 4'b0100 : 4'b0110;
											assign node1501 = (inp[7]) ? 4'b0100 : node1502;
												assign node1502 = (inp[15]) ? node1504 : 4'b0110;
													assign node1504 = (inp[1]) ? node1506 : 4'b0110;
														assign node1506 = (inp[11]) ? 4'b0100 : 4'b0110;
										assign node1510 = (inp[9]) ? node1516 : node1511;
											assign node1511 = (inp[15]) ? node1513 : 4'b0100;
												assign node1513 = (inp[7]) ? 4'b0110 : 4'b0100;
											assign node1516 = (inp[15]) ? node1520 : node1517;
												assign node1517 = (inp[7]) ? 4'b0000 : 4'b0010;
												assign node1520 = (inp[11]) ? node1522 : 4'b0010;
													assign node1522 = (inp[1]) ? 4'b0000 : 4'b0010;

endmodule