module dtc_split5_bm73 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node66;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node215;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node263;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node281;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node312;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node321;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node364;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node368;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node409;
	wire [3-1:0] node412;
	wire [3-1:0] node414;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node427;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node451;
	wire [3-1:0] node452;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node477;
	wire [3-1:0] node480;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node488;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node517;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node529;
	wire [3-1:0] node531;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node537;
	wire [3-1:0] node539;
	wire [3-1:0] node542;
	wire [3-1:0] node544;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node559;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node568;
	wire [3-1:0] node570;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node583;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node593;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node621;
	wire [3-1:0] node624;
	wire [3-1:0] node625;
	wire [3-1:0] node627;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node638;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node647;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node670;
	wire [3-1:0] node672;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node680;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node687;
	wire [3-1:0] node688;
	wire [3-1:0] node690;
	wire [3-1:0] node692;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node702;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node731;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node741;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node754;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node765;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node771;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node780;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node787;
	wire [3-1:0] node789;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node794;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node801;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node807;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node824;
	wire [3-1:0] node827;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node845;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node853;
	wire [3-1:0] node856;
	wire [3-1:0] node857;
	wire [3-1:0] node859;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node881;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node888;
	wire [3-1:0] node891;
	wire [3-1:0] node893;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node917;
	wire [3-1:0] node919;
	wire [3-1:0] node922;
	wire [3-1:0] node923;
	wire [3-1:0] node924;
	wire [3-1:0] node925;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node933;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node945;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node950;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node956;
	wire [3-1:0] node959;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node969;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node975;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node982;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node989;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node995;
	wire [3-1:0] node999;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1013;
	wire [3-1:0] node1016;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1027;
	wire [3-1:0] node1031;
	wire [3-1:0] node1032;
	wire [3-1:0] node1035;
	wire [3-1:0] node1037;
	wire [3-1:0] node1040;
	wire [3-1:0] node1041;
	wire [3-1:0] node1043;

	assign outp = (inp[9]) ? node298 : node1;
		assign node1 = (inp[6]) ? node219 : node2;
			assign node2 = (inp[3]) ? node156 : node3;
				assign node3 = (inp[10]) ? node95 : node4;
					assign node4 = (inp[7]) ? node36 : node5;
						assign node5 = (inp[4]) ? node21 : node6;
							assign node6 = (inp[11]) ? node14 : node7;
								assign node7 = (inp[8]) ? node11 : node8;
									assign node8 = (inp[5]) ? 3'b001 : 3'b101;
									assign node11 = (inp[5]) ? 3'b110 : 3'b001;
								assign node14 = (inp[5]) ? node18 : node15;
									assign node15 = (inp[8]) ? 3'b101 : 3'b011;
									assign node18 = (inp[8]) ? 3'b001 : 3'b101;
							assign node21 = (inp[5]) ? node29 : node22;
								assign node22 = (inp[8]) ? node26 : node23;
									assign node23 = (inp[11]) ? 3'b001 : 3'b110;
									assign node26 = (inp[11]) ? 3'b110 : 3'b010;
								assign node29 = (inp[8]) ? node33 : node30;
									assign node30 = (inp[11]) ? 3'b110 : 3'b010;
									assign node33 = (inp[11]) ? 3'b010 : 3'b100;
						assign node36 = (inp[4]) ? node74 : node37;
							assign node37 = (inp[1]) ? node53 : node38;
								assign node38 = (inp[5]) ? node46 : node39;
									assign node39 = (inp[11]) ? node43 : node40;
										assign node40 = (inp[8]) ? 3'b010 : 3'b110;
										assign node43 = (inp[8]) ? 3'b110 : 3'b001;
									assign node46 = (inp[8]) ? node50 : node47;
										assign node47 = (inp[11]) ? 3'b110 : 3'b010;
										assign node50 = (inp[11]) ? 3'b010 : 3'b100;
								assign node53 = (inp[8]) ? node63 : node54;
									assign node54 = (inp[0]) ? node56 : 3'b110;
										assign node56 = (inp[5]) ? node60 : node57;
											assign node57 = (inp[11]) ? 3'b001 : 3'b110;
											assign node60 = (inp[11]) ? 3'b110 : 3'b010;
									assign node63 = (inp[2]) ? node69 : node64;
										assign node64 = (inp[11]) ? node66 : 3'b010;
											assign node66 = (inp[5]) ? 3'b010 : 3'b110;
										assign node69 = (inp[5]) ? 3'b100 : node70;
											assign node70 = (inp[11]) ? 3'b110 : 3'b010;
							assign node74 = (inp[11]) ? node80 : node75;
								assign node75 = (inp[5]) ? 3'b000 : node76;
									assign node76 = (inp[8]) ? 3'b000 : 3'b100;
								assign node80 = (inp[2]) ? node88 : node81;
									assign node81 = (inp[8]) ? node85 : node82;
										assign node82 = (inp[5]) ? 3'b100 : 3'b010;
										assign node85 = (inp[5]) ? 3'b000 : 3'b100;
									assign node88 = (inp[0]) ? node90 : 3'b100;
										assign node90 = (inp[5]) ? 3'b100 : node91;
											assign node91 = (inp[8]) ? 3'b100 : 3'b010;
					assign node95 = (inp[7]) ? node125 : node96;
						assign node96 = (inp[4]) ? node110 : node97;
							assign node97 = (inp[11]) ? node105 : node98;
								assign node98 = (inp[8]) ? node102 : node99;
									assign node99 = (inp[5]) ? 3'b011 : 3'b111;
									assign node102 = (inp[5]) ? 3'b101 : 3'b011;
								assign node105 = (inp[8]) ? node107 : 3'b111;
									assign node107 = (inp[5]) ? 3'b011 : 3'b111;
							assign node110 = (inp[11]) ? node118 : node111;
								assign node111 = (inp[5]) ? node115 : node112;
									assign node112 = (inp[8]) ? 3'b001 : 3'b101;
									assign node115 = (inp[8]) ? 3'b110 : 3'b001;
								assign node118 = (inp[5]) ? node122 : node119;
									assign node119 = (inp[8]) ? 3'b101 : 3'b011;
									assign node122 = (inp[8]) ? 3'b001 : 3'b101;
						assign node125 = (inp[4]) ? node141 : node126;
							assign node126 = (inp[5]) ? node134 : node127;
								assign node127 = (inp[11]) ? node131 : node128;
									assign node128 = (inp[8]) ? 3'b001 : 3'b101;
									assign node131 = (inp[8]) ? 3'b101 : 3'b011;
								assign node134 = (inp[11]) ? node138 : node135;
									assign node135 = (inp[8]) ? 3'b110 : 3'b001;
									assign node138 = (inp[8]) ? 3'b001 : 3'b101;
							assign node141 = (inp[8]) ? node149 : node142;
								assign node142 = (inp[5]) ? node146 : node143;
									assign node143 = (inp[11]) ? 3'b001 : 3'b110;
									assign node146 = (inp[11]) ? 3'b110 : 3'b010;
								assign node149 = (inp[5]) ? node153 : node150;
									assign node150 = (inp[11]) ? 3'b110 : 3'b010;
									assign node153 = (inp[11]) ? 3'b010 : 3'b100;
				assign node156 = (inp[10]) ? node174 : node157;
					assign node157 = (inp[4]) ? 3'b000 : node158;
						assign node158 = (inp[7]) ? 3'b000 : node159;
							assign node159 = (inp[5]) ? node167 : node160;
								assign node160 = (inp[8]) ? node164 : node161;
									assign node161 = (inp[11]) ? 3'b010 : 3'b100;
									assign node164 = (inp[11]) ? 3'b100 : 3'b000;
								assign node167 = (inp[11]) ? node169 : 3'b000;
									assign node169 = (inp[8]) ? 3'b000 : 3'b100;
					assign node174 = (inp[7]) ? node204 : node175;
						assign node175 = (inp[4]) ? node191 : node176;
							assign node176 = (inp[11]) ? node184 : node177;
								assign node177 = (inp[5]) ? node181 : node178;
									assign node178 = (inp[8]) ? 3'b010 : 3'b110;
									assign node181 = (inp[8]) ? 3'b100 : 3'b010;
								assign node184 = (inp[8]) ? node188 : node185;
									assign node185 = (inp[5]) ? 3'b110 : 3'b001;
									assign node188 = (inp[5]) ? 3'b010 : 3'b110;
							assign node191 = (inp[5]) ? node199 : node192;
								assign node192 = (inp[8]) ? node196 : node193;
									assign node193 = (inp[11]) ? 3'b010 : 3'b100;
									assign node196 = (inp[11]) ? 3'b100 : 3'b000;
								assign node199 = (inp[11]) ? node201 : 3'b000;
									assign node201 = (inp[8]) ? 3'b000 : 3'b100;
						assign node204 = (inp[4]) ? 3'b000 : node205;
							assign node205 = (inp[5]) ? node213 : node206;
								assign node206 = (inp[11]) ? node210 : node207;
									assign node207 = (inp[8]) ? 3'b000 : 3'b100;
									assign node210 = (inp[8]) ? 3'b100 : 3'b010;
								assign node213 = (inp[11]) ? node215 : 3'b000;
									assign node215 = (inp[8]) ? 3'b000 : 3'b100;
			assign node219 = (inp[3]) ? 3'b000 : node220;
				assign node220 = (inp[10]) ? node238 : node221;
					assign node221 = (inp[7]) ? 3'b000 : node222;
						assign node222 = (inp[4]) ? 3'b000 : node223;
							assign node223 = (inp[8]) ? node231 : node224;
								assign node224 = (inp[11]) ? node228 : node225;
									assign node225 = (inp[5]) ? 3'b000 : 3'b100;
									assign node228 = (inp[5]) ? 3'b100 : 3'b010;
								assign node231 = (inp[11]) ? node233 : 3'b000;
									assign node233 = (inp[5]) ? 3'b000 : 3'b100;
					assign node238 = (inp[7]) ? node266 : node239;
						assign node239 = (inp[4]) ? node253 : node240;
							assign node240 = (inp[8]) ? node248 : node241;
								assign node241 = (inp[11]) ? node245 : node242;
									assign node242 = (inp[5]) ? 3'b010 : 3'b110;
									assign node245 = (inp[5]) ? 3'b110 : 3'b001;
								assign node248 = (inp[5]) ? 3'b010 : node249;
									assign node249 = (inp[11]) ? 3'b110 : 3'b010;
							assign node253 = (inp[8]) ? node261 : node254;
								assign node254 = (inp[11]) ? node258 : node255;
									assign node255 = (inp[5]) ? 3'b000 : 3'b100;
									assign node258 = (inp[5]) ? 3'b100 : 3'b010;
								assign node261 = (inp[11]) ? node263 : 3'b000;
									assign node263 = (inp[5]) ? 3'b000 : 3'b100;
						assign node266 = (inp[4]) ? node288 : node267;
							assign node267 = (inp[11]) ? node273 : node268;
								assign node268 = (inp[5]) ? 3'b000 : node269;
									assign node269 = (inp[8]) ? 3'b000 : 3'b100;
								assign node273 = (inp[5]) ? node281 : node274;
									assign node274 = (inp[8]) ? node276 : 3'b010;
										assign node276 = (inp[0]) ? 3'b100 : node277;
											assign node277 = (inp[1]) ? 3'b100 : 3'b000;
									assign node281 = (inp[8]) ? node283 : 3'b100;
										assign node283 = (inp[0]) ? 3'b000 : node284;
											assign node284 = (inp[2]) ? 3'b000 : 3'b100;
							assign node288 = (inp[8]) ? 3'b000 : node289;
								assign node289 = (inp[11]) ? node291 : 3'b000;
									assign node291 = (inp[2]) ? 3'b000 : node292;
										assign node292 = (inp[1]) ? 3'b000 : 3'b100;
		assign node298 = (inp[3]) ? node650 : node299;
			assign node299 = (inp[6]) ? node387 : node300;
				assign node300 = (inp[7]) ? node316 : node301;
					assign node301 = (inp[4]) ? node303 : 3'b111;
						assign node303 = (inp[10]) ? 3'b111 : node304;
							assign node304 = (inp[8]) ? node306 : 3'b111;
								assign node306 = (inp[5]) ? node310 : node307;
									assign node307 = (inp[11]) ? 3'b111 : 3'b011;
									assign node310 = (inp[11]) ? node312 : 3'b101;
										assign node312 = (inp[2]) ? 3'b011 : 3'b111;
					assign node316 = (inp[10]) ? node364 : node317;
						assign node317 = (inp[4]) ? node335 : node318;
							assign node318 = (inp[8]) ? node324 : node319;
								assign node319 = (inp[5]) ? node321 : 3'b111;
									assign node321 = (inp[11]) ? 3'b111 : 3'b011;
								assign node324 = (inp[11]) ? node328 : node325;
									assign node325 = (inp[5]) ? 3'b101 : 3'b011;
									assign node328 = (inp[5]) ? node330 : 3'b111;
										assign node330 = (inp[0]) ? 3'b011 : node331;
											assign node331 = (inp[1]) ? 3'b011 : 3'b011;
							assign node335 = (inp[0]) ? node357 : node336;
								assign node336 = (inp[8]) ? node348 : node337;
									assign node337 = (inp[11]) ? node341 : node338;
										assign node338 = (inp[5]) ? 3'b001 : 3'b101;
										assign node341 = (inp[5]) ? node345 : node342;
											assign node342 = (inp[2]) ? 3'b011 : 3'b011;
											assign node345 = (inp[2]) ? 3'b101 : 3'b011;
									assign node348 = (inp[5]) ? node352 : node349;
										assign node349 = (inp[11]) ? 3'b101 : 3'b001;
										assign node352 = (inp[11]) ? node354 : 3'b110;
											assign node354 = (inp[1]) ? 3'b001 : 3'b101;
								assign node357 = (inp[11]) ? 3'b101 : node358;
									assign node358 = (inp[2]) ? 3'b001 : node359;
										assign node359 = (inp[8]) ? 3'b001 : 3'b101;
						assign node364 = (inp[4]) ? node366 : 3'b111;
							assign node366 = (inp[5]) ? node372 : node367;
								assign node367 = (inp[11]) ? 3'b111 : node368;
									assign node368 = (inp[8]) ? 3'b011 : 3'b111;
								assign node372 = (inp[8]) ? node380 : node373;
									assign node373 = (inp[11]) ? 3'b111 : node374;
										assign node374 = (inp[0]) ? 3'b011 : node375;
											assign node375 = (inp[2]) ? 3'b011 : 3'b111;
									assign node380 = (inp[11]) ? 3'b011 : node381;
										assign node381 = (inp[0]) ? 3'b101 : node382;
											assign node382 = (inp[2]) ? 3'b101 : 3'b011;
				assign node387 = (inp[10]) ? node507 : node388;
					assign node388 = (inp[7]) ? node446 : node389;
						assign node389 = (inp[4]) ? node417 : node390;
							assign node390 = (inp[8]) ? node402 : node391;
								assign node391 = (inp[11]) ? node395 : node392;
									assign node392 = (inp[5]) ? 3'b001 : 3'b101;
									assign node395 = (inp[5]) ? node397 : 3'b011;
										assign node397 = (inp[1]) ? 3'b101 : node398;
											assign node398 = (inp[0]) ? 3'b101 : 3'b011;
								assign node402 = (inp[5]) ? node412 : node403;
									assign node403 = (inp[11]) ? node409 : node404;
										assign node404 = (inp[2]) ? 3'b001 : node405;
											assign node405 = (inp[0]) ? 3'b001 : 3'b101;
										assign node409 = (inp[1]) ? 3'b101 : 3'b011;
									assign node412 = (inp[11]) ? node414 : 3'b110;
										assign node414 = (inp[0]) ? 3'b001 : 3'b101;
							assign node417 = (inp[11]) ? node431 : node418;
								assign node418 = (inp[8]) ? node424 : node419;
									assign node419 = (inp[5]) ? node421 : 3'b110;
										assign node421 = (inp[0]) ? 3'b010 : 3'b110;
									assign node424 = (inp[5]) ? node426 : 3'b010;
										assign node426 = (inp[1]) ? 3'b100 : node427;
											assign node427 = (inp[0]) ? 3'b100 : 3'b010;
								assign node431 = (inp[0]) ? node437 : node432;
									assign node432 = (inp[5]) ? node434 : 3'b001;
										assign node434 = (inp[8]) ? 3'b110 : 3'b001;
									assign node437 = (inp[2]) ? node443 : node438;
										assign node438 = (inp[5]) ? node440 : 3'b110;
											assign node440 = (inp[8]) ? 3'b010 : 3'b110;
										assign node443 = (inp[5]) ? 3'b010 : 3'b001;
						assign node446 = (inp[4]) ? node480 : node447;
							assign node447 = (inp[11]) ? node465 : node448;
								assign node448 = (inp[8]) ? node456 : node449;
									assign node449 = (inp[5]) ? node451 : 3'b110;
										assign node451 = (inp[1]) ? 3'b010 : node452;
											assign node452 = (inp[0]) ? 3'b010 : 3'b110;
									assign node456 = (inp[5]) ? node462 : node457;
										assign node457 = (inp[0]) ? 3'b010 : node458;
											assign node458 = (inp[1]) ? 3'b010 : 3'b110;
										assign node462 = (inp[0]) ? 3'b100 : 3'b010;
								assign node465 = (inp[0]) ? node475 : node466;
									assign node466 = (inp[5]) ? node472 : node467;
										assign node467 = (inp[8]) ? 3'b001 : node468;
											assign node468 = (inp[2]) ? 3'b001 : 3'b101;
										assign node472 = (inp[8]) ? 3'b110 : 3'b001;
									assign node475 = (inp[5]) ? node477 : 3'b110;
										assign node477 = (inp[8]) ? 3'b010 : 3'b110;
							assign node480 = (inp[11]) ? node496 : node481;
								assign node481 = (inp[0]) ? 3'b000 : node482;
									assign node482 = (inp[2]) ? node488 : node483;
										assign node483 = (inp[8]) ? node485 : 3'b100;
											assign node485 = (inp[5]) ? 3'b000 : 3'b100;
										assign node488 = (inp[5]) ? node492 : node489;
											assign node489 = (inp[1]) ? 3'b100 : 3'b010;
											assign node492 = (inp[1]) ? 3'b000 : 3'b100;
								assign node496 = (inp[0]) ? node502 : node497;
									assign node497 = (inp[8]) ? 3'b010 : node498;
										assign node498 = (inp[5]) ? 3'b010 : 3'b110;
									assign node502 = (inp[8]) ? 3'b100 : node503;
										assign node503 = (inp[1]) ? 3'b010 : 3'b100;
					assign node507 = (inp[7]) ? node573 : node508;
						assign node508 = (inp[4]) ? node534 : node509;
							assign node509 = (inp[11]) ? node527 : node510;
								assign node510 = (inp[1]) ? node514 : node511;
									assign node511 = (inp[0]) ? 3'b101 : 3'b111;
									assign node514 = (inp[8]) ? node520 : node515;
										assign node515 = (inp[5]) ? node517 : 3'b111;
											assign node517 = (inp[0]) ? 3'b011 : 3'b111;
										assign node520 = (inp[0]) ? node524 : node521;
											assign node521 = (inp[5]) ? 3'b011 : 3'b111;
											assign node524 = (inp[5]) ? 3'b101 : 3'b011;
								assign node527 = (inp[8]) ? node529 : 3'b111;
									assign node529 = (inp[0]) ? node531 : 3'b111;
										assign node531 = (inp[5]) ? 3'b011 : 3'b111;
							assign node534 = (inp[11]) ? node552 : node535;
								assign node535 = (inp[0]) ? node547 : node536;
									assign node536 = (inp[1]) ? node542 : node537;
										assign node537 = (inp[8]) ? node539 : 3'b101;
											assign node539 = (inp[5]) ? 3'b001 : 3'b101;
										assign node542 = (inp[8]) ? node544 : 3'b011;
											assign node544 = (inp[5]) ? 3'b001 : 3'b101;
									assign node547 = (inp[5]) ? 3'b110 : node548;
										assign node548 = (inp[8]) ? 3'b001 : 3'b101;
								assign node552 = (inp[5]) ? node564 : node553;
									assign node553 = (inp[2]) ? node559 : node554;
										assign node554 = (inp[0]) ? 3'b011 : node555;
											assign node555 = (inp[8]) ? 3'b011 : 3'b111;
										assign node559 = (inp[8]) ? node561 : 3'b011;
											assign node561 = (inp[0]) ? 3'b101 : 3'b011;
									assign node564 = (inp[8]) ? node568 : node565;
										assign node565 = (inp[0]) ? 3'b101 : 3'b011;
										assign node568 = (inp[2]) ? node570 : 3'b101;
											assign node570 = (inp[0]) ? 3'b001 : 3'b101;
						assign node573 = (inp[4]) ? node617 : node574;
							assign node574 = (inp[11]) ? node596 : node575;
								assign node575 = (inp[1]) ? node583 : node576;
									assign node576 = (inp[5]) ? node578 : 3'b101;
										assign node578 = (inp[0]) ? 3'b001 : node579;
											assign node579 = (inp[8]) ? 3'b001 : 3'b101;
									assign node583 = (inp[0]) ? node591 : node584;
										assign node584 = (inp[5]) ? node588 : node585;
											assign node585 = (inp[8]) ? 3'b101 : 3'b011;
											assign node588 = (inp[8]) ? 3'b001 : 3'b101;
										assign node591 = (inp[5]) ? node593 : 3'b001;
											assign node593 = (inp[8]) ? 3'b110 : 3'b001;
								assign node596 = (inp[2]) ? node604 : node597;
									assign node597 = (inp[8]) ? 3'b011 : node598;
										assign node598 = (inp[5]) ? 3'b011 : node599;
											assign node599 = (inp[0]) ? 3'b011 : 3'b111;
									assign node604 = (inp[8]) ? node610 : node605;
										assign node605 = (inp[5]) ? node607 : 3'b011;
											assign node607 = (inp[0]) ? 3'b001 : 3'b011;
										assign node610 = (inp[5]) ? node614 : node611;
											assign node611 = (inp[0]) ? 3'b101 : 3'b011;
											assign node614 = (inp[0]) ? 3'b001 : 3'b101;
							assign node617 = (inp[8]) ? node631 : node618;
								assign node618 = (inp[0]) ? node624 : node619;
									assign node619 = (inp[11]) ? node621 : 3'b001;
										assign node621 = (inp[5]) ? 3'b001 : 3'b101;
									assign node624 = (inp[1]) ? 3'b110 : node625;
										assign node625 = (inp[11]) ? node627 : 3'b110;
											assign node627 = (inp[5]) ? 3'b001 : 3'b101;
								assign node631 = (inp[5]) ? node641 : node632;
									assign node632 = (inp[11]) ? node636 : node633;
										assign node633 = (inp[2]) ? 3'b110 : 3'b010;
										assign node636 = (inp[2]) ? node638 : 3'b001;
											assign node638 = (inp[1]) ? 3'b110 : 3'b001;
									assign node641 = (inp[0]) ? node645 : node642;
										assign node642 = (inp[11]) ? 3'b110 : 3'b010;
										assign node645 = (inp[11]) ? node647 : 3'b100;
											assign node647 = (inp[1]) ? 3'b010 : 3'b110;
			assign node650 = (inp[6]) ? node896 : node651;
				assign node651 = (inp[10]) ? node769 : node652;
					assign node652 = (inp[7]) ? node702 : node653;
						assign node653 = (inp[4]) ? node675 : node654;
							assign node654 = (inp[11]) ? node662 : node655;
								assign node655 = (inp[8]) ? node659 : node656;
									assign node656 = (inp[5]) ? 3'b001 : 3'b101;
									assign node659 = (inp[5]) ? 3'b110 : 3'b001;
								assign node662 = (inp[5]) ? node670 : node663;
									assign node663 = (inp[8]) ? node665 : 3'b011;
										assign node665 = (inp[0]) ? 3'b101 : node666;
											assign node666 = (inp[1]) ? 3'b101 : 3'b001;
									assign node670 = (inp[8]) ? node672 : 3'b101;
										assign node672 = (inp[2]) ? 3'b001 : 3'b101;
							assign node675 = (inp[11]) ? node687 : node676;
								assign node676 = (inp[8]) ? node680 : node677;
									assign node677 = (inp[5]) ? 3'b010 : 3'b110;
									assign node680 = (inp[5]) ? node682 : 3'b010;
										assign node682 = (inp[0]) ? 3'b100 : node683;
											assign node683 = (inp[1]) ? 3'b100 : 3'b010;
								assign node687 = (inp[5]) ? node695 : node688;
									assign node688 = (inp[8]) ? node690 : 3'b001;
										assign node690 = (inp[2]) ? node692 : 3'b110;
											assign node692 = (inp[1]) ? 3'b110 : 3'b001;
									assign node695 = (inp[0]) ? 3'b110 : node696;
										assign node696 = (inp[2]) ? 3'b110 : node697;
											assign node697 = (inp[1]) ? 3'b010 : 3'b001;
						assign node702 = (inp[4]) ? node744 : node703;
							assign node703 = (inp[1]) ? node729 : node704;
								assign node704 = (inp[2]) ? node714 : node705;
									assign node705 = (inp[11]) ? node709 : node706;
										assign node706 = (inp[0]) ? 3'b100 : 3'b110;
										assign node709 = (inp[5]) ? node711 : 3'b110;
											assign node711 = (inp[0]) ? 3'b010 : 3'b110;
									assign node714 = (inp[11]) ? node722 : node715;
										assign node715 = (inp[5]) ? node719 : node716;
											assign node716 = (inp[8]) ? 3'b010 : 3'b110;
											assign node719 = (inp[8]) ? 3'b100 : 3'b010;
										assign node722 = (inp[5]) ? node726 : node723;
											assign node723 = (inp[0]) ? 3'b001 : 3'b001;
											assign node726 = (inp[0]) ? 3'b010 : 3'b001;
								assign node729 = (inp[11]) ? node735 : node730;
									assign node730 = (inp[5]) ? 3'b010 : node731;
										assign node731 = (inp[8]) ? 3'b010 : 3'b110;
									assign node735 = (inp[5]) ? node739 : node736;
										assign node736 = (inp[8]) ? 3'b110 : 3'b001;
										assign node739 = (inp[8]) ? node741 : 3'b110;
											assign node741 = (inp[0]) ? 3'b010 : 3'b110;
							assign node744 = (inp[11]) ? node754 : node745;
								assign node745 = (inp[5]) ? 3'b000 : node746;
									assign node746 = (inp[8]) ? 3'b000 : node747;
										assign node747 = (inp[1]) ? 3'b100 : node748;
											assign node748 = (inp[2]) ? 3'b100 : 3'b010;
								assign node754 = (inp[5]) ? node762 : node755;
									assign node755 = (inp[1]) ? 3'b010 : node756;
										assign node756 = (inp[0]) ? 3'b100 : node757;
											assign node757 = (inp[8]) ? 3'b010 : 3'b110;
									assign node762 = (inp[1]) ? 3'b100 : node763;
										assign node763 = (inp[8]) ? node765 : 3'b010;
											assign node765 = (inp[2]) ? 3'b000 : 3'b100;
					assign node769 = (inp[7]) ? node827 : node770;
						assign node770 = (inp[4]) ? node792 : node771;
							assign node771 = (inp[11]) ? node787 : node772;
								assign node772 = (inp[8]) ? node780 : node773;
									assign node773 = (inp[5]) ? node775 : 3'b111;
										assign node775 = (inp[1]) ? 3'b011 : node776;
											assign node776 = (inp[0]) ? 3'b011 : 3'b111;
									assign node780 = (inp[5]) ? node782 : 3'b011;
										assign node782 = (inp[0]) ? 3'b101 : node783;
											assign node783 = (inp[2]) ? 3'b101 : 3'b011;
								assign node787 = (inp[8]) ? node789 : 3'b111;
									assign node789 = (inp[0]) ? 3'b011 : 3'b111;
							assign node792 = (inp[5]) ? node810 : node793;
								assign node793 = (inp[11]) ? node801 : node794;
									assign node794 = (inp[2]) ? 3'b101 : node795;
										assign node795 = (inp[8]) ? 3'b001 : node796;
											assign node796 = (inp[0]) ? 3'b101 : 3'b001;
									assign node801 = (inp[0]) ? node807 : node802;
										assign node802 = (inp[8]) ? 3'b011 : node803;
											assign node803 = (inp[2]) ? 3'b011 : 3'b111;
										assign node807 = (inp[1]) ? 3'b101 : 3'b011;
								assign node810 = (inp[11]) ? node820 : node811;
									assign node811 = (inp[0]) ? node817 : node812;
										assign node812 = (inp[2]) ? node814 : 3'b001;
											assign node814 = (inp[8]) ? 3'b000 : 3'b001;
										assign node817 = (inp[8]) ? 3'b110 : 3'b001;
									assign node820 = (inp[8]) ? node824 : node821;
										assign node821 = (inp[0]) ? 3'b101 : 3'b011;
										assign node824 = (inp[0]) ? 3'b001 : 3'b101;
						assign node827 = (inp[4]) ? node863 : node828;
							assign node828 = (inp[11]) ? node848 : node829;
								assign node829 = (inp[5]) ? node841 : node830;
									assign node830 = (inp[1]) ? node836 : node831;
										assign node831 = (inp[8]) ? 3'b101 : node832;
											assign node832 = (inp[0]) ? 3'b101 : 3'b011;
										assign node836 = (inp[2]) ? 3'b001 : node837;
											assign node837 = (inp[0]) ? 3'b001 : 3'b101;
									assign node841 = (inp[8]) ? node845 : node842;
										assign node842 = (inp[0]) ? 3'b001 : 3'b101;
										assign node845 = (inp[0]) ? 3'b110 : 3'b001;
								assign node848 = (inp[0]) ? node856 : node849;
									assign node849 = (inp[5]) ? node853 : node850;
										assign node850 = (inp[8]) ? 3'b011 : 3'b111;
										assign node853 = (inp[1]) ? 3'b101 : 3'b011;
									assign node856 = (inp[2]) ? 3'b101 : node857;
										assign node857 = (inp[8]) ? node859 : 3'b011;
											assign node859 = (inp[1]) ? 3'b001 : 3'b101;
							assign node863 = (inp[11]) ? node877 : node864;
								assign node864 = (inp[0]) ? node870 : node865;
									assign node865 = (inp[8]) ? node867 : 3'b110;
										assign node867 = (inp[5]) ? 3'b010 : 3'b110;
									assign node870 = (inp[8]) ? node874 : node871;
										assign node871 = (inp[5]) ? 3'b010 : 3'b110;
										assign node874 = (inp[5]) ? 3'b100 : 3'b010;
								assign node877 = (inp[8]) ? node885 : node878;
									assign node878 = (inp[5]) ? 3'b001 : node879;
										assign node879 = (inp[0]) ? node881 : 3'b101;
											assign node881 = (inp[1]) ? 3'b001 : 3'b001;
									assign node885 = (inp[5]) ? node891 : node886;
										assign node886 = (inp[0]) ? node888 : 3'b001;
											assign node888 = (inp[1]) ? 3'b110 : 3'b000;
										assign node891 = (inp[1]) ? node893 : 3'b110;
											assign node893 = (inp[0]) ? 3'b010 : 3'b110;
				assign node896 = (inp[10]) ? node942 : node897;
					assign node897 = (inp[4]) ? node931 : node898;
						assign node898 = (inp[7]) ? node922 : node899;
							assign node899 = (inp[11]) ? node909 : node900;
								assign node900 = (inp[0]) ? node904 : node901;
									assign node901 = (inp[5]) ? 3'b000 : 3'b010;
									assign node904 = (inp[8]) ? 3'b000 : node905;
										assign node905 = (inp[5]) ? 3'b000 : 3'b100;
								assign node909 = (inp[5]) ? node917 : node910;
									assign node910 = (inp[8]) ? node914 : node911;
										assign node911 = (inp[1]) ? 3'b010 : 3'b110;
										assign node914 = (inp[0]) ? 3'b100 : 3'b010;
									assign node917 = (inp[8]) ? node919 : 3'b100;
										assign node919 = (inp[0]) ? 3'b000 : 3'b100;
							assign node922 = (inp[8]) ? 3'b000 : node923;
								assign node923 = (inp[5]) ? 3'b000 : node924;
									assign node924 = (inp[0]) ? 3'b000 : node925;
										assign node925 = (inp[11]) ? 3'b100 : 3'b000;
						assign node931 = (inp[0]) ? 3'b000 : node932;
							assign node932 = (inp[8]) ? 3'b000 : node933;
								assign node933 = (inp[7]) ? 3'b000 : node934;
									assign node934 = (inp[2]) ? 3'b000 : node935;
										assign node935 = (inp[11]) ? 3'b100 : 3'b000;
					assign node942 = (inp[4]) ? node1006 : node943;
						assign node943 = (inp[7]) ? node985 : node944;
							assign node944 = (inp[11]) ? node962 : node945;
								assign node945 = (inp[0]) ? node953 : node946;
									assign node946 = (inp[5]) ? node950 : node947;
										assign node947 = (inp[8]) ? 3'b110 : 3'b001;
										assign node950 = (inp[8]) ? 3'b010 : 3'b110;
									assign node953 = (inp[5]) ? node959 : node954;
										assign node954 = (inp[2]) ? node956 : 3'b110;
											assign node956 = (inp[8]) ? 3'b010 : 3'b110;
										assign node959 = (inp[8]) ? 3'b100 : 3'b010;
								assign node962 = (inp[1]) ? node972 : node963;
									assign node963 = (inp[8]) ? node969 : node964;
										assign node964 = (inp[5]) ? 3'b001 : node965;
											assign node965 = (inp[0]) ? 3'b001 : 3'b101;
										assign node969 = (inp[5]) ? 3'b110 : 3'b001;
									assign node972 = (inp[5]) ? node978 : node973;
										assign node973 = (inp[8]) ? node975 : 3'b001;
											assign node975 = (inp[0]) ? 3'b110 : 3'b001;
										assign node978 = (inp[0]) ? node982 : node979;
											assign node979 = (inp[8]) ? 3'b110 : 3'b001;
											assign node982 = (inp[8]) ? 3'b010 : 3'b110;
							assign node985 = (inp[11]) ? node999 : node986;
								assign node986 = (inp[8]) ? node992 : node987;
									assign node987 = (inp[5]) ? node989 : 3'b010;
										assign node989 = (inp[0]) ? 3'b000 : 3'b100;
									assign node992 = (inp[5]) ? 3'b000 : node993;
										assign node993 = (inp[0]) ? node995 : 3'b100;
											assign node995 = (inp[1]) ? 3'b000 : 3'b100;
								assign node999 = (inp[5]) ? node1003 : node1000;
									assign node1000 = (inp[8]) ? 3'b010 : 3'b110;
									assign node1003 = (inp[8]) ? 3'b100 : 3'b010;
						assign node1006 = (inp[7]) ? node1040 : node1007;
							assign node1007 = (inp[5]) ? node1023 : node1008;
								assign node1008 = (inp[11]) ? node1016 : node1009;
									assign node1009 = (inp[0]) ? node1013 : node1010;
										assign node1010 = (inp[8]) ? 3'b100 : 3'b010;
										assign node1013 = (inp[8]) ? 3'b000 : 3'b100;
									assign node1016 = (inp[2]) ? node1018 : 3'b110;
										assign node1018 = (inp[0]) ? 3'b010 : node1019;
											assign node1019 = (inp[8]) ? 3'b010 : 3'b110;
								assign node1023 = (inp[11]) ? node1031 : node1024;
									assign node1024 = (inp[8]) ? 3'b000 : node1025;
										assign node1025 = (inp[0]) ? node1027 : 3'b100;
											assign node1027 = (inp[1]) ? 3'b000 : 3'b000;
									assign node1031 = (inp[8]) ? node1035 : node1032;
										assign node1032 = (inp[0]) ? 3'b100 : 3'b010;
										assign node1035 = (inp[2]) ? node1037 : 3'b100;
											assign node1037 = (inp[1]) ? 3'b000 : 3'b100;
							assign node1040 = (inp[8]) ? 3'b000 : node1041;
								assign node1041 = (inp[11]) ? node1043 : 3'b000;
									assign node1043 = (inp[5]) ? 3'b000 : 3'b100;

endmodule