module dtc_split25_bm99 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node26;
	wire [3-1:0] node32;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node137;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node141;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node188;

	assign outp = (inp[3]) ? node152 : node1;
		assign node1 = (inp[9]) ? node55 : node2;
			assign node2 = (inp[4]) ? node32 : node3;
				assign node3 = (inp[0]) ? node11 : node4;
					assign node4 = (inp[6]) ? 3'b000 : node5;
						assign node5 = (inp[5]) ? node7 : 3'b001;
							assign node7 = (inp[1]) ? 3'b001 : 3'b000;
					assign node11 = (inp[6]) ? 3'b001 : node12;
						assign node12 = (inp[5]) ? node22 : node13;
							assign node13 = (inp[1]) ? 3'b000 : node14;
								assign node14 = (inp[10]) ? node18 : node15;
									assign node15 = (inp[11]) ? 3'b000 : 3'b001;
									assign node18 = (inp[11]) ? 3'b001 : 3'b000;
							assign node22 = (inp[1]) ? 3'b001 : node23;
								assign node23 = (inp[10]) ? 3'b000 : node24;
									assign node24 = (inp[11]) ? node26 : 3'b000;
										assign node26 = (inp[2]) ? 3'b000 : 3'b001;
				assign node32 = (inp[0]) ? node34 : 3'b000;
					assign node34 = (inp[1]) ? node50 : node35;
						assign node35 = (inp[5]) ? node43 : node36;
							assign node36 = (inp[10]) ? node38 : 3'b000;
								assign node38 = (inp[2]) ? node40 : 3'b000;
									assign node40 = (inp[11]) ? 3'b000 : 3'b001;
							assign node43 = (inp[6]) ? 3'b001 : node44;
								assign node44 = (inp[7]) ? node46 : 3'b000;
									assign node46 = (inp[10]) ? 3'b001 : 3'b000;
						assign node50 = (inp[5]) ? 3'b000 : node51;
							assign node51 = (inp[6]) ? 3'b000 : 3'b001;
			assign node55 = (inp[6]) ? node113 : node56;
				assign node56 = (inp[4]) ? node88 : node57;
					assign node57 = (inp[0]) ? node67 : node58;
						assign node58 = (inp[1]) ? node64 : node59;
							assign node59 = (inp[5]) ? 3'b100 : node60;
								assign node60 = (inp[7]) ? 3'b110 : 3'b010;
							assign node64 = (inp[5]) ? 3'b010 : 3'b110;
						assign node67 = (inp[5]) ? node77 : node68;
							assign node68 = (inp[7]) ? node74 : node69;
								assign node69 = (inp[10]) ? node71 : 3'b001;
									assign node71 = (inp[1]) ? 3'b001 : 3'b110;
								assign node74 = (inp[11]) ? 3'b101 : 3'b001;
							assign node77 = (inp[1]) ? 3'b110 : node78;
								assign node78 = (inp[2]) ? node84 : node79;
									assign node79 = (inp[7]) ? node81 : 3'b001;
										assign node81 = (inp[11]) ? 3'b110 : 3'b001;
									assign node84 = (inp[8]) ? 3'b110 : 3'b001;
					assign node88 = (inp[0]) ? node98 : node89;
						assign node89 = (inp[2]) ? node91 : 3'b000;
							assign node91 = (inp[10]) ? node93 : 3'b000;
								assign node93 = (inp[5]) ? 3'b000 : node94;
									assign node94 = (inp[7]) ? 3'b000 : 3'b100;
						assign node98 = (inp[5]) ? node106 : node99;
							assign node99 = (inp[1]) ? 3'b010 : node100;
								assign node100 = (inp[10]) ? node102 : 3'b100;
									assign node102 = (inp[2]) ? 3'b010 : 3'b100;
							assign node106 = (inp[1]) ? 3'b100 : node107;
								assign node107 = (inp[10]) ? node109 : 3'b100;
									assign node109 = (inp[7]) ? 3'b010 : 3'b100;
				assign node113 = (inp[0]) ? node123 : node114;
					assign node114 = (inp[11]) ? node116 : 3'b001;
						assign node116 = (inp[4]) ? 3'b001 : node117;
							assign node117 = (inp[7]) ? node119 : 3'b001;
								assign node119 = (inp[2]) ? 3'b011 : 3'b001;
					assign node123 = (inp[4]) ? node137 : node124;
						assign node124 = (inp[5]) ? 3'b011 : node125;
							assign node125 = (inp[1]) ? 3'b111 : node126;
								assign node126 = (inp[8]) ? 3'b011 : node127;
									assign node127 = (inp[11]) ? node129 : 3'b111;
										assign node129 = (inp[10]) ? node131 : 3'b011;
											assign node131 = (inp[2]) ? 3'b111 : 3'b011;
						assign node137 = (inp[5]) ? node145 : node138;
							assign node138 = (inp[1]) ? 3'b101 : node139;
								assign node139 = (inp[8]) ? node141 : 3'b001;
									assign node141 = (inp[10]) ? 3'b101 : 3'b001;
							assign node145 = (inp[1]) ? 3'b001 : node146;
								assign node146 = (inp[10]) ? node148 : 3'b010;
									assign node148 = (inp[7]) ? 3'b110 : 3'b010;
		assign node152 = (inp[6]) ? node154 : 3'b000;
			assign node154 = (inp[0]) ? node170 : node155;
				assign node155 = (inp[9]) ? node167 : node156;
					assign node156 = (inp[4]) ? node158 : 3'b000;
						assign node158 = (inp[10]) ? node160 : 3'b010;
							assign node160 = (inp[5]) ? node164 : node161;
								assign node161 = (inp[2]) ? 3'b100 : 3'b010;
								assign node164 = (inp[1]) ? 3'b100 : 3'b010;
					assign node167 = (inp[4]) ? 3'b000 : 3'b100;
				assign node170 = (inp[4]) ? node174 : node171;
					assign node171 = (inp[9]) ? 3'b010 : 3'b001;
					assign node174 = (inp[9]) ? node186 : node175;
						assign node175 = (inp[10]) ? node181 : node176;
							assign node176 = (inp[7]) ? 3'b110 : node177;
								assign node177 = (inp[1]) ? 3'b110 : 3'b010;
							assign node181 = (inp[1]) ? node183 : 3'b010;
								assign node183 = (inp[7]) ? 3'b010 : 3'b110;
						assign node186 = (inp[11]) ? 3'b000 : node187;
							assign node187 = (inp[10]) ? 3'b000 : node188;
								assign node188 = (inp[7]) ? 3'b100 : 3'b000;

endmodule