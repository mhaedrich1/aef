module dtc_split33_bm26 (
	input  wire [15-1:0] inp,
	output wire [15-1:0] outp
);

	wire [15-1:0] node1;
	wire [15-1:0] node2;
	wire [15-1:0] node3;
	wire [15-1:0] node4;
	wire [15-1:0] node5;
	wire [15-1:0] node6;
	wire [15-1:0] node7;
	wire [15-1:0] node8;
	wire [15-1:0] node9;
	wire [15-1:0] node10;
	wire [15-1:0] node11;
	wire [15-1:0] node12;
	wire [15-1:0] node13;
	wire [15-1:0] node16;
	wire [15-1:0] node19;
	wire [15-1:0] node21;
	wire [15-1:0] node24;
	wire [15-1:0] node25;
	wire [15-1:0] node26;
	wire [15-1:0] node28;
	wire [15-1:0] node33;
	wire [15-1:0] node34;
	wire [15-1:0] node36;
	wire [15-1:0] node37;
	wire [15-1:0] node41;
	wire [15-1:0] node43;
	wire [15-1:0] node46;
	wire [15-1:0] node47;
	wire [15-1:0] node48;
	wire [15-1:0] node51;
	wire [15-1:0] node52;
	wire [15-1:0] node53;
	wire [15-1:0] node55;
	wire [15-1:0] node59;
	wire [15-1:0] node62;
	wire [15-1:0] node63;
	wire [15-1:0] node64;
	wire [15-1:0] node65;
	wire [15-1:0] node67;
	wire [15-1:0] node71;
	wire [15-1:0] node74;
	wire [15-1:0] node76;
	wire [15-1:0] node78;
	wire [15-1:0] node81;
	wire [15-1:0] node82;
	wire [15-1:0] node83;
	wire [15-1:0] node84;
	wire [15-1:0] node85;
	wire [15-1:0] node86;
	wire [15-1:0] node91;
	wire [15-1:0] node92;
	wire [15-1:0] node93;
	wire [15-1:0] node95;
	wire [15-1:0] node100;
	wire [15-1:0] node102;
	wire [15-1:0] node103;
	wire [15-1:0] node107;
	wire [15-1:0] node108;
	wire [15-1:0] node109;
	wire [15-1:0] node111;
	wire [15-1:0] node113;
	wire [15-1:0] node116;
	wire [15-1:0] node117;
	wire [15-1:0] node119;
	wire [15-1:0] node122;
	wire [15-1:0] node124;
	wire [15-1:0] node127;
	wire [15-1:0] node129;
	wire [15-1:0] node130;
	wire [15-1:0] node131;
	wire [15-1:0] node132;
	wire [15-1:0] node136;
	wire [15-1:0] node137;
	wire [15-1:0] node142;
	wire [15-1:0] node143;
	wire [15-1:0] node144;
	wire [15-1:0] node145;
	wire [15-1:0] node146;
	wire [15-1:0] node147;
	wire [15-1:0] node150;
	wire [15-1:0] node153;
	wire [15-1:0] node154;
	wire [15-1:0] node157;
	wire [15-1:0] node160;
	wire [15-1:0] node161;
	wire [15-1:0] node162;
	wire [15-1:0] node165;
	wire [15-1:0] node166;
	wire [15-1:0] node168;
	wire [15-1:0] node172;
	wire [15-1:0] node174;
	wire [15-1:0] node177;
	wire [15-1:0] node178;
	wire [15-1:0] node179;
	wire [15-1:0] node181;
	wire [15-1:0] node183;
	wire [15-1:0] node186;
	wire [15-1:0] node189;
	wire [15-1:0] node190;
	wire [15-1:0] node192;
	wire [15-1:0] node196;
	wire [15-1:0] node197;
	wire [15-1:0] node198;
	wire [15-1:0] node199;
	wire [15-1:0] node202;
	wire [15-1:0] node203;
	wire [15-1:0] node205;
	wire [15-1:0] node207;
	wire [15-1:0] node210;
	wire [15-1:0] node213;
	wire [15-1:0] node214;
	wire [15-1:0] node215;
	wire [15-1:0] node220;
	wire [15-1:0] node221;
	wire [15-1:0] node222;
	wire [15-1:0] node223;
	wire [15-1:0] node226;
	wire [15-1:0] node230;
	wire [15-1:0] node231;
	wire [15-1:0] node232;
	wire [15-1:0] node235;
	wire [15-1:0] node236;
	wire [15-1:0] node241;
	wire [15-1:0] node242;
	wire [15-1:0] node243;
	wire [15-1:0] node244;
	wire [15-1:0] node245;
	wire [15-1:0] node246;
	wire [15-1:0] node247;
	wire [15-1:0] node250;
	wire [15-1:0] node253;
	wire [15-1:0] node255;
	wire [15-1:0] node256;
	wire [15-1:0] node257;
	wire [15-1:0] node260;
	wire [15-1:0] node264;
	wire [15-1:0] node265;
	wire [15-1:0] node266;
	wire [15-1:0] node269;
	wire [15-1:0] node272;
	wire [15-1:0] node274;
	wire [15-1:0] node277;
	wire [15-1:0] node278;
	wire [15-1:0] node279;
	wire [15-1:0] node280;
	wire [15-1:0] node281;
	wire [15-1:0] node285;
	wire [15-1:0] node288;
	wire [15-1:0] node289;
	wire [15-1:0] node292;
	wire [15-1:0] node295;
	wire [15-1:0] node296;
	wire [15-1:0] node297;
	wire [15-1:0] node301;
	wire [15-1:0] node302;
	wire [15-1:0] node306;
	wire [15-1:0] node307;
	wire [15-1:0] node308;
	wire [15-1:0] node309;
	wire [15-1:0] node311;
	wire [15-1:0] node314;
	wire [15-1:0] node315;
	wire [15-1:0] node317;
	wire [15-1:0] node318;
	wire [15-1:0] node323;
	wire [15-1:0] node324;
	wire [15-1:0] node325;
	wire [15-1:0] node328;
	wire [15-1:0] node330;
	wire [15-1:0] node333;
	wire [15-1:0] node335;
	wire [15-1:0] node338;
	wire [15-1:0] node339;
	wire [15-1:0] node340;
	wire [15-1:0] node342;
	wire [15-1:0] node344;
	wire [15-1:0] node347;
	wire [15-1:0] node348;
	wire [15-1:0] node350;
	wire [15-1:0] node354;
	wire [15-1:0] node355;
	wire [15-1:0] node357;
	wire [15-1:0] node359;
	wire [15-1:0] node362;
	wire [15-1:0] node364;
	wire [15-1:0] node366;
	wire [15-1:0] node369;
	wire [15-1:0] node370;
	wire [15-1:0] node371;
	wire [15-1:0] node372;
	wire [15-1:0] node373;
	wire [15-1:0] node374;
	wire [15-1:0] node375;
	wire [15-1:0] node378;
	wire [15-1:0] node379;
	wire [15-1:0] node384;
	wire [15-1:0] node385;
	wire [15-1:0] node389;
	wire [15-1:0] node390;
	wire [15-1:0] node391;
	wire [15-1:0] node392;
	wire [15-1:0] node396;
	wire [15-1:0] node398;
	wire [15-1:0] node399;
	wire [15-1:0] node403;
	wire [15-1:0] node405;
	wire [15-1:0] node406;
	wire [15-1:0] node410;
	wire [15-1:0] node411;
	wire [15-1:0] node412;
	wire [15-1:0] node414;
	wire [15-1:0] node417;
	wire [15-1:0] node418;
	wire [15-1:0] node422;
	wire [15-1:0] node423;
	wire [15-1:0] node426;
	wire [15-1:0] node427;
	wire [15-1:0] node430;
	wire [15-1:0] node433;
	wire [15-1:0] node434;
	wire [15-1:0] node435;
	wire [15-1:0] node436;
	wire [15-1:0] node439;
	wire [15-1:0] node442;
	wire [15-1:0] node443;
	wire [15-1:0] node444;
	wire [15-1:0] node447;
	wire [15-1:0] node450;
	wire [15-1:0] node451;
	wire [15-1:0] node452;
	wire [15-1:0] node454;
	wire [15-1:0] node459;
	wire [15-1:0] node460;
	wire [15-1:0] node461;
	wire [15-1:0] node462;
	wire [15-1:0] node463;
	wire [15-1:0] node468;
	wire [15-1:0] node469;
	wire [15-1:0] node470;
	wire [15-1:0] node472;
	wire [15-1:0] node476;
	wire [15-1:0] node477;
	wire [15-1:0] node478;
	wire [15-1:0] node482;
	wire [15-1:0] node483;
	wire [15-1:0] node487;
	wire [15-1:0] node488;
	wire [15-1:0] node489;
	wire [15-1:0] node491;
	wire [15-1:0] node495;
	wire [15-1:0] node497;
	wire [15-1:0] node499;
	wire [15-1:0] node502;
	wire [15-1:0] node503;
	wire [15-1:0] node504;
	wire [15-1:0] node505;
	wire [15-1:0] node506;
	wire [15-1:0] node507;
	wire [15-1:0] node509;
	wire [15-1:0] node510;
	wire [15-1:0] node511;
	wire [15-1:0] node516;
	wire [15-1:0] node517;
	wire [15-1:0] node519;
	wire [15-1:0] node522;
	wire [15-1:0] node525;
	wire [15-1:0] node526;
	wire [15-1:0] node527;
	wire [15-1:0] node529;
	wire [15-1:0] node532;
	wire [15-1:0] node533;
	wire [15-1:0] node534;
	wire [15-1:0] node535;
	wire [15-1:0] node540;
	wire [15-1:0] node543;
	wire [15-1:0] node544;
	wire [15-1:0] node545;
	wire [15-1:0] node546;
	wire [15-1:0] node551;
	wire [15-1:0] node552;
	wire [15-1:0] node556;
	wire [15-1:0] node557;
	wire [15-1:0] node558;
	wire [15-1:0] node559;
	wire [15-1:0] node560;
	wire [15-1:0] node564;
	wire [15-1:0] node565;
	wire [15-1:0] node568;
	wire [15-1:0] node571;
	wire [15-1:0] node572;
	wire [15-1:0] node573;
	wire [15-1:0] node575;
	wire [15-1:0] node578;
	wire [15-1:0] node579;
	wire [15-1:0] node580;
	wire [15-1:0] node584;
	wire [15-1:0] node587;
	wire [15-1:0] node589;
	wire [15-1:0] node591;
	wire [15-1:0] node594;
	wire [15-1:0] node595;
	wire [15-1:0] node596;
	wire [15-1:0] node597;
	wire [15-1:0] node600;
	wire [15-1:0] node601;
	wire [15-1:0] node605;
	wire [15-1:0] node606;
	wire [15-1:0] node609;
	wire [15-1:0] node612;
	wire [15-1:0] node613;
	wire [15-1:0] node615;
	wire [15-1:0] node618;
	wire [15-1:0] node619;
	wire [15-1:0] node623;
	wire [15-1:0] node624;
	wire [15-1:0] node625;
	wire [15-1:0] node626;
	wire [15-1:0] node627;
	wire [15-1:0] node628;
	wire [15-1:0] node631;
	wire [15-1:0] node633;
	wire [15-1:0] node637;
	wire [15-1:0] node638;
	wire [15-1:0] node640;
	wire [15-1:0] node643;
	wire [15-1:0] node645;
	wire [15-1:0] node648;
	wire [15-1:0] node649;
	wire [15-1:0] node650;
	wire [15-1:0] node651;
	wire [15-1:0] node655;
	wire [15-1:0] node656;
	wire [15-1:0] node660;
	wire [15-1:0] node662;
	wire [15-1:0] node665;
	wire [15-1:0] node666;
	wire [15-1:0] node667;
	wire [15-1:0] node668;
	wire [15-1:0] node670;
	wire [15-1:0] node672;
	wire [15-1:0] node675;
	wire [15-1:0] node676;
	wire [15-1:0] node677;
	wire [15-1:0] node679;
	wire [15-1:0] node683;
	wire [15-1:0] node685;
	wire [15-1:0] node688;
	wire [15-1:0] node690;
	wire [15-1:0] node691;
	wire [15-1:0] node692;
	wire [15-1:0] node693;
	wire [15-1:0] node698;
	wire [15-1:0] node701;
	wire [15-1:0] node702;
	wire [15-1:0] node703;
	wire [15-1:0] node704;
	wire [15-1:0] node708;
	wire [15-1:0] node711;
	wire [15-1:0] node712;
	wire [15-1:0] node713;
	wire [15-1:0] node715;
	wire [15-1:0] node718;
	wire [15-1:0] node720;
	wire [15-1:0] node723;
	wire [15-1:0] node726;
	wire [15-1:0] node727;
	wire [15-1:0] node728;
	wire [15-1:0] node729;
	wire [15-1:0] node730;
	wire [15-1:0] node731;
	wire [15-1:0] node732;
	wire [15-1:0] node734;
	wire [15-1:0] node738;
	wire [15-1:0] node739;
	wire [15-1:0] node743;
	wire [15-1:0] node744;
	wire [15-1:0] node746;
	wire [15-1:0] node747;
	wire [15-1:0] node748;
	wire [15-1:0] node753;
	wire [15-1:0] node754;
	wire [15-1:0] node757;
	wire [15-1:0] node760;
	wire [15-1:0] node761;
	wire [15-1:0] node763;
	wire [15-1:0] node764;
	wire [15-1:0] node766;
	wire [15-1:0] node769;
	wire [15-1:0] node770;
	wire [15-1:0] node771;
	wire [15-1:0] node775;
	wire [15-1:0] node778;
	wire [15-1:0] node779;
	wire [15-1:0] node780;
	wire [15-1:0] node784;
	wire [15-1:0] node787;
	wire [15-1:0] node788;
	wire [15-1:0] node789;
	wire [15-1:0] node790;
	wire [15-1:0] node791;
	wire [15-1:0] node792;
	wire [15-1:0] node796;
	wire [15-1:0] node797;
	wire [15-1:0] node801;
	wire [15-1:0] node802;
	wire [15-1:0] node804;
	wire [15-1:0] node808;
	wire [15-1:0] node809;
	wire [15-1:0] node810;
	wire [15-1:0] node813;
	wire [15-1:0] node815;
	wire [15-1:0] node818;
	wire [15-1:0] node819;
	wire [15-1:0] node820;
	wire [15-1:0] node825;
	wire [15-1:0] node826;
	wire [15-1:0] node827;
	wire [15-1:0] node828;
	wire [15-1:0] node829;
	wire [15-1:0] node833;
	wire [15-1:0] node834;
	wire [15-1:0] node836;
	wire [15-1:0] node840;
	wire [15-1:0] node842;
	wire [15-1:0] node844;
	wire [15-1:0] node847;
	wire [15-1:0] node848;
	wire [15-1:0] node849;
	wire [15-1:0] node851;
	wire [15-1:0] node854;
	wire [15-1:0] node855;
	wire [15-1:0] node858;
	wire [15-1:0] node861;
	wire [15-1:0] node863;
	wire [15-1:0] node866;
	wire [15-1:0] node867;
	wire [15-1:0] node868;
	wire [15-1:0] node869;
	wire [15-1:0] node870;
	wire [15-1:0] node873;
	wire [15-1:0] node876;
	wire [15-1:0] node877;
	wire [15-1:0] node878;
	wire [15-1:0] node881;
	wire [15-1:0] node883;
	wire [15-1:0] node886;
	wire [15-1:0] node888;
	wire [15-1:0] node891;
	wire [15-1:0] node892;
	wire [15-1:0] node893;
	wire [15-1:0] node894;
	wire [15-1:0] node895;
	wire [15-1:0] node899;
	wire [15-1:0] node900;
	wire [15-1:0] node902;
	wire [15-1:0] node906;
	wire [15-1:0] node907;
	wire [15-1:0] node909;
	wire [15-1:0] node912;
	wire [15-1:0] node914;
	wire [15-1:0] node917;
	wire [15-1:0] node918;
	wire [15-1:0] node919;
	wire [15-1:0] node920;
	wire [15-1:0] node924;
	wire [15-1:0] node926;
	wire [15-1:0] node929;
	wire [15-1:0] node930;
	wire [15-1:0] node931;
	wire [15-1:0] node935;
	wire [15-1:0] node938;
	wire [15-1:0] node939;
	wire [15-1:0] node940;
	wire [15-1:0] node941;
	wire [15-1:0] node942;
	wire [15-1:0] node944;
	wire [15-1:0] node945;
	wire [15-1:0] node949;
	wire [15-1:0] node952;
	wire [15-1:0] node953;
	wire [15-1:0] node956;
	wire [15-1:0] node959;
	wire [15-1:0] node960;
	wire [15-1:0] node962;
	wire [15-1:0] node965;
	wire [15-1:0] node966;
	wire [15-1:0] node969;
	wire [15-1:0] node972;
	wire [15-1:0] node973;
	wire [15-1:0] node975;
	wire [15-1:0] node977;
	wire [15-1:0] node979;
	wire [15-1:0] node982;
	wire [15-1:0] node983;
	wire [15-1:0] node984;
	wire [15-1:0] node986;
	wire [15-1:0] node990;
	wire [15-1:0] node991;
	wire [15-1:0] node995;
	wire [15-1:0] node996;
	wire [15-1:0] node997;
	wire [15-1:0] node998;
	wire [15-1:0] node999;
	wire [15-1:0] node1000;
	wire [15-1:0] node1001;
	wire [15-1:0] node1002;
	wire [15-1:0] node1003;
	wire [15-1:0] node1004;
	wire [15-1:0] node1007;
	wire [15-1:0] node1010;
	wire [15-1:0] node1011;
	wire [15-1:0] node1013;
	wire [15-1:0] node1017;
	wire [15-1:0] node1018;
	wire [15-1:0] node1019;
	wire [15-1:0] node1021;
	wire [15-1:0] node1024;
	wire [15-1:0] node1025;
	wire [15-1:0] node1029;
	wire [15-1:0] node1031;
	wire [15-1:0] node1032;
	wire [15-1:0] node1036;
	wire [15-1:0] node1037;
	wire [15-1:0] node1039;
	wire [15-1:0] node1041;
	wire [15-1:0] node1044;
	wire [15-1:0] node1045;
	wire [15-1:0] node1049;
	wire [15-1:0] node1050;
	wire [15-1:0] node1051;
	wire [15-1:0] node1052;
	wire [15-1:0] node1053;
	wire [15-1:0] node1057;
	wire [15-1:0] node1060;
	wire [15-1:0] node1061;
	wire [15-1:0] node1063;
	wire [15-1:0] node1067;
	wire [15-1:0] node1068;
	wire [15-1:0] node1069;
	wire [15-1:0] node1071;
	wire [15-1:0] node1072;
	wire [15-1:0] node1076;
	wire [15-1:0] node1077;
	wire [15-1:0] node1081;
	wire [15-1:0] node1082;
	wire [15-1:0] node1083;
	wire [15-1:0] node1087;
	wire [15-1:0] node1090;
	wire [15-1:0] node1091;
	wire [15-1:0] node1092;
	wire [15-1:0] node1093;
	wire [15-1:0] node1094;
	wire [15-1:0] node1096;
	wire [15-1:0] node1097;
	wire [15-1:0] node1101;
	wire [15-1:0] node1103;
	wire [15-1:0] node1106;
	wire [15-1:0] node1107;
	wire [15-1:0] node1109;
	wire [15-1:0] node1112;
	wire [15-1:0] node1113;
	wire [15-1:0] node1115;
	wire [15-1:0] node1119;
	wire [15-1:0] node1120;
	wire [15-1:0] node1121;
	wire [15-1:0] node1122;
	wire [15-1:0] node1126;
	wire [15-1:0] node1128;
	wire [15-1:0] node1131;
	wire [15-1:0] node1132;
	wire [15-1:0] node1133;
	wire [15-1:0] node1135;
	wire [15-1:0] node1140;
	wire [15-1:0] node1141;
	wire [15-1:0] node1142;
	wire [15-1:0] node1143;
	wire [15-1:0] node1144;
	wire [15-1:0] node1148;
	wire [15-1:0] node1151;
	wire [15-1:0] node1152;
	wire [15-1:0] node1153;
	wire [15-1:0] node1158;
	wire [15-1:0] node1159;
	wire [15-1:0] node1160;
	wire [15-1:0] node1161;
	wire [15-1:0] node1163;
	wire [15-1:0] node1166;
	wire [15-1:0] node1167;
	wire [15-1:0] node1171;
	wire [15-1:0] node1174;
	wire [15-1:0] node1176;
	wire [15-1:0] node1177;
	wire [15-1:0] node1181;
	wire [15-1:0] node1182;
	wire [15-1:0] node1183;
	wire [15-1:0] node1184;
	wire [15-1:0] node1186;
	wire [15-1:0] node1187;
	wire [15-1:0] node1189;
	wire [15-1:0] node1192;
	wire [15-1:0] node1193;
	wire [15-1:0] node1194;
	wire [15-1:0] node1199;
	wire [15-1:0] node1200;
	wire [15-1:0] node1201;
	wire [15-1:0] node1204;
	wire [15-1:0] node1207;
	wire [15-1:0] node1209;
	wire [15-1:0] node1212;
	wire [15-1:0] node1213;
	wire [15-1:0] node1214;
	wire [15-1:0] node1215;
	wire [15-1:0] node1218;
	wire [15-1:0] node1222;
	wire [15-1:0] node1223;
	wire [15-1:0] node1224;
	wire [15-1:0] node1227;
	wire [15-1:0] node1229;
	wire [15-1:0] node1232;
	wire [15-1:0] node1233;
	wire [15-1:0] node1236;
	wire [15-1:0] node1239;
	wire [15-1:0] node1240;
	wire [15-1:0] node1241;
	wire [15-1:0] node1242;
	wire [15-1:0] node1244;
	wire [15-1:0] node1247;
	wire [15-1:0] node1248;
	wire [15-1:0] node1252;
	wire [15-1:0] node1253;
	wire [15-1:0] node1254;
	wire [15-1:0] node1255;
	wire [15-1:0] node1259;
	wire [15-1:0] node1260;
	wire [15-1:0] node1264;
	wire [15-1:0] node1265;
	wire [15-1:0] node1267;
	wire [15-1:0] node1271;
	wire [15-1:0] node1272;
	wire [15-1:0] node1273;
	wire [15-1:0] node1274;
	wire [15-1:0] node1275;
	wire [15-1:0] node1279;
	wire [15-1:0] node1280;
	wire [15-1:0] node1282;
	wire [15-1:0] node1286;
	wire [15-1:0] node1288;
	wire [15-1:0] node1291;
	wire [15-1:0] node1292;
	wire [15-1:0] node1293;
	wire [15-1:0] node1294;
	wire [15-1:0] node1299;
	wire [15-1:0] node1300;
	wire [15-1:0] node1302;
	wire [15-1:0] node1303;
	wire [15-1:0] node1307;
	wire [15-1:0] node1310;
	wire [15-1:0] node1311;
	wire [15-1:0] node1312;
	wire [15-1:0] node1313;
	wire [15-1:0] node1314;
	wire [15-1:0] node1315;
	wire [15-1:0] node1316;
	wire [15-1:0] node1319;
	wire [15-1:0] node1321;
	wire [15-1:0] node1324;
	wire [15-1:0] node1325;
	wire [15-1:0] node1327;
	wire [15-1:0] node1331;
	wire [15-1:0] node1332;
	wire [15-1:0] node1333;
	wire [15-1:0] node1335;
	wire [15-1:0] node1336;
	wire [15-1:0] node1341;
	wire [15-1:0] node1342;
	wire [15-1:0] node1345;
	wire [15-1:0] node1346;
	wire [15-1:0] node1350;
	wire [15-1:0] node1351;
	wire [15-1:0] node1352;
	wire [15-1:0] node1353;
	wire [15-1:0] node1356;
	wire [15-1:0] node1359;
	wire [15-1:0] node1360;
	wire [15-1:0] node1364;
	wire [15-1:0] node1365;
	wire [15-1:0] node1366;
	wire [15-1:0] node1367;
	wire [15-1:0] node1368;
	wire [15-1:0] node1373;
	wire [15-1:0] node1376;
	wire [15-1:0] node1379;
	wire [15-1:0] node1380;
	wire [15-1:0] node1381;
	wire [15-1:0] node1382;
	wire [15-1:0] node1385;
	wire [15-1:0] node1388;
	wire [15-1:0] node1389;
	wire [15-1:0] node1390;
	wire [15-1:0] node1392;
	wire [15-1:0] node1393;
	wire [15-1:0] node1398;
	wire [15-1:0] node1400;
	wire [15-1:0] node1401;
	wire [15-1:0] node1405;
	wire [15-1:0] node1406;
	wire [15-1:0] node1408;
	wire [15-1:0] node1409;
	wire [15-1:0] node1412;
	wire [15-1:0] node1413;
	wire [15-1:0] node1415;
	wire [15-1:0] node1419;
	wire [15-1:0] node1420;
	wire [15-1:0] node1421;
	wire [15-1:0] node1424;
	wire [15-1:0] node1426;
	wire [15-1:0] node1429;
	wire [15-1:0] node1430;
	wire [15-1:0] node1434;
	wire [15-1:0] node1435;
	wire [15-1:0] node1436;
	wire [15-1:0] node1437;
	wire [15-1:0] node1438;
	wire [15-1:0] node1441;
	wire [15-1:0] node1442;
	wire [15-1:0] node1444;
	wire [15-1:0] node1448;
	wire [15-1:0] node1449;
	wire [15-1:0] node1450;
	wire [15-1:0] node1451;
	wire [15-1:0] node1455;
	wire [15-1:0] node1458;
	wire [15-1:0] node1459;
	wire [15-1:0] node1460;
	wire [15-1:0] node1462;
	wire [15-1:0] node1466;
	wire [15-1:0] node1467;
	wire [15-1:0] node1471;
	wire [15-1:0] node1472;
	wire [15-1:0] node1473;
	wire [15-1:0] node1474;
	wire [15-1:0] node1475;
	wire [15-1:0] node1479;
	wire [15-1:0] node1481;
	wire [15-1:0] node1484;
	wire [15-1:0] node1485;
	wire [15-1:0] node1486;
	wire [15-1:0] node1491;
	wire [15-1:0] node1492;
	wire [15-1:0] node1493;
	wire [15-1:0] node1494;
	wire [15-1:0] node1496;
	wire [15-1:0] node1500;
	wire [15-1:0] node1503;
	wire [15-1:0] node1504;
	wire [15-1:0] node1505;
	wire [15-1:0] node1507;
	wire [15-1:0] node1511;
	wire [15-1:0] node1514;
	wire [15-1:0] node1515;
	wire [15-1:0] node1516;
	wire [15-1:0] node1517;
	wire [15-1:0] node1518;
	wire [15-1:0] node1521;
	wire [15-1:0] node1525;
	wire [15-1:0] node1526;
	wire [15-1:0] node1527;
	wire [15-1:0] node1530;
	wire [15-1:0] node1532;
	wire [15-1:0] node1535;
	wire [15-1:0] node1536;
	wire [15-1:0] node1537;
	wire [15-1:0] node1542;
	wire [15-1:0] node1543;
	wire [15-1:0] node1544;
	wire [15-1:0] node1545;
	wire [15-1:0] node1548;
	wire [15-1:0] node1550;
	wire [15-1:0] node1553;
	wire [15-1:0] node1554;
	wire [15-1:0] node1555;
	wire [15-1:0] node1559;
	wire [15-1:0] node1560;
	wire [15-1:0] node1564;
	wire [15-1:0] node1565;
	wire [15-1:0] node1566;
	wire [15-1:0] node1567;
	wire [15-1:0] node1570;
	wire [15-1:0] node1572;
	wire [15-1:0] node1575;
	wire [15-1:0] node1578;
	wire [15-1:0] node1579;
	wire [15-1:0] node1580;
	wire [15-1:0] node1584;
	wire [15-1:0] node1585;
	wire [15-1:0] node1589;
	wire [15-1:0] node1590;
	wire [15-1:0] node1591;
	wire [15-1:0] node1592;
	wire [15-1:0] node1593;
	wire [15-1:0] node1594;
	wire [15-1:0] node1595;
	wire [15-1:0] node1596;
	wire [15-1:0] node1597;
	wire [15-1:0] node1602;
	wire [15-1:0] node1603;
	wire [15-1:0] node1605;
	wire [15-1:0] node1606;
	wire [15-1:0] node1611;
	wire [15-1:0] node1612;
	wire [15-1:0] node1613;
	wire [15-1:0] node1616;
	wire [15-1:0] node1619;
	wire [15-1:0] node1620;
	wire [15-1:0] node1623;
	wire [15-1:0] node1624;
	wire [15-1:0] node1626;
	wire [15-1:0] node1630;
	wire [15-1:0] node1631;
	wire [15-1:0] node1632;
	wire [15-1:0] node1634;
	wire [15-1:0] node1637;
	wire [15-1:0] node1638;
	wire [15-1:0] node1641;
	wire [15-1:0] node1644;
	wire [15-1:0] node1645;
	wire [15-1:0] node1647;
	wire [15-1:0] node1649;
	wire [15-1:0] node1650;
	wire [15-1:0] node1655;
	wire [15-1:0] node1656;
	wire [15-1:0] node1657;
	wire [15-1:0] node1658;
	wire [15-1:0] node1659;
	wire [15-1:0] node1661;
	wire [15-1:0] node1665;
	wire [15-1:0] node1666;
	wire [15-1:0] node1670;
	wire [15-1:0] node1671;
	wire [15-1:0] node1673;
	wire [15-1:0] node1676;
	wire [15-1:0] node1677;
	wire [15-1:0] node1681;
	wire [15-1:0] node1682;
	wire [15-1:0] node1683;
	wire [15-1:0] node1684;
	wire [15-1:0] node1687;
	wire [15-1:0] node1690;
	wire [15-1:0] node1692;
	wire [15-1:0] node1693;
	wire [15-1:0] node1695;
	wire [15-1:0] node1699;
	wire [15-1:0] node1700;
	wire [15-1:0] node1701;
	wire [15-1:0] node1704;
	wire [15-1:0] node1705;
	wire [15-1:0] node1707;
	wire [15-1:0] node1711;
	wire [15-1:0] node1712;
	wire [15-1:0] node1713;
	wire [15-1:0] node1715;
	wire [15-1:0] node1720;
	wire [15-1:0] node1721;
	wire [15-1:0] node1722;
	wire [15-1:0] node1723;
	wire [15-1:0] node1724;
	wire [15-1:0] node1725;
	wire [15-1:0] node1727;
	wire [15-1:0] node1728;
	wire [15-1:0] node1732;
	wire [15-1:0] node1735;
	wire [15-1:0] node1736;
	wire [15-1:0] node1740;
	wire [15-1:0] node1741;
	wire [15-1:0] node1742;
	wire [15-1:0] node1743;
	wire [15-1:0] node1747;
	wire [15-1:0] node1750;
	wire [15-1:0] node1753;
	wire [15-1:0] node1754;
	wire [15-1:0] node1755;
	wire [15-1:0] node1758;
	wire [15-1:0] node1759;
	wire [15-1:0] node1763;
	wire [15-1:0] node1764;
	wire [15-1:0] node1765;
	wire [15-1:0] node1768;
	wire [15-1:0] node1769;
	wire [15-1:0] node1773;
	wire [15-1:0] node1775;
	wire [15-1:0] node1778;
	wire [15-1:0] node1779;
	wire [15-1:0] node1780;
	wire [15-1:0] node1781;
	wire [15-1:0] node1782;
	wire [15-1:0] node1783;
	wire [15-1:0] node1788;
	wire [15-1:0] node1789;
	wire [15-1:0] node1793;
	wire [15-1:0] node1794;
	wire [15-1:0] node1795;
	wire [15-1:0] node1798;
	wire [15-1:0] node1801;
	wire [15-1:0] node1802;
	wire [15-1:0] node1806;
	wire [15-1:0] node1807;
	wire [15-1:0] node1809;
	wire [15-1:0] node1811;
	wire [15-1:0] node1812;
	wire [15-1:0] node1816;
	wire [15-1:0] node1817;
	wire [15-1:0] node1819;
	wire [15-1:0] node1820;
	wire [15-1:0] node1824;
	wire [15-1:0] node1826;
	wire [15-1:0] node1827;
	wire [15-1:0] node1829;
	wire [15-1:0] node1833;
	wire [15-1:0] node1834;
	wire [15-1:0] node1835;
	wire [15-1:0] node1836;
	wire [15-1:0] node1837;
	wire [15-1:0] node1838;
	wire [15-1:0] node1839;
	wire [15-1:0] node1840;
	wire [15-1:0] node1845;
	wire [15-1:0] node1847;
	wire [15-1:0] node1848;
	wire [15-1:0] node1852;
	wire [15-1:0] node1853;
	wire [15-1:0] node1854;
	wire [15-1:0] node1858;
	wire [15-1:0] node1859;
	wire [15-1:0] node1861;
	wire [15-1:0] node1864;
	wire [15-1:0] node1865;
	wire [15-1:0] node1866;
	wire [15-1:0] node1870;
	wire [15-1:0] node1873;
	wire [15-1:0] node1874;
	wire [15-1:0] node1875;
	wire [15-1:0] node1876;
	wire [15-1:0] node1878;
	wire [15-1:0] node1882;
	wire [15-1:0] node1883;
	wire [15-1:0] node1887;
	wire [15-1:0] node1888;
	wire [15-1:0] node1890;
	wire [15-1:0] node1893;
	wire [15-1:0] node1895;
	wire [15-1:0] node1898;
	wire [15-1:0] node1899;
	wire [15-1:0] node1900;
	wire [15-1:0] node1901;
	wire [15-1:0] node1902;
	wire [15-1:0] node1906;
	wire [15-1:0] node1907;
	wire [15-1:0] node1909;
	wire [15-1:0] node1912;
	wire [15-1:0] node1915;
	wire [15-1:0] node1916;
	wire [15-1:0] node1917;
	wire [15-1:0] node1920;
	wire [15-1:0] node1921;
	wire [15-1:0] node1923;
	wire [15-1:0] node1927;
	wire [15-1:0] node1929;
	wire [15-1:0] node1932;
	wire [15-1:0] node1933;
	wire [15-1:0] node1934;
	wire [15-1:0] node1935;
	wire [15-1:0] node1939;
	wire [15-1:0] node1940;
	wire [15-1:0] node1944;
	wire [15-1:0] node1945;
	wire [15-1:0] node1946;
	wire [15-1:0] node1950;
	wire [15-1:0] node1953;
	wire [15-1:0] node1954;
	wire [15-1:0] node1955;
	wire [15-1:0] node1956;
	wire [15-1:0] node1957;
	wire [15-1:0] node1958;
	wire [15-1:0] node1962;
	wire [15-1:0] node1963;
	wire [15-1:0] node1965;
	wire [15-1:0] node1969;
	wire [15-1:0] node1970;
	wire [15-1:0] node1971;
	wire [15-1:0] node1973;
	wire [15-1:0] node1976;
	wire [15-1:0] node1979;
	wire [15-1:0] node1980;
	wire [15-1:0] node1983;
	wire [15-1:0] node1985;
	wire [15-1:0] node1988;
	wire [15-1:0] node1989;
	wire [15-1:0] node1990;
	wire [15-1:0] node1992;
	wire [15-1:0] node1994;
	wire [15-1:0] node1997;
	wire [15-1:0] node1998;
	wire [15-1:0] node2000;
	wire [15-1:0] node2003;
	wire [15-1:0] node2005;
	wire [15-1:0] node2008;
	wire [15-1:0] node2009;
	wire [15-1:0] node2010;
	wire [15-1:0] node2011;
	wire [15-1:0] node2015;
	wire [15-1:0] node2018;
	wire [15-1:0] node2020;
	wire [15-1:0] node2021;
	wire [15-1:0] node2023;
	wire [15-1:0] node2026;
	wire [15-1:0] node2029;
	wire [15-1:0] node2030;
	wire [15-1:0] node2031;
	wire [15-1:0] node2032;
	wire [15-1:0] node2033;
	wire [15-1:0] node2037;
	wire [15-1:0] node2039;
	wire [15-1:0] node2042;
	wire [15-1:0] node2043;
	wire [15-1:0] node2045;
	wire [15-1:0] node2046;
	wire [15-1:0] node2050;
	wire [15-1:0] node2051;
	wire [15-1:0] node2052;
	wire [15-1:0] node2057;
	wire [15-1:0] node2058;
	wire [15-1:0] node2059;
	wire [15-1:0] node2061;
	wire [15-1:0] node2062;
	wire [15-1:0] node2066;
	wire [15-1:0] node2067;
	wire [15-1:0] node2068;
	wire [15-1:0] node2072;
	wire [15-1:0] node2073;
	wire [15-1:0] node2075;
	wire [15-1:0] node2079;
	wire [15-1:0] node2080;
	wire [15-1:0] node2081;
	wire [15-1:0] node2084;
	wire [15-1:0] node2087;
	wire [15-1:0] node2089;
	wire [15-1:0] node2090;
	wire [15-1:0] node2092;
	wire [15-1:0] node2095;
	wire [15-1:0] node2098;
	wire [15-1:0] node2099;
	wire [15-1:0] node2100;
	wire [15-1:0] node2101;
	wire [15-1:0] node2102;
	wire [15-1:0] node2103;
	wire [15-1:0] node2104;
	wire [15-1:0] node2105;
	wire [15-1:0] node2106;
	wire [15-1:0] node2108;
	wire [15-1:0] node2111;
	wire [15-1:0] node2112;
	wire [15-1:0] node2114;
	wire [15-1:0] node2117;
	wire [15-1:0] node2119;
	wire [15-1:0] node2122;
	wire [15-1:0] node2123;
	wire [15-1:0] node2124;
	wire [15-1:0] node2127;
	wire [15-1:0] node2130;
	wire [15-1:0] node2131;
	wire [15-1:0] node2133;
	wire [15-1:0] node2137;
	wire [15-1:0] node2138;
	wire [15-1:0] node2139;
	wire [15-1:0] node2140;
	wire [15-1:0] node2143;
	wire [15-1:0] node2146;
	wire [15-1:0] node2147;
	wire [15-1:0] node2150;
	wire [15-1:0] node2152;
	wire [15-1:0] node2155;
	wire [15-1:0] node2156;
	wire [15-1:0] node2157;
	wire [15-1:0] node2158;
	wire [15-1:0] node2163;
	wire [15-1:0] node2164;
	wire [15-1:0] node2165;
	wire [15-1:0] node2169;
	wire [15-1:0] node2172;
	wire [15-1:0] node2173;
	wire [15-1:0] node2174;
	wire [15-1:0] node2175;
	wire [15-1:0] node2176;
	wire [15-1:0] node2178;
	wire [15-1:0] node2182;
	wire [15-1:0] node2183;
	wire [15-1:0] node2185;
	wire [15-1:0] node2188;
	wire [15-1:0] node2191;
	wire [15-1:0] node2192;
	wire [15-1:0] node2193;
	wire [15-1:0] node2196;
	wire [15-1:0] node2197;
	wire [15-1:0] node2199;
	wire [15-1:0] node2203;
	wire [15-1:0] node2204;
	wire [15-1:0] node2205;
	wire [15-1:0] node2210;
	wire [15-1:0] node2211;
	wire [15-1:0] node2212;
	wire [15-1:0] node2215;
	wire [15-1:0] node2216;
	wire [15-1:0] node2217;
	wire [15-1:0] node2219;
	wire [15-1:0] node2223;
	wire [15-1:0] node2224;
	wire [15-1:0] node2228;
	wire [15-1:0] node2229;
	wire [15-1:0] node2230;
	wire [15-1:0] node2232;
	wire [15-1:0] node2235;
	wire [15-1:0] node2238;
	wire [15-1:0] node2239;
	wire [15-1:0] node2240;
	wire [15-1:0] node2244;
	wire [15-1:0] node2247;
	wire [15-1:0] node2248;
	wire [15-1:0] node2249;
	wire [15-1:0] node2250;
	wire [15-1:0] node2251;
	wire [15-1:0] node2254;
	wire [15-1:0] node2255;
	wire [15-1:0] node2256;
	wire [15-1:0] node2259;
	wire [15-1:0] node2260;
	wire [15-1:0] node2264;
	wire [15-1:0] node2266;
	wire [15-1:0] node2269;
	wire [15-1:0] node2270;
	wire [15-1:0] node2271;
	wire [15-1:0] node2275;
	wire [15-1:0] node2276;
	wire [15-1:0] node2277;
	wire [15-1:0] node2279;
	wire [15-1:0] node2283;
	wire [15-1:0] node2286;
	wire [15-1:0] node2287;
	wire [15-1:0] node2288;
	wire [15-1:0] node2290;
	wire [15-1:0] node2291;
	wire [15-1:0] node2293;
	wire [15-1:0] node2296;
	wire [15-1:0] node2300;
	wire [15-1:0] node2301;
	wire [15-1:0] node2303;
	wire [15-1:0] node2305;
	wire [15-1:0] node2308;
	wire [15-1:0] node2309;
	wire [15-1:0] node2310;
	wire [15-1:0] node2315;
	wire [15-1:0] node2316;
	wire [15-1:0] node2317;
	wire [15-1:0] node2318;
	wire [15-1:0] node2320;
	wire [15-1:0] node2321;
	wire [15-1:0] node2325;
	wire [15-1:0] node2326;
	wire [15-1:0] node2329;
	wire [15-1:0] node2332;
	wire [15-1:0] node2333;
	wire [15-1:0] node2335;
	wire [15-1:0] node2336;
	wire [15-1:0] node2340;
	wire [15-1:0] node2341;
	wire [15-1:0] node2344;
	wire [15-1:0] node2345;
	wire [15-1:0] node2348;
	wire [15-1:0] node2351;
	wire [15-1:0] node2352;
	wire [15-1:0] node2354;
	wire [15-1:0] node2355;
	wire [15-1:0] node2359;
	wire [15-1:0] node2360;
	wire [15-1:0] node2362;
	wire [15-1:0] node2364;
	wire [15-1:0] node2365;
	wire [15-1:0] node2369;
	wire [15-1:0] node2372;
	wire [15-1:0] node2373;
	wire [15-1:0] node2374;
	wire [15-1:0] node2375;
	wire [15-1:0] node2376;
	wire [15-1:0] node2377;
	wire [15-1:0] node2380;
	wire [15-1:0] node2381;
	wire [15-1:0] node2384;
	wire [15-1:0] node2387;
	wire [15-1:0] node2389;
	wire [15-1:0] node2390;
	wire [15-1:0] node2394;
	wire [15-1:0] node2395;
	wire [15-1:0] node2396;
	wire [15-1:0] node2397;
	wire [15-1:0] node2398;
	wire [15-1:0] node2402;
	wire [15-1:0] node2404;
	wire [15-1:0] node2407;
	wire [15-1:0] node2408;
	wire [15-1:0] node2409;
	wire [15-1:0] node2411;
	wire [15-1:0] node2416;
	wire [15-1:0] node2417;
	wire [15-1:0] node2419;
	wire [15-1:0] node2422;
	wire [15-1:0] node2423;
	wire [15-1:0] node2426;
	wire [15-1:0] node2427;
	wire [15-1:0] node2429;
	wire [15-1:0] node2433;
	wire [15-1:0] node2434;
	wire [15-1:0] node2435;
	wire [15-1:0] node2436;
	wire [15-1:0] node2437;
	wire [15-1:0] node2438;
	wire [15-1:0] node2440;
	wire [15-1:0] node2445;
	wire [15-1:0] node2446;
	wire [15-1:0] node2447;
	wire [15-1:0] node2452;
	wire [15-1:0] node2453;
	wire [15-1:0] node2455;
	wire [15-1:0] node2458;
	wire [15-1:0] node2459;
	wire [15-1:0] node2462;
	wire [15-1:0] node2465;
	wire [15-1:0] node2466;
	wire [15-1:0] node2467;
	wire [15-1:0] node2469;
	wire [15-1:0] node2470;
	wire [15-1:0] node2474;
	wire [15-1:0] node2475;
	wire [15-1:0] node2478;
	wire [15-1:0] node2480;
	wire [15-1:0] node2483;
	wire [15-1:0] node2484;
	wire [15-1:0] node2485;
	wire [15-1:0] node2488;
	wire [15-1:0] node2490;
	wire [15-1:0] node2493;
	wire [15-1:0] node2494;
	wire [15-1:0] node2495;
	wire [15-1:0] node2500;
	wire [15-1:0] node2501;
	wire [15-1:0] node2502;
	wire [15-1:0] node2503;
	wire [15-1:0] node2504;
	wire [15-1:0] node2506;
	wire [15-1:0] node2507;
	wire [15-1:0] node2511;
	wire [15-1:0] node2513;
	wire [15-1:0] node2514;
	wire [15-1:0] node2515;
	wire [15-1:0] node2520;
	wire [15-1:0] node2521;
	wire [15-1:0] node2522;
	wire [15-1:0] node2523;
	wire [15-1:0] node2528;
	wire [15-1:0] node2529;
	wire [15-1:0] node2533;
	wire [15-1:0] node2534;
	wire [15-1:0] node2535;
	wire [15-1:0] node2536;
	wire [15-1:0] node2538;
	wire [15-1:0] node2542;
	wire [15-1:0] node2543;
	wire [15-1:0] node2544;
	wire [15-1:0] node2546;
	wire [15-1:0] node2550;
	wire [15-1:0] node2553;
	wire [15-1:0] node2554;
	wire [15-1:0] node2555;
	wire [15-1:0] node2556;
	wire [15-1:0] node2560;
	wire [15-1:0] node2561;
	wire [15-1:0] node2563;
	wire [15-1:0] node2567;
	wire [15-1:0] node2568;
	wire [15-1:0] node2571;
	wire [15-1:0] node2574;
	wire [15-1:0] node2575;
	wire [15-1:0] node2576;
	wire [15-1:0] node2577;
	wire [15-1:0] node2578;
	wire [15-1:0] node2581;
	wire [15-1:0] node2584;
	wire [15-1:0] node2585;
	wire [15-1:0] node2586;
	wire [15-1:0] node2588;
	wire [15-1:0] node2593;
	wire [15-1:0] node2594;
	wire [15-1:0] node2595;
	wire [15-1:0] node2598;
	wire [15-1:0] node2600;
	wire [15-1:0] node2601;
	wire [15-1:0] node2605;
	wire [15-1:0] node2606;
	wire [15-1:0] node2609;
	wire [15-1:0] node2611;
	wire [15-1:0] node2614;
	wire [15-1:0] node2615;
	wire [15-1:0] node2616;
	wire [15-1:0] node2618;
	wire [15-1:0] node2619;
	wire [15-1:0] node2620;
	wire [15-1:0] node2625;
	wire [15-1:0] node2626;
	wire [15-1:0] node2629;
	wire [15-1:0] node2631;
	wire [15-1:0] node2633;
	wire [15-1:0] node2636;
	wire [15-1:0] node2638;
	wire [15-1:0] node2639;
	wire [15-1:0] node2641;
	wire [15-1:0] node2642;
	wire [15-1:0] node2646;
	wire [15-1:0] node2649;
	wire [15-1:0] node2650;
	wire [15-1:0] node2651;
	wire [15-1:0] node2652;
	wire [15-1:0] node2653;
	wire [15-1:0] node2654;
	wire [15-1:0] node2655;
	wire [15-1:0] node2656;
	wire [15-1:0] node2659;
	wire [15-1:0] node2662;
	wire [15-1:0] node2663;
	wire [15-1:0] node2667;
	wire [15-1:0] node2668;
	wire [15-1:0] node2670;
	wire [15-1:0] node2673;
	wire [15-1:0] node2674;
	wire [15-1:0] node2675;
	wire [15-1:0] node2680;
	wire [15-1:0] node2681;
	wire [15-1:0] node2682;
	wire [15-1:0] node2683;
	wire [15-1:0] node2687;
	wire [15-1:0] node2689;
	wire [15-1:0] node2692;
	wire [15-1:0] node2693;
	wire [15-1:0] node2695;
	wire [15-1:0] node2698;
	wire [15-1:0] node2699;
	wire [15-1:0] node2703;
	wire [15-1:0] node2704;
	wire [15-1:0] node2705;
	wire [15-1:0] node2706;
	wire [15-1:0] node2707;
	wire [15-1:0] node2709;
	wire [15-1:0] node2712;
	wire [15-1:0] node2713;
	wire [15-1:0] node2715;
	wire [15-1:0] node2719;
	wire [15-1:0] node2720;
	wire [15-1:0] node2723;
	wire [15-1:0] node2726;
	wire [15-1:0] node2727;
	wire [15-1:0] node2728;
	wire [15-1:0] node2729;
	wire [15-1:0] node2733;
	wire [15-1:0] node2736;
	wire [15-1:0] node2738;
	wire [15-1:0] node2739;
	wire [15-1:0] node2742;
	wire [15-1:0] node2743;
	wire [15-1:0] node2747;
	wire [15-1:0] node2748;
	wire [15-1:0] node2749;
	wire [15-1:0] node2750;
	wire [15-1:0] node2753;
	wire [15-1:0] node2755;
	wire [15-1:0] node2759;
	wire [15-1:0] node2760;
	wire [15-1:0] node2761;
	wire [15-1:0] node2762;
	wire [15-1:0] node2766;
	wire [15-1:0] node2767;
	wire [15-1:0] node2769;
	wire [15-1:0] node2773;
	wire [15-1:0] node2776;
	wire [15-1:0] node2777;
	wire [15-1:0] node2778;
	wire [15-1:0] node2779;
	wire [15-1:0] node2780;
	wire [15-1:0] node2781;
	wire [15-1:0] node2782;
	wire [15-1:0] node2787;
	wire [15-1:0] node2789;
	wire [15-1:0] node2792;
	wire [15-1:0] node2794;
	wire [15-1:0] node2795;
	wire [15-1:0] node2797;
	wire [15-1:0] node2798;
	wire [15-1:0] node2802;
	wire [15-1:0] node2804;
	wire [15-1:0] node2807;
	wire [15-1:0] node2808;
	wire [15-1:0] node2809;
	wire [15-1:0] node2810;
	wire [15-1:0] node2814;
	wire [15-1:0] node2815;
	wire [15-1:0] node2818;
	wire [15-1:0] node2820;
	wire [15-1:0] node2823;
	wire [15-1:0] node2824;
	wire [15-1:0] node2827;
	wire [15-1:0] node2829;
	wire [15-1:0] node2831;
	wire [15-1:0] node2832;
	wire [15-1:0] node2836;
	wire [15-1:0] node2837;
	wire [15-1:0] node2838;
	wire [15-1:0] node2839;
	wire [15-1:0] node2841;
	wire [15-1:0] node2843;
	wire [15-1:0] node2844;
	wire [15-1:0] node2848;
	wire [15-1:0] node2849;
	wire [15-1:0] node2852;
	wire [15-1:0] node2853;
	wire [15-1:0] node2857;
	wire [15-1:0] node2858;
	wire [15-1:0] node2859;
	wire [15-1:0] node2862;
	wire [15-1:0] node2864;
	wire [15-1:0] node2867;
	wire [15-1:0] node2868;
	wire [15-1:0] node2871;
	wire [15-1:0] node2874;
	wire [15-1:0] node2875;
	wire [15-1:0] node2877;
	wire [15-1:0] node2878;
	wire [15-1:0] node2882;
	wire [15-1:0] node2883;
	wire [15-1:0] node2885;
	wire [15-1:0] node2886;
	wire [15-1:0] node2890;
	wire [15-1:0] node2891;
	wire [15-1:0] node2894;
	wire [15-1:0] node2897;
	wire [15-1:0] node2898;
	wire [15-1:0] node2899;
	wire [15-1:0] node2900;
	wire [15-1:0] node2901;
	wire [15-1:0] node2902;
	wire [15-1:0] node2903;
	wire [15-1:0] node2907;
	wire [15-1:0] node2908;
	wire [15-1:0] node2911;
	wire [15-1:0] node2914;
	wire [15-1:0] node2916;
	wire [15-1:0] node2917;
	wire [15-1:0] node2921;
	wire [15-1:0] node2922;
	wire [15-1:0] node2923;
	wire [15-1:0] node2924;
	wire [15-1:0] node2927;
	wire [15-1:0] node2929;
	wire [15-1:0] node2930;
	wire [15-1:0] node2934;
	wire [15-1:0] node2935;
	wire [15-1:0] node2938;
	wire [15-1:0] node2941;
	wire [15-1:0] node2942;
	wire [15-1:0] node2944;
	wire [15-1:0] node2945;
	wire [15-1:0] node2949;
	wire [15-1:0] node2951;
	wire [15-1:0] node2954;
	wire [15-1:0] node2955;
	wire [15-1:0] node2956;
	wire [15-1:0] node2957;
	wire [15-1:0] node2959;
	wire [15-1:0] node2960;
	wire [15-1:0] node2964;
	wire [15-1:0] node2965;
	wire [15-1:0] node2969;
	wire [15-1:0] node2970;
	wire [15-1:0] node2971;
	wire [15-1:0] node2973;
	wire [15-1:0] node2975;
	wire [15-1:0] node2979;
	wire [15-1:0] node2980;
	wire [15-1:0] node2982;
	wire [15-1:0] node2983;
	wire [15-1:0] node2988;
	wire [15-1:0] node2989;
	wire [15-1:0] node2990;
	wire [15-1:0] node2992;
	wire [15-1:0] node2993;
	wire [15-1:0] node2995;
	wire [15-1:0] node2998;
	wire [15-1:0] node3001;
	wire [15-1:0] node3002;
	wire [15-1:0] node3003;
	wire [15-1:0] node3008;
	wire [15-1:0] node3010;
	wire [15-1:0] node3011;
	wire [15-1:0] node3012;
	wire [15-1:0] node3017;
	wire [15-1:0] node3018;
	wire [15-1:0] node3019;
	wire [15-1:0] node3020;
	wire [15-1:0] node3021;
	wire [15-1:0] node3024;
	wire [15-1:0] node3027;
	wire [15-1:0] node3028;
	wire [15-1:0] node3029;
	wire [15-1:0] node3030;
	wire [15-1:0] node3034;
	wire [15-1:0] node3036;
	wire [15-1:0] node3040;
	wire [15-1:0] node3041;
	wire [15-1:0] node3042;
	wire [15-1:0] node3043;
	wire [15-1:0] node3046;
	wire [15-1:0] node3048;
	wire [15-1:0] node3049;
	wire [15-1:0] node3053;
	wire [15-1:0] node3054;
	wire [15-1:0] node3058;
	wire [15-1:0] node3060;
	wire [15-1:0] node3061;
	wire [15-1:0] node3064;
	wire [15-1:0] node3067;
	wire [15-1:0] node3068;
	wire [15-1:0] node3069;
	wire [15-1:0] node3070;
	wire [15-1:0] node3071;
	wire [15-1:0] node3075;
	wire [15-1:0] node3077;
	wire [15-1:0] node3078;
	wire [15-1:0] node3079;
	wire [15-1:0] node3084;
	wire [15-1:0] node3085;
	wire [15-1:0] node3087;
	wire [15-1:0] node3088;
	wire [15-1:0] node3089;
	wire [15-1:0] node3094;
	wire [15-1:0] node3095;
	wire [15-1:0] node3098;
	wire [15-1:0] node3101;
	wire [15-1:0] node3102;
	wire [15-1:0] node3103;
	wire [15-1:0] node3104;
	wire [15-1:0] node3107;
	wire [15-1:0] node3110;
	wire [15-1:0] node3111;
	wire [15-1:0] node3112;
	wire [15-1:0] node3115;
	wire [15-1:0] node3117;
	wire [15-1:0] node3120;
	wire [15-1:0] node3122;
	wire [15-1:0] node3124;
	wire [15-1:0] node3127;
	wire [15-1:0] node3128;
	wire [15-1:0] node3131;
	wire [15-1:0] node3133;
	wire [15-1:0] node3135;
	wire [15-1:0] node3138;
	wire [15-1:0] node3139;
	wire [15-1:0] node3140;
	wire [15-1:0] node3141;
	wire [15-1:0] node3142;
	wire [15-1:0] node3143;
	wire [15-1:0] node3144;
	wire [15-1:0] node3145;
	wire [15-1:0] node3146;
	wire [15-1:0] node3147;
	wire [15-1:0] node3152;
	wire [15-1:0] node3153;
	wire [15-1:0] node3154;
	wire [15-1:0] node3158;
	wire [15-1:0] node3159;
	wire [15-1:0] node3163;
	wire [15-1:0] node3164;
	wire [15-1:0] node3165;
	wire [15-1:0] node3169;
	wire [15-1:0] node3170;
	wire [15-1:0] node3174;
	wire [15-1:0] node3175;
	wire [15-1:0] node3176;
	wire [15-1:0] node3178;
	wire [15-1:0] node3181;
	wire [15-1:0] node3184;
	wire [15-1:0] node3185;
	wire [15-1:0] node3187;
	wire [15-1:0] node3190;
	wire [15-1:0] node3191;
	wire [15-1:0] node3194;
	wire [15-1:0] node3197;
	wire [15-1:0] node3198;
	wire [15-1:0] node3199;
	wire [15-1:0] node3200;
	wire [15-1:0] node3201;
	wire [15-1:0] node3205;
	wire [15-1:0] node3208;
	wire [15-1:0] node3209;
	wire [15-1:0] node3210;
	wire [15-1:0] node3211;
	wire [15-1:0] node3216;
	wire [15-1:0] node3217;
	wire [15-1:0] node3219;
	wire [15-1:0] node3223;
	wire [15-1:0] node3224;
	wire [15-1:0] node3225;
	wire [15-1:0] node3226;
	wire [15-1:0] node3228;
	wire [15-1:0] node3231;
	wire [15-1:0] node3233;
	wire [15-1:0] node3236;
	wire [15-1:0] node3237;
	wire [15-1:0] node3239;
	wire [15-1:0] node3240;
	wire [15-1:0] node3244;
	wire [15-1:0] node3247;
	wire [15-1:0] node3248;
	wire [15-1:0] node3250;
	wire [15-1:0] node3251;
	wire [15-1:0] node3255;
	wire [15-1:0] node3257;
	wire [15-1:0] node3260;
	wire [15-1:0] node3261;
	wire [15-1:0] node3262;
	wire [15-1:0] node3263;
	wire [15-1:0] node3264;
	wire [15-1:0] node3265;
	wire [15-1:0] node3269;
	wire [15-1:0] node3271;
	wire [15-1:0] node3274;
	wire [15-1:0] node3275;
	wire [15-1:0] node3276;
	wire [15-1:0] node3279;
	wire [15-1:0] node3281;
	wire [15-1:0] node3282;
	wire [15-1:0] node3287;
	wire [15-1:0] node3288;
	wire [15-1:0] node3289;
	wire [15-1:0] node3291;
	wire [15-1:0] node3294;
	wire [15-1:0] node3296;
	wire [15-1:0] node3297;
	wire [15-1:0] node3301;
	wire [15-1:0] node3302;
	wire [15-1:0] node3303;
	wire [15-1:0] node3305;
	wire [15-1:0] node3310;
	wire [15-1:0] node3311;
	wire [15-1:0] node3312;
	wire [15-1:0] node3313;
	wire [15-1:0] node3314;
	wire [15-1:0] node3317;
	wire [15-1:0] node3320;
	wire [15-1:0] node3321;
	wire [15-1:0] node3325;
	wire [15-1:0] node3326;
	wire [15-1:0] node3328;
	wire [15-1:0] node3330;
	wire [15-1:0] node3331;
	wire [15-1:0] node3335;
	wire [15-1:0] node3336;
	wire [15-1:0] node3340;
	wire [15-1:0] node3341;
	wire [15-1:0] node3342;
	wire [15-1:0] node3344;
	wire [15-1:0] node3348;
	wire [15-1:0] node3349;
	wire [15-1:0] node3350;
	wire [15-1:0] node3351;
	wire [15-1:0] node3356;
	wire [15-1:0] node3357;
	wire [15-1:0] node3358;
	wire [15-1:0] node3362;
	wire [15-1:0] node3363;
	wire [15-1:0] node3367;
	wire [15-1:0] node3368;
	wire [15-1:0] node3369;
	wire [15-1:0] node3370;
	wire [15-1:0] node3371;
	wire [15-1:0] node3372;
	wire [15-1:0] node3373;
	wire [15-1:0] node3377;
	wire [15-1:0] node3379;
	wire [15-1:0] node3380;
	wire [15-1:0] node3384;
	wire [15-1:0] node3385;
	wire [15-1:0] node3386;
	wire [15-1:0] node3388;
	wire [15-1:0] node3389;
	wire [15-1:0] node3393;
	wire [15-1:0] node3395;
	wire [15-1:0] node3398;
	wire [15-1:0] node3399;
	wire [15-1:0] node3402;
	wire [15-1:0] node3404;
	wire [15-1:0] node3407;
	wire [15-1:0] node3408;
	wire [15-1:0] node3409;
	wire [15-1:0] node3410;
	wire [15-1:0] node3413;
	wire [15-1:0] node3414;
	wire [15-1:0] node3416;
	wire [15-1:0] node3420;
	wire [15-1:0] node3421;
	wire [15-1:0] node3424;
	wire [15-1:0] node3427;
	wire [15-1:0] node3428;
	wire [15-1:0] node3429;
	wire [15-1:0] node3431;
	wire [15-1:0] node3432;
	wire [15-1:0] node3436;
	wire [15-1:0] node3438;
	wire [15-1:0] node3441;
	wire [15-1:0] node3442;
	wire [15-1:0] node3444;
	wire [15-1:0] node3446;
	wire [15-1:0] node3450;
	wire [15-1:0] node3451;
	wire [15-1:0] node3452;
	wire [15-1:0] node3453;
	wire [15-1:0] node3455;
	wire [15-1:0] node3458;
	wire [15-1:0] node3459;
	wire [15-1:0] node3460;
	wire [15-1:0] node3465;
	wire [15-1:0] node3466;
	wire [15-1:0] node3467;
	wire [15-1:0] node3470;
	wire [15-1:0] node3473;
	wire [15-1:0] node3474;
	wire [15-1:0] node3477;
	wire [15-1:0] node3480;
	wire [15-1:0] node3481;
	wire [15-1:0] node3482;
	wire [15-1:0] node3484;
	wire [15-1:0] node3486;
	wire [15-1:0] node3487;
	wire [15-1:0] node3491;
	wire [15-1:0] node3492;
	wire [15-1:0] node3493;
	wire [15-1:0] node3497;
	wire [15-1:0] node3499;
	wire [15-1:0] node3502;
	wire [15-1:0] node3503;
	wire [15-1:0] node3504;
	wire [15-1:0] node3508;
	wire [15-1:0] node3511;
	wire [15-1:0] node3512;
	wire [15-1:0] node3513;
	wire [15-1:0] node3514;
	wire [15-1:0] node3515;
	wire [15-1:0] node3516;
	wire [15-1:0] node3517;
	wire [15-1:0] node3521;
	wire [15-1:0] node3524;
	wire [15-1:0] node3526;
	wire [15-1:0] node3528;
	wire [15-1:0] node3531;
	wire [15-1:0] node3532;
	wire [15-1:0] node3535;
	wire [15-1:0] node3536;
	wire [15-1:0] node3537;
	wire [15-1:0] node3539;
	wire [15-1:0] node3544;
	wire [15-1:0] node3545;
	wire [15-1:0] node3546;
	wire [15-1:0] node3549;
	wire [15-1:0] node3550;
	wire [15-1:0] node3553;
	wire [15-1:0] node3555;
	wire [15-1:0] node3558;
	wire [15-1:0] node3559;
	wire [15-1:0] node3560;
	wire [15-1:0] node3564;
	wire [15-1:0] node3566;
	wire [15-1:0] node3567;
	wire [15-1:0] node3571;
	wire [15-1:0] node3572;
	wire [15-1:0] node3573;
	wire [15-1:0] node3574;
	wire [15-1:0] node3577;
	wire [15-1:0] node3578;
	wire [15-1:0] node3580;
	wire [15-1:0] node3583;
	wire [15-1:0] node3584;
	wire [15-1:0] node3585;
	wire [15-1:0] node3590;
	wire [15-1:0] node3591;
	wire [15-1:0] node3592;
	wire [15-1:0] node3595;
	wire [15-1:0] node3598;
	wire [15-1:0] node3599;
	wire [15-1:0] node3601;
	wire [15-1:0] node3604;
	wire [15-1:0] node3605;
	wire [15-1:0] node3608;
	wire [15-1:0] node3611;
	wire [15-1:0] node3612;
	wire [15-1:0] node3613;
	wire [15-1:0] node3614;
	wire [15-1:0] node3617;
	wire [15-1:0] node3618;
	wire [15-1:0] node3620;
	wire [15-1:0] node3624;
	wire [15-1:0] node3625;
	wire [15-1:0] node3626;
	wire [15-1:0] node3630;
	wire [15-1:0] node3633;
	wire [15-1:0] node3634;
	wire [15-1:0] node3636;
	wire [15-1:0] node3639;
	wire [15-1:0] node3640;
	wire [15-1:0] node3644;
	wire [15-1:0] node3645;
	wire [15-1:0] node3646;
	wire [15-1:0] node3647;
	wire [15-1:0] node3648;
	wire [15-1:0] node3649;
	wire [15-1:0] node3650;
	wire [15-1:0] node3653;
	wire [15-1:0] node3654;
	wire [15-1:0] node3655;
	wire [15-1:0] node3657;
	wire [15-1:0] node3662;
	wire [15-1:0] node3664;
	wire [15-1:0] node3665;
	wire [15-1:0] node3669;
	wire [15-1:0] node3670;
	wire [15-1:0] node3671;
	wire [15-1:0] node3672;
	wire [15-1:0] node3674;
	wire [15-1:0] node3678;
	wire [15-1:0] node3679;
	wire [15-1:0] node3680;
	wire [15-1:0] node3682;
	wire [15-1:0] node3686;
	wire [15-1:0] node3689;
	wire [15-1:0] node3690;
	wire [15-1:0] node3691;
	wire [15-1:0] node3693;
	wire [15-1:0] node3696;
	wire [15-1:0] node3698;
	wire [15-1:0] node3701;
	wire [15-1:0] node3703;
	wire [15-1:0] node3705;
	wire [15-1:0] node3708;
	wire [15-1:0] node3709;
	wire [15-1:0] node3710;
	wire [15-1:0] node3711;
	wire [15-1:0] node3712;
	wire [15-1:0] node3715;
	wire [15-1:0] node3717;
	wire [15-1:0] node3720;
	wire [15-1:0] node3723;
	wire [15-1:0] node3725;
	wire [15-1:0] node3726;
	wire [15-1:0] node3728;
	wire [15-1:0] node3731;
	wire [15-1:0] node3732;
	wire [15-1:0] node3736;
	wire [15-1:0] node3737;
	wire [15-1:0] node3738;
	wire [15-1:0] node3739;
	wire [15-1:0] node3740;
	wire [15-1:0] node3742;
	wire [15-1:0] node3747;
	wire [15-1:0] node3748;
	wire [15-1:0] node3751;
	wire [15-1:0] node3754;
	wire [15-1:0] node3755;
	wire [15-1:0] node3756;
	wire [15-1:0] node3759;
	wire [15-1:0] node3761;
	wire [15-1:0] node3764;
	wire [15-1:0] node3766;
	wire [15-1:0] node3769;
	wire [15-1:0] node3770;
	wire [15-1:0] node3771;
	wire [15-1:0] node3772;
	wire [15-1:0] node3773;
	wire [15-1:0] node3774;
	wire [15-1:0] node3777;
	wire [15-1:0] node3779;
	wire [15-1:0] node3782;
	wire [15-1:0] node3783;
	wire [15-1:0] node3787;
	wire [15-1:0] node3788;
	wire [15-1:0] node3789;
	wire [15-1:0] node3792;
	wire [15-1:0] node3793;
	wire [15-1:0] node3797;
	wire [15-1:0] node3800;
	wire [15-1:0] node3801;
	wire [15-1:0] node3802;
	wire [15-1:0] node3803;
	wire [15-1:0] node3807;
	wire [15-1:0] node3808;
	wire [15-1:0] node3810;
	wire [15-1:0] node3811;
	wire [15-1:0] node3815;
	wire [15-1:0] node3817;
	wire [15-1:0] node3820;
	wire [15-1:0] node3821;
	wire [15-1:0] node3823;
	wire [15-1:0] node3825;
	wire [15-1:0] node3826;
	wire [15-1:0] node3830;
	wire [15-1:0] node3831;
	wire [15-1:0] node3834;
	wire [15-1:0] node3835;
	wire [15-1:0] node3839;
	wire [15-1:0] node3840;
	wire [15-1:0] node3841;
	wire [15-1:0] node3842;
	wire [15-1:0] node3844;
	wire [15-1:0] node3848;
	wire [15-1:0] node3849;
	wire [15-1:0] node3850;
	wire [15-1:0] node3853;
	wire [15-1:0] node3856;
	wire [15-1:0] node3858;
	wire [15-1:0] node3861;
	wire [15-1:0] node3862;
	wire [15-1:0] node3863;
	wire [15-1:0] node3865;
	wire [15-1:0] node3866;
	wire [15-1:0] node3868;
	wire [15-1:0] node3872;
	wire [15-1:0] node3873;
	wire [15-1:0] node3874;
	wire [15-1:0] node3878;
	wire [15-1:0] node3881;
	wire [15-1:0] node3882;
	wire [15-1:0] node3883;
	wire [15-1:0] node3887;
	wire [15-1:0] node3890;
	wire [15-1:0] node3891;
	wire [15-1:0] node3892;
	wire [15-1:0] node3893;
	wire [15-1:0] node3894;
	wire [15-1:0] node3895;
	wire [15-1:0] node3896;
	wire [15-1:0] node3897;
	wire [15-1:0] node3901;
	wire [15-1:0] node3904;
	wire [15-1:0] node3906;
	wire [15-1:0] node3909;
	wire [15-1:0] node3910;
	wire [15-1:0] node3911;
	wire [15-1:0] node3915;
	wire [15-1:0] node3916;
	wire [15-1:0] node3920;
	wire [15-1:0] node3921;
	wire [15-1:0] node3922;
	wire [15-1:0] node3924;
	wire [15-1:0] node3925;
	wire [15-1:0] node3929;
	wire [15-1:0] node3930;
	wire [15-1:0] node3934;
	wire [15-1:0] node3935;
	wire [15-1:0] node3936;
	wire [15-1:0] node3939;
	wire [15-1:0] node3942;
	wire [15-1:0] node3943;
	wire [15-1:0] node3946;
	wire [15-1:0] node3947;
	wire [15-1:0] node3951;
	wire [15-1:0] node3952;
	wire [15-1:0] node3953;
	wire [15-1:0] node3954;
	wire [15-1:0] node3955;
	wire [15-1:0] node3956;
	wire [15-1:0] node3958;
	wire [15-1:0] node3963;
	wire [15-1:0] node3964;
	wire [15-1:0] node3967;
	wire [15-1:0] node3969;
	wire [15-1:0] node3972;
	wire [15-1:0] node3973;
	wire [15-1:0] node3974;
	wire [15-1:0] node3975;
	wire [15-1:0] node3979;
	wire [15-1:0] node3980;
	wire [15-1:0] node3984;
	wire [15-1:0] node3985;
	wire [15-1:0] node3989;
	wire [15-1:0] node3990;
	wire [15-1:0] node3991;
	wire [15-1:0] node3993;
	wire [15-1:0] node3995;
	wire [15-1:0] node3998;
	wire [15-1:0] node3999;
	wire [15-1:0] node4001;
	wire [15-1:0] node4002;
	wire [15-1:0] node4006;
	wire [15-1:0] node4007;
	wire [15-1:0] node4008;
	wire [15-1:0] node4012;
	wire [15-1:0] node4013;
	wire [15-1:0] node4017;
	wire [15-1:0] node4018;
	wire [15-1:0] node4020;
	wire [15-1:0] node4022;
	wire [15-1:0] node4024;
	wire [15-1:0] node4027;
	wire [15-1:0] node4029;
	wire [15-1:0] node4030;
	wire [15-1:0] node4032;
	wire [15-1:0] node4035;
	wire [15-1:0] node4037;
	wire [15-1:0] node4040;
	wire [15-1:0] node4041;
	wire [15-1:0] node4042;
	wire [15-1:0] node4043;
	wire [15-1:0] node4044;
	wire [15-1:0] node4046;
	wire [15-1:0] node4047;
	wire [15-1:0] node4048;
	wire [15-1:0] node4053;
	wire [15-1:0] node4054;
	wire [15-1:0] node4055;
	wire [15-1:0] node4060;
	wire [15-1:0] node4061;
	wire [15-1:0] node4062;
	wire [15-1:0] node4065;
	wire [15-1:0] node4068;
	wire [15-1:0] node4069;
	wire [15-1:0] node4070;
	wire [15-1:0] node4072;
	wire [15-1:0] node4075;
	wire [15-1:0] node4077;
	wire [15-1:0] node4080;
	wire [15-1:0] node4081;
	wire [15-1:0] node4084;
	wire [15-1:0] node4087;
	wire [15-1:0] node4088;
	wire [15-1:0] node4089;
	wire [15-1:0] node4091;
	wire [15-1:0] node4092;
	wire [15-1:0] node4097;
	wire [15-1:0] node4098;
	wire [15-1:0] node4100;
	wire [15-1:0] node4102;
	wire [15-1:0] node4105;
	wire [15-1:0] node4106;
	wire [15-1:0] node4107;
	wire [15-1:0] node4111;
	wire [15-1:0] node4113;
	wire [15-1:0] node4116;
	wire [15-1:0] node4117;
	wire [15-1:0] node4118;
	wire [15-1:0] node4119;
	wire [15-1:0] node4120;
	wire [15-1:0] node4124;
	wire [15-1:0] node4126;
	wire [15-1:0] node4128;
	wire [15-1:0] node4131;
	wire [15-1:0] node4132;
	wire [15-1:0] node4133;
	wire [15-1:0] node4134;
	wire [15-1:0] node4138;
	wire [15-1:0] node4141;
	wire [15-1:0] node4142;
	wire [15-1:0] node4145;
	wire [15-1:0] node4147;
	wire [15-1:0] node4150;
	wire [15-1:0] node4151;
	wire [15-1:0] node4152;
	wire [15-1:0] node4154;
	wire [15-1:0] node4156;
	wire [15-1:0] node4159;
	wire [15-1:0] node4161;
	wire [15-1:0] node4163;
	wire [15-1:0] node4166;
	wire [15-1:0] node4167;
	wire [15-1:0] node4169;
	wire [15-1:0] node4170;
	wire [15-1:0] node4174;
	wire [15-1:0] node4175;
	wire [15-1:0] node4177;
	wire [15-1:0] node4181;
	wire [15-1:0] node4182;
	wire [15-1:0] node4183;
	wire [15-1:0] node4184;
	wire [15-1:0] node4185;
	wire [15-1:0] node4186;
	wire [15-1:0] node4187;
	wire [15-1:0] node4188;
	wire [15-1:0] node4189;
	wire [15-1:0] node4190;
	wire [15-1:0] node4192;
	wire [15-1:0] node4195;
	wire [15-1:0] node4196;
	wire [15-1:0] node4197;
	wire [15-1:0] node4200;
	wire [15-1:0] node4203;
	wire [15-1:0] node4206;
	wire [15-1:0] node4207;
	wire [15-1:0] node4208;
	wire [15-1:0] node4211;
	wire [15-1:0] node4212;
	wire [15-1:0] node4213;
	wire [15-1:0] node4216;
	wire [15-1:0] node4219;
	wire [15-1:0] node4220;
	wire [15-1:0] node4224;
	wire [15-1:0] node4225;
	wire [15-1:0] node4228;
	wire [15-1:0] node4231;
	wire [15-1:0] node4232;
	wire [15-1:0] node4233;
	wire [15-1:0] node4234;
	wire [15-1:0] node4236;
	wire [15-1:0] node4237;
	wire [15-1:0] node4242;
	wire [15-1:0] node4243;
	wire [15-1:0] node4246;
	wire [15-1:0] node4249;
	wire [15-1:0] node4250;
	wire [15-1:0] node4252;
	wire [15-1:0] node4255;
	wire [15-1:0] node4256;
	wire [15-1:0] node4260;
	wire [15-1:0] node4261;
	wire [15-1:0] node4262;
	wire [15-1:0] node4263;
	wire [15-1:0] node4264;
	wire [15-1:0] node4267;
	wire [15-1:0] node4269;
	wire [15-1:0] node4273;
	wire [15-1:0] node4274;
	wire [15-1:0] node4275;
	wire [15-1:0] node4276;
	wire [15-1:0] node4280;
	wire [15-1:0] node4282;
	wire [15-1:0] node4285;
	wire [15-1:0] node4286;
	wire [15-1:0] node4290;
	wire [15-1:0] node4291;
	wire [15-1:0] node4292;
	wire [15-1:0] node4293;
	wire [15-1:0] node4295;
	wire [15-1:0] node4298;
	wire [15-1:0] node4300;
	wire [15-1:0] node4301;
	wire [15-1:0] node4305;
	wire [15-1:0] node4308;
	wire [15-1:0] node4309;
	wire [15-1:0] node4312;
	wire [15-1:0] node4313;
	wire [15-1:0] node4314;
	wire [15-1:0] node4316;
	wire [15-1:0] node4321;
	wire [15-1:0] node4322;
	wire [15-1:0] node4323;
	wire [15-1:0] node4324;
	wire [15-1:0] node4325;
	wire [15-1:0] node4326;
	wire [15-1:0] node4330;
	wire [15-1:0] node4331;
	wire [15-1:0] node4333;
	wire [15-1:0] node4334;
	wire [15-1:0] node4339;
	wire [15-1:0] node4340;
	wire [15-1:0] node4341;
	wire [15-1:0] node4342;
	wire [15-1:0] node4347;
	wire [15-1:0] node4348;
	wire [15-1:0] node4352;
	wire [15-1:0] node4353;
	wire [15-1:0] node4354;
	wire [15-1:0] node4355;
	wire [15-1:0] node4356;
	wire [15-1:0] node4358;
	wire [15-1:0] node4362;
	wire [15-1:0] node4365;
	wire [15-1:0] node4366;
	wire [15-1:0] node4370;
	wire [15-1:0] node4371;
	wire [15-1:0] node4372;
	wire [15-1:0] node4375;
	wire [15-1:0] node4377;
	wire [15-1:0] node4380;
	wire [15-1:0] node4382;
	wire [15-1:0] node4385;
	wire [15-1:0] node4386;
	wire [15-1:0] node4387;
	wire [15-1:0] node4388;
	wire [15-1:0] node4389;
	wire [15-1:0] node4391;
	wire [15-1:0] node4395;
	wire [15-1:0] node4396;
	wire [15-1:0] node4399;
	wire [15-1:0] node4402;
	wire [15-1:0] node4403;
	wire [15-1:0] node4404;
	wire [15-1:0] node4407;
	wire [15-1:0] node4409;
	wire [15-1:0] node4410;
	wire [15-1:0] node4415;
	wire [15-1:0] node4416;
	wire [15-1:0] node4417;
	wire [15-1:0] node4419;
	wire [15-1:0] node4422;
	wire [15-1:0] node4423;
	wire [15-1:0] node4424;
	wire [15-1:0] node4428;
	wire [15-1:0] node4430;
	wire [15-1:0] node4433;
	wire [15-1:0] node4435;
	wire [15-1:0] node4438;
	wire [15-1:0] node4439;
	wire [15-1:0] node4440;
	wire [15-1:0] node4441;
	wire [15-1:0] node4442;
	wire [15-1:0] node4443;
	wire [15-1:0] node4445;
	wire [15-1:0] node4447;
	wire [15-1:0] node4450;
	wire [15-1:0] node4451;
	wire [15-1:0] node4455;
	wire [15-1:0] node4456;
	wire [15-1:0] node4458;
	wire [15-1:0] node4461;
	wire [15-1:0] node4462;
	wire [15-1:0] node4464;
	wire [15-1:0] node4468;
	wire [15-1:0] node4469;
	wire [15-1:0] node4470;
	wire [15-1:0] node4471;
	wire [15-1:0] node4472;
	wire [15-1:0] node4476;
	wire [15-1:0] node4479;
	wire [15-1:0] node4480;
	wire [15-1:0] node4483;
	wire [15-1:0] node4485;
	wire [15-1:0] node4486;
	wire [15-1:0] node4490;
	wire [15-1:0] node4491;
	wire [15-1:0] node4492;
	wire [15-1:0] node4495;
	wire [15-1:0] node4498;
	wire [15-1:0] node4499;
	wire [15-1:0] node4502;
	wire [15-1:0] node4504;
	wire [15-1:0] node4506;
	wire [15-1:0] node4509;
	wire [15-1:0] node4510;
	wire [15-1:0] node4511;
	wire [15-1:0] node4513;
	wire [15-1:0] node4514;
	wire [15-1:0] node4515;
	wire [15-1:0] node4517;
	wire [15-1:0] node4520;
	wire [15-1:0] node4521;
	wire [15-1:0] node4526;
	wire [15-1:0] node4527;
	wire [15-1:0] node4529;
	wire [15-1:0] node4531;
	wire [15-1:0] node4534;
	wire [15-1:0] node4535;
	wire [15-1:0] node4536;
	wire [15-1:0] node4538;
	wire [15-1:0] node4542;
	wire [15-1:0] node4544;
	wire [15-1:0] node4547;
	wire [15-1:0] node4548;
	wire [15-1:0] node4549;
	wire [15-1:0] node4551;
	wire [15-1:0] node4553;
	wire [15-1:0] node4554;
	wire [15-1:0] node4558;
	wire [15-1:0] node4559;
	wire [15-1:0] node4563;
	wire [15-1:0] node4564;
	wire [15-1:0] node4565;
	wire [15-1:0] node4566;
	wire [15-1:0] node4568;
	wire [15-1:0] node4572;
	wire [15-1:0] node4575;
	wire [15-1:0] node4576;
	wire [15-1:0] node4577;
	wire [15-1:0] node4581;
	wire [15-1:0] node4584;
	wire [15-1:0] node4585;
	wire [15-1:0] node4586;
	wire [15-1:0] node4587;
	wire [15-1:0] node4588;
	wire [15-1:0] node4590;
	wire [15-1:0] node4592;
	wire [15-1:0] node4595;
	wire [15-1:0] node4597;
	wire [15-1:0] node4599;
	wire [15-1:0] node4602;
	wire [15-1:0] node4603;
	wire [15-1:0] node4604;
	wire [15-1:0] node4605;
	wire [15-1:0] node4609;
	wire [15-1:0] node4612;
	wire [15-1:0] node4613;
	wire [15-1:0] node4615;
	wire [15-1:0] node4616;
	wire [15-1:0] node4620;
	wire [15-1:0] node4622;
	wire [15-1:0] node4625;
	wire [15-1:0] node4626;
	wire [15-1:0] node4627;
	wire [15-1:0] node4629;
	wire [15-1:0] node4632;
	wire [15-1:0] node4633;
	wire [15-1:0] node4634;
	wire [15-1:0] node4636;
	wire [15-1:0] node4639;
	wire [15-1:0] node4642;
	wire [15-1:0] node4644;
	wire [15-1:0] node4647;
	wire [15-1:0] node4648;
	wire [15-1:0] node4651;
	wire [15-1:0] node4653;
	wire [15-1:0] node4656;
	wire [15-1:0] node4657;
	wire [15-1:0] node4658;
	wire [15-1:0] node4659;
	wire [15-1:0] node4660;
	wire [15-1:0] node4663;
	wire [15-1:0] node4665;
	wire [15-1:0] node4666;
	wire [15-1:0] node4670;
	wire [15-1:0] node4671;
	wire [15-1:0] node4672;
	wire [15-1:0] node4675;
	wire [15-1:0] node4678;
	wire [15-1:0] node4681;
	wire [15-1:0] node4682;
	wire [15-1:0] node4684;
	wire [15-1:0] node4688;
	wire [15-1:0] node4689;
	wire [15-1:0] node4690;
	wire [15-1:0] node4693;
	wire [15-1:0] node4694;
	wire [15-1:0] node4696;
	wire [15-1:0] node4700;
	wire [15-1:0] node4701;
	wire [15-1:0] node4704;
	wire [15-1:0] node4705;
	wire [15-1:0] node4707;
	wire [15-1:0] node4711;
	wire [15-1:0] node4712;
	wire [15-1:0] node4713;
	wire [15-1:0] node4714;
	wire [15-1:0] node4715;
	wire [15-1:0] node4716;
	wire [15-1:0] node4717;
	wire [15-1:0] node4718;
	wire [15-1:0] node4719;
	wire [15-1:0] node4723;
	wire [15-1:0] node4725;
	wire [15-1:0] node4728;
	wire [15-1:0] node4729;
	wire [15-1:0] node4730;
	wire [15-1:0] node4735;
	wire [15-1:0] node4736;
	wire [15-1:0] node4737;
	wire [15-1:0] node4741;
	wire [15-1:0] node4742;
	wire [15-1:0] node4743;
	wire [15-1:0] node4745;
	wire [15-1:0] node4750;
	wire [15-1:0] node4751;
	wire [15-1:0] node4752;
	wire [15-1:0] node4753;
	wire [15-1:0] node4754;
	wire [15-1:0] node4759;
	wire [15-1:0] node4760;
	wire [15-1:0] node4763;
	wire [15-1:0] node4766;
	wire [15-1:0] node4767;
	wire [15-1:0] node4768;
	wire [15-1:0] node4771;
	wire [15-1:0] node4773;
	wire [15-1:0] node4776;
	wire [15-1:0] node4777;
	wire [15-1:0] node4781;
	wire [15-1:0] node4782;
	wire [15-1:0] node4783;
	wire [15-1:0] node4784;
	wire [15-1:0] node4786;
	wire [15-1:0] node4789;
	wire [15-1:0] node4791;
	wire [15-1:0] node4794;
	wire [15-1:0] node4796;
	wire [15-1:0] node4797;
	wire [15-1:0] node4800;
	wire [15-1:0] node4803;
	wire [15-1:0] node4804;
	wire [15-1:0] node4805;
	wire [15-1:0] node4806;
	wire [15-1:0] node4808;
	wire [15-1:0] node4809;
	wire [15-1:0] node4813;
	wire [15-1:0] node4816;
	wire [15-1:0] node4817;
	wire [15-1:0] node4818;
	wire [15-1:0] node4822;
	wire [15-1:0] node4825;
	wire [15-1:0] node4826;
	wire [15-1:0] node4828;
	wire [15-1:0] node4831;
	wire [15-1:0] node4832;
	wire [15-1:0] node4833;
	wire [15-1:0] node4838;
	wire [15-1:0] node4839;
	wire [15-1:0] node4840;
	wire [15-1:0] node4841;
	wire [15-1:0] node4842;
	wire [15-1:0] node4844;
	wire [15-1:0] node4846;
	wire [15-1:0] node4849;
	wire [15-1:0] node4850;
	wire [15-1:0] node4853;
	wire [15-1:0] node4854;
	wire [15-1:0] node4858;
	wire [15-1:0] node4859;
	wire [15-1:0] node4861;
	wire [15-1:0] node4862;
	wire [15-1:0] node4866;
	wire [15-1:0] node4867;
	wire [15-1:0] node4869;
	wire [15-1:0] node4870;
	wire [15-1:0] node4874;
	wire [15-1:0] node4877;
	wire [15-1:0] node4878;
	wire [15-1:0] node4879;
	wire [15-1:0] node4881;
	wire [15-1:0] node4884;
	wire [15-1:0] node4886;
	wire [15-1:0] node4889;
	wire [15-1:0] node4891;
	wire [15-1:0] node4893;
	wire [15-1:0] node4896;
	wire [15-1:0] node4897;
	wire [15-1:0] node4898;
	wire [15-1:0] node4899;
	wire [15-1:0] node4900;
	wire [15-1:0] node4903;
	wire [15-1:0] node4906;
	wire [15-1:0] node4907;
	wire [15-1:0] node4910;
	wire [15-1:0] node4913;
	wire [15-1:0] node4914;
	wire [15-1:0] node4916;
	wire [15-1:0] node4918;
	wire [15-1:0] node4921;
	wire [15-1:0] node4923;
	wire [15-1:0] node4926;
	wire [15-1:0] node4927;
	wire [15-1:0] node4928;
	wire [15-1:0] node4930;
	wire [15-1:0] node4931;
	wire [15-1:0] node4935;
	wire [15-1:0] node4936;
	wire [15-1:0] node4937;
	wire [15-1:0] node4938;
	wire [15-1:0] node4941;
	wire [15-1:0] node4945;
	wire [15-1:0] node4947;
	wire [15-1:0] node4948;
	wire [15-1:0] node4951;
	wire [15-1:0] node4954;
	wire [15-1:0] node4955;
	wire [15-1:0] node4957;
	wire [15-1:0] node4960;
	wire [15-1:0] node4961;
	wire [15-1:0] node4963;
	wire [15-1:0] node4967;
	wire [15-1:0] node4968;
	wire [15-1:0] node4969;
	wire [15-1:0] node4970;
	wire [15-1:0] node4971;
	wire [15-1:0] node4972;
	wire [15-1:0] node4974;
	wire [15-1:0] node4976;
	wire [15-1:0] node4979;
	wire [15-1:0] node4980;
	wire [15-1:0] node4982;
	wire [15-1:0] node4983;
	wire [15-1:0] node4988;
	wire [15-1:0] node4990;
	wire [15-1:0] node4991;
	wire [15-1:0] node4993;
	wire [15-1:0] node4994;
	wire [15-1:0] node4999;
	wire [15-1:0] node5000;
	wire [15-1:0] node5001;
	wire [15-1:0] node5004;
	wire [15-1:0] node5005;
	wire [15-1:0] node5009;
	wire [15-1:0] node5010;
	wire [15-1:0] node5012;
	wire [15-1:0] node5014;
	wire [15-1:0] node5017;
	wire [15-1:0] node5019;
	wire [15-1:0] node5020;
	wire [15-1:0] node5024;
	wire [15-1:0] node5025;
	wire [15-1:0] node5026;
	wire [15-1:0] node5027;
	wire [15-1:0] node5029;
	wire [15-1:0] node5032;
	wire [15-1:0] node5034;
	wire [15-1:0] node5035;
	wire [15-1:0] node5039;
	wire [15-1:0] node5040;
	wire [15-1:0] node5042;
	wire [15-1:0] node5044;
	wire [15-1:0] node5047;
	wire [15-1:0] node5048;
	wire [15-1:0] node5052;
	wire [15-1:0] node5053;
	wire [15-1:0] node5054;
	wire [15-1:0] node5055;
	wire [15-1:0] node5056;
	wire [15-1:0] node5057;
	wire [15-1:0] node5062;
	wire [15-1:0] node5065;
	wire [15-1:0] node5066;
	wire [15-1:0] node5069;
	wire [15-1:0] node5070;
	wire [15-1:0] node5074;
	wire [15-1:0] node5075;
	wire [15-1:0] node5078;
	wire [15-1:0] node5080;
	wire [15-1:0] node5081;
	wire [15-1:0] node5085;
	wire [15-1:0] node5086;
	wire [15-1:0] node5087;
	wire [15-1:0] node5088;
	wire [15-1:0] node5089;
	wire [15-1:0] node5092;
	wire [15-1:0] node5095;
	wire [15-1:0] node5096;
	wire [15-1:0] node5098;
	wire [15-1:0] node5100;
	wire [15-1:0] node5103;
	wire [15-1:0] node5104;
	wire [15-1:0] node5105;
	wire [15-1:0] node5110;
	wire [15-1:0] node5111;
	wire [15-1:0] node5112;
	wire [15-1:0] node5113;
	wire [15-1:0] node5114;
	wire [15-1:0] node5118;
	wire [15-1:0] node5121;
	wire [15-1:0] node5122;
	wire [15-1:0] node5125;
	wire [15-1:0] node5127;
	wire [15-1:0] node5128;
	wire [15-1:0] node5132;
	wire [15-1:0] node5133;
	wire [15-1:0] node5134;
	wire [15-1:0] node5136;
	wire [15-1:0] node5139;
	wire [15-1:0] node5142;
	wire [15-1:0] node5143;
	wire [15-1:0] node5147;
	wire [15-1:0] node5148;
	wire [15-1:0] node5149;
	wire [15-1:0] node5150;
	wire [15-1:0] node5151;
	wire [15-1:0] node5155;
	wire [15-1:0] node5156;
	wire [15-1:0] node5157;
	wire [15-1:0] node5158;
	wire [15-1:0] node5162;
	wire [15-1:0] node5165;
	wire [15-1:0] node5168;
	wire [15-1:0] node5169;
	wire [15-1:0] node5170;
	wire [15-1:0] node5173;
	wire [15-1:0] node5176;
	wire [15-1:0] node5177;
	wire [15-1:0] node5178;
	wire [15-1:0] node5182;
	wire [15-1:0] node5183;
	wire [15-1:0] node5187;
	wire [15-1:0] node5188;
	wire [15-1:0] node5189;
	wire [15-1:0] node5191;
	wire [15-1:0] node5194;
	wire [15-1:0] node5196;
	wire [15-1:0] node5197;
	wire [15-1:0] node5201;
	wire [15-1:0] node5202;
	wire [15-1:0] node5203;
	wire [15-1:0] node5205;
	wire [15-1:0] node5207;
	wire [15-1:0] node5211;
	wire [15-1:0] node5212;
	wire [15-1:0] node5215;
	wire [15-1:0] node5216;
	wire [15-1:0] node5218;
	wire [15-1:0] node5222;
	wire [15-1:0] node5223;
	wire [15-1:0] node5224;
	wire [15-1:0] node5225;
	wire [15-1:0] node5226;
	wire [15-1:0] node5227;
	wire [15-1:0] node5228;
	wire [15-1:0] node5229;
	wire [15-1:0] node5230;
	wire [15-1:0] node5231;
	wire [15-1:0] node5235;
	wire [15-1:0] node5237;
	wire [15-1:0] node5240;
	wire [15-1:0] node5241;
	wire [15-1:0] node5244;
	wire [15-1:0] node5247;
	wire [15-1:0] node5249;
	wire [15-1:0] node5250;
	wire [15-1:0] node5251;
	wire [15-1:0] node5254;
	wire [15-1:0] node5255;
	wire [15-1:0] node5259;
	wire [15-1:0] node5261;
	wire [15-1:0] node5264;
	wire [15-1:0] node5265;
	wire [15-1:0] node5266;
	wire [15-1:0] node5267;
	wire [15-1:0] node5271;
	wire [15-1:0] node5272;
	wire [15-1:0] node5274;
	wire [15-1:0] node5275;
	wire [15-1:0] node5279;
	wire [15-1:0] node5281;
	wire [15-1:0] node5282;
	wire [15-1:0] node5286;
	wire [15-1:0] node5287;
	wire [15-1:0] node5288;
	wire [15-1:0] node5291;
	wire [15-1:0] node5294;
	wire [15-1:0] node5295;
	wire [15-1:0] node5298;
	wire [15-1:0] node5301;
	wire [15-1:0] node5302;
	wire [15-1:0] node5303;
	wire [15-1:0] node5304;
	wire [15-1:0] node5306;
	wire [15-1:0] node5309;
	wire [15-1:0] node5311;
	wire [15-1:0] node5314;
	wire [15-1:0] node5315;
	wire [15-1:0] node5317;
	wire [15-1:0] node5320;
	wire [15-1:0] node5321;
	wire [15-1:0] node5325;
	wire [15-1:0] node5326;
	wire [15-1:0] node5327;
	wire [15-1:0] node5328;
	wire [15-1:0] node5331;
	wire [15-1:0] node5334;
	wire [15-1:0] node5335;
	wire [15-1:0] node5339;
	wire [15-1:0] node5340;
	wire [15-1:0] node5343;
	wire [15-1:0] node5344;
	wire [15-1:0] node5346;
	wire [15-1:0] node5350;
	wire [15-1:0] node5351;
	wire [15-1:0] node5352;
	wire [15-1:0] node5353;
	wire [15-1:0] node5354;
	wire [15-1:0] node5355;
	wire [15-1:0] node5356;
	wire [15-1:0] node5358;
	wire [15-1:0] node5363;
	wire [15-1:0] node5364;
	wire [15-1:0] node5368;
	wire [15-1:0] node5369;
	wire [15-1:0] node5370;
	wire [15-1:0] node5373;
	wire [15-1:0] node5375;
	wire [15-1:0] node5378;
	wire [15-1:0] node5379;
	wire [15-1:0] node5380;
	wire [15-1:0] node5382;
	wire [15-1:0] node5387;
	wire [15-1:0] node5388;
	wire [15-1:0] node5389;
	wire [15-1:0] node5390;
	wire [15-1:0] node5391;
	wire [15-1:0] node5392;
	wire [15-1:0] node5397;
	wire [15-1:0] node5400;
	wire [15-1:0] node5401;
	wire [15-1:0] node5402;
	wire [15-1:0] node5404;
	wire [15-1:0] node5408;
	wire [15-1:0] node5411;
	wire [15-1:0] node5412;
	wire [15-1:0] node5414;
	wire [15-1:0] node5417;
	wire [15-1:0] node5418;
	wire [15-1:0] node5422;
	wire [15-1:0] node5423;
	wire [15-1:0] node5424;
	wire [15-1:0] node5425;
	wire [15-1:0] node5428;
	wire [15-1:0] node5429;
	wire [15-1:0] node5430;
	wire [15-1:0] node5435;
	wire [15-1:0] node5436;
	wire [15-1:0] node5437;
	wire [15-1:0] node5441;
	wire [15-1:0] node5444;
	wire [15-1:0] node5445;
	wire [15-1:0] node5446;
	wire [15-1:0] node5447;
	wire [15-1:0] node5450;
	wire [15-1:0] node5453;
	wire [15-1:0] node5454;
	wire [15-1:0] node5455;
	wire [15-1:0] node5459;
	wire [15-1:0] node5462;
	wire [15-1:0] node5463;
	wire [15-1:0] node5465;
	wire [15-1:0] node5467;
	wire [15-1:0] node5470;
	wire [15-1:0] node5472;
	wire [15-1:0] node5473;
	wire [15-1:0] node5477;
	wire [15-1:0] node5478;
	wire [15-1:0] node5479;
	wire [15-1:0] node5480;
	wire [15-1:0] node5481;
	wire [15-1:0] node5482;
	wire [15-1:0] node5483;
	wire [15-1:0] node5485;
	wire [15-1:0] node5488;
	wire [15-1:0] node5491;
	wire [15-1:0] node5493;
	wire [15-1:0] node5494;
	wire [15-1:0] node5498;
	wire [15-1:0] node5499;
	wire [15-1:0] node5500;
	wire [15-1:0] node5501;
	wire [15-1:0] node5503;
	wire [15-1:0] node5507;
	wire [15-1:0] node5510;
	wire [15-1:0] node5513;
	wire [15-1:0] node5514;
	wire [15-1:0] node5515;
	wire [15-1:0] node5517;
	wire [15-1:0] node5520;
	wire [15-1:0] node5521;
	wire [15-1:0] node5525;
	wire [15-1:0] node5526;
	wire [15-1:0] node5527;
	wire [15-1:0] node5529;
	wire [15-1:0] node5530;
	wire [15-1:0] node5534;
	wire [15-1:0] node5536;
	wire [15-1:0] node5537;
	wire [15-1:0] node5542;
	wire [15-1:0] node5543;
	wire [15-1:0] node5544;
	wire [15-1:0] node5545;
	wire [15-1:0] node5548;
	wire [15-1:0] node5551;
	wire [15-1:0] node5552;
	wire [15-1:0] node5553;
	wire [15-1:0] node5555;
	wire [15-1:0] node5559;
	wire [15-1:0] node5560;
	wire [15-1:0] node5562;
	wire [15-1:0] node5563;
	wire [15-1:0] node5567;
	wire [15-1:0] node5570;
	wire [15-1:0] node5571;
	wire [15-1:0] node5572;
	wire [15-1:0] node5573;
	wire [15-1:0] node5574;
	wire [15-1:0] node5578;
	wire [15-1:0] node5581;
	wire [15-1:0] node5582;
	wire [15-1:0] node5586;
	wire [15-1:0] node5587;
	wire [15-1:0] node5588;
	wire [15-1:0] node5589;
	wire [15-1:0] node5591;
	wire [15-1:0] node5596;
	wire [15-1:0] node5597;
	wire [15-1:0] node5600;
	wire [15-1:0] node5603;
	wire [15-1:0] node5604;
	wire [15-1:0] node5605;
	wire [15-1:0] node5606;
	wire [15-1:0] node5607;
	wire [15-1:0] node5608;
	wire [15-1:0] node5610;
	wire [15-1:0] node5611;
	wire [15-1:0] node5615;
	wire [15-1:0] node5618;
	wire [15-1:0] node5619;
	wire [15-1:0] node5623;
	wire [15-1:0] node5624;
	wire [15-1:0] node5625;
	wire [15-1:0] node5626;
	wire [15-1:0] node5630;
	wire [15-1:0] node5633;
	wire [15-1:0] node5634;
	wire [15-1:0] node5638;
	wire [15-1:0] node5639;
	wire [15-1:0] node5640;
	wire [15-1:0] node5641;
	wire [15-1:0] node5642;
	wire [15-1:0] node5647;
	wire [15-1:0] node5648;
	wire [15-1:0] node5651;
	wire [15-1:0] node5652;
	wire [15-1:0] node5654;
	wire [15-1:0] node5658;
	wire [15-1:0] node5659;
	wire [15-1:0] node5660;
	wire [15-1:0] node5664;
	wire [15-1:0] node5666;
	wire [15-1:0] node5667;
	wire [15-1:0] node5670;
	wire [15-1:0] node5673;
	wire [15-1:0] node5674;
	wire [15-1:0] node5675;
	wire [15-1:0] node5676;
	wire [15-1:0] node5677;
	wire [15-1:0] node5680;
	wire [15-1:0] node5682;
	wire [15-1:0] node5685;
	wire [15-1:0] node5686;
	wire [15-1:0] node5689;
	wire [15-1:0] node5692;
	wire [15-1:0] node5693;
	wire [15-1:0] node5695;
	wire [15-1:0] node5698;
	wire [15-1:0] node5699;
	wire [15-1:0] node5700;
	wire [15-1:0] node5704;
	wire [15-1:0] node5706;
	wire [15-1:0] node5709;
	wire [15-1:0] node5710;
	wire [15-1:0] node5711;
	wire [15-1:0] node5713;
	wire [15-1:0] node5715;
	wire [15-1:0] node5718;
	wire [15-1:0] node5720;
	wire [15-1:0] node5723;
	wire [15-1:0] node5724;
	wire [15-1:0] node5726;
	wire [15-1:0] node5729;
	wire [15-1:0] node5730;
	wire [15-1:0] node5733;
	wire [15-1:0] node5734;
	wire [15-1:0] node5736;
	wire [15-1:0] node5740;
	wire [15-1:0] node5741;
	wire [15-1:0] node5742;
	wire [15-1:0] node5743;
	wire [15-1:0] node5744;
	wire [15-1:0] node5745;
	wire [15-1:0] node5746;
	wire [15-1:0] node5747;
	wire [15-1:0] node5751;
	wire [15-1:0] node5754;
	wire [15-1:0] node5755;
	wire [15-1:0] node5756;
	wire [15-1:0] node5761;
	wire [15-1:0] node5762;
	wire [15-1:0] node5763;
	wire [15-1:0] node5764;
	wire [15-1:0] node5768;
	wire [15-1:0] node5769;
	wire [15-1:0] node5773;
	wire [15-1:0] node5774;
	wire [15-1:0] node5776;
	wire [15-1:0] node5779;
	wire [15-1:0] node5780;
	wire [15-1:0] node5784;
	wire [15-1:0] node5785;
	wire [15-1:0] node5786;
	wire [15-1:0] node5787;
	wire [15-1:0] node5788;
	wire [15-1:0] node5790;
	wire [15-1:0] node5793;
	wire [15-1:0] node5794;
	wire [15-1:0] node5795;
	wire [15-1:0] node5800;
	wire [15-1:0] node5802;
	wire [15-1:0] node5805;
	wire [15-1:0] node5806;
	wire [15-1:0] node5807;
	wire [15-1:0] node5809;
	wire [15-1:0] node5811;
	wire [15-1:0] node5815;
	wire [15-1:0] node5816;
	wire [15-1:0] node5819;
	wire [15-1:0] node5821;
	wire [15-1:0] node5824;
	wire [15-1:0] node5825;
	wire [15-1:0] node5826;
	wire [15-1:0] node5829;
	wire [15-1:0] node5830;
	wire [15-1:0] node5833;
	wire [15-1:0] node5835;
	wire [15-1:0] node5838;
	wire [15-1:0] node5840;
	wire [15-1:0] node5841;
	wire [15-1:0] node5843;
	wire [15-1:0] node5846;
	wire [15-1:0] node5848;
	wire [15-1:0] node5851;
	wire [15-1:0] node5852;
	wire [15-1:0] node5853;
	wire [15-1:0] node5854;
	wire [15-1:0] node5855;
	wire [15-1:0] node5857;
	wire [15-1:0] node5858;
	wire [15-1:0] node5862;
	wire [15-1:0] node5863;
	wire [15-1:0] node5864;
	wire [15-1:0] node5868;
	wire [15-1:0] node5871;
	wire [15-1:0] node5872;
	wire [15-1:0] node5874;
	wire [15-1:0] node5876;
	wire [15-1:0] node5879;
	wire [15-1:0] node5880;
	wire [15-1:0] node5882;
	wire [15-1:0] node5883;
	wire [15-1:0] node5887;
	wire [15-1:0] node5889;
	wire [15-1:0] node5892;
	wire [15-1:0] node5893;
	wire [15-1:0] node5894;
	wire [15-1:0] node5895;
	wire [15-1:0] node5898;
	wire [15-1:0] node5901;
	wire [15-1:0] node5902;
	wire [15-1:0] node5906;
	wire [15-1:0] node5907;
	wire [15-1:0] node5909;
	wire [15-1:0] node5912;
	wire [15-1:0] node5913;
	wire [15-1:0] node5914;
	wire [15-1:0] node5918;
	wire [15-1:0] node5921;
	wire [15-1:0] node5922;
	wire [15-1:0] node5923;
	wire [15-1:0] node5924;
	wire [15-1:0] node5925;
	wire [15-1:0] node5929;
	wire [15-1:0] node5930;
	wire [15-1:0] node5933;
	wire [15-1:0] node5935;
	wire [15-1:0] node5938;
	wire [15-1:0] node5939;
	wire [15-1:0] node5940;
	wire [15-1:0] node5942;
	wire [15-1:0] node5945;
	wire [15-1:0] node5948;
	wire [15-1:0] node5949;
	wire [15-1:0] node5950;
	wire [15-1:0] node5954;
	wire [15-1:0] node5957;
	wire [15-1:0] node5958;
	wire [15-1:0] node5959;
	wire [15-1:0] node5960;
	wire [15-1:0] node5963;
	wire [15-1:0] node5966;
	wire [15-1:0] node5967;
	wire [15-1:0] node5971;
	wire [15-1:0] node5972;
	wire [15-1:0] node5973;
	wire [15-1:0] node5974;
	wire [15-1:0] node5976;
	wire [15-1:0] node5980;
	wire [15-1:0] node5982;
	wire [15-1:0] node5985;
	wire [15-1:0] node5986;
	wire [15-1:0] node5990;
	wire [15-1:0] node5991;
	wire [15-1:0] node5992;
	wire [15-1:0] node5993;
	wire [15-1:0] node5994;
	wire [15-1:0] node5995;
	wire [15-1:0] node5997;
	wire [15-1:0] node6000;
	wire [15-1:0] node6003;
	wire [15-1:0] node6004;
	wire [15-1:0] node6007;
	wire [15-1:0] node6008;
	wire [15-1:0] node6012;
	wire [15-1:0] node6013;
	wire [15-1:0] node6014;
	wire [15-1:0] node6015;
	wire [15-1:0] node6018;
	wire [15-1:0] node6021;
	wire [15-1:0] node6022;
	wire [15-1:0] node6023;
	wire [15-1:0] node6027;
	wire [15-1:0] node6030;
	wire [15-1:0] node6032;
	wire [15-1:0] node6033;
	wire [15-1:0] node6036;
	wire [15-1:0] node6039;
	wire [15-1:0] node6040;
	wire [15-1:0] node6041;
	wire [15-1:0] node6042;
	wire [15-1:0] node6043;
	wire [15-1:0] node6046;
	wire [15-1:0] node6048;
	wire [15-1:0] node6051;
	wire [15-1:0] node6052;
	wire [15-1:0] node6054;
	wire [15-1:0] node6055;
	wire [15-1:0] node6059;
	wire [15-1:0] node6061;
	wire [15-1:0] node6064;
	wire [15-1:0] node6065;
	wire [15-1:0] node6066;
	wire [15-1:0] node6069;
	wire [15-1:0] node6072;
	wire [15-1:0] node6073;
	wire [15-1:0] node6074;
	wire [15-1:0] node6078;
	wire [15-1:0] node6079;
	wire [15-1:0] node6083;
	wire [15-1:0] node6084;
	wire [15-1:0] node6086;
	wire [15-1:0] node6087;
	wire [15-1:0] node6091;
	wire [15-1:0] node6092;
	wire [15-1:0] node6093;
	wire [15-1:0] node6095;
	wire [15-1:0] node6099;
	wire [15-1:0] node6101;
	wire [15-1:0] node6104;
	wire [15-1:0] node6105;
	wire [15-1:0] node6106;
	wire [15-1:0] node6107;
	wire [15-1:0] node6108;
	wire [15-1:0] node6111;
	wire [15-1:0] node6112;
	wire [15-1:0] node6115;
	wire [15-1:0] node6118;
	wire [15-1:0] node6119;
	wire [15-1:0] node6121;
	wire [15-1:0] node6124;
	wire [15-1:0] node6126;
	wire [15-1:0] node6129;
	wire [15-1:0] node6130;
	wire [15-1:0] node6131;
	wire [15-1:0] node6134;
	wire [15-1:0] node6135;
	wire [15-1:0] node6136;
	wire [15-1:0] node6140;
	wire [15-1:0] node6143;
	wire [15-1:0] node6144;
	wire [15-1:0] node6146;
	wire [15-1:0] node6149;
	wire [15-1:0] node6151;
	wire [15-1:0] node6154;
	wire [15-1:0] node6155;
	wire [15-1:0] node6156;
	wire [15-1:0] node6157;
	wire [15-1:0] node6159;
	wire [15-1:0] node6162;
	wire [15-1:0] node6163;
	wire [15-1:0] node6167;
	wire [15-1:0] node6168;
	wire [15-1:0] node6170;
	wire [15-1:0] node6171;
	wire [15-1:0] node6173;
	wire [15-1:0] node6177;
	wire [15-1:0] node6178;
	wire [15-1:0] node6181;
	wire [15-1:0] node6183;
	wire [15-1:0] node6186;
	wire [15-1:0] node6187;
	wire [15-1:0] node6188;
	wire [15-1:0] node6189;
	wire [15-1:0] node6190;
	wire [15-1:0] node6194;
	wire [15-1:0] node6196;
	wire [15-1:0] node6200;
	wire [15-1:0] node6201;
	wire [15-1:0] node6202;
	wire [15-1:0] node6203;
	wire [15-1:0] node6207;
	wire [15-1:0] node6210;
	wire [15-1:0] node6211;
	wire [15-1:0] node6214;
	wire [15-1:0] node6216;
	wire [15-1:0] node6219;
	wire [15-1:0] node6220;
	wire [15-1:0] node6221;
	wire [15-1:0] node6222;
	wire [15-1:0] node6223;
	wire [15-1:0] node6224;
	wire [15-1:0] node6225;
	wire [15-1:0] node6226;
	wire [15-1:0] node6228;
	wire [15-1:0] node6229;
	wire [15-1:0] node6230;
	wire [15-1:0] node6234;
	wire [15-1:0] node6237;
	wire [15-1:0] node6238;
	wire [15-1:0] node6239;
	wire [15-1:0] node6243;
	wire [15-1:0] node6245;
	wire [15-1:0] node6248;
	wire [15-1:0] node6249;
	wire [15-1:0] node6250;
	wire [15-1:0] node6253;
	wire [15-1:0] node6254;
	wire [15-1:0] node6257;
	wire [15-1:0] node6260;
	wire [15-1:0] node6262;
	wire [15-1:0] node6263;
	wire [15-1:0] node6264;
	wire [15-1:0] node6266;
	wire [15-1:0] node6270;
	wire [15-1:0] node6273;
	wire [15-1:0] node6274;
	wire [15-1:0] node6275;
	wire [15-1:0] node6277;
	wire [15-1:0] node6278;
	wire [15-1:0] node6282;
	wire [15-1:0] node6283;
	wire [15-1:0] node6286;
	wire [15-1:0] node6287;
	wire [15-1:0] node6289;
	wire [15-1:0] node6290;
	wire [15-1:0] node6295;
	wire [15-1:0] node6296;
	wire [15-1:0] node6297;
	wire [15-1:0] node6298;
	wire [15-1:0] node6302;
	wire [15-1:0] node6303;
	wire [15-1:0] node6306;
	wire [15-1:0] node6308;
	wire [15-1:0] node6311;
	wire [15-1:0] node6312;
	wire [15-1:0] node6314;
	wire [15-1:0] node6316;
	wire [15-1:0] node6319;
	wire [15-1:0] node6320;
	wire [15-1:0] node6322;
	wire [15-1:0] node6326;
	wire [15-1:0] node6327;
	wire [15-1:0] node6328;
	wire [15-1:0] node6329;
	wire [15-1:0] node6330;
	wire [15-1:0] node6331;
	wire [15-1:0] node6333;
	wire [15-1:0] node6336;
	wire [15-1:0] node6337;
	wire [15-1:0] node6339;
	wire [15-1:0] node6343;
	wire [15-1:0] node6344;
	wire [15-1:0] node6345;
	wire [15-1:0] node6347;
	wire [15-1:0] node6350;
	wire [15-1:0] node6353;
	wire [15-1:0] node6356;
	wire [15-1:0] node6357;
	wire [15-1:0] node6358;
	wire [15-1:0] node6361;
	wire [15-1:0] node6363;
	wire [15-1:0] node6366;
	wire [15-1:0] node6368;
	wire [15-1:0] node6369;
	wire [15-1:0] node6371;
	wire [15-1:0] node6375;
	wire [15-1:0] node6376;
	wire [15-1:0] node6377;
	wire [15-1:0] node6378;
	wire [15-1:0] node6381;
	wire [15-1:0] node6384;
	wire [15-1:0] node6386;
	wire [15-1:0] node6389;
	wire [15-1:0] node6390;
	wire [15-1:0] node6391;
	wire [15-1:0] node6395;
	wire [15-1:0] node6397;
	wire [15-1:0] node6398;
	wire [15-1:0] node6402;
	wire [15-1:0] node6403;
	wire [15-1:0] node6404;
	wire [15-1:0] node6406;
	wire [15-1:0] node6408;
	wire [15-1:0] node6411;
	wire [15-1:0] node6413;
	wire [15-1:0] node6414;
	wire [15-1:0] node6415;
	wire [15-1:0] node6420;
	wire [15-1:0] node6421;
	wire [15-1:0] node6422;
	wire [15-1:0] node6424;
	wire [15-1:0] node6427;
	wire [15-1:0] node6428;
	wire [15-1:0] node6432;
	wire [15-1:0] node6433;
	wire [15-1:0] node6435;
	wire [15-1:0] node6437;
	wire [15-1:0] node6438;
	wire [15-1:0] node6442;
	wire [15-1:0] node6443;
	wire [15-1:0] node6447;
	wire [15-1:0] node6448;
	wire [15-1:0] node6449;
	wire [15-1:0] node6450;
	wire [15-1:0] node6451;
	wire [15-1:0] node6452;
	wire [15-1:0] node6453;
	wire [15-1:0] node6456;
	wire [15-1:0] node6457;
	wire [15-1:0] node6459;
	wire [15-1:0] node6462;
	wire [15-1:0] node6463;
	wire [15-1:0] node6467;
	wire [15-1:0] node6468;
	wire [15-1:0] node6472;
	wire [15-1:0] node6473;
	wire [15-1:0] node6474;
	wire [15-1:0] node6475;
	wire [15-1:0] node6479;
	wire [15-1:0] node6482;
	wire [15-1:0] node6484;
	wire [15-1:0] node6487;
	wire [15-1:0] node6488;
	wire [15-1:0] node6489;
	wire [15-1:0] node6490;
	wire [15-1:0] node6493;
	wire [15-1:0] node6496;
	wire [15-1:0] node6498;
	wire [15-1:0] node6501;
	wire [15-1:0] node6502;
	wire [15-1:0] node6503;
	wire [15-1:0] node6506;
	wire [15-1:0] node6507;
	wire [15-1:0] node6511;
	wire [15-1:0] node6512;
	wire [15-1:0] node6516;
	wire [15-1:0] node6517;
	wire [15-1:0] node6518;
	wire [15-1:0] node6519;
	wire [15-1:0] node6520;
	wire [15-1:0] node6522;
	wire [15-1:0] node6526;
	wire [15-1:0] node6527;
	wire [15-1:0] node6529;
	wire [15-1:0] node6532;
	wire [15-1:0] node6534;
	wire [15-1:0] node6535;
	wire [15-1:0] node6539;
	wire [15-1:0] node6540;
	wire [15-1:0] node6541;
	wire [15-1:0] node6543;
	wire [15-1:0] node6546;
	wire [15-1:0] node6548;
	wire [15-1:0] node6551;
	wire [15-1:0] node6552;
	wire [15-1:0] node6553;
	wire [15-1:0] node6555;
	wire [15-1:0] node6559;
	wire [15-1:0] node6561;
	wire [15-1:0] node6564;
	wire [15-1:0] node6565;
	wire [15-1:0] node6566;
	wire [15-1:0] node6569;
	wire [15-1:0] node6570;
	wire [15-1:0] node6571;
	wire [15-1:0] node6573;
	wire [15-1:0] node6578;
	wire [15-1:0] node6579;
	wire [15-1:0] node6580;
	wire [15-1:0] node6581;
	wire [15-1:0] node6585;
	wire [15-1:0] node6586;
	wire [15-1:0] node6590;
	wire [15-1:0] node6593;
	wire [15-1:0] node6594;
	wire [15-1:0] node6595;
	wire [15-1:0] node6596;
	wire [15-1:0] node6597;
	wire [15-1:0] node6599;
	wire [15-1:0] node6602;
	wire [15-1:0] node6603;
	wire [15-1:0] node6604;
	wire [15-1:0] node6608;
	wire [15-1:0] node6611;
	wire [15-1:0] node6612;
	wire [15-1:0] node6614;
	wire [15-1:0] node6615;
	wire [15-1:0] node6617;
	wire [15-1:0] node6620;
	wire [15-1:0] node6623;
	wire [15-1:0] node6624;
	wire [15-1:0] node6627;
	wire [15-1:0] node6629;
	wire [15-1:0] node6632;
	wire [15-1:0] node6633;
	wire [15-1:0] node6634;
	wire [15-1:0] node6635;
	wire [15-1:0] node6637;
	wire [15-1:0] node6641;
	wire [15-1:0] node6642;
	wire [15-1:0] node6643;
	wire [15-1:0] node6647;
	wire [15-1:0] node6650;
	wire [15-1:0] node6652;
	wire [15-1:0] node6653;
	wire [15-1:0] node6654;
	wire [15-1:0] node6657;
	wire [15-1:0] node6659;
	wire [15-1:0] node6663;
	wire [15-1:0] node6664;
	wire [15-1:0] node6665;
	wire [15-1:0] node6666;
	wire [15-1:0] node6667;
	wire [15-1:0] node6670;
	wire [15-1:0] node6673;
	wire [15-1:0] node6674;
	wire [15-1:0] node6678;
	wire [15-1:0] node6679;
	wire [15-1:0] node6683;
	wire [15-1:0] node6684;
	wire [15-1:0] node6685;
	wire [15-1:0] node6686;
	wire [15-1:0] node6690;
	wire [15-1:0] node6692;
	wire [15-1:0] node6695;
	wire [15-1:0] node6696;
	wire [15-1:0] node6697;
	wire [15-1:0] node6700;
	wire [15-1:0] node6703;
	wire [15-1:0] node6704;
	wire [15-1:0] node6708;
	wire [15-1:0] node6709;
	wire [15-1:0] node6710;
	wire [15-1:0] node6711;
	wire [15-1:0] node6712;
	wire [15-1:0] node6713;
	wire [15-1:0] node6714;
	wire [15-1:0] node6715;
	wire [15-1:0] node6717;
	wire [15-1:0] node6720;
	wire [15-1:0] node6723;
	wire [15-1:0] node6724;
	wire [15-1:0] node6725;
	wire [15-1:0] node6727;
	wire [15-1:0] node6731;
	wire [15-1:0] node6734;
	wire [15-1:0] node6735;
	wire [15-1:0] node6737;
	wire [15-1:0] node6741;
	wire [15-1:0] node6742;
	wire [15-1:0] node6743;
	wire [15-1:0] node6744;
	wire [15-1:0] node6746;
	wire [15-1:0] node6749;
	wire [15-1:0] node6751;
	wire [15-1:0] node6754;
	wire [15-1:0] node6755;
	wire [15-1:0] node6757;
	wire [15-1:0] node6758;
	wire [15-1:0] node6763;
	wire [15-1:0] node6764;
	wire [15-1:0] node6766;
	wire [15-1:0] node6769;
	wire [15-1:0] node6770;
	wire [15-1:0] node6774;
	wire [15-1:0] node6775;
	wire [15-1:0] node6776;
	wire [15-1:0] node6777;
	wire [15-1:0] node6778;
	wire [15-1:0] node6780;
	wire [15-1:0] node6784;
	wire [15-1:0] node6785;
	wire [15-1:0] node6789;
	wire [15-1:0] node6790;
	wire [15-1:0] node6792;
	wire [15-1:0] node6796;
	wire [15-1:0] node6797;
	wire [15-1:0] node6798;
	wire [15-1:0] node6799;
	wire [15-1:0] node6802;
	wire [15-1:0] node6805;
	wire [15-1:0] node6807;
	wire [15-1:0] node6810;
	wire [15-1:0] node6812;
	wire [15-1:0] node6813;
	wire [15-1:0] node6816;
	wire [15-1:0] node6817;
	wire [15-1:0] node6819;
	wire [15-1:0] node6823;
	wire [15-1:0] node6824;
	wire [15-1:0] node6825;
	wire [15-1:0] node6826;
	wire [15-1:0] node6827;
	wire [15-1:0] node6828;
	wire [15-1:0] node6831;
	wire [15-1:0] node6832;
	wire [15-1:0] node6836;
	wire [15-1:0] node6837;
	wire [15-1:0] node6841;
	wire [15-1:0] node6842;
	wire [15-1:0] node6843;
	wire [15-1:0] node6845;
	wire [15-1:0] node6847;
	wire [15-1:0] node6850;
	wire [15-1:0] node6851;
	wire [15-1:0] node6855;
	wire [15-1:0] node6857;
	wire [15-1:0] node6859;
	wire [15-1:0] node6862;
	wire [15-1:0] node6863;
	wire [15-1:0] node6864;
	wire [15-1:0] node6866;
	wire [15-1:0] node6867;
	wire [15-1:0] node6871;
	wire [15-1:0] node6872;
	wire [15-1:0] node6873;
	wire [15-1:0] node6877;
	wire [15-1:0] node6880;
	wire [15-1:0] node6881;
	wire [15-1:0] node6882;
	wire [15-1:0] node6885;
	wire [15-1:0] node6886;
	wire [15-1:0] node6888;
	wire [15-1:0] node6892;
	wire [15-1:0] node6893;
	wire [15-1:0] node6897;
	wire [15-1:0] node6898;
	wire [15-1:0] node6899;
	wire [15-1:0] node6900;
	wire [15-1:0] node6901;
	wire [15-1:0] node6902;
	wire [15-1:0] node6904;
	wire [15-1:0] node6908;
	wire [15-1:0] node6911;
	wire [15-1:0] node6912;
	wire [15-1:0] node6915;
	wire [15-1:0] node6918;
	wire [15-1:0] node6919;
	wire [15-1:0] node6920;
	wire [15-1:0] node6921;
	wire [15-1:0] node6925;
	wire [15-1:0] node6928;
	wire [15-1:0] node6929;
	wire [15-1:0] node6930;
	wire [15-1:0] node6934;
	wire [15-1:0] node6936;
	wire [15-1:0] node6939;
	wire [15-1:0] node6940;
	wire [15-1:0] node6941;
	wire [15-1:0] node6942;
	wire [15-1:0] node6945;
	wire [15-1:0] node6946;
	wire [15-1:0] node6948;
	wire [15-1:0] node6952;
	wire [15-1:0] node6953;
	wire [15-1:0] node6954;
	wire [15-1:0] node6958;
	wire [15-1:0] node6959;
	wire [15-1:0] node6961;
	wire [15-1:0] node6965;
	wire [15-1:0] node6966;
	wire [15-1:0] node6968;
	wire [15-1:0] node6971;
	wire [15-1:0] node6974;
	wire [15-1:0] node6975;
	wire [15-1:0] node6976;
	wire [15-1:0] node6977;
	wire [15-1:0] node6978;
	wire [15-1:0] node6979;
	wire [15-1:0] node6981;
	wire [15-1:0] node6983;
	wire [15-1:0] node6984;
	wire [15-1:0] node6988;
	wire [15-1:0] node6989;
	wire [15-1:0] node6990;
	wire [15-1:0] node6994;
	wire [15-1:0] node6997;
	wire [15-1:0] node6998;
	wire [15-1:0] node6999;
	wire [15-1:0] node7002;
	wire [15-1:0] node7004;
	wire [15-1:0] node7007;
	wire [15-1:0] node7008;
	wire [15-1:0] node7009;
	wire [15-1:0] node7011;
	wire [15-1:0] node7015;
	wire [15-1:0] node7018;
	wire [15-1:0] node7019;
	wire [15-1:0] node7020;
	wire [15-1:0] node7022;
	wire [15-1:0] node7024;
	wire [15-1:0] node7027;
	wire [15-1:0] node7028;
	wire [15-1:0] node7029;
	wire [15-1:0] node7034;
	wire [15-1:0] node7035;
	wire [15-1:0] node7036;
	wire [15-1:0] node7039;
	wire [15-1:0] node7042;
	wire [15-1:0] node7043;
	wire [15-1:0] node7046;
	wire [15-1:0] node7048;
	wire [15-1:0] node7051;
	wire [15-1:0] node7052;
	wire [15-1:0] node7053;
	wire [15-1:0] node7054;
	wire [15-1:0] node7055;
	wire [15-1:0] node7059;
	wire [15-1:0] node7060;
	wire [15-1:0] node7063;
	wire [15-1:0] node7066;
	wire [15-1:0] node7067;
	wire [15-1:0] node7069;
	wire [15-1:0] node7072;
	wire [15-1:0] node7073;
	wire [15-1:0] node7075;
	wire [15-1:0] node7076;
	wire [15-1:0] node7080;
	wire [15-1:0] node7083;
	wire [15-1:0] node7084;
	wire [15-1:0] node7085;
	wire [15-1:0] node7088;
	wire [15-1:0] node7089;
	wire [15-1:0] node7093;
	wire [15-1:0] node7094;
	wire [15-1:0] node7096;
	wire [15-1:0] node7099;
	wire [15-1:0] node7101;
	wire [15-1:0] node7103;
	wire [15-1:0] node7104;
	wire [15-1:0] node7108;
	wire [15-1:0] node7109;
	wire [15-1:0] node7110;
	wire [15-1:0] node7111;
	wire [15-1:0] node7112;
	wire [15-1:0] node7113;
	wire [15-1:0] node7117;
	wire [15-1:0] node7118;
	wire [15-1:0] node7121;
	wire [15-1:0] node7124;
	wire [15-1:0] node7125;
	wire [15-1:0] node7127;
	wire [15-1:0] node7130;
	wire [15-1:0] node7131;
	wire [15-1:0] node7132;
	wire [15-1:0] node7137;
	wire [15-1:0] node7138;
	wire [15-1:0] node7139;
	wire [15-1:0] node7140;
	wire [15-1:0] node7142;
	wire [15-1:0] node7146;
	wire [15-1:0] node7147;
	wire [15-1:0] node7148;
	wire [15-1:0] node7150;
	wire [15-1:0] node7154;
	wire [15-1:0] node7157;
	wire [15-1:0] node7158;
	wire [15-1:0] node7160;
	wire [15-1:0] node7161;
	wire [15-1:0] node7164;
	wire [15-1:0] node7168;
	wire [15-1:0] node7169;
	wire [15-1:0] node7170;
	wire [15-1:0] node7171;
	wire [15-1:0] node7172;
	wire [15-1:0] node7176;
	wire [15-1:0] node7177;
	wire [15-1:0] node7178;
	wire [15-1:0] node7180;
	wire [15-1:0] node7184;
	wire [15-1:0] node7187;
	wire [15-1:0] node7188;
	wire [15-1:0] node7189;
	wire [15-1:0] node7192;
	wire [15-1:0] node7194;
	wire [15-1:0] node7197;
	wire [15-1:0] node7198;
	wire [15-1:0] node7202;
	wire [15-1:0] node7203;
	wire [15-1:0] node7204;
	wire [15-1:0] node7206;
	wire [15-1:0] node7208;
	wire [15-1:0] node7211;
	wire [15-1:0] node7212;
	wire [15-1:0] node7215;
	wire [15-1:0] node7218;
	wire [15-1:0] node7219;
	wire [15-1:0] node7221;
	wire [15-1:0] node7223;
	wire [15-1:0] node7226;
	wire [15-1:0] node7227;
	wire [15-1:0] node7230;
	wire [15-1:0] node7233;
	wire [15-1:0] node7234;
	wire [15-1:0] node7235;
	wire [15-1:0] node7236;
	wire [15-1:0] node7237;
	wire [15-1:0] node7238;
	wire [15-1:0] node7239;
	wire [15-1:0] node7240;
	wire [15-1:0] node7241;
	wire [15-1:0] node7243;
	wire [15-1:0] node7246;
	wire [15-1:0] node7247;
	wire [15-1:0] node7251;
	wire [15-1:0] node7253;
	wire [15-1:0] node7255;
	wire [15-1:0] node7258;
	wire [15-1:0] node7259;
	wire [15-1:0] node7260;
	wire [15-1:0] node7262;
	wire [15-1:0] node7263;
	wire [15-1:0] node7268;
	wire [15-1:0] node7269;
	wire [15-1:0] node7270;
	wire [15-1:0] node7272;
	wire [15-1:0] node7277;
	wire [15-1:0] node7278;
	wire [15-1:0] node7279;
	wire [15-1:0] node7281;
	wire [15-1:0] node7284;
	wire [15-1:0] node7285;
	wire [15-1:0] node7286;
	wire [15-1:0] node7288;
	wire [15-1:0] node7292;
	wire [15-1:0] node7293;
	wire [15-1:0] node7295;
	wire [15-1:0] node7299;
	wire [15-1:0] node7300;
	wire [15-1:0] node7304;
	wire [15-1:0] node7305;
	wire [15-1:0] node7306;
	wire [15-1:0] node7307;
	wire [15-1:0] node7310;
	wire [15-1:0] node7311;
	wire [15-1:0] node7313;
	wire [15-1:0] node7314;
	wire [15-1:0] node7319;
	wire [15-1:0] node7320;
	wire [15-1:0] node7321;
	wire [15-1:0] node7323;
	wire [15-1:0] node7326;
	wire [15-1:0] node7327;
	wire [15-1:0] node7328;
	wire [15-1:0] node7333;
	wire [15-1:0] node7334;
	wire [15-1:0] node7337;
	wire [15-1:0] node7339;
	wire [15-1:0] node7341;
	wire [15-1:0] node7344;
	wire [15-1:0] node7345;
	wire [15-1:0] node7347;
	wire [15-1:0] node7348;
	wire [15-1:0] node7350;
	wire [15-1:0] node7353;
	wire [15-1:0] node7354;
	wire [15-1:0] node7355;
	wire [15-1:0] node7360;
	wire [15-1:0] node7363;
	wire [15-1:0] node7364;
	wire [15-1:0] node7365;
	wire [15-1:0] node7366;
	wire [15-1:0] node7367;
	wire [15-1:0] node7368;
	wire [15-1:0] node7369;
	wire [15-1:0] node7373;
	wire [15-1:0] node7376;
	wire [15-1:0] node7377;
	wire [15-1:0] node7379;
	wire [15-1:0] node7382;
	wire [15-1:0] node7384;
	wire [15-1:0] node7387;
	wire [15-1:0] node7388;
	wire [15-1:0] node7389;
	wire [15-1:0] node7392;
	wire [15-1:0] node7395;
	wire [15-1:0] node7396;
	wire [15-1:0] node7400;
	wire [15-1:0] node7401;
	wire [15-1:0] node7402;
	wire [15-1:0] node7403;
	wire [15-1:0] node7405;
	wire [15-1:0] node7407;
	wire [15-1:0] node7411;
	wire [15-1:0] node7413;
	wire [15-1:0] node7416;
	wire [15-1:0] node7417;
	wire [15-1:0] node7419;
	wire [15-1:0] node7422;
	wire [15-1:0] node7424;
	wire [15-1:0] node7427;
	wire [15-1:0] node7428;
	wire [15-1:0] node7429;
	wire [15-1:0] node7431;
	wire [15-1:0] node7432;
	wire [15-1:0] node7435;
	wire [15-1:0] node7438;
	wire [15-1:0] node7439;
	wire [15-1:0] node7441;
	wire [15-1:0] node7443;
	wire [15-1:0] node7444;
	wire [15-1:0] node7448;
	wire [15-1:0] node7449;
	wire [15-1:0] node7450;
	wire [15-1:0] node7455;
	wire [15-1:0] node7456;
	wire [15-1:0] node7457;
	wire [15-1:0] node7458;
	wire [15-1:0] node7461;
	wire [15-1:0] node7462;
	wire [15-1:0] node7466;
	wire [15-1:0] node7469;
	wire [15-1:0] node7470;
	wire [15-1:0] node7472;
	wire [15-1:0] node7474;
	wire [15-1:0] node7477;
	wire [15-1:0] node7479;
	wire [15-1:0] node7482;
	wire [15-1:0] node7483;
	wire [15-1:0] node7484;
	wire [15-1:0] node7485;
	wire [15-1:0] node7486;
	wire [15-1:0] node7487;
	wire [15-1:0] node7488;
	wire [15-1:0] node7492;
	wire [15-1:0] node7494;
	wire [15-1:0] node7495;
	wire [15-1:0] node7496;
	wire [15-1:0] node7501;
	wire [15-1:0] node7502;
	wire [15-1:0] node7503;
	wire [15-1:0] node7504;
	wire [15-1:0] node7506;
	wire [15-1:0] node7510;
	wire [15-1:0] node7511;
	wire [15-1:0] node7513;
	wire [15-1:0] node7517;
	wire [15-1:0] node7518;
	wire [15-1:0] node7521;
	wire [15-1:0] node7523;
	wire [15-1:0] node7525;
	wire [15-1:0] node7528;
	wire [15-1:0] node7529;
	wire [15-1:0] node7530;
	wire [15-1:0] node7532;
	wire [15-1:0] node7535;
	wire [15-1:0] node7536;
	wire [15-1:0] node7539;
	wire [15-1:0] node7540;
	wire [15-1:0] node7544;
	wire [15-1:0] node7545;
	wire [15-1:0] node7547;
	wire [15-1:0] node7551;
	wire [15-1:0] node7552;
	wire [15-1:0] node7553;
	wire [15-1:0] node7554;
	wire [15-1:0] node7556;
	wire [15-1:0] node7559;
	wire [15-1:0] node7560;
	wire [15-1:0] node7561;
	wire [15-1:0] node7565;
	wire [15-1:0] node7566;
	wire [15-1:0] node7568;
	wire [15-1:0] node7572;
	wire [15-1:0] node7574;
	wire [15-1:0] node7575;
	wire [15-1:0] node7576;
	wire [15-1:0] node7581;
	wire [15-1:0] node7582;
	wire [15-1:0] node7583;
	wire [15-1:0] node7584;
	wire [15-1:0] node7586;
	wire [15-1:0] node7589;
	wire [15-1:0] node7591;
	wire [15-1:0] node7593;
	wire [15-1:0] node7597;
	wire [15-1:0] node7598;
	wire [15-1:0] node7599;
	wire [15-1:0] node7603;
	wire [15-1:0] node7605;
	wire [15-1:0] node7608;
	wire [15-1:0] node7609;
	wire [15-1:0] node7610;
	wire [15-1:0] node7611;
	wire [15-1:0] node7612;
	wire [15-1:0] node7614;
	wire [15-1:0] node7617;
	wire [15-1:0] node7619;
	wire [15-1:0] node7620;
	wire [15-1:0] node7624;
	wire [15-1:0] node7625;
	wire [15-1:0] node7626;
	wire [15-1:0] node7627;
	wire [15-1:0] node7628;
	wire [15-1:0] node7632;
	wire [15-1:0] node7634;
	wire [15-1:0] node7638;
	wire [15-1:0] node7639;
	wire [15-1:0] node7642;
	wire [15-1:0] node7645;
	wire [15-1:0] node7646;
	wire [15-1:0] node7647;
	wire [15-1:0] node7650;
	wire [15-1:0] node7651;
	wire [15-1:0] node7653;
	wire [15-1:0] node7654;
	wire [15-1:0] node7657;
	wire [15-1:0] node7660;
	wire [15-1:0] node7661;
	wire [15-1:0] node7665;
	wire [15-1:0] node7666;
	wire [15-1:0] node7669;
	wire [15-1:0] node7670;
	wire [15-1:0] node7671;
	wire [15-1:0] node7673;
	wire [15-1:0] node7677;
	wire [15-1:0] node7679;
	wire [15-1:0] node7682;
	wire [15-1:0] node7683;
	wire [15-1:0] node7684;
	wire [15-1:0] node7685;
	wire [15-1:0] node7686;
	wire [15-1:0] node7691;
	wire [15-1:0] node7692;
	wire [15-1:0] node7693;
	wire [15-1:0] node7695;
	wire [15-1:0] node7698;
	wire [15-1:0] node7701;
	wire [15-1:0] node7702;
	wire [15-1:0] node7706;
	wire [15-1:0] node7707;
	wire [15-1:0] node7708;
	wire [15-1:0] node7709;
	wire [15-1:0] node7712;
	wire [15-1:0] node7713;
	wire [15-1:0] node7715;
	wire [15-1:0] node7719;
	wire [15-1:0] node7720;
	wire [15-1:0] node7722;
	wire [15-1:0] node7726;
	wire [15-1:0] node7728;
	wire [15-1:0] node7729;
	wire [15-1:0] node7730;
	wire [15-1:0] node7734;
	wire [15-1:0] node7735;
	wire [15-1:0] node7739;
	wire [15-1:0] node7740;
	wire [15-1:0] node7741;
	wire [15-1:0] node7742;
	wire [15-1:0] node7743;
	wire [15-1:0] node7744;
	wire [15-1:0] node7745;
	wire [15-1:0] node7746;
	wire [15-1:0] node7748;
	wire [15-1:0] node7752;
	wire [15-1:0] node7754;
	wire [15-1:0] node7757;
	wire [15-1:0] node7758;
	wire [15-1:0] node7759;
	wire [15-1:0] node7761;
	wire [15-1:0] node7764;
	wire [15-1:0] node7766;
	wire [15-1:0] node7769;
	wire [15-1:0] node7772;
	wire [15-1:0] node7773;
	wire [15-1:0] node7774;
	wire [15-1:0] node7775;
	wire [15-1:0] node7779;
	wire [15-1:0] node7780;
	wire [15-1:0] node7783;
	wire [15-1:0] node7786;
	wire [15-1:0] node7787;
	wire [15-1:0] node7790;
	wire [15-1:0] node7792;
	wire [15-1:0] node7794;
	wire [15-1:0] node7797;
	wire [15-1:0] node7798;
	wire [15-1:0] node7799;
	wire [15-1:0] node7800;
	wire [15-1:0] node7802;
	wire [15-1:0] node7804;
	wire [15-1:0] node7805;
	wire [15-1:0] node7809;
	wire [15-1:0] node7810;
	wire [15-1:0] node7811;
	wire [15-1:0] node7816;
	wire [15-1:0] node7818;
	wire [15-1:0] node7819;
	wire [15-1:0] node7821;
	wire [15-1:0] node7822;
	wire [15-1:0] node7826;
	wire [15-1:0] node7829;
	wire [15-1:0] node7830;
	wire [15-1:0] node7831;
	wire [15-1:0] node7834;
	wire [15-1:0] node7835;
	wire [15-1:0] node7839;
	wire [15-1:0] node7840;
	wire [15-1:0] node7841;
	wire [15-1:0] node7844;
	wire [15-1:0] node7846;
	wire [15-1:0] node7849;
	wire [15-1:0] node7850;
	wire [15-1:0] node7854;
	wire [15-1:0] node7855;
	wire [15-1:0] node7856;
	wire [15-1:0] node7857;
	wire [15-1:0] node7858;
	wire [15-1:0] node7859;
	wire [15-1:0] node7862;
	wire [15-1:0] node7865;
	wire [15-1:0] node7866;
	wire [15-1:0] node7870;
	wire [15-1:0] node7871;
	wire [15-1:0] node7872;
	wire [15-1:0] node7874;
	wire [15-1:0] node7878;
	wire [15-1:0] node7879;
	wire [15-1:0] node7881;
	wire [15-1:0] node7882;
	wire [15-1:0] node7886;
	wire [15-1:0] node7887;
	wire [15-1:0] node7891;
	wire [15-1:0] node7892;
	wire [15-1:0] node7893;
	wire [15-1:0] node7895;
	wire [15-1:0] node7899;
	wire [15-1:0] node7900;
	wire [15-1:0] node7901;
	wire [15-1:0] node7904;
	wire [15-1:0] node7907;
	wire [15-1:0] node7908;
	wire [15-1:0] node7912;
	wire [15-1:0] node7913;
	wire [15-1:0] node7914;
	wire [15-1:0] node7915;
	wire [15-1:0] node7916;
	wire [15-1:0] node7920;
	wire [15-1:0] node7921;
	wire [15-1:0] node7923;
	wire [15-1:0] node7926;
	wire [15-1:0] node7929;
	wire [15-1:0] node7930;
	wire [15-1:0] node7932;
	wire [15-1:0] node7935;
	wire [15-1:0] node7936;
	wire [15-1:0] node7937;
	wire [15-1:0] node7939;
	wire [15-1:0] node7943;
	wire [15-1:0] node7946;
	wire [15-1:0] node7947;
	wire [15-1:0] node7948;
	wire [15-1:0] node7949;
	wire [15-1:0] node7952;
	wire [15-1:0] node7955;
	wire [15-1:0] node7957;
	wire [15-1:0] node7960;
	wire [15-1:0] node7961;
	wire [15-1:0] node7963;
	wire [15-1:0] node7964;
	wire [15-1:0] node7966;
	wire [15-1:0] node7970;
	wire [15-1:0] node7971;
	wire [15-1:0] node7973;
	wire [15-1:0] node7974;
	wire [15-1:0] node7978;
	wire [15-1:0] node7981;
	wire [15-1:0] node7982;
	wire [15-1:0] node7983;
	wire [15-1:0] node7984;
	wire [15-1:0] node7985;
	wire [15-1:0] node7986;
	wire [15-1:0] node7987;
	wire [15-1:0] node7988;
	wire [15-1:0] node7993;
	wire [15-1:0] node7994;
	wire [15-1:0] node7998;
	wire [15-1:0] node7999;
	wire [15-1:0] node8000;
	wire [15-1:0] node8004;
	wire [15-1:0] node8007;
	wire [15-1:0] node8008;
	wire [15-1:0] node8010;
	wire [15-1:0] node8011;
	wire [15-1:0] node8012;
	wire [15-1:0] node8014;
	wire [15-1:0] node8018;
	wire [15-1:0] node8021;
	wire [15-1:0] node8023;
	wire [15-1:0] node8024;
	wire [15-1:0] node8027;
	wire [15-1:0] node8030;
	wire [15-1:0] node8031;
	wire [15-1:0] node8032;
	wire [15-1:0] node8034;
	wire [15-1:0] node8035;
	wire [15-1:0] node8037;
	wire [15-1:0] node8038;
	wire [15-1:0] node8043;
	wire [15-1:0] node8044;
	wire [15-1:0] node8045;
	wire [15-1:0] node8048;
	wire [15-1:0] node8050;
	wire [15-1:0] node8051;
	wire [15-1:0] node8055;
	wire [15-1:0] node8056;
	wire [15-1:0] node8059;
	wire [15-1:0] node8061;
	wire [15-1:0] node8064;
	wire [15-1:0] node8065;
	wire [15-1:0] node8066;
	wire [15-1:0] node8068;
	wire [15-1:0] node8071;
	wire [15-1:0] node8073;
	wire [15-1:0] node8076;
	wire [15-1:0] node8077;
	wire [15-1:0] node8079;
	wire [15-1:0] node8081;
	wire [15-1:0] node8085;
	wire [15-1:0] node8086;
	wire [15-1:0] node8087;
	wire [15-1:0] node8088;
	wire [15-1:0] node8089;
	wire [15-1:0] node8090;
	wire [15-1:0] node8094;
	wire [15-1:0] node8095;
	wire [15-1:0] node8097;
	wire [15-1:0] node8100;
	wire [15-1:0] node8102;
	wire [15-1:0] node8105;
	wire [15-1:0] node8106;
	wire [15-1:0] node8107;
	wire [15-1:0] node8111;
	wire [15-1:0] node8112;
	wire [15-1:0] node8114;
	wire [15-1:0] node8117;
	wire [15-1:0] node8119;
	wire [15-1:0] node8122;
	wire [15-1:0] node8123;
	wire [15-1:0] node8124;
	wire [15-1:0] node8125;
	wire [15-1:0] node8129;
	wire [15-1:0] node8130;
	wire [15-1:0] node8131;
	wire [15-1:0] node8135;
	wire [15-1:0] node8138;
	wire [15-1:0] node8139;
	wire [15-1:0] node8140;
	wire [15-1:0] node8143;
	wire [15-1:0] node8145;
	wire [15-1:0] node8148;
	wire [15-1:0] node8149;
	wire [15-1:0] node8151;
	wire [15-1:0] node8153;
	wire [15-1:0] node8156;
	wire [15-1:0] node8157;
	wire [15-1:0] node8158;
	wire [15-1:0] node8163;
	wire [15-1:0] node8164;
	wire [15-1:0] node8165;
	wire [15-1:0] node8166;
	wire [15-1:0] node8168;
	wire [15-1:0] node8170;
	wire [15-1:0] node8173;
	wire [15-1:0] node8174;
	wire [15-1:0] node8178;
	wire [15-1:0] node8179;
	wire [15-1:0] node8181;
	wire [15-1:0] node8184;
	wire [15-1:0] node8185;
	wire [15-1:0] node8186;
	wire [15-1:0] node8191;
	wire [15-1:0] node8192;
	wire [15-1:0] node8193;
	wire [15-1:0] node8194;
	wire [15-1:0] node8195;
	wire [15-1:0] node8199;
	wire [15-1:0] node8202;
	wire [15-1:0] node8203;
	wire [15-1:0] node8204;
	wire [15-1:0] node8208;
	wire [15-1:0] node8211;
	wire [15-1:0] node8212;
	wire [15-1:0] node8213;
	wire [15-1:0] node8216;
	wire [15-1:0] node8218;
	wire [15-1:0] node8219;
	wire [15-1:0] node8223;
	wire [15-1:0] node8224;
	wire [15-1:0] node8226;
	wire [15-1:0] node8227;
	wire [15-1:0] node8231;
	wire [15-1:0] node8233;
	wire [15-1:0] node8235;
	wire [15-1:0] node8238;
	wire [15-1:0] node8239;
	wire [15-1:0] node8240;
	wire [15-1:0] node8241;
	wire [15-1:0] node8242;
	wire [15-1:0] node8243;
	wire [15-1:0] node8244;
	wire [15-1:0] node8245;
	wire [15-1:0] node8246;
	wire [15-1:0] node8247;
	wire [15-1:0] node8248;
	wire [15-1:0] node8249;
	wire [15-1:0] node8252;
	wire [15-1:0] node8255;
	wire [15-1:0] node8256;
	wire [15-1:0] node8259;
	wire [15-1:0] node8260;
	wire [15-1:0] node8261;
	wire [15-1:0] node8266;
	wire [15-1:0] node8267;
	wire [15-1:0] node8268;
	wire [15-1:0] node8269;
	wire [15-1:0] node8273;
	wire [15-1:0] node8276;
	wire [15-1:0] node8278;
	wire [15-1:0] node8281;
	wire [15-1:0] node8282;
	wire [15-1:0] node8283;
	wire [15-1:0] node8284;
	wire [15-1:0] node8286;
	wire [15-1:0] node8287;
	wire [15-1:0] node8292;
	wire [15-1:0] node8293;
	wire [15-1:0] node8296;
	wire [15-1:0] node8298;
	wire [15-1:0] node8301;
	wire [15-1:0] node8303;
	wire [15-1:0] node8304;
	wire [15-1:0] node8305;
	wire [15-1:0] node8308;
	wire [15-1:0] node8309;
	wire [15-1:0] node8314;
	wire [15-1:0] node8315;
	wire [15-1:0] node8316;
	wire [15-1:0] node8317;
	wire [15-1:0] node8318;
	wire [15-1:0] node8321;
	wire [15-1:0] node8323;
	wire [15-1:0] node8326;
	wire [15-1:0] node8327;
	wire [15-1:0] node8331;
	wire [15-1:0] node8332;
	wire [15-1:0] node8333;
	wire [15-1:0] node8335;
	wire [15-1:0] node8338;
	wire [15-1:0] node8341;
	wire [15-1:0] node8342;
	wire [15-1:0] node8343;
	wire [15-1:0] node8347;
	wire [15-1:0] node8350;
	wire [15-1:0] node8351;
	wire [15-1:0] node8352;
	wire [15-1:0] node8355;
	wire [15-1:0] node8356;
	wire [15-1:0] node8359;
	wire [15-1:0] node8362;
	wire [15-1:0] node8363;
	wire [15-1:0] node8365;
	wire [15-1:0] node8368;
	wire [15-1:0] node8369;
	wire [15-1:0] node8371;
	wire [15-1:0] node8373;
	wire [15-1:0] node8376;
	wire [15-1:0] node8377;
	wire [15-1:0] node8381;
	wire [15-1:0] node8382;
	wire [15-1:0] node8383;
	wire [15-1:0] node8384;
	wire [15-1:0] node8385;
	wire [15-1:0] node8387;
	wire [15-1:0] node8389;
	wire [15-1:0] node8392;
	wire [15-1:0] node8393;
	wire [15-1:0] node8396;
	wire [15-1:0] node8399;
	wire [15-1:0] node8400;
	wire [15-1:0] node8401;
	wire [15-1:0] node8404;
	wire [15-1:0] node8407;
	wire [15-1:0] node8408;
	wire [15-1:0] node8410;
	wire [15-1:0] node8411;
	wire [15-1:0] node8415;
	wire [15-1:0] node8418;
	wire [15-1:0] node8419;
	wire [15-1:0] node8420;
	wire [15-1:0] node8421;
	wire [15-1:0] node8424;
	wire [15-1:0] node8427;
	wire [15-1:0] node8428;
	wire [15-1:0] node8430;
	wire [15-1:0] node8431;
	wire [15-1:0] node8435;
	wire [15-1:0] node8438;
	wire [15-1:0] node8439;
	wire [15-1:0] node8440;
	wire [15-1:0] node8441;
	wire [15-1:0] node8445;
	wire [15-1:0] node8448;
	wire [15-1:0] node8449;
	wire [15-1:0] node8453;
	wire [15-1:0] node8454;
	wire [15-1:0] node8455;
	wire [15-1:0] node8456;
	wire [15-1:0] node8457;
	wire [15-1:0] node8460;
	wire [15-1:0] node8461;
	wire [15-1:0] node8463;
	wire [15-1:0] node8467;
	wire [15-1:0] node8468;
	wire [15-1:0] node8469;
	wire [15-1:0] node8474;
	wire [15-1:0] node8475;
	wire [15-1:0] node8477;
	wire [15-1:0] node8479;
	wire [15-1:0] node8482;
	wire [15-1:0] node8483;
	wire [15-1:0] node8484;
	wire [15-1:0] node8486;
	wire [15-1:0] node8490;
	wire [15-1:0] node8493;
	wire [15-1:0] node8494;
	wire [15-1:0] node8495;
	wire [15-1:0] node8496;
	wire [15-1:0] node8497;
	wire [15-1:0] node8501;
	wire [15-1:0] node8503;
	wire [15-1:0] node8504;
	wire [15-1:0] node8508;
	wire [15-1:0] node8509;
	wire [15-1:0] node8513;
	wire [15-1:0] node8514;
	wire [15-1:0] node8517;
	wire [15-1:0] node8518;
	wire [15-1:0] node8519;
	wire [15-1:0] node8522;
	wire [15-1:0] node8523;
	wire [15-1:0] node8528;
	wire [15-1:0] node8529;
	wire [15-1:0] node8530;
	wire [15-1:0] node8531;
	wire [15-1:0] node8532;
	wire [15-1:0] node8533;
	wire [15-1:0] node8534;
	wire [15-1:0] node8535;
	wire [15-1:0] node8539;
	wire [15-1:0] node8540;
	wire [15-1:0] node8543;
	wire [15-1:0] node8544;
	wire [15-1:0] node8548;
	wire [15-1:0] node8549;
	wire [15-1:0] node8553;
	wire [15-1:0] node8554;
	wire [15-1:0] node8556;
	wire [15-1:0] node8557;
	wire [15-1:0] node8561;
	wire [15-1:0] node8562;
	wire [15-1:0] node8564;
	wire [15-1:0] node8567;
	wire [15-1:0] node8568;
	wire [15-1:0] node8572;
	wire [15-1:0] node8573;
	wire [15-1:0] node8574;
	wire [15-1:0] node8576;
	wire [15-1:0] node8579;
	wire [15-1:0] node8581;
	wire [15-1:0] node8584;
	wire [15-1:0] node8585;
	wire [15-1:0] node8586;
	wire [15-1:0] node8589;
	wire [15-1:0] node8592;
	wire [15-1:0] node8593;
	wire [15-1:0] node8597;
	wire [15-1:0] node8598;
	wire [15-1:0] node8599;
	wire [15-1:0] node8601;
	wire [15-1:0] node8602;
	wire [15-1:0] node8604;
	wire [15-1:0] node8605;
	wire [15-1:0] node8609;
	wire [15-1:0] node8612;
	wire [15-1:0] node8613;
	wire [15-1:0] node8614;
	wire [15-1:0] node8617;
	wire [15-1:0] node8618;
	wire [15-1:0] node8619;
	wire [15-1:0] node8622;
	wire [15-1:0] node8626;
	wire [15-1:0] node8627;
	wire [15-1:0] node8629;
	wire [15-1:0] node8632;
	wire [15-1:0] node8634;
	wire [15-1:0] node8637;
	wire [15-1:0] node8638;
	wire [15-1:0] node8639;
	wire [15-1:0] node8642;
	wire [15-1:0] node8643;
	wire [15-1:0] node8644;
	wire [15-1:0] node8648;
	wire [15-1:0] node8649;
	wire [15-1:0] node8653;
	wire [15-1:0] node8654;
	wire [15-1:0] node8655;
	wire [15-1:0] node8656;
	wire [15-1:0] node8660;
	wire [15-1:0] node8661;
	wire [15-1:0] node8665;
	wire [15-1:0] node8666;
	wire [15-1:0] node8668;
	wire [15-1:0] node8672;
	wire [15-1:0] node8673;
	wire [15-1:0] node8674;
	wire [15-1:0] node8675;
	wire [15-1:0] node8676;
	wire [15-1:0] node8678;
	wire [15-1:0] node8680;
	wire [15-1:0] node8683;
	wire [15-1:0] node8685;
	wire [15-1:0] node8688;
	wire [15-1:0] node8689;
	wire [15-1:0] node8691;
	wire [15-1:0] node8693;
	wire [15-1:0] node8696;
	wire [15-1:0] node8699;
	wire [15-1:0] node8700;
	wire [15-1:0] node8701;
	wire [15-1:0] node8702;
	wire [15-1:0] node8705;
	wire [15-1:0] node8707;
	wire [15-1:0] node8710;
	wire [15-1:0] node8711;
	wire [15-1:0] node8714;
	wire [15-1:0] node8715;
	wire [15-1:0] node8717;
	wire [15-1:0] node8721;
	wire [15-1:0] node8722;
	wire [15-1:0] node8723;
	wire [15-1:0] node8726;
	wire [15-1:0] node8729;
	wire [15-1:0] node8730;
	wire [15-1:0] node8734;
	wire [15-1:0] node8735;
	wire [15-1:0] node8736;
	wire [15-1:0] node8737;
	wire [15-1:0] node8739;
	wire [15-1:0] node8742;
	wire [15-1:0] node8743;
	wire [15-1:0] node8747;
	wire [15-1:0] node8748;
	wire [15-1:0] node8750;
	wire [15-1:0] node8753;
	wire [15-1:0] node8754;
	wire [15-1:0] node8757;
	wire [15-1:0] node8759;
	wire [15-1:0] node8762;
	wire [15-1:0] node8763;
	wire [15-1:0] node8764;
	wire [15-1:0] node8765;
	wire [15-1:0] node8769;
	wire [15-1:0] node8770;
	wire [15-1:0] node8773;
	wire [15-1:0] node8776;
	wire [15-1:0] node8777;
	wire [15-1:0] node8779;
	wire [15-1:0] node8782;
	wire [15-1:0] node8783;
	wire [15-1:0] node8785;
	wire [15-1:0] node8789;
	wire [15-1:0] node8790;
	wire [15-1:0] node8791;
	wire [15-1:0] node8792;
	wire [15-1:0] node8793;
	wire [15-1:0] node8794;
	wire [15-1:0] node8795;
	wire [15-1:0] node8796;
	wire [15-1:0] node8797;
	wire [15-1:0] node8799;
	wire [15-1:0] node8802;
	wire [15-1:0] node8804;
	wire [15-1:0] node8807;
	wire [15-1:0] node8810;
	wire [15-1:0] node8811;
	wire [15-1:0] node8814;
	wire [15-1:0] node8817;
	wire [15-1:0] node8818;
	wire [15-1:0] node8820;
	wire [15-1:0] node8823;
	wire [15-1:0] node8824;
	wire [15-1:0] node8826;
	wire [15-1:0] node8829;
	wire [15-1:0] node8832;
	wire [15-1:0] node8833;
	wire [15-1:0] node8834;
	wire [15-1:0] node8835;
	wire [15-1:0] node8839;
	wire [15-1:0] node8842;
	wire [15-1:0] node8843;
	wire [15-1:0] node8844;
	wire [15-1:0] node8845;
	wire [15-1:0] node8847;
	wire [15-1:0] node8852;
	wire [15-1:0] node8853;
	wire [15-1:0] node8857;
	wire [15-1:0] node8858;
	wire [15-1:0] node8859;
	wire [15-1:0] node8860;
	wire [15-1:0] node8861;
	wire [15-1:0] node8862;
	wire [15-1:0] node8866;
	wire [15-1:0] node8867;
	wire [15-1:0] node8869;
	wire [15-1:0] node8873;
	wire [15-1:0] node8874;
	wire [15-1:0] node8877;
	wire [15-1:0] node8880;
	wire [15-1:0] node8881;
	wire [15-1:0] node8883;
	wire [15-1:0] node8885;
	wire [15-1:0] node8888;
	wire [15-1:0] node8891;
	wire [15-1:0] node8892;
	wire [15-1:0] node8893;
	wire [15-1:0] node8894;
	wire [15-1:0] node8898;
	wire [15-1:0] node8899;
	wire [15-1:0] node8901;
	wire [15-1:0] node8902;
	wire [15-1:0] node8906;
	wire [15-1:0] node8907;
	wire [15-1:0] node8911;
	wire [15-1:0] node8912;
	wire [15-1:0] node8913;
	wire [15-1:0] node8916;
	wire [15-1:0] node8917;
	wire [15-1:0] node8920;
	wire [15-1:0] node8921;
	wire [15-1:0] node8925;
	wire [15-1:0] node8926;
	wire [15-1:0] node8930;
	wire [15-1:0] node8931;
	wire [15-1:0] node8932;
	wire [15-1:0] node8933;
	wire [15-1:0] node8934;
	wire [15-1:0] node8936;
	wire [15-1:0] node8939;
	wire [15-1:0] node8940;
	wire [15-1:0] node8942;
	wire [15-1:0] node8943;
	wire [15-1:0] node8948;
	wire [15-1:0] node8949;
	wire [15-1:0] node8950;
	wire [15-1:0] node8951;
	wire [15-1:0] node8955;
	wire [15-1:0] node8958;
	wire [15-1:0] node8959;
	wire [15-1:0] node8962;
	wire [15-1:0] node8964;
	wire [15-1:0] node8967;
	wire [15-1:0] node8968;
	wire [15-1:0] node8969;
	wire [15-1:0] node8971;
	wire [15-1:0] node8973;
	wire [15-1:0] node8976;
	wire [15-1:0] node8977;
	wire [15-1:0] node8979;
	wire [15-1:0] node8983;
	wire [15-1:0] node8984;
	wire [15-1:0] node8985;
	wire [15-1:0] node8989;
	wire [15-1:0] node8990;
	wire [15-1:0] node8994;
	wire [15-1:0] node8995;
	wire [15-1:0] node8996;
	wire [15-1:0] node8997;
	wire [15-1:0] node8998;
	wire [15-1:0] node8999;
	wire [15-1:0] node9003;
	wire [15-1:0] node9005;
	wire [15-1:0] node9006;
	wire [15-1:0] node9010;
	wire [15-1:0] node9011;
	wire [15-1:0] node9014;
	wire [15-1:0] node9017;
	wire [15-1:0] node9018;
	wire [15-1:0] node9019;
	wire [15-1:0] node9020;
	wire [15-1:0] node9025;
	wire [15-1:0] node9026;
	wire [15-1:0] node9029;
	wire [15-1:0] node9032;
	wire [15-1:0] node9033;
	wire [15-1:0] node9034;
	wire [15-1:0] node9035;
	wire [15-1:0] node9037;
	wire [15-1:0] node9038;
	wire [15-1:0] node9042;
	wire [15-1:0] node9043;
	wire [15-1:0] node9045;
	wire [15-1:0] node9049;
	wire [15-1:0] node9051;
	wire [15-1:0] node9054;
	wire [15-1:0] node9055;
	wire [15-1:0] node9056;
	wire [15-1:0] node9058;
	wire [15-1:0] node9061;
	wire [15-1:0] node9062;
	wire [15-1:0] node9066;
	wire [15-1:0] node9067;
	wire [15-1:0] node9068;
	wire [15-1:0] node9072;
	wire [15-1:0] node9074;
	wire [15-1:0] node9077;
	wire [15-1:0] node9078;
	wire [15-1:0] node9079;
	wire [15-1:0] node9080;
	wire [15-1:0] node9081;
	wire [15-1:0] node9082;
	wire [15-1:0] node9083;
	wire [15-1:0] node9086;
	wire [15-1:0] node9089;
	wire [15-1:0] node9091;
	wire [15-1:0] node9092;
	wire [15-1:0] node9093;
	wire [15-1:0] node9097;
	wire [15-1:0] node9100;
	wire [15-1:0] node9101;
	wire [15-1:0] node9102;
	wire [15-1:0] node9105;
	wire [15-1:0] node9108;
	wire [15-1:0] node9109;
	wire [15-1:0] node9113;
	wire [15-1:0] node9114;
	wire [15-1:0] node9115;
	wire [15-1:0] node9116;
	wire [15-1:0] node9119;
	wire [15-1:0] node9122;
	wire [15-1:0] node9123;
	wire [15-1:0] node9125;
	wire [15-1:0] node9128;
	wire [15-1:0] node9130;
	wire [15-1:0] node9131;
	wire [15-1:0] node9135;
	wire [15-1:0] node9136;
	wire [15-1:0] node9138;
	wire [15-1:0] node9140;
	wire [15-1:0] node9143;
	wire [15-1:0] node9144;
	wire [15-1:0] node9148;
	wire [15-1:0] node9149;
	wire [15-1:0] node9150;
	wire [15-1:0] node9151;
	wire [15-1:0] node9152;
	wire [15-1:0] node9155;
	wire [15-1:0] node9158;
	wire [15-1:0] node9159;
	wire [15-1:0] node9162;
	wire [15-1:0] node9163;
	wire [15-1:0] node9165;
	wire [15-1:0] node9169;
	wire [15-1:0] node9170;
	wire [15-1:0] node9171;
	wire [15-1:0] node9174;
	wire [15-1:0] node9177;
	wire [15-1:0] node9179;
	wire [15-1:0] node9182;
	wire [15-1:0] node9183;
	wire [15-1:0] node9184;
	wire [15-1:0] node9185;
	wire [15-1:0] node9188;
	wire [15-1:0] node9189;
	wire [15-1:0] node9191;
	wire [15-1:0] node9195;
	wire [15-1:0] node9198;
	wire [15-1:0] node9199;
	wire [15-1:0] node9200;
	wire [15-1:0] node9203;
	wire [15-1:0] node9204;
	wire [15-1:0] node9206;
	wire [15-1:0] node9210;
	wire [15-1:0] node9211;
	wire [15-1:0] node9212;
	wire [15-1:0] node9216;
	wire [15-1:0] node9219;
	wire [15-1:0] node9220;
	wire [15-1:0] node9221;
	wire [15-1:0] node9222;
	wire [15-1:0] node9223;
	wire [15-1:0] node9226;
	wire [15-1:0] node9227;
	wire [15-1:0] node9231;
	wire [15-1:0] node9233;
	wire [15-1:0] node9234;
	wire [15-1:0] node9236;
	wire [15-1:0] node9239;
	wire [15-1:0] node9242;
	wire [15-1:0] node9243;
	wire [15-1:0] node9244;
	wire [15-1:0] node9245;
	wire [15-1:0] node9246;
	wire [15-1:0] node9250;
	wire [15-1:0] node9253;
	wire [15-1:0] node9254;
	wire [15-1:0] node9258;
	wire [15-1:0] node9259;
	wire [15-1:0] node9260;
	wire [15-1:0] node9263;
	wire [15-1:0] node9266;
	wire [15-1:0] node9268;
	wire [15-1:0] node9271;
	wire [15-1:0] node9272;
	wire [15-1:0] node9273;
	wire [15-1:0] node9274;
	wire [15-1:0] node9276;
	wire [15-1:0] node9279;
	wire [15-1:0] node9280;
	wire [15-1:0] node9281;
	wire [15-1:0] node9286;
	wire [15-1:0] node9287;
	wire [15-1:0] node9289;
	wire [15-1:0] node9292;
	wire [15-1:0] node9294;
	wire [15-1:0] node9297;
	wire [15-1:0] node9298;
	wire [15-1:0] node9299;
	wire [15-1:0] node9301;
	wire [15-1:0] node9304;
	wire [15-1:0] node9305;
	wire [15-1:0] node9307;
	wire [15-1:0] node9310;
	wire [15-1:0] node9311;
	wire [15-1:0] node9312;
	wire [15-1:0] node9316;
	wire [15-1:0] node9319;
	wire [15-1:0] node9320;
	wire [15-1:0] node9321;
	wire [15-1:0] node9322;
	wire [15-1:0] node9326;
	wire [15-1:0] node9329;
	wire [15-1:0] node9330;
	wire [15-1:0] node9331;
	wire [15-1:0] node9334;
	wire [15-1:0] node9336;
	wire [15-1:0] node9339;
	wire [15-1:0] node9340;
	wire [15-1:0] node9344;
	wire [15-1:0] node9345;
	wire [15-1:0] node9346;
	wire [15-1:0] node9347;
	wire [15-1:0] node9348;
	wire [15-1:0] node9349;
	wire [15-1:0] node9350;
	wire [15-1:0] node9351;
	wire [15-1:0] node9353;
	wire [15-1:0] node9354;
	wire [15-1:0] node9358;
	wire [15-1:0] node9359;
	wire [15-1:0] node9360;
	wire [15-1:0] node9361;
	wire [15-1:0] node9367;
	wire [15-1:0] node9368;
	wire [15-1:0] node9369;
	wire [15-1:0] node9370;
	wire [15-1:0] node9373;
	wire [15-1:0] node9374;
	wire [15-1:0] node9379;
	wire [15-1:0] node9380;
	wire [15-1:0] node9384;
	wire [15-1:0] node9385;
	wire [15-1:0] node9386;
	wire [15-1:0] node9387;
	wire [15-1:0] node9390;
	wire [15-1:0] node9392;
	wire [15-1:0] node9393;
	wire [15-1:0] node9397;
	wire [15-1:0] node9398;
	wire [15-1:0] node9401;
	wire [15-1:0] node9403;
	wire [15-1:0] node9406;
	wire [15-1:0] node9407;
	wire [15-1:0] node9408;
	wire [15-1:0] node9409;
	wire [15-1:0] node9414;
	wire [15-1:0] node9415;
	wire [15-1:0] node9416;
	wire [15-1:0] node9421;
	wire [15-1:0] node9422;
	wire [15-1:0] node9423;
	wire [15-1:0] node9424;
	wire [15-1:0] node9426;
	wire [15-1:0] node9428;
	wire [15-1:0] node9431;
	wire [15-1:0] node9432;
	wire [15-1:0] node9435;
	wire [15-1:0] node9437;
	wire [15-1:0] node9438;
	wire [15-1:0] node9442;
	wire [15-1:0] node9443;
	wire [15-1:0] node9444;
	wire [15-1:0] node9445;
	wire [15-1:0] node9450;
	wire [15-1:0] node9451;
	wire [15-1:0] node9454;
	wire [15-1:0] node9457;
	wire [15-1:0] node9458;
	wire [15-1:0] node9459;
	wire [15-1:0] node9460;
	wire [15-1:0] node9464;
	wire [15-1:0] node9465;
	wire [15-1:0] node9466;
	wire [15-1:0] node9471;
	wire [15-1:0] node9472;
	wire [15-1:0] node9474;
	wire [15-1:0] node9477;
	wire [15-1:0] node9478;
	wire [15-1:0] node9481;
	wire [15-1:0] node9483;
	wire [15-1:0] node9486;
	wire [15-1:0] node9487;
	wire [15-1:0] node9488;
	wire [15-1:0] node9489;
	wire [15-1:0] node9490;
	wire [15-1:0] node9491;
	wire [15-1:0] node9492;
	wire [15-1:0] node9494;
	wire [15-1:0] node9499;
	wire [15-1:0] node9501;
	wire [15-1:0] node9502;
	wire [15-1:0] node9506;
	wire [15-1:0] node9508;
	wire [15-1:0] node9510;
	wire [15-1:0] node9511;
	wire [15-1:0] node9512;
	wire [15-1:0] node9517;
	wire [15-1:0] node9518;
	wire [15-1:0] node9519;
	wire [15-1:0] node9520;
	wire [15-1:0] node9525;
	wire [15-1:0] node9527;
	wire [15-1:0] node9528;
	wire [15-1:0] node9530;
	wire [15-1:0] node9534;
	wire [15-1:0] node9535;
	wire [15-1:0] node9536;
	wire [15-1:0] node9537;
	wire [15-1:0] node9539;
	wire [15-1:0] node9541;
	wire [15-1:0] node9542;
	wire [15-1:0] node9546;
	wire [15-1:0] node9549;
	wire [15-1:0] node9550;
	wire [15-1:0] node9551;
	wire [15-1:0] node9552;
	wire [15-1:0] node9556;
	wire [15-1:0] node9559;
	wire [15-1:0] node9560;
	wire [15-1:0] node9561;
	wire [15-1:0] node9565;
	wire [15-1:0] node9567;
	wire [15-1:0] node9568;
	wire [15-1:0] node9572;
	wire [15-1:0] node9573;
	wire [15-1:0] node9574;
	wire [15-1:0] node9576;
	wire [15-1:0] node9580;
	wire [15-1:0] node9581;
	wire [15-1:0] node9582;
	wire [15-1:0] node9583;
	wire [15-1:0] node9587;
	wire [15-1:0] node9590;
	wire [15-1:0] node9592;
	wire [15-1:0] node9594;
	wire [15-1:0] node9597;
	wire [15-1:0] node9598;
	wire [15-1:0] node9599;
	wire [15-1:0] node9600;
	wire [15-1:0] node9601;
	wire [15-1:0] node9602;
	wire [15-1:0] node9603;
	wire [15-1:0] node9605;
	wire [15-1:0] node9606;
	wire [15-1:0] node9610;
	wire [15-1:0] node9612;
	wire [15-1:0] node9615;
	wire [15-1:0] node9616;
	wire [15-1:0] node9619;
	wire [15-1:0] node9622;
	wire [15-1:0] node9623;
	wire [15-1:0] node9624;
	wire [15-1:0] node9627;
	wire [15-1:0] node9629;
	wire [15-1:0] node9632;
	wire [15-1:0] node9633;
	wire [15-1:0] node9634;
	wire [15-1:0] node9639;
	wire [15-1:0] node9640;
	wire [15-1:0] node9641;
	wire [15-1:0] node9643;
	wire [15-1:0] node9645;
	wire [15-1:0] node9648;
	wire [15-1:0] node9649;
	wire [15-1:0] node9650;
	wire [15-1:0] node9655;
	wire [15-1:0] node9656;
	wire [15-1:0] node9658;
	wire [15-1:0] node9661;
	wire [15-1:0] node9662;
	wire [15-1:0] node9663;
	wire [15-1:0] node9667;
	wire [15-1:0] node9670;
	wire [15-1:0] node9671;
	wire [15-1:0] node9672;
	wire [15-1:0] node9673;
	wire [15-1:0] node9674;
	wire [15-1:0] node9676;
	wire [15-1:0] node9679;
	wire [15-1:0] node9682;
	wire [15-1:0] node9683;
	wire [15-1:0] node9687;
	wire [15-1:0] node9688;
	wire [15-1:0] node9690;
	wire [15-1:0] node9693;
	wire [15-1:0] node9695;
	wire [15-1:0] node9697;
	wire [15-1:0] node9700;
	wire [15-1:0] node9701;
	wire [15-1:0] node9702;
	wire [15-1:0] node9703;
	wire [15-1:0] node9704;
	wire [15-1:0] node9708;
	wire [15-1:0] node9709;
	wire [15-1:0] node9713;
	wire [15-1:0] node9716;
	wire [15-1:0] node9717;
	wire [15-1:0] node9718;
	wire [15-1:0] node9721;
	wire [15-1:0] node9722;
	wire [15-1:0] node9726;
	wire [15-1:0] node9728;
	wire [15-1:0] node9731;
	wire [15-1:0] node9732;
	wire [15-1:0] node9733;
	wire [15-1:0] node9734;
	wire [15-1:0] node9735;
	wire [15-1:0] node9736;
	wire [15-1:0] node9737;
	wire [15-1:0] node9742;
	wire [15-1:0] node9743;
	wire [15-1:0] node9746;
	wire [15-1:0] node9748;
	wire [15-1:0] node9751;
	wire [15-1:0] node9752;
	wire [15-1:0] node9753;
	wire [15-1:0] node9756;
	wire [15-1:0] node9758;
	wire [15-1:0] node9761;
	wire [15-1:0] node9762;
	wire [15-1:0] node9763;
	wire [15-1:0] node9768;
	wire [15-1:0] node9769;
	wire [15-1:0] node9771;
	wire [15-1:0] node9772;
	wire [15-1:0] node9776;
	wire [15-1:0] node9777;
	wire [15-1:0] node9778;
	wire [15-1:0] node9781;
	wire [15-1:0] node9782;
	wire [15-1:0] node9786;
	wire [15-1:0] node9788;
	wire [15-1:0] node9789;
	wire [15-1:0] node9793;
	wire [15-1:0] node9794;
	wire [15-1:0] node9795;
	wire [15-1:0] node9796;
	wire [15-1:0] node9797;
	wire [15-1:0] node9800;
	wire [15-1:0] node9801;
	wire [15-1:0] node9803;
	wire [15-1:0] node9806;
	wire [15-1:0] node9808;
	wire [15-1:0] node9811;
	wire [15-1:0] node9812;
	wire [15-1:0] node9815;
	wire [15-1:0] node9817;
	wire [15-1:0] node9818;
	wire [15-1:0] node9822;
	wire [15-1:0] node9823;
	wire [15-1:0] node9825;
	wire [15-1:0] node9827;
	wire [15-1:0] node9830;
	wire [15-1:0] node9832;
	wire [15-1:0] node9835;
	wire [15-1:0] node9836;
	wire [15-1:0] node9837;
	wire [15-1:0] node9839;
	wire [15-1:0] node9842;
	wire [15-1:0] node9843;
	wire [15-1:0] node9844;
	wire [15-1:0] node9848;
	wire [15-1:0] node9849;
	wire [15-1:0] node9853;
	wire [15-1:0] node9854;
	wire [15-1:0] node9855;
	wire [15-1:0] node9859;
	wire [15-1:0] node9860;
	wire [15-1:0] node9863;
	wire [15-1:0] node9865;
	wire [15-1:0] node9867;
	wire [15-1:0] node9870;
	wire [15-1:0] node9871;
	wire [15-1:0] node9872;
	wire [15-1:0] node9873;
	wire [15-1:0] node9874;
	wire [15-1:0] node9875;
	wire [15-1:0] node9876;
	wire [15-1:0] node9877;
	wire [15-1:0] node9878;
	wire [15-1:0] node9882;
	wire [15-1:0] node9884;
	wire [15-1:0] node9887;
	wire [15-1:0] node9888;
	wire [15-1:0] node9891;
	wire [15-1:0] node9894;
	wire [15-1:0] node9895;
	wire [15-1:0] node9896;
	wire [15-1:0] node9897;
	wire [15-1:0] node9901;
	wire [15-1:0] node9904;
	wire [15-1:0] node9905;
	wire [15-1:0] node9906;
	wire [15-1:0] node9911;
	wire [15-1:0] node9912;
	wire [15-1:0] node9913;
	wire [15-1:0] node9914;
	wire [15-1:0] node9917;
	wire [15-1:0] node9918;
	wire [15-1:0] node9919;
	wire [15-1:0] node9922;
	wire [15-1:0] node9926;
	wire [15-1:0] node9927;
	wire [15-1:0] node9928;
	wire [15-1:0] node9930;
	wire [15-1:0] node9933;
	wire [15-1:0] node9934;
	wire [15-1:0] node9938;
	wire [15-1:0] node9941;
	wire [15-1:0] node9942;
	wire [15-1:0] node9944;
	wire [15-1:0] node9945;
	wire [15-1:0] node9947;
	wire [15-1:0] node9951;
	wire [15-1:0] node9952;
	wire [15-1:0] node9953;
	wire [15-1:0] node9955;
	wire [15-1:0] node9958;
	wire [15-1:0] node9961;
	wire [15-1:0] node9964;
	wire [15-1:0] node9965;
	wire [15-1:0] node9966;
	wire [15-1:0] node9967;
	wire [15-1:0] node9970;
	wire [15-1:0] node9973;
	wire [15-1:0] node9974;
	wire [15-1:0] node9975;
	wire [15-1:0] node9976;
	wire [15-1:0] node9980;
	wire [15-1:0] node9982;
	wire [15-1:0] node9983;
	wire [15-1:0] node9987;
	wire [15-1:0] node9988;
	wire [15-1:0] node9990;
	wire [15-1:0] node9991;
	wire [15-1:0] node9995;
	wire [15-1:0] node9998;
	wire [15-1:0] node9999;
	wire [15-1:0] node10000;
	wire [15-1:0] node10001;
	wire [15-1:0] node10002;
	wire [15-1:0] node10006;
	wire [15-1:0] node10007;
	wire [15-1:0] node10012;
	wire [15-1:0] node10013;
	wire [15-1:0] node10016;
	wire [15-1:0] node10017;
	wire [15-1:0] node10018;
	wire [15-1:0] node10020;
	wire [15-1:0] node10024;
	wire [15-1:0] node10025;
	wire [15-1:0] node10026;
	wire [15-1:0] node10031;
	wire [15-1:0] node10032;
	wire [15-1:0] node10033;
	wire [15-1:0] node10034;
	wire [15-1:0] node10035;
	wire [15-1:0] node10036;
	wire [15-1:0] node10039;
	wire [15-1:0] node10042;
	wire [15-1:0] node10043;
	wire [15-1:0] node10047;
	wire [15-1:0] node10048;
	wire [15-1:0] node10051;
	wire [15-1:0] node10052;
	wire [15-1:0] node10054;
	wire [15-1:0] node10058;
	wire [15-1:0] node10059;
	wire [15-1:0] node10060;
	wire [15-1:0] node10062;
	wire [15-1:0] node10065;
	wire [15-1:0] node10067;
	wire [15-1:0] node10068;
	wire [15-1:0] node10072;
	wire [15-1:0] node10073;
	wire [15-1:0] node10074;
	wire [15-1:0] node10075;
	wire [15-1:0] node10077;
	wire [15-1:0] node10081;
	wire [15-1:0] node10084;
	wire [15-1:0] node10085;
	wire [15-1:0] node10086;
	wire [15-1:0] node10091;
	wire [15-1:0] node10092;
	wire [15-1:0] node10093;
	wire [15-1:0] node10094;
	wire [15-1:0] node10095;
	wire [15-1:0] node10096;
	wire [15-1:0] node10101;
	wire [15-1:0] node10102;
	wire [15-1:0] node10106;
	wire [15-1:0] node10108;
	wire [15-1:0] node10110;
	wire [15-1:0] node10113;
	wire [15-1:0] node10114;
	wire [15-1:0] node10115;
	wire [15-1:0] node10116;
	wire [15-1:0] node10119;
	wire [15-1:0] node10122;
	wire [15-1:0] node10123;
	wire [15-1:0] node10124;
	wire [15-1:0] node10128;
	wire [15-1:0] node10131;
	wire [15-1:0] node10132;
	wire [15-1:0] node10133;
	wire [15-1:0] node10136;
	wire [15-1:0] node10138;
	wire [15-1:0] node10140;
	wire [15-1:0] node10143;
	wire [15-1:0] node10144;
	wire [15-1:0] node10146;
	wire [15-1:0] node10147;
	wire [15-1:0] node10151;
	wire [15-1:0] node10154;
	wire [15-1:0] node10155;
	wire [15-1:0] node10156;
	wire [15-1:0] node10157;
	wire [15-1:0] node10158;
	wire [15-1:0] node10159;
	wire [15-1:0] node10161;
	wire [15-1:0] node10162;
	wire [15-1:0] node10164;
	wire [15-1:0] node10169;
	wire [15-1:0] node10170;
	wire [15-1:0] node10171;
	wire [15-1:0] node10173;
	wire [15-1:0] node10174;
	wire [15-1:0] node10178;
	wire [15-1:0] node10181;
	wire [15-1:0] node10182;
	wire [15-1:0] node10185;
	wire [15-1:0] node10188;
	wire [15-1:0] node10189;
	wire [15-1:0] node10190;
	wire [15-1:0] node10191;
	wire [15-1:0] node10193;
	wire [15-1:0] node10194;
	wire [15-1:0] node10199;
	wire [15-1:0] node10200;
	wire [15-1:0] node10204;
	wire [15-1:0] node10205;
	wire [15-1:0] node10207;
	wire [15-1:0] node10209;
	wire [15-1:0] node10210;
	wire [15-1:0] node10214;
	wire [15-1:0] node10216;
	wire [15-1:0] node10217;
	wire [15-1:0] node10221;
	wire [15-1:0] node10222;
	wire [15-1:0] node10223;
	wire [15-1:0] node10224;
	wire [15-1:0] node10226;
	wire [15-1:0] node10227;
	wire [15-1:0] node10228;
	wire [15-1:0] node10233;
	wire [15-1:0] node10234;
	wire [15-1:0] node10237;
	wire [15-1:0] node10239;
	wire [15-1:0] node10242;
	wire [15-1:0] node10243;
	wire [15-1:0] node10245;
	wire [15-1:0] node10248;
	wire [15-1:0] node10249;
	wire [15-1:0] node10251;
	wire [15-1:0] node10255;
	wire [15-1:0] node10256;
	wire [15-1:0] node10257;
	wire [15-1:0] node10259;
	wire [15-1:0] node10261;
	wire [15-1:0] node10262;
	wire [15-1:0] node10266;
	wire [15-1:0] node10267;
	wire [15-1:0] node10271;
	wire [15-1:0] node10272;
	wire [15-1:0] node10273;
	wire [15-1:0] node10276;
	wire [15-1:0] node10279;
	wire [15-1:0] node10280;
	wire [15-1:0] node10282;
	wire [15-1:0] node10286;
	wire [15-1:0] node10287;
	wire [15-1:0] node10288;
	wire [15-1:0] node10289;
	wire [15-1:0] node10290;
	wire [15-1:0] node10291;
	wire [15-1:0] node10295;
	wire [15-1:0] node10296;
	wire [15-1:0] node10298;
	wire [15-1:0] node10301;
	wire [15-1:0] node10302;
	wire [15-1:0] node10306;
	wire [15-1:0] node10307;
	wire [15-1:0] node10308;
	wire [15-1:0] node10311;
	wire [15-1:0] node10314;
	wire [15-1:0] node10315;
	wire [15-1:0] node10317;
	wire [15-1:0] node10320;
	wire [15-1:0] node10323;
	wire [15-1:0] node10324;
	wire [15-1:0] node10325;
	wire [15-1:0] node10326;
	wire [15-1:0] node10330;
	wire [15-1:0] node10332;
	wire [15-1:0] node10335;
	wire [15-1:0] node10336;
	wire [15-1:0] node10337;
	wire [15-1:0] node10339;
	wire [15-1:0] node10343;
	wire [15-1:0] node10345;
	wire [15-1:0] node10348;
	wire [15-1:0] node10349;
	wire [15-1:0] node10350;
	wire [15-1:0] node10351;
	wire [15-1:0] node10352;
	wire [15-1:0] node10356;
	wire [15-1:0] node10357;
	wire [15-1:0] node10361;
	wire [15-1:0] node10362;
	wire [15-1:0] node10365;
	wire [15-1:0] node10366;
	wire [15-1:0] node10367;
	wire [15-1:0] node10371;
	wire [15-1:0] node10374;
	wire [15-1:0] node10375;
	wire [15-1:0] node10376;
	wire [15-1:0] node10377;
	wire [15-1:0] node10379;
	wire [15-1:0] node10380;
	wire [15-1:0] node10384;
	wire [15-1:0] node10387;
	wire [15-1:0] node10388;
	wire [15-1:0] node10391;
	wire [15-1:0] node10394;
	wire [15-1:0] node10395;
	wire [15-1:0] node10396;
	wire [15-1:0] node10397;
	wire [15-1:0] node10401;
	wire [15-1:0] node10403;
	wire [15-1:0] node10404;
	wire [15-1:0] node10408;
	wire [15-1:0] node10409;
	wire [15-1:0] node10412;
	wire [15-1:0] node10414;
	wire [15-1:0] node10415;
	wire [15-1:0] node10419;
	wire [15-1:0] node10420;
	wire [15-1:0] node10421;
	wire [15-1:0] node10422;
	wire [15-1:0] node10423;
	wire [15-1:0] node10424;
	wire [15-1:0] node10425;
	wire [15-1:0] node10426;
	wire [15-1:0] node10427;
	wire [15-1:0] node10428;
	wire [15-1:0] node10430;
	wire [15-1:0] node10431;
	wire [15-1:0] node10435;
	wire [15-1:0] node10438;
	wire [15-1:0] node10440;
	wire [15-1:0] node10443;
	wire [15-1:0] node10444;
	wire [15-1:0] node10445;
	wire [15-1:0] node10449;
	wire [15-1:0] node10450;
	wire [15-1:0] node10452;
	wire [15-1:0] node10453;
	wire [15-1:0] node10457;
	wire [15-1:0] node10458;
	wire [15-1:0] node10459;
	wire [15-1:0] node10464;
	wire [15-1:0] node10465;
	wire [15-1:0] node10466;
	wire [15-1:0] node10467;
	wire [15-1:0] node10470;
	wire [15-1:0] node10471;
	wire [15-1:0] node10475;
	wire [15-1:0] node10477;
	wire [15-1:0] node10480;
	wire [15-1:0] node10481;
	wire [15-1:0] node10482;
	wire [15-1:0] node10485;
	wire [15-1:0] node10488;
	wire [15-1:0] node10490;
	wire [15-1:0] node10493;
	wire [15-1:0] node10494;
	wire [15-1:0] node10495;
	wire [15-1:0] node10496;
	wire [15-1:0] node10497;
	wire [15-1:0] node10498;
	wire [15-1:0] node10500;
	wire [15-1:0] node10504;
	wire [15-1:0] node10507;
	wire [15-1:0] node10509;
	wire [15-1:0] node10510;
	wire [15-1:0] node10513;
	wire [15-1:0] node10514;
	wire [15-1:0] node10518;
	wire [15-1:0] node10519;
	wire [15-1:0] node10520;
	wire [15-1:0] node10523;
	wire [15-1:0] node10526;
	wire [15-1:0] node10527;
	wire [15-1:0] node10528;
	wire [15-1:0] node10531;
	wire [15-1:0] node10533;
	wire [15-1:0] node10537;
	wire [15-1:0] node10538;
	wire [15-1:0] node10539;
	wire [15-1:0] node10541;
	wire [15-1:0] node10544;
	wire [15-1:0] node10546;
	wire [15-1:0] node10547;
	wire [15-1:0] node10551;
	wire [15-1:0] node10553;
	wire [15-1:0] node10554;
	wire [15-1:0] node10556;
	wire [15-1:0] node10557;
	wire [15-1:0] node10561;
	wire [15-1:0] node10564;
	wire [15-1:0] node10565;
	wire [15-1:0] node10566;
	wire [15-1:0] node10567;
	wire [15-1:0] node10568;
	wire [15-1:0] node10570;
	wire [15-1:0] node10573;
	wire [15-1:0] node10574;
	wire [15-1:0] node10577;
	wire [15-1:0] node10579;
	wire [15-1:0] node10582;
	wire [15-1:0] node10583;
	wire [15-1:0] node10586;
	wire [15-1:0] node10587;
	wire [15-1:0] node10589;
	wire [15-1:0] node10593;
	wire [15-1:0] node10594;
	wire [15-1:0] node10595;
	wire [15-1:0] node10596;
	wire [15-1:0] node10599;
	wire [15-1:0] node10602;
	wire [15-1:0] node10604;
	wire [15-1:0] node10605;
	wire [15-1:0] node10606;
	wire [15-1:0] node10610;
	wire [15-1:0] node10613;
	wire [15-1:0] node10614;
	wire [15-1:0] node10615;
	wire [15-1:0] node10616;
	wire [15-1:0] node10619;
	wire [15-1:0] node10622;
	wire [15-1:0] node10624;
	wire [15-1:0] node10627;
	wire [15-1:0] node10628;
	wire [15-1:0] node10630;
	wire [15-1:0] node10631;
	wire [15-1:0] node10635;
	wire [15-1:0] node10636;
	wire [15-1:0] node10640;
	wire [15-1:0] node10641;
	wire [15-1:0] node10642;
	wire [15-1:0] node10643;
	wire [15-1:0] node10644;
	wire [15-1:0] node10648;
	wire [15-1:0] node10649;
	wire [15-1:0] node10652;
	wire [15-1:0] node10655;
	wire [15-1:0] node10656;
	wire [15-1:0] node10657;
	wire [15-1:0] node10658;
	wire [15-1:0] node10662;
	wire [15-1:0] node10664;
	wire [15-1:0] node10667;
	wire [15-1:0] node10669;
	wire [15-1:0] node10672;
	wire [15-1:0] node10673;
	wire [15-1:0] node10674;
	wire [15-1:0] node10676;
	wire [15-1:0] node10679;
	wire [15-1:0] node10681;
	wire [15-1:0] node10683;
	wire [15-1:0] node10686;
	wire [15-1:0] node10687;
	wire [15-1:0] node10689;
	wire [15-1:0] node10691;
	wire [15-1:0] node10694;
	wire [15-1:0] node10696;
	wire [15-1:0] node10699;
	wire [15-1:0] node10700;
	wire [15-1:0] node10701;
	wire [15-1:0] node10702;
	wire [15-1:0] node10703;
	wire [15-1:0] node10704;
	wire [15-1:0] node10705;
	wire [15-1:0] node10709;
	wire [15-1:0] node10710;
	wire [15-1:0] node10714;
	wire [15-1:0] node10715;
	wire [15-1:0] node10716;
	wire [15-1:0] node10717;
	wire [15-1:0] node10719;
	wire [15-1:0] node10723;
	wire [15-1:0] node10724;
	wire [15-1:0] node10728;
	wire [15-1:0] node10731;
	wire [15-1:0] node10732;
	wire [15-1:0] node10733;
	wire [15-1:0] node10735;
	wire [15-1:0] node10738;
	wire [15-1:0] node10739;
	wire [15-1:0] node10743;
	wire [15-1:0] node10744;
	wire [15-1:0] node10745;
	wire [15-1:0] node10746;
	wire [15-1:0] node10750;
	wire [15-1:0] node10751;
	wire [15-1:0] node10754;
	wire [15-1:0] node10755;
	wire [15-1:0] node10759;
	wire [15-1:0] node10760;
	wire [15-1:0] node10762;
	wire [15-1:0] node10766;
	wire [15-1:0] node10767;
	wire [15-1:0] node10768;
	wire [15-1:0] node10769;
	wire [15-1:0] node10770;
	wire [15-1:0] node10771;
	wire [15-1:0] node10775;
	wire [15-1:0] node10778;
	wire [15-1:0] node10779;
	wire [15-1:0] node10783;
	wire [15-1:0] node10784;
	wire [15-1:0] node10785;
	wire [15-1:0] node10788;
	wire [15-1:0] node10790;
	wire [15-1:0] node10793;
	wire [15-1:0] node10794;
	wire [15-1:0] node10798;
	wire [15-1:0] node10799;
	wire [15-1:0] node10800;
	wire [15-1:0] node10802;
	wire [15-1:0] node10804;
	wire [15-1:0] node10805;
	wire [15-1:0] node10809;
	wire [15-1:0] node10810;
	wire [15-1:0] node10814;
	wire [15-1:0] node10815;
	wire [15-1:0] node10816;
	wire [15-1:0] node10817;
	wire [15-1:0] node10821;
	wire [15-1:0] node10823;
	wire [15-1:0] node10826;
	wire [15-1:0] node10827;
	wire [15-1:0] node10830;
	wire [15-1:0] node10833;
	wire [15-1:0] node10834;
	wire [15-1:0] node10835;
	wire [15-1:0] node10836;
	wire [15-1:0] node10837;
	wire [15-1:0] node10838;
	wire [15-1:0] node10841;
	wire [15-1:0] node10845;
	wire [15-1:0] node10846;
	wire [15-1:0] node10847;
	wire [15-1:0] node10849;
	wire [15-1:0] node10853;
	wire [15-1:0] node10854;
	wire [15-1:0] node10855;
	wire [15-1:0] node10860;
	wire [15-1:0] node10861;
	wire [15-1:0] node10862;
	wire [15-1:0] node10863;
	wire [15-1:0] node10866;
	wire [15-1:0] node10867;
	wire [15-1:0] node10871;
	wire [15-1:0] node10872;
	wire [15-1:0] node10873;
	wire [15-1:0] node10877;
	wire [15-1:0] node10879;
	wire [15-1:0] node10882;
	wire [15-1:0] node10883;
	wire [15-1:0] node10885;
	wire [15-1:0] node10888;
	wire [15-1:0] node10890;
	wire [15-1:0] node10892;
	wire [15-1:0] node10895;
	wire [15-1:0] node10896;
	wire [15-1:0] node10897;
	wire [15-1:0] node10898;
	wire [15-1:0] node10899;
	wire [15-1:0] node10902;
	wire [15-1:0] node10905;
	wire [15-1:0] node10906;
	wire [15-1:0] node10907;
	wire [15-1:0] node10909;
	wire [15-1:0] node10913;
	wire [15-1:0] node10914;
	wire [15-1:0] node10918;
	wire [15-1:0] node10919;
	wire [15-1:0] node10921;
	wire [15-1:0] node10922;
	wire [15-1:0] node10924;
	wire [15-1:0] node10927;
	wire [15-1:0] node10928;
	wire [15-1:0] node10932;
	wire [15-1:0] node10934;
	wire [15-1:0] node10937;
	wire [15-1:0] node10938;
	wire [15-1:0] node10939;
	wire [15-1:0] node10940;
	wire [15-1:0] node10941;
	wire [15-1:0] node10945;
	wire [15-1:0] node10948;
	wire [15-1:0] node10949;
	wire [15-1:0] node10952;
	wire [15-1:0] node10953;
	wire [15-1:0] node10957;
	wire [15-1:0] node10958;
	wire [15-1:0] node10960;
	wire [15-1:0] node10962;
	wire [15-1:0] node10963;
	wire [15-1:0] node10967;
	wire [15-1:0] node10968;
	wire [15-1:0] node10971;
	wire [15-1:0] node10974;
	wire [15-1:0] node10975;
	wire [15-1:0] node10976;
	wire [15-1:0] node10977;
	wire [15-1:0] node10978;
	wire [15-1:0] node10979;
	wire [15-1:0] node10980;
	wire [15-1:0] node10981;
	wire [15-1:0] node10984;
	wire [15-1:0] node10987;
	wire [15-1:0] node10988;
	wire [15-1:0] node10989;
	wire [15-1:0] node10991;
	wire [15-1:0] node10995;
	wire [15-1:0] node10998;
	wire [15-1:0] node10999;
	wire [15-1:0] node11001;
	wire [15-1:0] node11005;
	wire [15-1:0] node11006;
	wire [15-1:0] node11007;
	wire [15-1:0] node11008;
	wire [15-1:0] node11009;
	wire [15-1:0] node11013;
	wire [15-1:0] node11016;
	wire [15-1:0] node11018;
	wire [15-1:0] node11020;
	wire [15-1:0] node11023;
	wire [15-1:0] node11024;
	wire [15-1:0] node11026;
	wire [15-1:0] node11029;
	wire [15-1:0] node11030;
	wire [15-1:0] node11034;
	wire [15-1:0] node11035;
	wire [15-1:0] node11036;
	wire [15-1:0] node11037;
	wire [15-1:0] node11041;
	wire [15-1:0] node11042;
	wire [15-1:0] node11043;
	wire [15-1:0] node11044;
	wire [15-1:0] node11046;
	wire [15-1:0] node11050;
	wire [15-1:0] node11053;
	wire [15-1:0] node11054;
	wire [15-1:0] node11056;
	wire [15-1:0] node11057;
	wire [15-1:0] node11062;
	wire [15-1:0] node11063;
	wire [15-1:0] node11064;
	wire [15-1:0] node11066;
	wire [15-1:0] node11067;
	wire [15-1:0] node11071;
	wire [15-1:0] node11074;
	wire [15-1:0] node11075;
	wire [15-1:0] node11076;
	wire [15-1:0] node11079;
	wire [15-1:0] node11082;
	wire [15-1:0] node11083;
	wire [15-1:0] node11084;
	wire [15-1:0] node11088;
	wire [15-1:0] node11090;
	wire [15-1:0] node11093;
	wire [15-1:0] node11094;
	wire [15-1:0] node11095;
	wire [15-1:0] node11096;
	wire [15-1:0] node11097;
	wire [15-1:0] node11099;
	wire [15-1:0] node11100;
	wire [15-1:0] node11104;
	wire [15-1:0] node11106;
	wire [15-1:0] node11109;
	wire [15-1:0] node11110;
	wire [15-1:0] node11112;
	wire [15-1:0] node11114;
	wire [15-1:0] node11117;
	wire [15-1:0] node11119;
	wire [15-1:0] node11122;
	wire [15-1:0] node11123;
	wire [15-1:0] node11124;
	wire [15-1:0] node11127;
	wire [15-1:0] node11128;
	wire [15-1:0] node11129;
	wire [15-1:0] node11131;
	wire [15-1:0] node11135;
	wire [15-1:0] node11138;
	wire [15-1:0] node11139;
	wire [15-1:0] node11141;
	wire [15-1:0] node11144;
	wire [15-1:0] node11146;
	wire [15-1:0] node11149;
	wire [15-1:0] node11150;
	wire [15-1:0] node11151;
	wire [15-1:0] node11152;
	wire [15-1:0] node11153;
	wire [15-1:0] node11157;
	wire [15-1:0] node11160;
	wire [15-1:0] node11161;
	wire [15-1:0] node11163;
	wire [15-1:0] node11166;
	wire [15-1:0] node11167;
	wire [15-1:0] node11170;
	wire [15-1:0] node11172;
	wire [15-1:0] node11175;
	wire [15-1:0] node11176;
	wire [15-1:0] node11177;
	wire [15-1:0] node11179;
	wire [15-1:0] node11181;
	wire [15-1:0] node11185;
	wire [15-1:0] node11186;
	wire [15-1:0] node11187;
	wire [15-1:0] node11190;
	wire [15-1:0] node11193;
	wire [15-1:0] node11194;
	wire [15-1:0] node11197;
	wire [15-1:0] node11199;
	wire [15-1:0] node11202;
	wire [15-1:0] node11203;
	wire [15-1:0] node11204;
	wire [15-1:0] node11205;
	wire [15-1:0] node11206;
	wire [15-1:0] node11207;
	wire [15-1:0] node11208;
	wire [15-1:0] node11211;
	wire [15-1:0] node11212;
	wire [15-1:0] node11214;
	wire [15-1:0] node11219;
	wire [15-1:0] node11220;
	wire [15-1:0] node11221;
	wire [15-1:0] node11224;
	wire [15-1:0] node11225;
	wire [15-1:0] node11229;
	wire [15-1:0] node11230;
	wire [15-1:0] node11232;
	wire [15-1:0] node11233;
	wire [15-1:0] node11238;
	wire [15-1:0] node11239;
	wire [15-1:0] node11241;
	wire [15-1:0] node11242;
	wire [15-1:0] node11243;
	wire [15-1:0] node11245;
	wire [15-1:0] node11250;
	wire [15-1:0] node11251;
	wire [15-1:0] node11252;
	wire [15-1:0] node11253;
	wire [15-1:0] node11257;
	wire [15-1:0] node11258;
	wire [15-1:0] node11260;
	wire [15-1:0] node11264;
	wire [15-1:0] node11265;
	wire [15-1:0] node11268;
	wire [15-1:0] node11270;
	wire [15-1:0] node11273;
	wire [15-1:0] node11274;
	wire [15-1:0] node11275;
	wire [15-1:0] node11276;
	wire [15-1:0] node11277;
	wire [15-1:0] node11278;
	wire [15-1:0] node11279;
	wire [15-1:0] node11285;
	wire [15-1:0] node11286;
	wire [15-1:0] node11287;
	wire [15-1:0] node11291;
	wire [15-1:0] node11294;
	wire [15-1:0] node11295;
	wire [15-1:0] node11296;
	wire [15-1:0] node11298;
	wire [15-1:0] node11300;
	wire [15-1:0] node11303;
	wire [15-1:0] node11304;
	wire [15-1:0] node11308;
	wire [15-1:0] node11309;
	wire [15-1:0] node11310;
	wire [15-1:0] node11314;
	wire [15-1:0] node11316;
	wire [15-1:0] node11319;
	wire [15-1:0] node11320;
	wire [15-1:0] node11321;
	wire [15-1:0] node11323;
	wire [15-1:0] node11326;
	wire [15-1:0] node11327;
	wire [15-1:0] node11328;
	wire [15-1:0] node11332;
	wire [15-1:0] node11333;
	wire [15-1:0] node11337;
	wire [15-1:0] node11338;
	wire [15-1:0] node11340;
	wire [15-1:0] node11343;
	wire [15-1:0] node11344;
	wire [15-1:0] node11347;
	wire [15-1:0] node11350;
	wire [15-1:0] node11351;
	wire [15-1:0] node11352;
	wire [15-1:0] node11353;
	wire [15-1:0] node11354;
	wire [15-1:0] node11356;
	wire [15-1:0] node11359;
	wire [15-1:0] node11360;
	wire [15-1:0] node11363;
	wire [15-1:0] node11366;
	wire [15-1:0] node11367;
	wire [15-1:0] node11368;
	wire [15-1:0] node11370;
	wire [15-1:0] node11371;
	wire [15-1:0] node11376;
	wire [15-1:0] node11378;
	wire [15-1:0] node11379;
	wire [15-1:0] node11383;
	wire [15-1:0] node11384;
	wire [15-1:0] node11385;
	wire [15-1:0] node11386;
	wire [15-1:0] node11391;
	wire [15-1:0] node11392;
	wire [15-1:0] node11394;
	wire [15-1:0] node11395;
	wire [15-1:0] node11397;
	wire [15-1:0] node11401;
	wire [15-1:0] node11402;
	wire [15-1:0] node11405;
	wire [15-1:0] node11408;
	wire [15-1:0] node11409;
	wire [15-1:0] node11410;
	wire [15-1:0] node11411;
	wire [15-1:0] node11413;
	wire [15-1:0] node11416;
	wire [15-1:0] node11417;
	wire [15-1:0] node11421;
	wire [15-1:0] node11422;
	wire [15-1:0] node11426;
	wire [15-1:0] node11427;
	wire [15-1:0] node11428;
	wire [15-1:0] node11429;
	wire [15-1:0] node11431;
	wire [15-1:0] node11433;
	wire [15-1:0] node11436;
	wire [15-1:0] node11437;
	wire [15-1:0] node11441;
	wire [15-1:0] node11442;
	wire [15-1:0] node11445;
	wire [15-1:0] node11448;
	wire [15-1:0] node11449;
	wire [15-1:0] node11450;
	wire [15-1:0] node11453;
	wire [15-1:0] node11456;
	wire [15-1:0] node11457;
	wire [15-1:0] node11458;
	wire [15-1:0] node11462;
	wire [15-1:0] node11465;
	wire [15-1:0] node11466;
	wire [15-1:0] node11467;
	wire [15-1:0] node11468;
	wire [15-1:0] node11469;
	wire [15-1:0] node11470;
	wire [15-1:0] node11471;
	wire [15-1:0] node11472;
	wire [15-1:0] node11473;
	wire [15-1:0] node11474;
	wire [15-1:0] node11479;
	wire [15-1:0] node11480;
	wire [15-1:0] node11484;
	wire [15-1:0] node11485;
	wire [15-1:0] node11486;
	wire [15-1:0] node11487;
	wire [15-1:0] node11489;
	wire [15-1:0] node11492;
	wire [15-1:0] node11493;
	wire [15-1:0] node11497;
	wire [15-1:0] node11500;
	wire [15-1:0] node11501;
	wire [15-1:0] node11505;
	wire [15-1:0] node11506;
	wire [15-1:0] node11507;
	wire [15-1:0] node11508;
	wire [15-1:0] node11512;
	wire [15-1:0] node11513;
	wire [15-1:0] node11515;
	wire [15-1:0] node11516;
	wire [15-1:0] node11521;
	wire [15-1:0] node11522;
	wire [15-1:0] node11523;
	wire [15-1:0] node11527;
	wire [15-1:0] node11529;
	wire [15-1:0] node11532;
	wire [15-1:0] node11533;
	wire [15-1:0] node11534;
	wire [15-1:0] node11535;
	wire [15-1:0] node11536;
	wire [15-1:0] node11538;
	wire [15-1:0] node11539;
	wire [15-1:0] node11544;
	wire [15-1:0] node11546;
	wire [15-1:0] node11547;
	wire [15-1:0] node11549;
	wire [15-1:0] node11553;
	wire [15-1:0] node11554;
	wire [15-1:0] node11555;
	wire [15-1:0] node11558;
	wire [15-1:0] node11560;
	wire [15-1:0] node11561;
	wire [15-1:0] node11565;
	wire [15-1:0] node11566;
	wire [15-1:0] node11567;
	wire [15-1:0] node11572;
	wire [15-1:0] node11573;
	wire [15-1:0] node11575;
	wire [15-1:0] node11576;
	wire [15-1:0] node11580;
	wire [15-1:0] node11581;
	wire [15-1:0] node11582;
	wire [15-1:0] node11584;
	wire [15-1:0] node11588;
	wire [15-1:0] node11589;
	wire [15-1:0] node11591;
	wire [15-1:0] node11594;
	wire [15-1:0] node11596;
	wire [15-1:0] node11599;
	wire [15-1:0] node11600;
	wire [15-1:0] node11601;
	wire [15-1:0] node11602;
	wire [15-1:0] node11603;
	wire [15-1:0] node11604;
	wire [15-1:0] node11606;
	wire [15-1:0] node11609;
	wire [15-1:0] node11612;
	wire [15-1:0] node11613;
	wire [15-1:0] node11616;
	wire [15-1:0] node11618;
	wire [15-1:0] node11619;
	wire [15-1:0] node11623;
	wire [15-1:0] node11624;
	wire [15-1:0] node11626;
	wire [15-1:0] node11628;
	wire [15-1:0] node11631;
	wire [15-1:0] node11632;
	wire [15-1:0] node11633;
	wire [15-1:0] node11635;
	wire [15-1:0] node11638;
	wire [15-1:0] node11639;
	wire [15-1:0] node11643;
	wire [15-1:0] node11646;
	wire [15-1:0] node11647;
	wire [15-1:0] node11648;
	wire [15-1:0] node11649;
	wire [15-1:0] node11653;
	wire [15-1:0] node11654;
	wire [15-1:0] node11657;
	wire [15-1:0] node11658;
	wire [15-1:0] node11660;
	wire [15-1:0] node11664;
	wire [15-1:0] node11665;
	wire [15-1:0] node11666;
	wire [15-1:0] node11669;
	wire [15-1:0] node11672;
	wire [15-1:0] node11675;
	wire [15-1:0] node11676;
	wire [15-1:0] node11677;
	wire [15-1:0] node11678;
	wire [15-1:0] node11679;
	wire [15-1:0] node11680;
	wire [15-1:0] node11684;
	wire [15-1:0] node11687;
	wire [15-1:0] node11688;
	wire [15-1:0] node11691;
	wire [15-1:0] node11694;
	wire [15-1:0] node11695;
	wire [15-1:0] node11697;
	wire [15-1:0] node11700;
	wire [15-1:0] node11703;
	wire [15-1:0] node11704;
	wire [15-1:0] node11705;
	wire [15-1:0] node11706;
	wire [15-1:0] node11707;
	wire [15-1:0] node11711;
	wire [15-1:0] node11714;
	wire [15-1:0] node11716;
	wire [15-1:0] node11719;
	wire [15-1:0] node11720;
	wire [15-1:0] node11721;
	wire [15-1:0] node11723;
	wire [15-1:0] node11727;
	wire [15-1:0] node11729;
	wire [15-1:0] node11732;
	wire [15-1:0] node11733;
	wire [15-1:0] node11734;
	wire [15-1:0] node11735;
	wire [15-1:0] node11736;
	wire [15-1:0] node11738;
	wire [15-1:0] node11739;
	wire [15-1:0] node11742;
	wire [15-1:0] node11744;
	wire [15-1:0] node11747;
	wire [15-1:0] node11748;
	wire [15-1:0] node11750;
	wire [15-1:0] node11751;
	wire [15-1:0] node11753;
	wire [15-1:0] node11757;
	wire [15-1:0] node11758;
	wire [15-1:0] node11759;
	wire [15-1:0] node11764;
	wire [15-1:0] node11765;
	wire [15-1:0] node11766;
	wire [15-1:0] node11767;
	wire [15-1:0] node11770;
	wire [15-1:0] node11773;
	wire [15-1:0] node11774;
	wire [15-1:0] node11778;
	wire [15-1:0] node11779;
	wire [15-1:0] node11781;
	wire [15-1:0] node11783;
	wire [15-1:0] node11786;
	wire [15-1:0] node11787;
	wire [15-1:0] node11789;
	wire [15-1:0] node11790;
	wire [15-1:0] node11794;
	wire [15-1:0] node11797;
	wire [15-1:0] node11798;
	wire [15-1:0] node11799;
	wire [15-1:0] node11800;
	wire [15-1:0] node11801;
	wire [15-1:0] node11805;
	wire [15-1:0] node11806;
	wire [15-1:0] node11809;
	wire [15-1:0] node11811;
	wire [15-1:0] node11814;
	wire [15-1:0] node11815;
	wire [15-1:0] node11816;
	wire [15-1:0] node11819;
	wire [15-1:0] node11821;
	wire [15-1:0] node11822;
	wire [15-1:0] node11826;
	wire [15-1:0] node11828;
	wire [15-1:0] node11831;
	wire [15-1:0] node11832;
	wire [15-1:0] node11833;
	wire [15-1:0] node11834;
	wire [15-1:0] node11837;
	wire [15-1:0] node11839;
	wire [15-1:0] node11842;
	wire [15-1:0] node11843;
	wire [15-1:0] node11845;
	wire [15-1:0] node11848;
	wire [15-1:0] node11850;
	wire [15-1:0] node11851;
	wire [15-1:0] node11855;
	wire [15-1:0] node11856;
	wire [15-1:0] node11857;
	wire [15-1:0] node11860;
	wire [15-1:0] node11862;
	wire [15-1:0] node11865;
	wire [15-1:0] node11866;
	wire [15-1:0] node11869;
	wire [15-1:0] node11872;
	wire [15-1:0] node11873;
	wire [15-1:0] node11874;
	wire [15-1:0] node11875;
	wire [15-1:0] node11876;
	wire [15-1:0] node11877;
	wire [15-1:0] node11878;
	wire [15-1:0] node11882;
	wire [15-1:0] node11885;
	wire [15-1:0] node11886;
	wire [15-1:0] node11888;
	wire [15-1:0] node11889;
	wire [15-1:0] node11893;
	wire [15-1:0] node11896;
	wire [15-1:0] node11897;
	wire [15-1:0] node11898;
	wire [15-1:0] node11901;
	wire [15-1:0] node11903;
	wire [15-1:0] node11906;
	wire [15-1:0] node11907;
	wire [15-1:0] node11910;
	wire [15-1:0] node11912;
	wire [15-1:0] node11915;
	wire [15-1:0] node11916;
	wire [15-1:0] node11918;
	wire [15-1:0] node11919;
	wire [15-1:0] node11921;
	wire [15-1:0] node11924;
	wire [15-1:0] node11925;
	wire [15-1:0] node11929;
	wire [15-1:0] node11930;
	wire [15-1:0] node11931;
	wire [15-1:0] node11932;
	wire [15-1:0] node11936;
	wire [15-1:0] node11937;
	wire [15-1:0] node11941;
	wire [15-1:0] node11942;
	wire [15-1:0] node11946;
	wire [15-1:0] node11947;
	wire [15-1:0] node11948;
	wire [15-1:0] node11949;
	wire [15-1:0] node11950;
	wire [15-1:0] node11951;
	wire [15-1:0] node11956;
	wire [15-1:0] node11957;
	wire [15-1:0] node11960;
	wire [15-1:0] node11963;
	wire [15-1:0] node11964;
	wire [15-1:0] node11965;
	wire [15-1:0] node11968;
	wire [15-1:0] node11969;
	wire [15-1:0] node11971;
	wire [15-1:0] node11975;
	wire [15-1:0] node11976;
	wire [15-1:0] node11980;
	wire [15-1:0] node11981;
	wire [15-1:0] node11982;
	wire [15-1:0] node11984;
	wire [15-1:0] node11986;
	wire [15-1:0] node11989;
	wire [15-1:0] node11992;
	wire [15-1:0] node11993;
	wire [15-1:0] node11995;
	wire [15-1:0] node11998;
	wire [15-1:0] node11999;
	wire [15-1:0] node12002;
	wire [15-1:0] node12004;
	wire [15-1:0] node12007;
	wire [15-1:0] node12008;
	wire [15-1:0] node12009;
	wire [15-1:0] node12010;
	wire [15-1:0] node12011;
	wire [15-1:0] node12012;
	wire [15-1:0] node12014;
	wire [15-1:0] node12015;
	wire [15-1:0] node12017;
	wire [15-1:0] node12018;
	wire [15-1:0] node12023;
	wire [15-1:0] node12024;
	wire [15-1:0] node12025;
	wire [15-1:0] node12026;
	wire [15-1:0] node12027;
	wire [15-1:0] node12032;
	wire [15-1:0] node12035;
	wire [15-1:0] node12037;
	wire [15-1:0] node12039;
	wire [15-1:0] node12041;
	wire [15-1:0] node12044;
	wire [15-1:0] node12045;
	wire [15-1:0] node12046;
	wire [15-1:0] node12047;
	wire [15-1:0] node12052;
	wire [15-1:0] node12053;
	wire [15-1:0] node12055;
	wire [15-1:0] node12058;
	wire [15-1:0] node12060;
	wire [15-1:0] node12063;
	wire [15-1:0] node12064;
	wire [15-1:0] node12065;
	wire [15-1:0] node12066;
	wire [15-1:0] node12067;
	wire [15-1:0] node12069;
	wire [15-1:0] node12072;
	wire [15-1:0] node12075;
	wire [15-1:0] node12076;
	wire [15-1:0] node12077;
	wire [15-1:0] node12082;
	wire [15-1:0] node12083;
	wire [15-1:0] node12084;
	wire [15-1:0] node12086;
	wire [15-1:0] node12088;
	wire [15-1:0] node12091;
	wire [15-1:0] node12094;
	wire [15-1:0] node12095;
	wire [15-1:0] node12096;
	wire [15-1:0] node12098;
	wire [15-1:0] node12102;
	wire [15-1:0] node12105;
	wire [15-1:0] node12106;
	wire [15-1:0] node12108;
	wire [15-1:0] node12109;
	wire [15-1:0] node12112;
	wire [15-1:0] node12113;
	wire [15-1:0] node12114;
	wire [15-1:0] node12119;
	wire [15-1:0] node12120;
	wire [15-1:0] node12121;
	wire [15-1:0] node12122;
	wire [15-1:0] node12126;
	wire [15-1:0] node12129;
	wire [15-1:0] node12131;
	wire [15-1:0] node12134;
	wire [15-1:0] node12135;
	wire [15-1:0] node12136;
	wire [15-1:0] node12137;
	wire [15-1:0] node12138;
	wire [15-1:0] node12139;
	wire [15-1:0] node12142;
	wire [15-1:0] node12145;
	wire [15-1:0] node12146;
	wire [15-1:0] node12149;
	wire [15-1:0] node12151;
	wire [15-1:0] node12154;
	wire [15-1:0] node12155;
	wire [15-1:0] node12156;
	wire [15-1:0] node12157;
	wire [15-1:0] node12162;
	wire [15-1:0] node12164;
	wire [15-1:0] node12167;
	wire [15-1:0] node12168;
	wire [15-1:0] node12169;
	wire [15-1:0] node12172;
	wire [15-1:0] node12173;
	wire [15-1:0] node12177;
	wire [15-1:0] node12178;
	wire [15-1:0] node12179;
	wire [15-1:0] node12182;
	wire [15-1:0] node12185;
	wire [15-1:0] node12186;
	wire [15-1:0] node12188;
	wire [15-1:0] node12189;
	wire [15-1:0] node12194;
	wire [15-1:0] node12195;
	wire [15-1:0] node12196;
	wire [15-1:0] node12197;
	wire [15-1:0] node12198;
	wire [15-1:0] node12200;
	wire [15-1:0] node12203;
	wire [15-1:0] node12205;
	wire [15-1:0] node12208;
	wire [15-1:0] node12209;
	wire [15-1:0] node12212;
	wire [15-1:0] node12215;
	wire [15-1:0] node12216;
	wire [15-1:0] node12218;
	wire [15-1:0] node12221;
	wire [15-1:0] node12222;
	wire [15-1:0] node12226;
	wire [15-1:0] node12227;
	wire [15-1:0] node12228;
	wire [15-1:0] node12229;
	wire [15-1:0] node12232;
	wire [15-1:0] node12235;
	wire [15-1:0] node12236;
	wire [15-1:0] node12237;
	wire [15-1:0] node12241;
	wire [15-1:0] node12242;
	wire [15-1:0] node12246;
	wire [15-1:0] node12247;
	wire [15-1:0] node12249;
	wire [15-1:0] node12251;
	wire [15-1:0] node12252;
	wire [15-1:0] node12256;
	wire [15-1:0] node12258;
	wire [15-1:0] node12260;
	wire [15-1:0] node12263;
	wire [15-1:0] node12264;
	wire [15-1:0] node12265;
	wire [15-1:0] node12266;
	wire [15-1:0] node12267;
	wire [15-1:0] node12268;
	wire [15-1:0] node12269;
	wire [15-1:0] node12270;
	wire [15-1:0] node12274;
	wire [15-1:0] node12276;
	wire [15-1:0] node12279;
	wire [15-1:0] node12282;
	wire [15-1:0] node12283;
	wire [15-1:0] node12286;
	wire [15-1:0] node12287;
	wire [15-1:0] node12291;
	wire [15-1:0] node12292;
	wire [15-1:0] node12293;
	wire [15-1:0] node12294;
	wire [15-1:0] node12295;
	wire [15-1:0] node12296;
	wire [15-1:0] node12301;
	wire [15-1:0] node12304;
	wire [15-1:0] node12305;
	wire [15-1:0] node12307;
	wire [15-1:0] node12308;
	wire [15-1:0] node12312;
	wire [15-1:0] node12315;
	wire [15-1:0] node12316;
	wire [15-1:0] node12317;
	wire [15-1:0] node12320;
	wire [15-1:0] node12322;
	wire [15-1:0] node12323;
	wire [15-1:0] node12327;
	wire [15-1:0] node12328;
	wire [15-1:0] node12331;
	wire [15-1:0] node12334;
	wire [15-1:0] node12335;
	wire [15-1:0] node12336;
	wire [15-1:0] node12337;
	wire [15-1:0] node12339;
	wire [15-1:0] node12342;
	wire [15-1:0] node12343;
	wire [15-1:0] node12346;
	wire [15-1:0] node12349;
	wire [15-1:0] node12351;
	wire [15-1:0] node12352;
	wire [15-1:0] node12354;
	wire [15-1:0] node12355;
	wire [15-1:0] node12358;
	wire [15-1:0] node12361;
	wire [15-1:0] node12364;
	wire [15-1:0] node12365;
	wire [15-1:0] node12366;
	wire [15-1:0] node12368;
	wire [15-1:0] node12370;
	wire [15-1:0] node12373;
	wire [15-1:0] node12376;
	wire [15-1:0] node12377;
	wire [15-1:0] node12380;
	wire [15-1:0] node12382;
	wire [15-1:0] node12383;
	wire [15-1:0] node12386;
	wire [15-1:0] node12389;
	wire [15-1:0] node12390;
	wire [15-1:0] node12391;
	wire [15-1:0] node12392;
	wire [15-1:0] node12393;
	wire [15-1:0] node12394;
	wire [15-1:0] node12395;
	wire [15-1:0] node12400;
	wire [15-1:0] node12401;
	wire [15-1:0] node12404;
	wire [15-1:0] node12405;
	wire [15-1:0] node12408;
	wire [15-1:0] node12411;
	wire [15-1:0] node12412;
	wire [15-1:0] node12414;
	wire [15-1:0] node12416;
	wire [15-1:0] node12417;
	wire [15-1:0] node12421;
	wire [15-1:0] node12422;
	wire [15-1:0] node12425;
	wire [15-1:0] node12428;
	wire [15-1:0] node12429;
	wire [15-1:0] node12430;
	wire [15-1:0] node12432;
	wire [15-1:0] node12433;
	wire [15-1:0] node12435;
	wire [15-1:0] node12439;
	wire [15-1:0] node12440;
	wire [15-1:0] node12443;
	wire [15-1:0] node12446;
	wire [15-1:0] node12448;
	wire [15-1:0] node12449;
	wire [15-1:0] node12453;
	wire [15-1:0] node12454;
	wire [15-1:0] node12455;
	wire [15-1:0] node12456;
	wire [15-1:0] node12459;
	wire [15-1:0] node12462;
	wire [15-1:0] node12463;
	wire [15-1:0] node12464;
	wire [15-1:0] node12468;
	wire [15-1:0] node12469;
	wire [15-1:0] node12472;
	wire [15-1:0] node12474;
	wire [15-1:0] node12476;
	wire [15-1:0] node12479;
	wire [15-1:0] node12480;
	wire [15-1:0] node12481;
	wire [15-1:0] node12482;
	wire [15-1:0] node12485;
	wire [15-1:0] node12487;
	wire [15-1:0] node12489;
	wire [15-1:0] node12492;
	wire [15-1:0] node12493;
	wire [15-1:0] node12495;
	wire [15-1:0] node12497;
	wire [15-1:0] node12501;
	wire [15-1:0] node12502;
	wire [15-1:0] node12505;
	wire [15-1:0] node12506;
	wire [15-1:0] node12507;
	wire [15-1:0] node12511;
	wire [15-1:0] node12512;
	wire [15-1:0] node12514;
	wire [15-1:0] node12518;
	wire [15-1:0] node12519;
	wire [15-1:0] node12520;
	wire [15-1:0] node12521;
	wire [15-1:0] node12522;
	wire [15-1:0] node12523;
	wire [15-1:0] node12524;
	wire [15-1:0] node12525;
	wire [15-1:0] node12526;
	wire [15-1:0] node12527;
	wire [15-1:0] node12528;
	wire [15-1:0] node12529;
	wire [15-1:0] node12532;
	wire [15-1:0] node12535;
	wire [15-1:0] node12538;
	wire [15-1:0] node12539;
	wire [15-1:0] node12541;
	wire [15-1:0] node12542;
	wire [15-1:0] node12546;
	wire [15-1:0] node12549;
	wire [15-1:0] node12550;
	wire [15-1:0] node12551;
	wire [15-1:0] node12556;
	wire [15-1:0] node12557;
	wire [15-1:0] node12558;
	wire [15-1:0] node12559;
	wire [15-1:0] node12563;
	wire [15-1:0] node12564;
	wire [15-1:0] node12565;
	wire [15-1:0] node12569;
	wire [15-1:0] node12572;
	wire [15-1:0] node12573;
	wire [15-1:0] node12574;
	wire [15-1:0] node12577;
	wire [15-1:0] node12581;
	wire [15-1:0] node12582;
	wire [15-1:0] node12583;
	wire [15-1:0] node12584;
	wire [15-1:0] node12585;
	wire [15-1:0] node12586;
	wire [15-1:0] node12587;
	wire [15-1:0] node12592;
	wire [15-1:0] node12595;
	wire [15-1:0] node12596;
	wire [15-1:0] node12597;
	wire [15-1:0] node12599;
	wire [15-1:0] node12603;
	wire [15-1:0] node12606;
	wire [15-1:0] node12607;
	wire [15-1:0] node12609;
	wire [15-1:0] node12612;
	wire [15-1:0] node12614;
	wire [15-1:0] node12617;
	wire [15-1:0] node12618;
	wire [15-1:0] node12619;
	wire [15-1:0] node12620;
	wire [15-1:0] node12623;
	wire [15-1:0] node12625;
	wire [15-1:0] node12626;
	wire [15-1:0] node12630;
	wire [15-1:0] node12631;
	wire [15-1:0] node12634;
	wire [15-1:0] node12637;
	wire [15-1:0] node12638;
	wire [15-1:0] node12639;
	wire [15-1:0] node12641;
	wire [15-1:0] node12644;
	wire [15-1:0] node12646;
	wire [15-1:0] node12649;
	wire [15-1:0] node12650;
	wire [15-1:0] node12654;
	wire [15-1:0] node12655;
	wire [15-1:0] node12656;
	wire [15-1:0] node12657;
	wire [15-1:0] node12658;
	wire [15-1:0] node12659;
	wire [15-1:0] node12661;
	wire [15-1:0] node12664;
	wire [15-1:0] node12667;
	wire [15-1:0] node12668;
	wire [15-1:0] node12670;
	wire [15-1:0] node12673;
	wire [15-1:0] node12674;
	wire [15-1:0] node12675;
	wire [15-1:0] node12680;
	wire [15-1:0] node12682;
	wire [15-1:0] node12683;
	wire [15-1:0] node12685;
	wire [15-1:0] node12688;
	wire [15-1:0] node12691;
	wire [15-1:0] node12692;
	wire [15-1:0] node12693;
	wire [15-1:0] node12696;
	wire [15-1:0] node12697;
	wire [15-1:0] node12701;
	wire [15-1:0] node12702;
	wire [15-1:0] node12704;
	wire [15-1:0] node12707;
	wire [15-1:0] node12708;
	wire [15-1:0] node12712;
	wire [15-1:0] node12713;
	wire [15-1:0] node12714;
	wire [15-1:0] node12715;
	wire [15-1:0] node12716;
	wire [15-1:0] node12717;
	wire [15-1:0] node12719;
	wire [15-1:0] node12723;
	wire [15-1:0] node12725;
	wire [15-1:0] node12728;
	wire [15-1:0] node12729;
	wire [15-1:0] node12733;
	wire [15-1:0] node12734;
	wire [15-1:0] node12735;
	wire [15-1:0] node12737;
	wire [15-1:0] node12741;
	wire [15-1:0] node12742;
	wire [15-1:0] node12743;
	wire [15-1:0] node12745;
	wire [15-1:0] node12750;
	wire [15-1:0] node12751;
	wire [15-1:0] node12752;
	wire [15-1:0] node12755;
	wire [15-1:0] node12756;
	wire [15-1:0] node12757;
	wire [15-1:0] node12762;
	wire [15-1:0] node12763;
	wire [15-1:0] node12766;
	wire [15-1:0] node12767;
	wire [15-1:0] node12768;
	wire [15-1:0] node12770;
	wire [15-1:0] node12775;
	wire [15-1:0] node12776;
	wire [15-1:0] node12777;
	wire [15-1:0] node12778;
	wire [15-1:0] node12779;
	wire [15-1:0] node12780;
	wire [15-1:0] node12782;
	wire [15-1:0] node12783;
	wire [15-1:0] node12788;
	wire [15-1:0] node12789;
	wire [15-1:0] node12792;
	wire [15-1:0] node12793;
	wire [15-1:0] node12797;
	wire [15-1:0] node12798;
	wire [15-1:0] node12799;
	wire [15-1:0] node12800;
	wire [15-1:0] node12801;
	wire [15-1:0] node12803;
	wire [15-1:0] node12807;
	wire [15-1:0] node12810;
	wire [15-1:0] node12811;
	wire [15-1:0] node12813;
	wire [15-1:0] node12814;
	wire [15-1:0] node12817;
	wire [15-1:0] node12821;
	wire [15-1:0] node12822;
	wire [15-1:0] node12825;
	wire [15-1:0] node12826;
	wire [15-1:0] node12827;
	wire [15-1:0] node12829;
	wire [15-1:0] node12834;
	wire [15-1:0] node12835;
	wire [15-1:0] node12836;
	wire [15-1:0] node12837;
	wire [15-1:0] node12838;
	wire [15-1:0] node12842;
	wire [15-1:0] node12843;
	wire [15-1:0] node12846;
	wire [15-1:0] node12849;
	wire [15-1:0] node12850;
	wire [15-1:0] node12851;
	wire [15-1:0] node12856;
	wire [15-1:0] node12857;
	wire [15-1:0] node12858;
	wire [15-1:0] node12859;
	wire [15-1:0] node12861;
	wire [15-1:0] node12865;
	wire [15-1:0] node12866;
	wire [15-1:0] node12868;
	wire [15-1:0] node12872;
	wire [15-1:0] node12873;
	wire [15-1:0] node12876;
	wire [15-1:0] node12877;
	wire [15-1:0] node12881;
	wire [15-1:0] node12882;
	wire [15-1:0] node12883;
	wire [15-1:0] node12884;
	wire [15-1:0] node12886;
	wire [15-1:0] node12887;
	wire [15-1:0] node12888;
	wire [15-1:0] node12889;
	wire [15-1:0] node12893;
	wire [15-1:0] node12896;
	wire [15-1:0] node12897;
	wire [15-1:0] node12901;
	wire [15-1:0] node12902;
	wire [15-1:0] node12904;
	wire [15-1:0] node12907;
	wire [15-1:0] node12908;
	wire [15-1:0] node12910;
	wire [15-1:0] node12914;
	wire [15-1:0] node12915;
	wire [15-1:0] node12916;
	wire [15-1:0] node12917;
	wire [15-1:0] node12919;
	wire [15-1:0] node12921;
	wire [15-1:0] node12924;
	wire [15-1:0] node12925;
	wire [15-1:0] node12927;
	wire [15-1:0] node12932;
	wire [15-1:0] node12933;
	wire [15-1:0] node12934;
	wire [15-1:0] node12935;
	wire [15-1:0] node12939;
	wire [15-1:0] node12941;
	wire [15-1:0] node12944;
	wire [15-1:0] node12945;
	wire [15-1:0] node12948;
	wire [15-1:0] node12951;
	wire [15-1:0] node12952;
	wire [15-1:0] node12953;
	wire [15-1:0] node12954;
	wire [15-1:0] node12955;
	wire [15-1:0] node12956;
	wire [15-1:0] node12960;
	wire [15-1:0] node12963;
	wire [15-1:0] node12964;
	wire [15-1:0] node12966;
	wire [15-1:0] node12969;
	wire [15-1:0] node12972;
	wire [15-1:0] node12973;
	wire [15-1:0] node12974;
	wire [15-1:0] node12976;
	wire [15-1:0] node12977;
	wire [15-1:0] node12982;
	wire [15-1:0] node12985;
	wire [15-1:0] node12986;
	wire [15-1:0] node12987;
	wire [15-1:0] node12988;
	wire [15-1:0] node12990;
	wire [15-1:0] node12993;
	wire [15-1:0] node12995;
	wire [15-1:0] node12998;
	wire [15-1:0] node13000;
	wire [15-1:0] node13003;
	wire [15-1:0] node13004;
	wire [15-1:0] node13005;
	wire [15-1:0] node13006;
	wire [15-1:0] node13010;
	wire [15-1:0] node13013;
	wire [15-1:0] node13014;
	wire [15-1:0] node13015;
	wire [15-1:0] node13019;
	wire [15-1:0] node13021;
	wire [15-1:0] node13024;
	wire [15-1:0] node13025;
	wire [15-1:0] node13026;
	wire [15-1:0] node13027;
	wire [15-1:0] node13028;
	wire [15-1:0] node13029;
	wire [15-1:0] node13030;
	wire [15-1:0] node13031;
	wire [15-1:0] node13035;
	wire [15-1:0] node13038;
	wire [15-1:0] node13039;
	wire [15-1:0] node13040;
	wire [15-1:0] node13041;
	wire [15-1:0] node13043;
	wire [15-1:0] node13047;
	wire [15-1:0] node13050;
	wire [15-1:0] node13051;
	wire [15-1:0] node13055;
	wire [15-1:0] node13056;
	wire [15-1:0] node13057;
	wire [15-1:0] node13058;
	wire [15-1:0] node13060;
	wire [15-1:0] node13061;
	wire [15-1:0] node13065;
	wire [15-1:0] node13067;
	wire [15-1:0] node13070;
	wire [15-1:0] node13071;
	wire [15-1:0] node13073;
	wire [15-1:0] node13076;
	wire [15-1:0] node13079;
	wire [15-1:0] node13080;
	wire [15-1:0] node13081;
	wire [15-1:0] node13082;
	wire [15-1:0] node13086;
	wire [15-1:0] node13089;
	wire [15-1:0] node13090;
	wire [15-1:0] node13094;
	wire [15-1:0] node13095;
	wire [15-1:0] node13096;
	wire [15-1:0] node13097;
	wire [15-1:0] node13100;
	wire [15-1:0] node13102;
	wire [15-1:0] node13103;
	wire [15-1:0] node13107;
	wire [15-1:0] node13108;
	wire [15-1:0] node13109;
	wire [15-1:0] node13113;
	wire [15-1:0] node13115;
	wire [15-1:0] node13118;
	wire [15-1:0] node13119;
	wire [15-1:0] node13120;
	wire [15-1:0] node13122;
	wire [15-1:0] node13125;
	wire [15-1:0] node13126;
	wire [15-1:0] node13129;
	wire [15-1:0] node13130;
	wire [15-1:0] node13134;
	wire [15-1:0] node13135;
	wire [15-1:0] node13137;
	wire [15-1:0] node13140;
	wire [15-1:0] node13141;
	wire [15-1:0] node13142;
	wire [15-1:0] node13146;
	wire [15-1:0] node13148;
	wire [15-1:0] node13151;
	wire [15-1:0] node13152;
	wire [15-1:0] node13153;
	wire [15-1:0] node13154;
	wire [15-1:0] node13155;
	wire [15-1:0] node13156;
	wire [15-1:0] node13157;
	wire [15-1:0] node13159;
	wire [15-1:0] node13163;
	wire [15-1:0] node13166;
	wire [15-1:0] node13167;
	wire [15-1:0] node13170;
	wire [15-1:0] node13173;
	wire [15-1:0] node13175;
	wire [15-1:0] node13176;
	wire [15-1:0] node13179;
	wire [15-1:0] node13182;
	wire [15-1:0] node13183;
	wire [15-1:0] node13184;
	wire [15-1:0] node13186;
	wire [15-1:0] node13188;
	wire [15-1:0] node13189;
	wire [15-1:0] node13193;
	wire [15-1:0] node13194;
	wire [15-1:0] node13195;
	wire [15-1:0] node13199;
	wire [15-1:0] node13202;
	wire [15-1:0] node13204;
	wire [15-1:0] node13207;
	wire [15-1:0] node13208;
	wire [15-1:0] node13209;
	wire [15-1:0] node13210;
	wire [15-1:0] node13211;
	wire [15-1:0] node13215;
	wire [15-1:0] node13216;
	wire [15-1:0] node13218;
	wire [15-1:0] node13222;
	wire [15-1:0] node13223;
	wire [15-1:0] node13224;
	wire [15-1:0] node13227;
	wire [15-1:0] node13229;
	wire [15-1:0] node13232;
	wire [15-1:0] node13233;
	wire [15-1:0] node13236;
	wire [15-1:0] node13239;
	wire [15-1:0] node13240;
	wire [15-1:0] node13241;
	wire [15-1:0] node13242;
	wire [15-1:0] node13245;
	wire [15-1:0] node13247;
	wire [15-1:0] node13248;
	wire [15-1:0] node13252;
	wire [15-1:0] node13253;
	wire [15-1:0] node13256;
	wire [15-1:0] node13259;
	wire [15-1:0] node13260;
	wire [15-1:0] node13262;
	wire [15-1:0] node13264;
	wire [15-1:0] node13267;
	wire [15-1:0] node13269;
	wire [15-1:0] node13272;
	wire [15-1:0] node13273;
	wire [15-1:0] node13274;
	wire [15-1:0] node13275;
	wire [15-1:0] node13276;
	wire [15-1:0] node13277;
	wire [15-1:0] node13278;
	wire [15-1:0] node13280;
	wire [15-1:0] node13283;
	wire [15-1:0] node13286;
	wire [15-1:0] node13287;
	wire [15-1:0] node13288;
	wire [15-1:0] node13290;
	wire [15-1:0] node13294;
	wire [15-1:0] node13296;
	wire [15-1:0] node13297;
	wire [15-1:0] node13301;
	wire [15-1:0] node13302;
	wire [15-1:0] node13303;
	wire [15-1:0] node13304;
	wire [15-1:0] node13306;
	wire [15-1:0] node13310;
	wire [15-1:0] node13313;
	wire [15-1:0] node13316;
	wire [15-1:0] node13317;
	wire [15-1:0] node13318;
	wire [15-1:0] node13319;
	wire [15-1:0] node13322;
	wire [15-1:0] node13323;
	wire [15-1:0] node13325;
	wire [15-1:0] node13328;
	wire [15-1:0] node13332;
	wire [15-1:0] node13333;
	wire [15-1:0] node13335;
	wire [15-1:0] node13338;
	wire [15-1:0] node13341;
	wire [15-1:0] node13342;
	wire [15-1:0] node13343;
	wire [15-1:0] node13344;
	wire [15-1:0] node13345;
	wire [15-1:0] node13349;
	wire [15-1:0] node13350;
	wire [15-1:0] node13354;
	wire [15-1:0] node13356;
	wire [15-1:0] node13357;
	wire [15-1:0] node13360;
	wire [15-1:0] node13363;
	wire [15-1:0] node13364;
	wire [15-1:0] node13365;
	wire [15-1:0] node13366;
	wire [15-1:0] node13369;
	wire [15-1:0] node13370;
	wire [15-1:0] node13372;
	wire [15-1:0] node13376;
	wire [15-1:0] node13377;
	wire [15-1:0] node13380;
	wire [15-1:0] node13382;
	wire [15-1:0] node13385;
	wire [15-1:0] node13386;
	wire [15-1:0] node13387;
	wire [15-1:0] node13390;
	wire [15-1:0] node13393;
	wire [15-1:0] node13394;
	wire [15-1:0] node13397;
	wire [15-1:0] node13400;
	wire [15-1:0] node13401;
	wire [15-1:0] node13402;
	wire [15-1:0] node13403;
	wire [15-1:0] node13404;
	wire [15-1:0] node13405;
	wire [15-1:0] node13409;
	wire [15-1:0] node13410;
	wire [15-1:0] node13413;
	wire [15-1:0] node13415;
	wire [15-1:0] node13418;
	wire [15-1:0] node13419;
	wire [15-1:0] node13421;
	wire [15-1:0] node13425;
	wire [15-1:0] node13426;
	wire [15-1:0] node13427;
	wire [15-1:0] node13428;
	wire [15-1:0] node13431;
	wire [15-1:0] node13432;
	wire [15-1:0] node13434;
	wire [15-1:0] node13438;
	wire [15-1:0] node13440;
	wire [15-1:0] node13443;
	wire [15-1:0] node13444;
	wire [15-1:0] node13445;
	wire [15-1:0] node13446;
	wire [15-1:0] node13448;
	wire [15-1:0] node13452;
	wire [15-1:0] node13454;
	wire [15-1:0] node13456;
	wire [15-1:0] node13459;
	wire [15-1:0] node13460;
	wire [15-1:0] node13463;
	wire [15-1:0] node13466;
	wire [15-1:0] node13467;
	wire [15-1:0] node13468;
	wire [15-1:0] node13469;
	wire [15-1:0] node13470;
	wire [15-1:0] node13473;
	wire [15-1:0] node13476;
	wire [15-1:0] node13477;
	wire [15-1:0] node13478;
	wire [15-1:0] node13480;
	wire [15-1:0] node13483;
	wire [15-1:0] node13485;
	wire [15-1:0] node13488;
	wire [15-1:0] node13490;
	wire [15-1:0] node13491;
	wire [15-1:0] node13495;
	wire [15-1:0] node13496;
	wire [15-1:0] node13497;
	wire [15-1:0] node13499;
	wire [15-1:0] node13501;
	wire [15-1:0] node13506;
	wire [15-1:0] node13507;
	wire [15-1:0] node13509;
	wire [15-1:0] node13510;
	wire [15-1:0] node13511;
	wire [15-1:0] node13516;
	wire [15-1:0] node13517;
	wire [15-1:0] node13518;
	wire [15-1:0] node13519;
	wire [15-1:0] node13523;
	wire [15-1:0] node13526;
	wire [15-1:0] node13528;
	wire [15-1:0] node13529;
	wire [15-1:0] node13531;
	wire [15-1:0] node13534;
	wire [15-1:0] node13536;
	wire [15-1:0] node13539;
	wire [15-1:0] node13540;
	wire [15-1:0] node13541;
	wire [15-1:0] node13542;
	wire [15-1:0] node13543;
	wire [15-1:0] node13544;
	wire [15-1:0] node13545;
	wire [15-1:0] node13546;
	wire [15-1:0] node13547;
	wire [15-1:0] node13548;
	wire [15-1:0] node13552;
	wire [15-1:0] node13555;
	wire [15-1:0] node13556;
	wire [15-1:0] node13558;
	wire [15-1:0] node13562;
	wire [15-1:0] node13563;
	wire [15-1:0] node13564;
	wire [15-1:0] node13567;
	wire [15-1:0] node13570;
	wire [15-1:0] node13571;
	wire [15-1:0] node13573;
	wire [15-1:0] node13574;
	wire [15-1:0] node13578;
	wire [15-1:0] node13581;
	wire [15-1:0] node13582;
	wire [15-1:0] node13583;
	wire [15-1:0] node13585;
	wire [15-1:0] node13586;
	wire [15-1:0] node13589;
	wire [15-1:0] node13590;
	wire [15-1:0] node13594;
	wire [15-1:0] node13596;
	wire [15-1:0] node13599;
	wire [15-1:0] node13600;
	wire [15-1:0] node13601;
	wire [15-1:0] node13602;
	wire [15-1:0] node13606;
	wire [15-1:0] node13609;
	wire [15-1:0] node13611;
	wire [15-1:0] node13612;
	wire [15-1:0] node13614;
	wire [15-1:0] node13618;
	wire [15-1:0] node13619;
	wire [15-1:0] node13620;
	wire [15-1:0] node13621;
	wire [15-1:0] node13622;
	wire [15-1:0] node13624;
	wire [15-1:0] node13628;
	wire [15-1:0] node13629;
	wire [15-1:0] node13630;
	wire [15-1:0] node13635;
	wire [15-1:0] node13636;
	wire [15-1:0] node13638;
	wire [15-1:0] node13639;
	wire [15-1:0] node13643;
	wire [15-1:0] node13646;
	wire [15-1:0] node13647;
	wire [15-1:0] node13648;
	wire [15-1:0] node13651;
	wire [15-1:0] node13652;
	wire [15-1:0] node13654;
	wire [15-1:0] node13657;
	wire [15-1:0] node13658;
	wire [15-1:0] node13659;
	wire [15-1:0] node13663;
	wire [15-1:0] node13666;
	wire [15-1:0] node13667;
	wire [15-1:0] node13670;
	wire [15-1:0] node13671;
	wire [15-1:0] node13673;
	wire [15-1:0] node13677;
	wire [15-1:0] node13678;
	wire [15-1:0] node13679;
	wire [15-1:0] node13680;
	wire [15-1:0] node13681;
	wire [15-1:0] node13682;
	wire [15-1:0] node13685;
	wire [15-1:0] node13688;
	wire [15-1:0] node13689;
	wire [15-1:0] node13691;
	wire [15-1:0] node13695;
	wire [15-1:0] node13696;
	wire [15-1:0] node13697;
	wire [15-1:0] node13698;
	wire [15-1:0] node13702;
	wire [15-1:0] node13705;
	wire [15-1:0] node13706;
	wire [15-1:0] node13708;
	wire [15-1:0] node13711;
	wire [15-1:0] node13714;
	wire [15-1:0] node13715;
	wire [15-1:0] node13716;
	wire [15-1:0] node13717;
	wire [15-1:0] node13718;
	wire [15-1:0] node13719;
	wire [15-1:0] node13724;
	wire [15-1:0] node13727;
	wire [15-1:0] node13728;
	wire [15-1:0] node13730;
	wire [15-1:0] node13732;
	wire [15-1:0] node13736;
	wire [15-1:0] node13737;
	wire [15-1:0] node13738;
	wire [15-1:0] node13742;
	wire [15-1:0] node13745;
	wire [15-1:0] node13746;
	wire [15-1:0] node13747;
	wire [15-1:0] node13748;
	wire [15-1:0] node13749;
	wire [15-1:0] node13751;
	wire [15-1:0] node13755;
	wire [15-1:0] node13756;
	wire [15-1:0] node13757;
	wire [15-1:0] node13761;
	wire [15-1:0] node13764;
	wire [15-1:0] node13765;
	wire [15-1:0] node13766;
	wire [15-1:0] node13767;
	wire [15-1:0] node13772;
	wire [15-1:0] node13773;
	wire [15-1:0] node13776;
	wire [15-1:0] node13778;
	wire [15-1:0] node13780;
	wire [15-1:0] node13783;
	wire [15-1:0] node13784;
	wire [15-1:0] node13785;
	wire [15-1:0] node13787;
	wire [15-1:0] node13790;
	wire [15-1:0] node13791;
	wire [15-1:0] node13794;
	wire [15-1:0] node13797;
	wire [15-1:0] node13798;
	wire [15-1:0] node13800;
	wire [15-1:0] node13801;
	wire [15-1:0] node13803;
	wire [15-1:0] node13807;
	wire [15-1:0] node13808;
	wire [15-1:0] node13812;
	wire [15-1:0] node13813;
	wire [15-1:0] node13814;
	wire [15-1:0] node13815;
	wire [15-1:0] node13816;
	wire [15-1:0] node13817;
	wire [15-1:0] node13819;
	wire [15-1:0] node13822;
	wire [15-1:0] node13823;
	wire [15-1:0] node13824;
	wire [15-1:0] node13826;
	wire [15-1:0] node13830;
	wire [15-1:0] node13833;
	wire [15-1:0] node13835;
	wire [15-1:0] node13836;
	wire [15-1:0] node13837;
	wire [15-1:0] node13838;
	wire [15-1:0] node13844;
	wire [15-1:0] node13845;
	wire [15-1:0] node13846;
	wire [15-1:0] node13847;
	wire [15-1:0] node13850;
	wire [15-1:0] node13852;
	wire [15-1:0] node13855;
	wire [15-1:0] node13856;
	wire [15-1:0] node13860;
	wire [15-1:0] node13861;
	wire [15-1:0] node13862;
	wire [15-1:0] node13866;
	wire [15-1:0] node13868;
	wire [15-1:0] node13871;
	wire [15-1:0] node13872;
	wire [15-1:0] node13873;
	wire [15-1:0] node13874;
	wire [15-1:0] node13875;
	wire [15-1:0] node13876;
	wire [15-1:0] node13880;
	wire [15-1:0] node13883;
	wire [15-1:0] node13884;
	wire [15-1:0] node13888;
	wire [15-1:0] node13889;
	wire [15-1:0] node13890;
	wire [15-1:0] node13891;
	wire [15-1:0] node13895;
	wire [15-1:0] node13898;
	wire [15-1:0] node13899;
	wire [15-1:0] node13900;
	wire [15-1:0] node13902;
	wire [15-1:0] node13906;
	wire [15-1:0] node13908;
	wire [15-1:0] node13911;
	wire [15-1:0] node13912;
	wire [15-1:0] node13913;
	wire [15-1:0] node13914;
	wire [15-1:0] node13915;
	wire [15-1:0] node13919;
	wire [15-1:0] node13922;
	wire [15-1:0] node13923;
	wire [15-1:0] node13926;
	wire [15-1:0] node13929;
	wire [15-1:0] node13930;
	wire [15-1:0] node13931;
	wire [15-1:0] node13935;
	wire [15-1:0] node13936;
	wire [15-1:0] node13937;
	wire [15-1:0] node13939;
	wire [15-1:0] node13944;
	wire [15-1:0] node13945;
	wire [15-1:0] node13946;
	wire [15-1:0] node13947;
	wire [15-1:0] node13948;
	wire [15-1:0] node13949;
	wire [15-1:0] node13952;
	wire [15-1:0] node13955;
	wire [15-1:0] node13956;
	wire [15-1:0] node13958;
	wire [15-1:0] node13961;
	wire [15-1:0] node13964;
	wire [15-1:0] node13965;
	wire [15-1:0] node13966;
	wire [15-1:0] node13967;
	wire [15-1:0] node13971;
	wire [15-1:0] node13974;
	wire [15-1:0] node13975;
	wire [15-1:0] node13978;
	wire [15-1:0] node13981;
	wire [15-1:0] node13982;
	wire [15-1:0] node13983;
	wire [15-1:0] node13984;
	wire [15-1:0] node13988;
	wire [15-1:0] node13989;
	wire [15-1:0] node13992;
	wire [15-1:0] node13993;
	wire [15-1:0] node13997;
	wire [15-1:0] node13998;
	wire [15-1:0] node13999;
	wire [15-1:0] node14001;
	wire [15-1:0] node14003;
	wire [15-1:0] node14007;
	wire [15-1:0] node14008;
	wire [15-1:0] node14011;
	wire [15-1:0] node14012;
	wire [15-1:0] node14014;
	wire [15-1:0] node14018;
	wire [15-1:0] node14019;
	wire [15-1:0] node14020;
	wire [15-1:0] node14023;
	wire [15-1:0] node14024;
	wire [15-1:0] node14026;
	wire [15-1:0] node14029;
	wire [15-1:0] node14030;
	wire [15-1:0] node14031;
	wire [15-1:0] node14036;
	wire [15-1:0] node14037;
	wire [15-1:0] node14038;
	wire [15-1:0] node14040;
	wire [15-1:0] node14043;
	wire [15-1:0] node14044;
	wire [15-1:0] node14047;
	wire [15-1:0] node14050;
	wire [15-1:0] node14051;
	wire [15-1:0] node14052;
	wire [15-1:0] node14055;
	wire [15-1:0] node14057;
	wire [15-1:0] node14060;
	wire [15-1:0] node14061;
	wire [15-1:0] node14064;
	wire [15-1:0] node14067;
	wire [15-1:0] node14068;
	wire [15-1:0] node14069;
	wire [15-1:0] node14070;
	wire [15-1:0] node14071;
	wire [15-1:0] node14072;
	wire [15-1:0] node14073;
	wire [15-1:0] node14076;
	wire [15-1:0] node14078;
	wire [15-1:0] node14081;
	wire [15-1:0] node14082;
	wire [15-1:0] node14083;
	wire [15-1:0] node14086;
	wire [15-1:0] node14087;
	wire [15-1:0] node14092;
	wire [15-1:0] node14093;
	wire [15-1:0] node14094;
	wire [15-1:0] node14096;
	wire [15-1:0] node14099;
	wire [15-1:0] node14101;
	wire [15-1:0] node14103;
	wire [15-1:0] node14106;
	wire [15-1:0] node14107;
	wire [15-1:0] node14108;
	wire [15-1:0] node14112;
	wire [15-1:0] node14114;
	wire [15-1:0] node14117;
	wire [15-1:0] node14118;
	wire [15-1:0] node14119;
	wire [15-1:0] node14120;
	wire [15-1:0] node14121;
	wire [15-1:0] node14125;
	wire [15-1:0] node14126;
	wire [15-1:0] node14129;
	wire [15-1:0] node14132;
	wire [15-1:0] node14133;
	wire [15-1:0] node14134;
	wire [15-1:0] node14138;
	wire [15-1:0] node14139;
	wire [15-1:0] node14141;
	wire [15-1:0] node14144;
	wire [15-1:0] node14145;
	wire [15-1:0] node14146;
	wire [15-1:0] node14150;
	wire [15-1:0] node14153;
	wire [15-1:0] node14154;
	wire [15-1:0] node14155;
	wire [15-1:0] node14156;
	wire [15-1:0] node14158;
	wire [15-1:0] node14159;
	wire [15-1:0] node14163;
	wire [15-1:0] node14164;
	wire [15-1:0] node14166;
	wire [15-1:0] node14170;
	wire [15-1:0] node14171;
	wire [15-1:0] node14174;
	wire [15-1:0] node14175;
	wire [15-1:0] node14177;
	wire [15-1:0] node14181;
	wire [15-1:0] node14182;
	wire [15-1:0] node14183;
	wire [15-1:0] node14186;
	wire [15-1:0] node14187;
	wire [15-1:0] node14191;
	wire [15-1:0] node14192;
	wire [15-1:0] node14193;
	wire [15-1:0] node14197;
	wire [15-1:0] node14200;
	wire [15-1:0] node14201;
	wire [15-1:0] node14202;
	wire [15-1:0] node14203;
	wire [15-1:0] node14204;
	wire [15-1:0] node14205;
	wire [15-1:0] node14206;
	wire [15-1:0] node14207;
	wire [15-1:0] node14211;
	wire [15-1:0] node14215;
	wire [15-1:0] node14217;
	wire [15-1:0] node14219;
	wire [15-1:0] node14222;
	wire [15-1:0] node14223;
	wire [15-1:0] node14224;
	wire [15-1:0] node14228;
	wire [15-1:0] node14229;
	wire [15-1:0] node14230;
	wire [15-1:0] node14234;
	wire [15-1:0] node14237;
	wire [15-1:0] node14238;
	wire [15-1:0] node14239;
	wire [15-1:0] node14240;
	wire [15-1:0] node14241;
	wire [15-1:0] node14245;
	wire [15-1:0] node14247;
	wire [15-1:0] node14248;
	wire [15-1:0] node14252;
	wire [15-1:0] node14253;
	wire [15-1:0] node14254;
	wire [15-1:0] node14258;
	wire [15-1:0] node14261;
	wire [15-1:0] node14262;
	wire [15-1:0] node14263;
	wire [15-1:0] node14266;
	wire [15-1:0] node14269;
	wire [15-1:0] node14270;
	wire [15-1:0] node14272;
	wire [15-1:0] node14275;
	wire [15-1:0] node14277;
	wire [15-1:0] node14280;
	wire [15-1:0] node14281;
	wire [15-1:0] node14282;
	wire [15-1:0] node14283;
	wire [15-1:0] node14285;
	wire [15-1:0] node14289;
	wire [15-1:0] node14290;
	wire [15-1:0] node14291;
	wire [15-1:0] node14294;
	wire [15-1:0] node14297;
	wire [15-1:0] node14298;
	wire [15-1:0] node14301;
	wire [15-1:0] node14304;
	wire [15-1:0] node14305;
	wire [15-1:0] node14306;
	wire [15-1:0] node14307;
	wire [15-1:0] node14310;
	wire [15-1:0] node14313;
	wire [15-1:0] node14314;
	wire [15-1:0] node14318;
	wire [15-1:0] node14319;
	wire [15-1:0] node14320;
	wire [15-1:0] node14323;
	wire [15-1:0] node14325;
	wire [15-1:0] node14328;
	wire [15-1:0] node14329;
	wire [15-1:0] node14332;
	wire [15-1:0] node14334;
	wire [15-1:0] node14337;
	wire [15-1:0] node14338;
	wire [15-1:0] node14339;
	wire [15-1:0] node14340;
	wire [15-1:0] node14341;
	wire [15-1:0] node14342;
	wire [15-1:0] node14343;
	wire [15-1:0] node14347;
	wire [15-1:0] node14348;
	wire [15-1:0] node14349;
	wire [15-1:0] node14353;
	wire [15-1:0] node14356;
	wire [15-1:0] node14357;
	wire [15-1:0] node14359;
	wire [15-1:0] node14362;
	wire [15-1:0] node14363;
	wire [15-1:0] node14364;
	wire [15-1:0] node14369;
	wire [15-1:0] node14370;
	wire [15-1:0] node14372;
	wire [15-1:0] node14373;
	wire [15-1:0] node14374;
	wire [15-1:0] node14379;
	wire [15-1:0] node14380;
	wire [15-1:0] node14382;
	wire [15-1:0] node14385;
	wire [15-1:0] node14386;
	wire [15-1:0] node14390;
	wire [15-1:0] node14391;
	wire [15-1:0] node14392;
	wire [15-1:0] node14393;
	wire [15-1:0] node14394;
	wire [15-1:0] node14397;
	wire [15-1:0] node14399;
	wire [15-1:0] node14400;
	wire [15-1:0] node14404;
	wire [15-1:0] node14405;
	wire [15-1:0] node14406;
	wire [15-1:0] node14411;
	wire [15-1:0] node14412;
	wire [15-1:0] node14413;
	wire [15-1:0] node14414;
	wire [15-1:0] node14418;
	wire [15-1:0] node14421;
	wire [15-1:0] node14424;
	wire [15-1:0] node14425;
	wire [15-1:0] node14426;
	wire [15-1:0] node14427;
	wire [15-1:0] node14430;
	wire [15-1:0] node14432;
	wire [15-1:0] node14435;
	wire [15-1:0] node14436;
	wire [15-1:0] node14439;
	wire [15-1:0] node14440;
	wire [15-1:0] node14443;
	wire [15-1:0] node14444;
	wire [15-1:0] node14448;
	wire [15-1:0] node14450;
	wire [15-1:0] node14451;
	wire [15-1:0] node14452;
	wire [15-1:0] node14456;
	wire [15-1:0] node14457;
	wire [15-1:0] node14459;
	wire [15-1:0] node14463;
	wire [15-1:0] node14464;
	wire [15-1:0] node14465;
	wire [15-1:0] node14466;
	wire [15-1:0] node14467;
	wire [15-1:0] node14468;
	wire [15-1:0] node14469;
	wire [15-1:0] node14471;
	wire [15-1:0] node14476;
	wire [15-1:0] node14477;
	wire [15-1:0] node14478;
	wire [15-1:0] node14480;
	wire [15-1:0] node14485;
	wire [15-1:0] node14486;
	wire [15-1:0] node14487;
	wire [15-1:0] node14490;
	wire [15-1:0] node14491;
	wire [15-1:0] node14492;
	wire [15-1:0] node14495;
	wire [15-1:0] node14499;
	wire [15-1:0] node14500;
	wire [15-1:0] node14501;
	wire [15-1:0] node14506;
	wire [15-1:0] node14507;
	wire [15-1:0] node14508;
	wire [15-1:0] node14510;
	wire [15-1:0] node14512;
	wire [15-1:0] node14515;
	wire [15-1:0] node14516;
	wire [15-1:0] node14517;
	wire [15-1:0] node14519;
	wire [15-1:0] node14523;
	wire [15-1:0] node14526;
	wire [15-1:0] node14527;
	wire [15-1:0] node14528;
	wire [15-1:0] node14531;
	wire [15-1:0] node14534;
	wire [15-1:0] node14536;
	wire [15-1:0] node14537;
	wire [15-1:0] node14541;
	wire [15-1:0] node14542;
	wire [15-1:0] node14543;
	wire [15-1:0] node14545;
	wire [15-1:0] node14547;
	wire [15-1:0] node14550;
	wire [15-1:0] node14552;
	wire [15-1:0] node14553;
	wire [15-1:0] node14554;
	wire [15-1:0] node14556;
	wire [15-1:0] node14559;
	wire [15-1:0] node14561;
	wire [15-1:0] node14565;
	wire [15-1:0] node14566;
	wire [15-1:0] node14567;
	wire [15-1:0] node14569;
	wire [15-1:0] node14571;
	wire [15-1:0] node14572;
	wire [15-1:0] node14576;
	wire [15-1:0] node14577;
	wire [15-1:0] node14578;
	wire [15-1:0] node14580;
	wire [15-1:0] node14584;
	wire [15-1:0] node14585;
	wire [15-1:0] node14587;
	wire [15-1:0] node14591;
	wire [15-1:0] node14593;
	wire [15-1:0] node14595;
	wire [15-1:0] node14597;
	wire [15-1:0] node14598;
	wire [15-1:0] node14602;
	wire [15-1:0] node14603;
	wire [15-1:0] node14604;
	wire [15-1:0] node14605;
	wire [15-1:0] node14606;
	wire [15-1:0] node14607;
	wire [15-1:0] node14608;
	wire [15-1:0] node14609;
	wire [15-1:0] node14610;
	wire [15-1:0] node14611;
	wire [15-1:0] node14612;
	wire [15-1:0] node14616;
	wire [15-1:0] node14619;
	wire [15-1:0] node14620;
	wire [15-1:0] node14621;
	wire [15-1:0] node14623;
	wire [15-1:0] node14627;
	wire [15-1:0] node14630;
	wire [15-1:0] node14631;
	wire [15-1:0] node14632;
	wire [15-1:0] node14635;
	wire [15-1:0] node14637;
	wire [15-1:0] node14640;
	wire [15-1:0] node14641;
	wire [15-1:0] node14642;
	wire [15-1:0] node14644;
	wire [15-1:0] node14648;
	wire [15-1:0] node14650;
	wire [15-1:0] node14653;
	wire [15-1:0] node14654;
	wire [15-1:0] node14655;
	wire [15-1:0] node14656;
	wire [15-1:0] node14660;
	wire [15-1:0] node14661;
	wire [15-1:0] node14663;
	wire [15-1:0] node14664;
	wire [15-1:0] node14669;
	wire [15-1:0] node14670;
	wire [15-1:0] node14671;
	wire [15-1:0] node14672;
	wire [15-1:0] node14677;
	wire [15-1:0] node14678;
	wire [15-1:0] node14681;
	wire [15-1:0] node14684;
	wire [15-1:0] node14685;
	wire [15-1:0] node14686;
	wire [15-1:0] node14687;
	wire [15-1:0] node14688;
	wire [15-1:0] node14691;
	wire [15-1:0] node14694;
	wire [15-1:0] node14696;
	wire [15-1:0] node14698;
	wire [15-1:0] node14701;
	wire [15-1:0] node14702;
	wire [15-1:0] node14703;
	wire [15-1:0] node14704;
	wire [15-1:0] node14708;
	wire [15-1:0] node14709;
	wire [15-1:0] node14711;
	wire [15-1:0] node14715;
	wire [15-1:0] node14717;
	wire [15-1:0] node14720;
	wire [15-1:0] node14721;
	wire [15-1:0] node14722;
	wire [15-1:0] node14724;
	wire [15-1:0] node14728;
	wire [15-1:0] node14729;
	wire [15-1:0] node14732;
	wire [15-1:0] node14735;
	wire [15-1:0] node14736;
	wire [15-1:0] node14737;
	wire [15-1:0] node14738;
	wire [15-1:0] node14739;
	wire [15-1:0] node14740;
	wire [15-1:0] node14743;
	wire [15-1:0] node14746;
	wire [15-1:0] node14747;
	wire [15-1:0] node14751;
	wire [15-1:0] node14752;
	wire [15-1:0] node14755;
	wire [15-1:0] node14756;
	wire [15-1:0] node14759;
	wire [15-1:0] node14762;
	wire [15-1:0] node14763;
	wire [15-1:0] node14764;
	wire [15-1:0] node14765;
	wire [15-1:0] node14768;
	wire [15-1:0] node14770;
	wire [15-1:0] node14774;
	wire [15-1:0] node14776;
	wire [15-1:0] node14777;
	wire [15-1:0] node14779;
	wire [15-1:0] node14782;
	wire [15-1:0] node14785;
	wire [15-1:0] node14786;
	wire [15-1:0] node14787;
	wire [15-1:0] node14788;
	wire [15-1:0] node14789;
	wire [15-1:0] node14793;
	wire [15-1:0] node14795;
	wire [15-1:0] node14798;
	wire [15-1:0] node14799;
	wire [15-1:0] node14800;
	wire [15-1:0] node14801;
	wire [15-1:0] node14805;
	wire [15-1:0] node14808;
	wire [15-1:0] node14809;
	wire [15-1:0] node14810;
	wire [15-1:0] node14814;
	wire [15-1:0] node14817;
	wire [15-1:0] node14818;
	wire [15-1:0] node14819;
	wire [15-1:0] node14821;
	wire [15-1:0] node14822;
	wire [15-1:0] node14826;
	wire [15-1:0] node14827;
	wire [15-1:0] node14828;
	wire [15-1:0] node14832;
	wire [15-1:0] node14835;
	wire [15-1:0] node14836;
	wire [15-1:0] node14837;
	wire [15-1:0] node14840;
	wire [15-1:0] node14841;
	wire [15-1:0] node14843;
	wire [15-1:0] node14847;
	wire [15-1:0] node14850;
	wire [15-1:0] node14851;
	wire [15-1:0] node14852;
	wire [15-1:0] node14853;
	wire [15-1:0] node14854;
	wire [15-1:0] node14855;
	wire [15-1:0] node14856;
	wire [15-1:0] node14858;
	wire [15-1:0] node14861;
	wire [15-1:0] node14864;
	wire [15-1:0] node14866;
	wire [15-1:0] node14868;
	wire [15-1:0] node14871;
	wire [15-1:0] node14872;
	wire [15-1:0] node14873;
	wire [15-1:0] node14875;
	wire [15-1:0] node14878;
	wire [15-1:0] node14880;
	wire [15-1:0] node14881;
	wire [15-1:0] node14885;
	wire [15-1:0] node14886;
	wire [15-1:0] node14890;
	wire [15-1:0] node14891;
	wire [15-1:0] node14892;
	wire [15-1:0] node14893;
	wire [15-1:0] node14895;
	wire [15-1:0] node14898;
	wire [15-1:0] node14899;
	wire [15-1:0] node14903;
	wire [15-1:0] node14904;
	wire [15-1:0] node14907;
	wire [15-1:0] node14909;
	wire [15-1:0] node14910;
	wire [15-1:0] node14914;
	wire [15-1:0] node14915;
	wire [15-1:0] node14918;
	wire [15-1:0] node14919;
	wire [15-1:0] node14921;
	wire [15-1:0] node14925;
	wire [15-1:0] node14926;
	wire [15-1:0] node14927;
	wire [15-1:0] node14928;
	wire [15-1:0] node14929;
	wire [15-1:0] node14933;
	wire [15-1:0] node14934;
	wire [15-1:0] node14937;
	wire [15-1:0] node14939;
	wire [15-1:0] node14942;
	wire [15-1:0] node14943;
	wire [15-1:0] node14945;
	wire [15-1:0] node14948;
	wire [15-1:0] node14949;
	wire [15-1:0] node14953;
	wire [15-1:0] node14954;
	wire [15-1:0] node14955;
	wire [15-1:0] node14956;
	wire [15-1:0] node14957;
	wire [15-1:0] node14959;
	wire [15-1:0] node14963;
	wire [15-1:0] node14964;
	wire [15-1:0] node14966;
	wire [15-1:0] node14970;
	wire [15-1:0] node14971;
	wire [15-1:0] node14974;
	wire [15-1:0] node14975;
	wire [15-1:0] node14979;
	wire [15-1:0] node14980;
	wire [15-1:0] node14981;
	wire [15-1:0] node14983;
	wire [15-1:0] node14985;
	wire [15-1:0] node14988;
	wire [15-1:0] node14989;
	wire [15-1:0] node14993;
	wire [15-1:0] node14994;
	wire [15-1:0] node14997;
	wire [15-1:0] node15000;
	wire [15-1:0] node15001;
	wire [15-1:0] node15002;
	wire [15-1:0] node15003;
	wire [15-1:0] node15004;
	wire [15-1:0] node15005;
	wire [15-1:0] node15009;
	wire [15-1:0] node15010;
	wire [15-1:0] node15011;
	wire [15-1:0] node15013;
	wire [15-1:0] node15017;
	wire [15-1:0] node15020;
	wire [15-1:0] node15021;
	wire [15-1:0] node15023;
	wire [15-1:0] node15025;
	wire [15-1:0] node15028;
	wire [15-1:0] node15029;
	wire [15-1:0] node15033;
	wire [15-1:0] node15034;
	wire [15-1:0] node15035;
	wire [15-1:0] node15036;
	wire [15-1:0] node15037;
	wire [15-1:0] node15040;
	wire [15-1:0] node15042;
	wire [15-1:0] node15045;
	wire [15-1:0] node15046;
	wire [15-1:0] node15050;
	wire [15-1:0] node15052;
	wire [15-1:0] node15053;
	wire [15-1:0] node15057;
	wire [15-1:0] node15058;
	wire [15-1:0] node15059;
	wire [15-1:0] node15062;
	wire [15-1:0] node15063;
	wire [15-1:0] node15067;
	wire [15-1:0] node15068;
	wire [15-1:0] node15072;
	wire [15-1:0] node15073;
	wire [15-1:0] node15074;
	wire [15-1:0] node15075;
	wire [15-1:0] node15078;
	wire [15-1:0] node15079;
	wire [15-1:0] node15080;
	wire [15-1:0] node15082;
	wire [15-1:0] node15086;
	wire [15-1:0] node15088;
	wire [15-1:0] node15091;
	wire [15-1:0] node15092;
	wire [15-1:0] node15093;
	wire [15-1:0] node15097;
	wire [15-1:0] node15098;
	wire [15-1:0] node15101;
	wire [15-1:0] node15103;
	wire [15-1:0] node15106;
	wire [15-1:0] node15107;
	wire [15-1:0] node15108;
	wire [15-1:0] node15110;
	wire [15-1:0] node15113;
	wire [15-1:0] node15114;
	wire [15-1:0] node15117;
	wire [15-1:0] node15119;
	wire [15-1:0] node15122;
	wire [15-1:0] node15123;
	wire [15-1:0] node15124;
	wire [15-1:0] node15125;
	wire [15-1:0] node15129;
	wire [15-1:0] node15132;
	wire [15-1:0] node15133;
	wire [15-1:0] node15135;
	wire [15-1:0] node15138;
	wire [15-1:0] node15140;
	wire [15-1:0] node15141;
	wire [15-1:0] node15145;
	wire [15-1:0] node15146;
	wire [15-1:0] node15147;
	wire [15-1:0] node15148;
	wire [15-1:0] node15149;
	wire [15-1:0] node15150;
	wire [15-1:0] node15152;
	wire [15-1:0] node15153;
	wire [15-1:0] node15157;
	wire [15-1:0] node15158;
	wire [15-1:0] node15159;
	wire [15-1:0] node15161;
	wire [15-1:0] node15163;
	wire [15-1:0] node15166;
	wire [15-1:0] node15168;
	wire [15-1:0] node15171;
	wire [15-1:0] node15172;
	wire [15-1:0] node15176;
	wire [15-1:0] node15177;
	wire [15-1:0] node15178;
	wire [15-1:0] node15179;
	wire [15-1:0] node15180;
	wire [15-1:0] node15182;
	wire [15-1:0] node15185;
	wire [15-1:0] node15187;
	wire [15-1:0] node15190;
	wire [15-1:0] node15192;
	wire [15-1:0] node15193;
	wire [15-1:0] node15197;
	wire [15-1:0] node15198;
	wire [15-1:0] node15201;
	wire [15-1:0] node15202;
	wire [15-1:0] node15206;
	wire [15-1:0] node15207;
	wire [15-1:0] node15208;
	wire [15-1:0] node15209;
	wire [15-1:0] node15211;
	wire [15-1:0] node15215;
	wire [15-1:0] node15218;
	wire [15-1:0] node15219;
	wire [15-1:0] node15220;
	wire [15-1:0] node15225;
	wire [15-1:0] node15226;
	wire [15-1:0] node15227;
	wire [15-1:0] node15228;
	wire [15-1:0] node15229;
	wire [15-1:0] node15233;
	wire [15-1:0] node15234;
	wire [15-1:0] node15238;
	wire [15-1:0] node15239;
	wire [15-1:0] node15240;
	wire [15-1:0] node15243;
	wire [15-1:0] node15246;
	wire [15-1:0] node15247;
	wire [15-1:0] node15251;
	wire [15-1:0] node15252;
	wire [15-1:0] node15253;
	wire [15-1:0] node15254;
	wire [15-1:0] node15258;
	wire [15-1:0] node15259;
	wire [15-1:0] node15261;
	wire [15-1:0] node15264;
	wire [15-1:0] node15265;
	wire [15-1:0] node15269;
	wire [15-1:0] node15270;
	wire [15-1:0] node15271;
	wire [15-1:0] node15274;
	wire [15-1:0] node15277;
	wire [15-1:0] node15280;
	wire [15-1:0] node15281;
	wire [15-1:0] node15282;
	wire [15-1:0] node15283;
	wire [15-1:0] node15284;
	wire [15-1:0] node15285;
	wire [15-1:0] node15289;
	wire [15-1:0] node15290;
	wire [15-1:0] node15291;
	wire [15-1:0] node15296;
	wire [15-1:0] node15297;
	wire [15-1:0] node15298;
	wire [15-1:0] node15299;
	wire [15-1:0] node15300;
	wire [15-1:0] node15304;
	wire [15-1:0] node15307;
	wire [15-1:0] node15308;
	wire [15-1:0] node15312;
	wire [15-1:0] node15314;
	wire [15-1:0] node15317;
	wire [15-1:0] node15318;
	wire [15-1:0] node15319;
	wire [15-1:0] node15320;
	wire [15-1:0] node15321;
	wire [15-1:0] node15325;
	wire [15-1:0] node15328;
	wire [15-1:0] node15329;
	wire [15-1:0] node15333;
	wire [15-1:0] node15334;
	wire [15-1:0] node15335;
	wire [15-1:0] node15338;
	wire [15-1:0] node15341;
	wire [15-1:0] node15342;
	wire [15-1:0] node15344;
	wire [15-1:0] node15345;
	wire [15-1:0] node15349;
	wire [15-1:0] node15352;
	wire [15-1:0] node15353;
	wire [15-1:0] node15354;
	wire [15-1:0] node15355;
	wire [15-1:0] node15357;
	wire [15-1:0] node15359;
	wire [15-1:0] node15362;
	wire [15-1:0] node15363;
	wire [15-1:0] node15364;
	wire [15-1:0] node15368;
	wire [15-1:0] node15371;
	wire [15-1:0] node15372;
	wire [15-1:0] node15373;
	wire [15-1:0] node15374;
	wire [15-1:0] node15378;
	wire [15-1:0] node15381;
	wire [15-1:0] node15382;
	wire [15-1:0] node15383;
	wire [15-1:0] node15387;
	wire [15-1:0] node15390;
	wire [15-1:0] node15391;
	wire [15-1:0] node15392;
	wire [15-1:0] node15393;
	wire [15-1:0] node15396;
	wire [15-1:0] node15399;
	wire [15-1:0] node15400;
	wire [15-1:0] node15404;
	wire [15-1:0] node15405;
	wire [15-1:0] node15406;
	wire [15-1:0] node15409;
	wire [15-1:0] node15412;
	wire [15-1:0] node15413;
	wire [15-1:0] node15414;
	wire [15-1:0] node15416;
	wire [15-1:0] node15420;
	wire [15-1:0] node15421;
	wire [15-1:0] node15424;
	wire [15-1:0] node15426;
	wire [15-1:0] node15429;
	wire [15-1:0] node15430;
	wire [15-1:0] node15431;
	wire [15-1:0] node15432;
	wire [15-1:0] node15433;
	wire [15-1:0] node15435;
	wire [15-1:0] node15436;
	wire [15-1:0] node15438;
	wire [15-1:0] node15439;
	wire [15-1:0] node15444;
	wire [15-1:0] node15445;
	wire [15-1:0] node15446;
	wire [15-1:0] node15447;
	wire [15-1:0] node15451;
	wire [15-1:0] node15452;
	wire [15-1:0] node15455;
	wire [15-1:0] node15456;
	wire [15-1:0] node15460;
	wire [15-1:0] node15461;
	wire [15-1:0] node15462;
	wire [15-1:0] node15466;
	wire [15-1:0] node15469;
	wire [15-1:0] node15470;
	wire [15-1:0] node15471;
	wire [15-1:0] node15472;
	wire [15-1:0] node15473;
	wire [15-1:0] node15478;
	wire [15-1:0] node15479;
	wire [15-1:0] node15482;
	wire [15-1:0] node15485;
	wire [15-1:0] node15486;
	wire [15-1:0] node15487;
	wire [15-1:0] node15488;
	wire [15-1:0] node15492;
	wire [15-1:0] node15495;
	wire [15-1:0] node15496;
	wire [15-1:0] node15499;
	wire [15-1:0] node15500;
	wire [15-1:0] node15504;
	wire [15-1:0] node15505;
	wire [15-1:0] node15506;
	wire [15-1:0] node15507;
	wire [15-1:0] node15508;
	wire [15-1:0] node15512;
	wire [15-1:0] node15513;
	wire [15-1:0] node15517;
	wire [15-1:0] node15518;
	wire [15-1:0] node15519;
	wire [15-1:0] node15522;
	wire [15-1:0] node15524;
	wire [15-1:0] node15525;
	wire [15-1:0] node15529;
	wire [15-1:0] node15530;
	wire [15-1:0] node15531;
	wire [15-1:0] node15533;
	wire [15-1:0] node15536;
	wire [15-1:0] node15539;
	wire [15-1:0] node15542;
	wire [15-1:0] node15543;
	wire [15-1:0] node15544;
	wire [15-1:0] node15546;
	wire [15-1:0] node15548;
	wire [15-1:0] node15549;
	wire [15-1:0] node15553;
	wire [15-1:0] node15554;
	wire [15-1:0] node15557;
	wire [15-1:0] node15560;
	wire [15-1:0] node15561;
	wire [15-1:0] node15562;
	wire [15-1:0] node15564;
	wire [15-1:0] node15566;
	wire [15-1:0] node15569;
	wire [15-1:0] node15572;
	wire [15-1:0] node15574;
	wire [15-1:0] node15577;
	wire [15-1:0] node15578;
	wire [15-1:0] node15579;
	wire [15-1:0] node15580;
	wire [15-1:0] node15581;
	wire [15-1:0] node15585;
	wire [15-1:0] node15587;
	wire [15-1:0] node15588;
	wire [15-1:0] node15589;
	wire [15-1:0] node15593;
	wire [15-1:0] node15596;
	wire [15-1:0] node15597;
	wire [15-1:0] node15598;
	wire [15-1:0] node15600;
	wire [15-1:0] node15603;
	wire [15-1:0] node15605;
	wire [15-1:0] node15608;
	wire [15-1:0] node15609;
	wire [15-1:0] node15612;
	wire [15-1:0] node15613;
	wire [15-1:0] node15616;
	wire [15-1:0] node15617;
	wire [15-1:0] node15619;
	wire [15-1:0] node15623;
	wire [15-1:0] node15624;
	wire [15-1:0] node15625;
	wire [15-1:0] node15626;
	wire [15-1:0] node15627;
	wire [15-1:0] node15629;
	wire [15-1:0] node15633;
	wire [15-1:0] node15634;
	wire [15-1:0] node15637;
	wire [15-1:0] node15638;
	wire [15-1:0] node15642;
	wire [15-1:0] node15643;
	wire [15-1:0] node15644;
	wire [15-1:0] node15647;
	wire [15-1:0] node15649;
	wire [15-1:0] node15652;
	wire [15-1:0] node15653;
	wire [15-1:0] node15656;
	wire [15-1:0] node15658;
	wire [15-1:0] node15661;
	wire [15-1:0] node15662;
	wire [15-1:0] node15663;
	wire [15-1:0] node15665;
	wire [15-1:0] node15666;
	wire [15-1:0] node15668;
	wire [15-1:0] node15672;
	wire [15-1:0] node15673;
	wire [15-1:0] node15677;
	wire [15-1:0] node15678;
	wire [15-1:0] node15680;
	wire [15-1:0] node15681;
	wire [15-1:0] node15685;
	wire [15-1:0] node15687;
	wire [15-1:0] node15690;
	wire [15-1:0] node15691;
	wire [15-1:0] node15692;
	wire [15-1:0] node15693;
	wire [15-1:0] node15694;
	wire [15-1:0] node15695;
	wire [15-1:0] node15696;
	wire [15-1:0] node15697;
	wire [15-1:0] node15698;
	wire [15-1:0] node15700;
	wire [15-1:0] node15701;
	wire [15-1:0] node15705;
	wire [15-1:0] node15708;
	wire [15-1:0] node15710;
	wire [15-1:0] node15713;
	wire [15-1:0] node15714;
	wire [15-1:0] node15715;
	wire [15-1:0] node15717;
	wire [15-1:0] node15718;
	wire [15-1:0] node15723;
	wire [15-1:0] node15724;
	wire [15-1:0] node15728;
	wire [15-1:0] node15729;
	wire [15-1:0] node15730;
	wire [15-1:0] node15732;
	wire [15-1:0] node15733;
	wire [15-1:0] node15737;
	wire [15-1:0] node15738;
	wire [15-1:0] node15741;
	wire [15-1:0] node15744;
	wire [15-1:0] node15747;
	wire [15-1:0] node15748;
	wire [15-1:0] node15749;
	wire [15-1:0] node15750;
	wire [15-1:0] node15753;
	wire [15-1:0] node15755;
	wire [15-1:0] node15758;
	wire [15-1:0] node15759;
	wire [15-1:0] node15760;
	wire [15-1:0] node15761;
	wire [15-1:0] node15766;
	wire [15-1:0] node15768;
	wire [15-1:0] node15771;
	wire [15-1:0] node15772;
	wire [15-1:0] node15773;
	wire [15-1:0] node15774;
	wire [15-1:0] node15777;
	wire [15-1:0] node15780;
	wire [15-1:0] node15783;
	wire [15-1:0] node15784;
	wire [15-1:0] node15786;
	wire [15-1:0] node15789;
	wire [15-1:0] node15792;
	wire [15-1:0] node15793;
	wire [15-1:0] node15794;
	wire [15-1:0] node15795;
	wire [15-1:0] node15796;
	wire [15-1:0] node15797;
	wire [15-1:0] node15800;
	wire [15-1:0] node15801;
	wire [15-1:0] node15803;
	wire [15-1:0] node15807;
	wire [15-1:0] node15808;
	wire [15-1:0] node15809;
	wire [15-1:0] node15814;
	wire [15-1:0] node15815;
	wire [15-1:0] node15816;
	wire [15-1:0] node15819;
	wire [15-1:0] node15822;
	wire [15-1:0] node15823;
	wire [15-1:0] node15825;
	wire [15-1:0] node15829;
	wire [15-1:0] node15830;
	wire [15-1:0] node15831;
	wire [15-1:0] node15832;
	wire [15-1:0] node15834;
	wire [15-1:0] node15835;
	wire [15-1:0] node15839;
	wire [15-1:0] node15840;
	wire [15-1:0] node15842;
	wire [15-1:0] node15846;
	wire [15-1:0] node15848;
	wire [15-1:0] node15849;
	wire [15-1:0] node15853;
	wire [15-1:0] node15854;
	wire [15-1:0] node15856;
	wire [15-1:0] node15859;
	wire [15-1:0] node15860;
	wire [15-1:0] node15862;
	wire [15-1:0] node15865;
	wire [15-1:0] node15868;
	wire [15-1:0] node15869;
	wire [15-1:0] node15870;
	wire [15-1:0] node15871;
	wire [15-1:0] node15872;
	wire [15-1:0] node15873;
	wire [15-1:0] node15875;
	wire [15-1:0] node15878;
	wire [15-1:0] node15880;
	wire [15-1:0] node15883;
	wire [15-1:0] node15885;
	wire [15-1:0] node15887;
	wire [15-1:0] node15890;
	wire [15-1:0] node15891;
	wire [15-1:0] node15893;
	wire [15-1:0] node15897;
	wire [15-1:0] node15898;
	wire [15-1:0] node15899;
	wire [15-1:0] node15901;
	wire [15-1:0] node15905;
	wire [15-1:0] node15907;
	wire [15-1:0] node15908;
	wire [15-1:0] node15912;
	wire [15-1:0] node15913;
	wire [15-1:0] node15914;
	wire [15-1:0] node15916;
	wire [15-1:0] node15920;
	wire [15-1:0] node15921;
	wire [15-1:0] node15923;
	wire [15-1:0] node15924;
	wire [15-1:0] node15928;
	wire [15-1:0] node15929;
	wire [15-1:0] node15931;
	wire [15-1:0] node15932;
	wire [15-1:0] node15937;
	wire [15-1:0] node15938;
	wire [15-1:0] node15939;
	wire [15-1:0] node15940;
	wire [15-1:0] node15941;
	wire [15-1:0] node15942;
	wire [15-1:0] node15945;
	wire [15-1:0] node15946;
	wire [15-1:0] node15949;
	wire [15-1:0] node15952;
	wire [15-1:0] node15953;
	wire [15-1:0] node15954;
	wire [15-1:0] node15957;
	wire [15-1:0] node15961;
	wire [15-1:0] node15962;
	wire [15-1:0] node15964;
	wire [15-1:0] node15965;
	wire [15-1:0] node15967;
	wire [15-1:0] node15968;
	wire [15-1:0] node15973;
	wire [15-1:0] node15974;
	wire [15-1:0] node15975;
	wire [15-1:0] node15977;
	wire [15-1:0] node15981;
	wire [15-1:0] node15982;
	wire [15-1:0] node15986;
	wire [15-1:0] node15987;
	wire [15-1:0] node15988;
	wire [15-1:0] node15989;
	wire [15-1:0] node15990;
	wire [15-1:0] node15992;
	wire [15-1:0] node15995;
	wire [15-1:0] node15996;
	wire [15-1:0] node15998;
	wire [15-1:0] node16002;
	wire [15-1:0] node16003;
	wire [15-1:0] node16004;
	wire [15-1:0] node16008;
	wire [15-1:0] node16011;
	wire [15-1:0] node16012;
	wire [15-1:0] node16013;
	wire [15-1:0] node16017;
	wire [15-1:0] node16018;
	wire [15-1:0] node16020;
	wire [15-1:0] node16021;
	wire [15-1:0] node16025;
	wire [15-1:0] node16028;
	wire [15-1:0] node16029;
	wire [15-1:0] node16030;
	wire [15-1:0] node16031;
	wire [15-1:0] node16034;
	wire [15-1:0] node16037;
	wire [15-1:0] node16039;
	wire [15-1:0] node16041;
	wire [15-1:0] node16044;
	wire [15-1:0] node16045;
	wire [15-1:0] node16046;
	wire [15-1:0] node16048;
	wire [15-1:0] node16050;
	wire [15-1:0] node16054;
	wire [15-1:0] node16056;
	wire [15-1:0] node16059;
	wire [15-1:0] node16060;
	wire [15-1:0] node16061;
	wire [15-1:0] node16062;
	wire [15-1:0] node16063;
	wire [15-1:0] node16066;
	wire [15-1:0] node16067;
	wire [15-1:0] node16068;
	wire [15-1:0] node16072;
	wire [15-1:0] node16075;
	wire [15-1:0] node16076;
	wire [15-1:0] node16077;
	wire [15-1:0] node16078;
	wire [15-1:0] node16080;
	wire [15-1:0] node16084;
	wire [15-1:0] node16085;
	wire [15-1:0] node16087;
	wire [15-1:0] node16091;
	wire [15-1:0] node16092;
	wire [15-1:0] node16095;
	wire [15-1:0] node16098;
	wire [15-1:0] node16099;
	wire [15-1:0] node16100;
	wire [15-1:0] node16101;
	wire [15-1:0] node16104;
	wire [15-1:0] node16107;
	wire [15-1:0] node16108;
	wire [15-1:0] node16109;
	wire [15-1:0] node16111;
	wire [15-1:0] node16115;
	wire [15-1:0] node16118;
	wire [15-1:0] node16119;
	wire [15-1:0] node16120;
	wire [15-1:0] node16123;
	wire [15-1:0] node16126;
	wire [15-1:0] node16127;
	wire [15-1:0] node16130;
	wire [15-1:0] node16131;
	wire [15-1:0] node16135;
	wire [15-1:0] node16136;
	wire [15-1:0] node16137;
	wire [15-1:0] node16138;
	wire [15-1:0] node16139;
	wire [15-1:0] node16142;
	wire [15-1:0] node16144;
	wire [15-1:0] node16147;
	wire [15-1:0] node16148;
	wire [15-1:0] node16151;
	wire [15-1:0] node16154;
	wire [15-1:0] node16155;
	wire [15-1:0] node16156;
	wire [15-1:0] node16157;
	wire [15-1:0] node16161;
	wire [15-1:0] node16163;
	wire [15-1:0] node16165;
	wire [15-1:0] node16168;
	wire [15-1:0] node16169;
	wire [15-1:0] node16171;
	wire [15-1:0] node16173;
	wire [15-1:0] node16177;
	wire [15-1:0] node16178;
	wire [15-1:0] node16179;
	wire [15-1:0] node16181;
	wire [15-1:0] node16184;
	wire [15-1:0] node16185;
	wire [15-1:0] node16186;
	wire [15-1:0] node16190;
	wire [15-1:0] node16193;
	wire [15-1:0] node16194;
	wire [15-1:0] node16196;
	wire [15-1:0] node16199;
	wire [15-1:0] node16200;
	wire [15-1:0] node16203;
	wire [15-1:0] node16206;
	wire [15-1:0] node16207;
	wire [15-1:0] node16208;
	wire [15-1:0] node16209;
	wire [15-1:0] node16210;
	wire [15-1:0] node16211;
	wire [15-1:0] node16213;
	wire [15-1:0] node16214;
	wire [15-1:0] node16216;
	wire [15-1:0] node16219;
	wire [15-1:0] node16220;
	wire [15-1:0] node16224;
	wire [15-1:0] node16225;
	wire [15-1:0] node16226;
	wire [15-1:0] node16229;
	wire [15-1:0] node16231;
	wire [15-1:0] node16234;
	wire [15-1:0] node16235;
	wire [15-1:0] node16238;
	wire [15-1:0] node16241;
	wire [15-1:0] node16242;
	wire [15-1:0] node16243;
	wire [15-1:0] node16245;
	wire [15-1:0] node16248;
	wire [15-1:0] node16249;
	wire [15-1:0] node16252;
	wire [15-1:0] node16255;
	wire [15-1:0] node16256;
	wire [15-1:0] node16258;
	wire [15-1:0] node16261;
	wire [15-1:0] node16262;
	wire [15-1:0] node16266;
	wire [15-1:0] node16267;
	wire [15-1:0] node16268;
	wire [15-1:0] node16269;
	wire [15-1:0] node16270;
	wire [15-1:0] node16271;
	wire [15-1:0] node16275;
	wire [15-1:0] node16277;
	wire [15-1:0] node16278;
	wire [15-1:0] node16282;
	wire [15-1:0] node16283;
	wire [15-1:0] node16285;
	wire [15-1:0] node16287;
	wire [15-1:0] node16290;
	wire [15-1:0] node16293;
	wire [15-1:0] node16294;
	wire [15-1:0] node16295;
	wire [15-1:0] node16297;
	wire [15-1:0] node16301;
	wire [15-1:0] node16302;
	wire [15-1:0] node16306;
	wire [15-1:0] node16307;
	wire [15-1:0] node16308;
	wire [15-1:0] node16310;
	wire [15-1:0] node16311;
	wire [15-1:0] node16313;
	wire [15-1:0] node16317;
	wire [15-1:0] node16318;
	wire [15-1:0] node16321;
	wire [15-1:0] node16322;
	wire [15-1:0] node16326;
	wire [15-1:0] node16327;
	wire [15-1:0] node16330;
	wire [15-1:0] node16333;
	wire [15-1:0] node16334;
	wire [15-1:0] node16335;
	wire [15-1:0] node16336;
	wire [15-1:0] node16337;
	wire [15-1:0] node16338;
	wire [15-1:0] node16341;
	wire [15-1:0] node16343;
	wire [15-1:0] node16346;
	wire [15-1:0] node16347;
	wire [15-1:0] node16349;
	wire [15-1:0] node16352;
	wire [15-1:0] node16355;
	wire [15-1:0] node16356;
	wire [15-1:0] node16357;
	wire [15-1:0] node16361;
	wire [15-1:0] node16362;
	wire [15-1:0] node16365;
	wire [15-1:0] node16368;
	wire [15-1:0] node16369;
	wire [15-1:0] node16370;
	wire [15-1:0] node16372;
	wire [15-1:0] node16373;
	wire [15-1:0] node16375;
	wire [15-1:0] node16379;
	wire [15-1:0] node16380;
	wire [15-1:0] node16382;
	wire [15-1:0] node16385;
	wire [15-1:0] node16387;
	wire [15-1:0] node16390;
	wire [15-1:0] node16391;
	wire [15-1:0] node16392;
	wire [15-1:0] node16395;
	wire [15-1:0] node16396;
	wire [15-1:0] node16400;
	wire [15-1:0] node16401;
	wire [15-1:0] node16404;
	wire [15-1:0] node16406;
	wire [15-1:0] node16407;
	wire [15-1:0] node16411;
	wire [15-1:0] node16412;
	wire [15-1:0] node16413;
	wire [15-1:0] node16414;
	wire [15-1:0] node16416;
	wire [15-1:0] node16419;
	wire [15-1:0] node16420;
	wire [15-1:0] node16421;
	wire [15-1:0] node16425;
	wire [15-1:0] node16428;
	wire [15-1:0] node16429;
	wire [15-1:0] node16430;
	wire [15-1:0] node16432;
	wire [15-1:0] node16434;
	wire [15-1:0] node16438;
	wire [15-1:0] node16439;
	wire [15-1:0] node16442;
	wire [15-1:0] node16443;
	wire [15-1:0] node16447;
	wire [15-1:0] node16448;
	wire [15-1:0] node16449;
	wire [15-1:0] node16451;
	wire [15-1:0] node16454;
	wire [15-1:0] node16455;
	wire [15-1:0] node16458;
	wire [15-1:0] node16460;
	wire [15-1:0] node16461;
	wire [15-1:0] node16465;
	wire [15-1:0] node16466;
	wire [15-1:0] node16467;
	wire [15-1:0] node16469;
	wire [15-1:0] node16473;
	wire [15-1:0] node16474;
	wire [15-1:0] node16475;
	wire [15-1:0] node16480;
	wire [15-1:0] node16481;
	wire [15-1:0] node16482;
	wire [15-1:0] node16483;
	wire [15-1:0] node16484;
	wire [15-1:0] node16486;
	wire [15-1:0] node16488;
	wire [15-1:0] node16491;
	wire [15-1:0] node16492;
	wire [15-1:0] node16493;
	wire [15-1:0] node16494;
	wire [15-1:0] node16498;
	wire [15-1:0] node16499;
	wire [15-1:0] node16503;
	wire [15-1:0] node16504;
	wire [15-1:0] node16508;
	wire [15-1:0] node16509;
	wire [15-1:0] node16510;
	wire [15-1:0] node16511;
	wire [15-1:0] node16514;
	wire [15-1:0] node16517;
	wire [15-1:0] node16518;
	wire [15-1:0] node16521;
	wire [15-1:0] node16522;
	wire [15-1:0] node16526;
	wire [15-1:0] node16527;
	wire [15-1:0] node16528;
	wire [15-1:0] node16529;
	wire [15-1:0] node16533;
	wire [15-1:0] node16536;
	wire [15-1:0] node16537;
	wire [15-1:0] node16538;
	wire [15-1:0] node16542;
	wire [15-1:0] node16545;
	wire [15-1:0] node16546;
	wire [15-1:0] node16547;
	wire [15-1:0] node16548;
	wire [15-1:0] node16549;
	wire [15-1:0] node16551;
	wire [15-1:0] node16555;
	wire [15-1:0] node16558;
	wire [15-1:0] node16559;
	wire [15-1:0] node16561;
	wire [15-1:0] node16563;
	wire [15-1:0] node16564;
	wire [15-1:0] node16568;
	wire [15-1:0] node16569;
	wire [15-1:0] node16573;
	wire [15-1:0] node16574;
	wire [15-1:0] node16575;
	wire [15-1:0] node16577;
	wire [15-1:0] node16580;
	wire [15-1:0] node16581;
	wire [15-1:0] node16584;
	wire [15-1:0] node16585;
	wire [15-1:0] node16589;
	wire [15-1:0] node16590;
	wire [15-1:0] node16591;
	wire [15-1:0] node16592;
	wire [15-1:0] node16597;
	wire [15-1:0] node16599;
	wire [15-1:0] node16600;
	wire [15-1:0] node16602;
	wire [15-1:0] node16605;
	wire [15-1:0] node16607;
	wire [15-1:0] node16610;
	wire [15-1:0] node16611;
	wire [15-1:0] node16612;
	wire [15-1:0] node16613;
	wire [15-1:0] node16614;
	wire [15-1:0] node16616;
	wire [15-1:0] node16618;
	wire [15-1:0] node16619;
	wire [15-1:0] node16623;
	wire [15-1:0] node16624;
	wire [15-1:0] node16627;
	wire [15-1:0] node16630;
	wire [15-1:0] node16631;
	wire [15-1:0] node16632;
	wire [15-1:0] node16636;
	wire [15-1:0] node16639;
	wire [15-1:0] node16640;
	wire [15-1:0] node16641;
	wire [15-1:0] node16644;
	wire [15-1:0] node16645;
	wire [15-1:0] node16647;
	wire [15-1:0] node16650;
	wire [15-1:0] node16652;
	wire [15-1:0] node16655;
	wire [15-1:0] node16656;
	wire [15-1:0] node16658;
	wire [15-1:0] node16661;
	wire [15-1:0] node16662;
	wire [15-1:0] node16663;
	wire [15-1:0] node16667;
	wire [15-1:0] node16670;
	wire [15-1:0] node16671;
	wire [15-1:0] node16672;
	wire [15-1:0] node16673;
	wire [15-1:0] node16675;
	wire [15-1:0] node16678;
	wire [15-1:0] node16679;
	wire [15-1:0] node16682;
	wire [15-1:0] node16685;
	wire [15-1:0] node16686;
	wire [15-1:0] node16688;
	wire [15-1:0] node16691;
	wire [15-1:0] node16692;
	wire [15-1:0] node16695;
	wire [15-1:0] node16697;
	wire [15-1:0] node16699;
	wire [15-1:0] node16702;
	wire [15-1:0] node16703;
	wire [15-1:0] node16704;
	wire [15-1:0] node16705;
	wire [15-1:0] node16708;
	wire [15-1:0] node16711;
	wire [15-1:0] node16712;
	wire [15-1:0] node16715;
	wire [15-1:0] node16717;
	wire [15-1:0] node16719;
	wire [15-1:0] node16722;
	wire [15-1:0] node16723;
	wire [15-1:0] node16725;
	wire [15-1:0] node16728;
	wire [15-1:0] node16729;
	wire [15-1:0] node16732;
	wire [15-1:0] node16733;

	assign outp = (inp[7]) ? node8238 : node1;
		assign node1 = (inp[12]) ? node4181 : node2;
			assign node2 = (inp[8]) ? node2098 : node3;
				assign node3 = (inp[9]) ? node995 : node4;
					assign node4 = (inp[14]) ? node502 : node5;
						assign node5 = (inp[10]) ? node241 : node6;
							assign node6 = (inp[1]) ? node142 : node7;
								assign node7 = (inp[13]) ? node81 : node8;
									assign node8 = (inp[2]) ? node46 : node9;
										assign node9 = (inp[11]) ? node33 : node10;
											assign node10 = (inp[6]) ? node24 : node11;
												assign node11 = (inp[4]) ? node19 : node12;
													assign node12 = (inp[5]) ? node16 : node13;
														assign node13 = (inp[3]) ? 15'b011111111111111 : 15'b111111111111111;
														assign node16 = (inp[3]) ? 15'b001111111111111 : 15'b011111111111111;
													assign node19 = (inp[3]) ? node21 : 15'b001111111111111;
														assign node21 = (inp[5]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node24 = (inp[5]) ? 15'b000111111111111 : node25;
													assign node25 = (inp[4]) ? 15'b000111111111111 : node26;
														assign node26 = (inp[3]) ? node28 : 15'b001111111111111;
															assign node28 = (inp[0]) ? 15'b000111111111111 : 15'b001111111111111;
											assign node33 = (inp[4]) ? node41 : node34;
												assign node34 = (inp[3]) ? node36 : 15'b001111111111111;
													assign node36 = (inp[0]) ? 15'b000011111111111 : node37;
														assign node37 = (inp[5]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node41 = (inp[6]) ? node43 : 15'b000111111111111;
													assign node43 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node46 = (inp[11]) ? node62 : node47;
											assign node47 = (inp[0]) ? node51 : node48;
												assign node48 = (inp[5]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node51 = (inp[4]) ? node59 : node52;
													assign node52 = (inp[3]) ? 15'b000011111111111 : node53;
														assign node53 = (inp[6]) ? node55 : 15'b000111111111111;
															assign node55 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node59 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node62 = (inp[4]) ? node74 : node63;
												assign node63 = (inp[0]) ? node71 : node64;
													assign node64 = (inp[5]) ? 15'b000011111111111 : node65;
														assign node65 = (inp[6]) ? node67 : 15'b000111111111111;
															assign node67 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node71 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node74 = (inp[0]) ? node76 : 15'b000001111111111;
													assign node76 = (inp[3]) ? node78 : 15'b000001111111111;
														assign node78 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node81 = (inp[6]) ? node107 : node82;
										assign node82 = (inp[4]) ? node100 : node83;
											assign node83 = (inp[2]) ? node91 : node84;
												assign node84 = (inp[5]) ? 15'b000111111111111 : node85;
													assign node85 = (inp[3]) ? 15'b000111111111111 : node86;
														assign node86 = (inp[0]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node91 = (inp[5]) ? 15'b000001111111111 : node92;
													assign node92 = (inp[3]) ? 15'b000011111111111 : node93;
														assign node93 = (inp[0]) ? node95 : 15'b000111111111111;
															assign node95 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node100 = (inp[3]) ? node102 : 15'b000011111111111;
												assign node102 = (inp[5]) ? 15'b000000111111111 : node103;
													assign node103 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node107 = (inp[4]) ? node127 : node108;
											assign node108 = (inp[2]) ? node116 : node109;
												assign node109 = (inp[5]) ? node111 : 15'b000111111111111;
													assign node111 = (inp[3]) ? node113 : 15'b000011111111111;
														assign node113 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node116 = (inp[11]) ? node122 : node117;
													assign node117 = (inp[0]) ? node119 : 15'b000011111111111;
														assign node119 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node122 = (inp[5]) ? node124 : 15'b000001111111111;
														assign node124 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node127 = (inp[11]) ? node129 : 15'b000001111111111;
												assign node129 = (inp[2]) ? 15'b000000011111111 : node130;
													assign node130 = (inp[3]) ? node136 : node131;
														assign node131 = (inp[5]) ? 15'b000001111111111 : node132;
															assign node132 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
														assign node136 = (inp[5]) ? 15'b000000111111111 : node137;
															assign node137 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
								assign node142 = (inp[2]) ? node196 : node143;
									assign node143 = (inp[0]) ? node177 : node144;
										assign node144 = (inp[5]) ? node160 : node145;
											assign node145 = (inp[3]) ? node153 : node146;
												assign node146 = (inp[6]) ? node150 : node147;
													assign node147 = (inp[4]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node150 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node153 = (inp[13]) ? node157 : node154;
													assign node154 = (inp[6]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node157 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node160 = (inp[3]) ? node172 : node161;
												assign node161 = (inp[4]) ? node165 : node162;
													assign node162 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node165 = (inp[6]) ? 15'b000001111111111 : node166;
														assign node166 = (inp[13]) ? node168 : 15'b000011111111111;
															assign node168 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node172 = (inp[13]) ? node174 : 15'b000001111111111;
													assign node174 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node177 = (inp[4]) ? node189 : node178;
											assign node178 = (inp[11]) ? node186 : node179;
												assign node179 = (inp[3]) ? node181 : 15'b000111111111111;
													assign node181 = (inp[5]) ? node183 : 15'b000111111111111;
														assign node183 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node186 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node189 = (inp[11]) ? 15'b000000111111111 : node190;
												assign node190 = (inp[6]) ? node192 : 15'b000001111111111;
													assign node192 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node196 = (inp[11]) ? node220 : node197;
										assign node197 = (inp[5]) ? node213 : node198;
											assign node198 = (inp[13]) ? node202 : node199;
												assign node199 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node202 = (inp[6]) ? node210 : node203;
													assign node203 = (inp[0]) ? node205 : 15'b000001111111111;
														assign node205 = (inp[3]) ? node207 : 15'b000001111111111;
															assign node207 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node210 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node213 = (inp[0]) ? 15'b000000111111111 : node214;
												assign node214 = (inp[6]) ? 15'b000000111111111 : node215;
													assign node215 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node220 = (inp[4]) ? node230 : node221;
											assign node221 = (inp[13]) ? 15'b000000111111111 : node222;
												assign node222 = (inp[3]) ? node226 : node223;
													assign node223 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node226 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node230 = (inp[0]) ? 15'b000000011111111 : node231;
												assign node231 = (inp[3]) ? node235 : node232;
													assign node232 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node235 = (inp[5]) ? 15'b000000011111111 : node236;
														assign node236 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
							assign node241 = (inp[11]) ? node369 : node242;
								assign node242 = (inp[6]) ? node306 : node243;
									assign node243 = (inp[2]) ? node277 : node244;
										assign node244 = (inp[3]) ? node264 : node245;
											assign node245 = (inp[4]) ? node253 : node246;
												assign node246 = (inp[13]) ? node250 : node247;
													assign node247 = (inp[5]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node250 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node253 = (inp[0]) ? node255 : 15'b000111111111111;
													assign node255 = (inp[1]) ? 15'b000001111111111 : node256;
														assign node256 = (inp[5]) ? node260 : node257;
															assign node257 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
															assign node260 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node264 = (inp[5]) ? node272 : node265;
												assign node265 = (inp[0]) ? node269 : node266;
													assign node266 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node269 = (inp[13]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node272 = (inp[1]) ? node274 : 15'b000001111111111;
													assign node274 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node277 = (inp[5]) ? node295 : node278;
											assign node278 = (inp[0]) ? node288 : node279;
												assign node279 = (inp[3]) ? node285 : node280;
													assign node280 = (inp[13]) ? 15'b000011111111111 : node281;
														assign node281 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node285 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node288 = (inp[3]) ? node292 : node289;
													assign node289 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node292 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node295 = (inp[4]) ? node301 : node296;
												assign node296 = (inp[1]) ? 15'b000001111111111 : node297;
													assign node297 = (inp[13]) ? 15'b000001111111111 : 15'b000111111111111;
												assign node301 = (inp[0]) ? 15'b000000111111111 : node302;
													assign node302 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node306 = (inp[0]) ? node338 : node307;
										assign node307 = (inp[5]) ? node323 : node308;
											assign node308 = (inp[4]) ? node314 : node309;
												assign node309 = (inp[1]) ? node311 : 15'b000111111111111;
													assign node311 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node314 = (inp[13]) ? 15'b000001111111111 : node315;
													assign node315 = (inp[1]) ? node317 : 15'b000011111111111;
														assign node317 = (inp[2]) ? 15'b000001111111111 : node318;
															assign node318 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node323 = (inp[13]) ? node333 : node324;
												assign node324 = (inp[4]) ? node328 : node325;
													assign node325 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node328 = (inp[3]) ? node330 : 15'b000001111111111;
														assign node330 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node333 = (inp[4]) ? node335 : 15'b000001111111111;
													assign node335 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node338 = (inp[4]) ? node354 : node339;
											assign node339 = (inp[5]) ? node347 : node340;
												assign node340 = (inp[13]) ? node342 : 15'b000001111111111;
													assign node342 = (inp[1]) ? node344 : 15'b000001111111111;
														assign node344 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node347 = (inp[3]) ? 15'b000000111111111 : node348;
													assign node348 = (inp[1]) ? node350 : 15'b000001111111111;
														assign node350 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node354 = (inp[2]) ? node362 : node355;
												assign node355 = (inp[3]) ? node357 : 15'b000000111111111;
													assign node357 = (inp[1]) ? node359 : 15'b000000111111111;
														assign node359 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node362 = (inp[1]) ? node364 : 15'b000000011111111;
													assign node364 = (inp[3]) ? node366 : 15'b000000011111111;
														assign node366 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node369 = (inp[3]) ? node433 : node370;
									assign node370 = (inp[5]) ? node410 : node371;
										assign node371 = (inp[6]) ? node389 : node372;
											assign node372 = (inp[4]) ? node384 : node373;
												assign node373 = (inp[13]) ? 15'b000011111111111 : node374;
													assign node374 = (inp[1]) ? node378 : node375;
														assign node375 = (inp[0]) ? 15'b000111111111111 : 15'b001111111111111;
														assign node378 = (inp[0]) ? 15'b000011111111111 : node379;
															assign node379 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node384 = (inp[2]) ? 15'b000001111111111 : node385;
													assign node385 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node389 = (inp[2]) ? node403 : node390;
												assign node390 = (inp[13]) ? node396 : node391;
													assign node391 = (inp[4]) ? 15'b000001111111111 : node392;
														assign node392 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node396 = (inp[0]) ? node398 : 15'b000001111111111;
														assign node398 = (inp[1]) ? 15'b000000111111111 : node399;
															assign node399 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node403 = (inp[0]) ? node405 : 15'b000000111111111;
													assign node405 = (inp[4]) ? 15'b000000111111111 : node406;
														assign node406 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node410 = (inp[13]) ? node422 : node411;
											assign node411 = (inp[4]) ? node417 : node412;
												assign node412 = (inp[0]) ? node414 : 15'b000011111111111;
													assign node414 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node417 = (inp[0]) ? 15'b000000111111111 : node418;
													assign node418 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node422 = (inp[4]) ? node426 : node423;
												assign node423 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node426 = (inp[0]) ? node430 : node427;
													assign node427 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node430 = (inp[6]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node433 = (inp[2]) ? node459 : node434;
										assign node434 = (inp[13]) ? node442 : node435;
											assign node435 = (inp[1]) ? node439 : node436;
												assign node436 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node439 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node442 = (inp[5]) ? node450 : node443;
												assign node443 = (inp[4]) ? node447 : node444;
													assign node444 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node447 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node450 = (inp[6]) ? 15'b000000001111111 : node451;
													assign node451 = (inp[4]) ? 15'b000000011111111 : node452;
														assign node452 = (inp[0]) ? node454 : 15'b000000111111111;
															assign node454 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node459 = (inp[4]) ? node487 : node460;
											assign node460 = (inp[0]) ? node468 : node461;
												assign node461 = (inp[1]) ? 15'b000000011111111 : node462;
													assign node462 = (inp[6]) ? 15'b000000111111111 : node463;
														assign node463 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node468 = (inp[5]) ? node476 : node469;
													assign node469 = (inp[1]) ? 15'b000000011111111 : node470;
														assign node470 = (inp[6]) ? node472 : 15'b000000111111111;
															assign node472 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node476 = (inp[13]) ? node482 : node477;
														assign node477 = (inp[1]) ? 15'b000000011111111 : node478;
															assign node478 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node482 = (inp[1]) ? 15'b000000001111111 : node483;
															assign node483 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node487 = (inp[5]) ? node495 : node488;
												assign node488 = (inp[1]) ? 15'b000000001111111 : node489;
													assign node489 = (inp[0]) ? node491 : 15'b000000111111111;
														assign node491 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node495 = (inp[0]) ? node497 : 15'b000000001111111;
													assign node497 = (inp[6]) ? node499 : 15'b000000001111111;
														assign node499 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node502 = (inp[2]) ? node726 : node503;
							assign node503 = (inp[13]) ? node623 : node504;
								assign node504 = (inp[10]) ? node556 : node505;
									assign node505 = (inp[1]) ? node525 : node506;
										assign node506 = (inp[11]) ? node516 : node507;
											assign node507 = (inp[6]) ? node509 : 15'b000111111111111;
												assign node509 = (inp[5]) ? 15'b000011111111111 : node510;
													assign node510 = (inp[4]) ? 15'b000011111111111 : node511;
														assign node511 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node516 = (inp[6]) ? node522 : node517;
												assign node517 = (inp[0]) ? node519 : 15'b000011111111111;
													assign node519 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node522 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node525 = (inp[11]) ? node543 : node526;
											assign node526 = (inp[3]) ? node532 : node527;
												assign node527 = (inp[6]) ? node529 : 15'b000011111111111;
													assign node529 = (inp[5]) ? 15'b000011111111111 : 15'b000001111111111;
												assign node532 = (inp[0]) ? node540 : node533;
													assign node533 = (inp[4]) ? 15'b000001111111111 : node534;
														assign node534 = (inp[6]) ? 15'b000011111111111 : node535;
															assign node535 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node540 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node543 = (inp[6]) ? node551 : node544;
												assign node544 = (inp[5]) ? 15'b000001111111111 : node545;
													assign node545 = (inp[0]) ? 15'b000001111111111 : node546;
														assign node546 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node551 = (inp[0]) ? 15'b000000011111111 : node552;
													assign node552 = (inp[3]) ? 15'b000001111111111 : 15'b000000111111111;
									assign node556 = (inp[0]) ? node594 : node557;
										assign node557 = (inp[3]) ? node571 : node558;
											assign node558 = (inp[11]) ? node564 : node559;
												assign node559 = (inp[5]) ? 15'b000011111111111 : node560;
													assign node560 = (inp[4]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node564 = (inp[4]) ? node568 : node565;
													assign node565 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node568 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node571 = (inp[1]) ? node587 : node572;
												assign node572 = (inp[11]) ? node578 : node573;
													assign node573 = (inp[4]) ? node575 : 15'b000011111111111;
														assign node575 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node578 = (inp[6]) ? node584 : node579;
														assign node579 = (inp[4]) ? 15'b000001111111111 : node580;
															assign node580 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
														assign node584 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node587 = (inp[6]) ? node589 : 15'b000000111111111;
													assign node589 = (inp[4]) ? node591 : 15'b000000111111111;
														assign node591 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node594 = (inp[11]) ? node612 : node595;
											assign node595 = (inp[5]) ? node605 : node596;
												assign node596 = (inp[3]) ? node600 : node597;
													assign node597 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node600 = (inp[6]) ? 15'b000000111111111 : node601;
														assign node601 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node605 = (inp[1]) ? node609 : node606;
													assign node606 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node609 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node612 = (inp[5]) ? node618 : node613;
												assign node613 = (inp[1]) ? node615 : 15'b000000111111111;
													assign node615 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node618 = (inp[6]) ? 15'b000000001111111 : node619;
													assign node619 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node623 = (inp[6]) ? node665 : node624;
									assign node624 = (inp[5]) ? node648 : node625;
										assign node625 = (inp[0]) ? node637 : node626;
											assign node626 = (inp[10]) ? 15'b000001111111111 : node627;
												assign node627 = (inp[3]) ? node631 : node628;
													assign node628 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node631 = (inp[4]) ? node633 : 15'b000011111111111;
														assign node633 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node637 = (inp[11]) ? node643 : node638;
												assign node638 = (inp[4]) ? node640 : 15'b000001111111111;
													assign node640 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node643 = (inp[1]) ? node645 : 15'b000001111111111;
													assign node645 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node648 = (inp[11]) ? node660 : node649;
											assign node649 = (inp[1]) ? node655 : node650;
												assign node650 = (inp[0]) ? 15'b000000111111111 : node651;
													assign node651 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node655 = (inp[4]) ? 15'b000000011111111 : node656;
													assign node656 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node660 = (inp[10]) ? node662 : 15'b000000011111111;
												assign node662 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node665 = (inp[1]) ? node701 : node666;
										assign node666 = (inp[11]) ? node688 : node667;
											assign node667 = (inp[4]) ? node675 : node668;
												assign node668 = (inp[10]) ? node670 : 15'b000001111111111;
													assign node670 = (inp[0]) ? node672 : 15'b000001111111111;
														assign node672 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node675 = (inp[10]) ? node683 : node676;
													assign node676 = (inp[0]) ? 15'b000000111111111 : node677;
														assign node677 = (inp[5]) ? node679 : 15'b000001111111111;
															assign node679 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node683 = (inp[3]) ? node685 : 15'b000000111111111;
														assign node685 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node688 = (inp[10]) ? node690 : 15'b000000111111111;
												assign node690 = (inp[0]) ? node698 : node691;
													assign node691 = (inp[3]) ? 15'b000000011111111 : node692;
														assign node692 = (inp[4]) ? 15'b000000111111111 : node693;
															assign node693 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node698 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node701 = (inp[3]) ? node711 : node702;
											assign node702 = (inp[10]) ? node708 : node703;
												assign node703 = (inp[4]) ? 15'b000000111111111 : node704;
													assign node704 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node708 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node711 = (inp[0]) ? node723 : node712;
												assign node712 = (inp[11]) ? node718 : node713;
													assign node713 = (inp[4]) ? node715 : 15'b000000111111111;
														assign node715 = (inp[10]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node718 = (inp[4]) ? node720 : 15'b000000011111111;
														assign node720 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node723 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node726 = (inp[3]) ? node866 : node727;
								assign node727 = (inp[11]) ? node787 : node728;
									assign node728 = (inp[6]) ? node760 : node729;
										assign node729 = (inp[4]) ? node743 : node730;
											assign node730 = (inp[10]) ? node738 : node731;
												assign node731 = (inp[1]) ? 15'b000011111111111 : node732;
													assign node732 = (inp[5]) ? node734 : 15'b000111111111111;
														assign node734 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node738 = (inp[5]) ? 15'b000001111111111 : node739;
													assign node739 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node743 = (inp[13]) ? node753 : node744;
												assign node744 = (inp[0]) ? node746 : 15'b000111111111111;
													assign node746 = (inp[5]) ? 15'b000000111111111 : node747;
														assign node747 = (inp[10]) ? 15'b000001111111111 : node748;
															assign node748 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node753 = (inp[0]) ? node757 : node754;
													assign node754 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node757 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node760 = (inp[10]) ? node778 : node761;
											assign node761 = (inp[4]) ? node763 : 15'b000001111111111;
												assign node763 = (inp[5]) ? node769 : node764;
													assign node764 = (inp[13]) ? node766 : 15'b000001111111111;
														assign node766 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node769 = (inp[13]) ? node775 : node770;
														assign node770 = (inp[1]) ? 15'b000000111111111 : node771;
															assign node771 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node775 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node778 = (inp[0]) ? node784 : node779;
												assign node779 = (inp[1]) ? 15'b000000111111111 : node780;
													assign node780 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node784 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node787 = (inp[13]) ? node825 : node788;
										assign node788 = (inp[4]) ? node808 : node789;
											assign node789 = (inp[6]) ? node801 : node790;
												assign node790 = (inp[5]) ? node796 : node791;
													assign node791 = (inp[0]) ? 15'b000011111111111 : node792;
														assign node792 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node796 = (inp[0]) ? 15'b000001111111111 : node797;
														assign node797 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node801 = (inp[0]) ? 15'b000000011111111 : node802;
													assign node802 = (inp[5]) ? node804 : 15'b000001111111111;
														assign node804 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node808 = (inp[1]) ? node818 : node809;
												assign node809 = (inp[0]) ? node813 : node810;
													assign node810 = (inp[6]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node813 = (inp[5]) ? node815 : 15'b000000111111111;
														assign node815 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node818 = (inp[0]) ? 15'b000000001111111 : node819;
													assign node819 = (inp[6]) ? 15'b000000011111111 : node820;
														assign node820 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node825 = (inp[5]) ? node847 : node826;
											assign node826 = (inp[4]) ? node840 : node827;
												assign node827 = (inp[6]) ? node833 : node828;
													assign node828 = (inp[0]) ? 15'b000000111111111 : node829;
														assign node829 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node833 = (inp[1]) ? 15'b000000011111111 : node834;
														assign node834 = (inp[0]) ? node836 : 15'b000000111111111;
															assign node836 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node840 = (inp[1]) ? node842 : 15'b000000011111111;
													assign node842 = (inp[0]) ? node844 : 15'b000000011111111;
														assign node844 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node847 = (inp[10]) ? node861 : node848;
												assign node848 = (inp[6]) ? node854 : node849;
													assign node849 = (inp[4]) ? node851 : 15'b000000011111111;
														assign node851 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node854 = (inp[4]) ? node858 : node855;
														assign node855 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node858 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node861 = (inp[6]) ? node863 : 15'b000000001111111;
													assign node863 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node866 = (inp[5]) ? node938 : node867;
									assign node867 = (inp[6]) ? node891 : node868;
										assign node868 = (inp[4]) ? node876 : node869;
											assign node869 = (inp[13]) ? node873 : node870;
												assign node870 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node873 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node876 = (inp[10]) ? node886 : node877;
												assign node877 = (inp[13]) ? node881 : node878;
													assign node878 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node881 = (inp[1]) ? node883 : 15'b000000111111111;
														assign node883 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node886 = (inp[13]) ? node888 : 15'b000000111111111;
													assign node888 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node891 = (inp[1]) ? node917 : node892;
											assign node892 = (inp[13]) ? node906 : node893;
												assign node893 = (inp[10]) ? node899 : node894;
													assign node894 = (inp[4]) ? 15'b000000111111111 : node895;
														assign node895 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node899 = (inp[11]) ? 15'b000000011111111 : node900;
														assign node900 = (inp[0]) ? node902 : 15'b000000111111111;
															assign node902 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node906 = (inp[11]) ? node912 : node907;
													assign node907 = (inp[10]) ? node909 : 15'b000000111111111;
														assign node909 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node912 = (inp[4]) ? node914 : 15'b000000011111111;
														assign node914 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node917 = (inp[11]) ? node929 : node918;
												assign node918 = (inp[13]) ? node924 : node919;
													assign node919 = (inp[4]) ? 15'b000000011111111 : node920;
														assign node920 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node924 = (inp[10]) ? node926 : 15'b000000011111111;
														assign node926 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node929 = (inp[10]) ? node935 : node930;
													assign node930 = (inp[0]) ? 15'b000000001111111 : node931;
														assign node931 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node935 = (inp[4]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node938 = (inp[6]) ? node972 : node939;
										assign node939 = (inp[10]) ? node959 : node940;
											assign node940 = (inp[13]) ? node952 : node941;
												assign node941 = (inp[11]) ? node949 : node942;
													assign node942 = (inp[4]) ? node944 : 15'b000001111111111;
														assign node944 = (inp[1]) ? 15'b000000111111111 : node945;
															assign node945 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node949 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node952 = (inp[1]) ? node956 : node953;
													assign node953 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node956 = (inp[11]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node959 = (inp[13]) ? node965 : node960;
												assign node960 = (inp[4]) ? node962 : 15'b000000111111111;
													assign node962 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node965 = (inp[11]) ? node969 : node966;
													assign node966 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node969 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node972 = (inp[0]) ? node982 : node973;
											assign node973 = (inp[10]) ? node975 : 15'b000000011111111;
												assign node975 = (inp[1]) ? node977 : 15'b000000011111111;
													assign node977 = (inp[11]) ? node979 : 15'b000000001111111;
														assign node979 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node982 = (inp[1]) ? node990 : node983;
												assign node983 = (inp[13]) ? 15'b000000001111111 : node984;
													assign node984 = (inp[10]) ? node986 : 15'b000000001111111;
														assign node986 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node990 = (inp[13]) ? 15'b000000000011111 : node991;
													assign node991 = (inp[11]) ? 15'b000000000011111 : 15'b000000001111111;
					assign node995 = (inp[4]) ? node1589 : node996;
						assign node996 = (inp[6]) ? node1310 : node997;
							assign node997 = (inp[5]) ? node1181 : node998;
								assign node998 = (inp[11]) ? node1090 : node999;
									assign node999 = (inp[13]) ? node1049 : node1000;
										assign node1000 = (inp[2]) ? node1036 : node1001;
											assign node1001 = (inp[0]) ? node1017 : node1002;
												assign node1002 = (inp[14]) ? node1010 : node1003;
													assign node1003 = (inp[1]) ? node1007 : node1004;
														assign node1004 = (inp[3]) ? 15'b001111111111111 : 15'b011111111111111;
														assign node1007 = (inp[3]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node1010 = (inp[3]) ? 15'b000011111111111 : node1011;
														assign node1011 = (inp[1]) ? node1013 : 15'b000111111111111;
															assign node1013 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node1017 = (inp[1]) ? node1029 : node1018;
													assign node1018 = (inp[3]) ? node1024 : node1019;
														assign node1019 = (inp[14]) ? node1021 : 15'b000111111111111;
															assign node1021 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
														assign node1024 = (inp[14]) ? 15'b000011111111111 : node1025;
															assign node1025 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1029 = (inp[3]) ? node1031 : 15'b000011111111111;
														assign node1031 = (inp[10]) ? 15'b000001111111111 : node1032;
															assign node1032 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1036 = (inp[1]) ? node1044 : node1037;
												assign node1037 = (inp[0]) ? node1039 : 15'b000111111111111;
													assign node1039 = (inp[10]) ? node1041 : 15'b000011111111111;
														assign node1041 = (inp[3]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node1044 = (inp[10]) ? 15'b000001111111111 : node1045;
													assign node1045 = (inp[3]) ? 15'b000001111111111 : 15'b000111111111111;
										assign node1049 = (inp[10]) ? node1067 : node1050;
											assign node1050 = (inp[3]) ? node1060 : node1051;
												assign node1051 = (inp[14]) ? node1057 : node1052;
													assign node1052 = (inp[2]) ? 15'b000011111111111 : node1053;
														assign node1053 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1057 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1060 = (inp[1]) ? 15'b000001111111111 : node1061;
													assign node1061 = (inp[2]) ? node1063 : 15'b000011111111111;
														assign node1063 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1067 = (inp[14]) ? node1081 : node1068;
												assign node1068 = (inp[1]) ? node1076 : node1069;
													assign node1069 = (inp[0]) ? node1071 : 15'b000011111111111;
														assign node1071 = (inp[2]) ? 15'b000001111111111 : node1072;
															assign node1072 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1076 = (inp[3]) ? 15'b000000111111111 : node1077;
														assign node1077 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1081 = (inp[3]) ? node1087 : node1082;
													assign node1082 = (inp[2]) ? 15'b000000111111111 : node1083;
														assign node1083 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1087 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1090 = (inp[13]) ? node1140 : node1091;
										assign node1091 = (inp[14]) ? node1119 : node1092;
											assign node1092 = (inp[3]) ? node1106 : node1093;
												assign node1093 = (inp[0]) ? node1101 : node1094;
													assign node1094 = (inp[1]) ? node1096 : 15'b000111111111111;
														assign node1096 = (inp[10]) ? 15'b000011111111111 : node1097;
															assign node1097 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1101 = (inp[10]) ? node1103 : 15'b000011111111111;
														assign node1103 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1106 = (inp[2]) ? node1112 : node1107;
													assign node1107 = (inp[1]) ? node1109 : 15'b000011111111111;
														assign node1109 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1112 = (inp[10]) ? 15'b000000111111111 : node1113;
														assign node1113 = (inp[1]) ? node1115 : 15'b000001111111111;
															assign node1115 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1119 = (inp[3]) ? node1131 : node1120;
												assign node1120 = (inp[0]) ? node1126 : node1121;
													assign node1121 = (inp[10]) ? 15'b000001111111111 : node1122;
														assign node1122 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1126 = (inp[2]) ? node1128 : 15'b000001111111111;
														assign node1128 = (inp[10]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node1131 = (inp[10]) ? 15'b000000111111111 : node1132;
													assign node1132 = (inp[0]) ? 15'b000000111111111 : node1133;
														assign node1133 = (inp[1]) ? node1135 : 15'b000001111111111;
															assign node1135 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node1140 = (inp[10]) ? node1158 : node1141;
											assign node1141 = (inp[1]) ? node1151 : node1142;
												assign node1142 = (inp[14]) ? node1148 : node1143;
													assign node1143 = (inp[3]) ? 15'b000001111111111 : node1144;
														assign node1144 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1148 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1151 = (inp[2]) ? 15'b000000111111111 : node1152;
													assign node1152 = (inp[3]) ? 15'b000000111111111 : node1153;
														assign node1153 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1158 = (inp[3]) ? node1174 : node1159;
												assign node1159 = (inp[0]) ? node1171 : node1160;
													assign node1160 = (inp[2]) ? node1166 : node1161;
														assign node1161 = (inp[1]) ? node1163 : 15'b000001111111111;
															assign node1163 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node1166 = (inp[14]) ? 15'b000000111111111 : node1167;
															assign node1167 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1171 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node1174 = (inp[0]) ? node1176 : 15'b000000011111111;
													assign node1176 = (inp[1]) ? 15'b000000000111111 : node1177;
														assign node1177 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node1181 = (inp[10]) ? node1239 : node1182;
									assign node1182 = (inp[13]) ? node1212 : node1183;
										assign node1183 = (inp[14]) ? node1199 : node1184;
											assign node1184 = (inp[3]) ? node1186 : 15'b000111111111111;
												assign node1186 = (inp[0]) ? node1192 : node1187;
													assign node1187 = (inp[1]) ? node1189 : 15'b000011111111111;
														assign node1189 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1192 = (inp[11]) ? 15'b000001111111111 : node1193;
														assign node1193 = (inp[2]) ? 15'b000001111111111 : node1194;
															assign node1194 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1199 = (inp[11]) ? node1207 : node1200;
												assign node1200 = (inp[1]) ? node1204 : node1201;
													assign node1201 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1204 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1207 = (inp[3]) ? node1209 : 15'b000001111111111;
													assign node1209 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1212 = (inp[3]) ? node1222 : node1213;
											assign node1213 = (inp[0]) ? 15'b000000111111111 : node1214;
												assign node1214 = (inp[11]) ? node1218 : node1215;
													assign node1215 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1218 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1222 = (inp[14]) ? node1232 : node1223;
												assign node1223 = (inp[0]) ? node1227 : node1224;
													assign node1224 = (inp[2]) ? 15'b000001111111111 : 15'b000000111111111;
													assign node1227 = (inp[1]) ? node1229 : 15'b000000111111111;
														assign node1229 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1232 = (inp[1]) ? node1236 : node1233;
													assign node1233 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1236 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1239 = (inp[1]) ? node1271 : node1240;
										assign node1240 = (inp[11]) ? node1252 : node1241;
											assign node1241 = (inp[0]) ? node1247 : node1242;
												assign node1242 = (inp[2]) ? node1244 : 15'b000011111111111;
													assign node1244 = (inp[14]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node1247 = (inp[13]) ? 15'b000000011111111 : node1248;
													assign node1248 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1252 = (inp[13]) ? node1264 : node1253;
												assign node1253 = (inp[3]) ? node1259 : node1254;
													assign node1254 = (inp[0]) ? 15'b000000111111111 : node1255;
														assign node1255 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1259 = (inp[0]) ? 15'b000000011111111 : node1260;
														assign node1260 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1264 = (inp[14]) ? 15'b000000011111111 : node1265;
													assign node1265 = (inp[2]) ? node1267 : 15'b000000111111111;
														assign node1267 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1271 = (inp[11]) ? node1291 : node1272;
											assign node1272 = (inp[2]) ? node1286 : node1273;
												assign node1273 = (inp[3]) ? node1279 : node1274;
													assign node1274 = (inp[13]) ? 15'b000000111111111 : node1275;
														assign node1275 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1279 = (inp[0]) ? 15'b000000011111111 : node1280;
														assign node1280 = (inp[13]) ? node1282 : 15'b000001111111111;
															assign node1282 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1286 = (inp[0]) ? node1288 : 15'b000000011111111;
													assign node1288 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1291 = (inp[13]) ? node1299 : node1292;
												assign node1292 = (inp[0]) ? 15'b000000011111111 : node1293;
													assign node1293 = (inp[2]) ? 15'b000000011111111 : node1294;
														assign node1294 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1299 = (inp[3]) ? node1307 : node1300;
													assign node1300 = (inp[2]) ? node1302 : 15'b000000011111111;
														assign node1302 = (inp[14]) ? 15'b000000001111111 : node1303;
															assign node1303 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1307 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node1310 = (inp[13]) ? node1434 : node1311;
								assign node1311 = (inp[14]) ? node1379 : node1312;
									assign node1312 = (inp[10]) ? node1350 : node1313;
										assign node1313 = (inp[3]) ? node1331 : node1314;
											assign node1314 = (inp[1]) ? node1324 : node1315;
												assign node1315 = (inp[2]) ? node1319 : node1316;
													assign node1316 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node1319 = (inp[5]) ? node1321 : 15'b000011111111111;
														assign node1321 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1324 = (inp[2]) ? 15'b000001111111111 : node1325;
													assign node1325 = (inp[0]) ? node1327 : 15'b000011111111111;
														assign node1327 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1331 = (inp[11]) ? node1341 : node1332;
												assign node1332 = (inp[0]) ? 15'b000001111111111 : node1333;
													assign node1333 = (inp[1]) ? node1335 : 15'b000111111111111;
														assign node1335 = (inp[5]) ? 15'b000001111111111 : node1336;
															assign node1336 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1341 = (inp[0]) ? node1345 : node1342;
													assign node1342 = (inp[2]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node1345 = (inp[1]) ? 15'b000000011111111 : node1346;
														assign node1346 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1350 = (inp[5]) ? node1364 : node1351;
											assign node1351 = (inp[3]) ? node1359 : node1352;
												assign node1352 = (inp[1]) ? node1356 : node1353;
													assign node1353 = (inp[2]) ? 15'b000011111111111 : 15'b000001111111111;
													assign node1356 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1359 = (inp[2]) ? 15'b000000111111111 : node1360;
													assign node1360 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1364 = (inp[2]) ? node1376 : node1365;
												assign node1365 = (inp[11]) ? node1373 : node1366;
													assign node1366 = (inp[0]) ? 15'b000000111111111 : node1367;
														assign node1367 = (inp[1]) ? 15'b000001111111111 : node1368;
															assign node1368 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1373 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1376 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node1379 = (inp[1]) ? node1405 : node1380;
										assign node1380 = (inp[0]) ? node1388 : node1381;
											assign node1381 = (inp[2]) ? node1385 : node1382;
												assign node1382 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1385 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1388 = (inp[10]) ? node1398 : node1389;
												assign node1389 = (inp[3]) ? 15'b000000011111111 : node1390;
													assign node1390 = (inp[11]) ? node1392 : 15'b000001111111111;
														assign node1392 = (inp[2]) ? 15'b000000111111111 : node1393;
															assign node1393 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1398 = (inp[11]) ? node1400 : 15'b000000011111111;
													assign node1400 = (inp[3]) ? 15'b000000001111111 : node1401;
														assign node1401 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1405 = (inp[0]) ? node1419 : node1406;
											assign node1406 = (inp[3]) ? node1408 : 15'b000000111111111;
												assign node1408 = (inp[11]) ? node1412 : node1409;
													assign node1409 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1412 = (inp[2]) ? 15'b000000001111111 : node1413;
														assign node1413 = (inp[10]) ? node1415 : 15'b000000011111111;
															assign node1415 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1419 = (inp[5]) ? node1429 : node1420;
												assign node1420 = (inp[11]) ? node1424 : node1421;
													assign node1421 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1424 = (inp[3]) ? node1426 : 15'b000000011111111;
														assign node1426 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1429 = (inp[10]) ? 15'b000000001111111 : node1430;
													assign node1430 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1434 = (inp[5]) ? node1514 : node1435;
									assign node1435 = (inp[11]) ? node1471 : node1436;
										assign node1436 = (inp[1]) ? node1448 : node1437;
											assign node1437 = (inp[2]) ? node1441 : node1438;
												assign node1438 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1441 = (inp[0]) ? 15'b000000111111111 : node1442;
													assign node1442 = (inp[10]) ? node1444 : 15'b000000111111111;
														assign node1444 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1448 = (inp[10]) ? node1458 : node1449;
												assign node1449 = (inp[3]) ? node1455 : node1450;
													assign node1450 = (inp[14]) ? 15'b000000111111111 : node1451;
														assign node1451 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1455 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1458 = (inp[2]) ? node1466 : node1459;
													assign node1459 = (inp[3]) ? 15'b000000011111111 : node1460;
														assign node1460 = (inp[14]) ? node1462 : 15'b000000111111111;
															assign node1462 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1466 = (inp[14]) ? 15'b000000001111111 : node1467;
														assign node1467 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1471 = (inp[2]) ? node1491 : node1472;
											assign node1472 = (inp[0]) ? node1484 : node1473;
												assign node1473 = (inp[10]) ? node1479 : node1474;
													assign node1474 = (inp[1]) ? 15'b000001111111111 : node1475;
														assign node1475 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1479 = (inp[1]) ? node1481 : 15'b000000111111111;
														assign node1481 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1484 = (inp[1]) ? 15'b000000001111111 : node1485;
													assign node1485 = (inp[14]) ? 15'b000000011111111 : node1486;
														assign node1486 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1491 = (inp[1]) ? node1503 : node1492;
												assign node1492 = (inp[0]) ? node1500 : node1493;
													assign node1493 = (inp[10]) ? 15'b000000011111111 : node1494;
														assign node1494 = (inp[14]) ? node1496 : 15'b000000111111111;
															assign node1496 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1500 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1503 = (inp[0]) ? node1511 : node1504;
													assign node1504 = (inp[14]) ? 15'b000000001111111 : node1505;
														assign node1505 = (inp[10]) ? node1507 : 15'b000000011111111;
															assign node1507 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1511 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1514 = (inp[3]) ? node1542 : node1515;
										assign node1515 = (inp[2]) ? node1525 : node1516;
											assign node1516 = (inp[0]) ? 15'b000000011111111 : node1517;
												assign node1517 = (inp[10]) ? node1521 : node1518;
													assign node1518 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1521 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1525 = (inp[1]) ? node1535 : node1526;
												assign node1526 = (inp[11]) ? node1530 : node1527;
													assign node1527 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1530 = (inp[10]) ? node1532 : 15'b000000011111111;
														assign node1532 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1535 = (inp[14]) ? 15'b000000001111111 : node1536;
													assign node1536 = (inp[0]) ? 15'b000000001111111 : node1537;
														assign node1537 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1542 = (inp[1]) ? node1564 : node1543;
											assign node1543 = (inp[2]) ? node1553 : node1544;
												assign node1544 = (inp[0]) ? node1548 : node1545;
													assign node1545 = (inp[14]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node1548 = (inp[14]) ? node1550 : 15'b000000011111111;
														assign node1550 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1553 = (inp[14]) ? node1559 : node1554;
													assign node1554 = (inp[0]) ? 15'b000000001111111 : node1555;
														assign node1555 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1559 = (inp[10]) ? 15'b000000000111111 : node1560;
														assign node1560 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1564 = (inp[0]) ? node1578 : node1565;
												assign node1565 = (inp[11]) ? node1575 : node1566;
													assign node1566 = (inp[10]) ? node1570 : node1567;
														assign node1567 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node1570 = (inp[2]) ? node1572 : 15'b000000001111111;
															assign node1572 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node1575 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1578 = (inp[14]) ? node1584 : node1579;
													assign node1579 = (inp[2]) ? 15'b000000000111111 : node1580;
														assign node1580 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node1584 = (inp[11]) ? 15'b000000000001111 : node1585;
														assign node1585 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node1589 = (inp[10]) ? node1833 : node1590;
							assign node1590 = (inp[0]) ? node1720 : node1591;
								assign node1591 = (inp[5]) ? node1655 : node1592;
									assign node1592 = (inp[11]) ? node1630 : node1593;
										assign node1593 = (inp[13]) ? node1611 : node1594;
											assign node1594 = (inp[1]) ? node1602 : node1595;
												assign node1595 = (inp[3]) ? 15'b000011111111111 : node1596;
													assign node1596 = (inp[2]) ? 15'b000011111111111 : node1597;
														assign node1597 = (inp[14]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node1602 = (inp[6]) ? 15'b000001111111111 : node1603;
													assign node1603 = (inp[3]) ? node1605 : 15'b000011111111111;
														assign node1605 = (inp[14]) ? 15'b000001111111111 : node1606;
															assign node1606 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node1611 = (inp[3]) ? node1619 : node1612;
												assign node1612 = (inp[14]) ? node1616 : node1613;
													assign node1613 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1616 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1619 = (inp[1]) ? node1623 : node1620;
													assign node1620 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1623 = (inp[2]) ? 15'b000000011111111 : node1624;
														assign node1624 = (inp[14]) ? node1626 : 15'b000000111111111;
															assign node1626 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1630 = (inp[3]) ? node1644 : node1631;
											assign node1631 = (inp[6]) ? node1637 : node1632;
												assign node1632 = (inp[13]) ? node1634 : 15'b000001111111111;
													assign node1634 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1637 = (inp[2]) ? node1641 : node1638;
													assign node1638 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1641 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1644 = (inp[14]) ? 15'b000000011111111 : node1645;
												assign node1645 = (inp[13]) ? node1647 : 15'b000000111111111;
													assign node1647 = (inp[6]) ? node1649 : 15'b000000111111111;
														assign node1649 = (inp[1]) ? 15'b000000011111111 : node1650;
															assign node1650 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node1655 = (inp[1]) ? node1681 : node1656;
										assign node1656 = (inp[2]) ? node1670 : node1657;
											assign node1657 = (inp[3]) ? node1665 : node1658;
												assign node1658 = (inp[13]) ? 15'b000001111111111 : node1659;
													assign node1659 = (inp[14]) ? node1661 : 15'b000011111111111;
														assign node1661 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node1665 = (inp[13]) ? 15'b000000111111111 : node1666;
													assign node1666 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1670 = (inp[13]) ? node1676 : node1671;
												assign node1671 = (inp[11]) ? node1673 : 15'b000001111111111;
													assign node1673 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1676 = (inp[3]) ? 15'b000000001111111 : node1677;
													assign node1677 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node1681 = (inp[3]) ? node1699 : node1682;
											assign node1682 = (inp[14]) ? node1690 : node1683;
												assign node1683 = (inp[11]) ? node1687 : node1684;
													assign node1684 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1687 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1690 = (inp[13]) ? node1692 : 15'b000000111111111;
													assign node1692 = (inp[11]) ? 15'b000000000111111 : node1693;
														assign node1693 = (inp[6]) ? node1695 : 15'b000000011111111;
															assign node1695 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1699 = (inp[11]) ? node1711 : node1700;
												assign node1700 = (inp[2]) ? node1704 : node1701;
													assign node1701 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1704 = (inp[14]) ? 15'b000000001111111 : node1705;
														assign node1705 = (inp[6]) ? node1707 : 15'b000000011111111;
															assign node1707 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1711 = (inp[13]) ? 15'b000000001111111 : node1712;
													assign node1712 = (inp[6]) ? 15'b000000001111111 : node1713;
														assign node1713 = (inp[14]) ? node1715 : 15'b000000011111111;
															assign node1715 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node1720 = (inp[14]) ? node1778 : node1721;
									assign node1721 = (inp[5]) ? node1753 : node1722;
										assign node1722 = (inp[1]) ? node1740 : node1723;
											assign node1723 = (inp[13]) ? node1735 : node1724;
												assign node1724 = (inp[6]) ? node1732 : node1725;
													assign node1725 = (inp[3]) ? node1727 : 15'b000011111111111;
														assign node1727 = (inp[11]) ? 15'b000001111111111 : node1728;
															assign node1728 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node1732 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1735 = (inp[3]) ? 15'b000000011111111 : node1736;
													assign node1736 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node1740 = (inp[2]) ? node1750 : node1741;
												assign node1741 = (inp[11]) ? node1747 : node1742;
													assign node1742 = (inp[3]) ? 15'b000000111111111 : node1743;
														assign node1743 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node1747 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1750 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1753 = (inp[11]) ? node1763 : node1754;
											assign node1754 = (inp[13]) ? node1758 : node1755;
												assign node1755 = (inp[3]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node1758 = (inp[6]) ? 15'b000000011111111 : node1759;
													assign node1759 = (inp[3]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node1763 = (inp[1]) ? node1773 : node1764;
												assign node1764 = (inp[3]) ? node1768 : node1765;
													assign node1765 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1768 = (inp[13]) ? 15'b000000001111111 : node1769;
														assign node1769 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1773 = (inp[2]) ? node1775 : 15'b000000001111111;
													assign node1775 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1778 = (inp[2]) ? node1806 : node1779;
										assign node1779 = (inp[13]) ? node1793 : node1780;
											assign node1780 = (inp[11]) ? node1788 : node1781;
												assign node1781 = (inp[6]) ? 15'b000000011111111 : node1782;
													assign node1782 = (inp[3]) ? 15'b000000111111111 : node1783;
														assign node1783 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1788 = (inp[6]) ? 15'b000000011111111 : node1789;
													assign node1789 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1793 = (inp[5]) ? node1801 : node1794;
												assign node1794 = (inp[11]) ? node1798 : node1795;
													assign node1795 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1798 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1801 = (inp[3]) ? 15'b000000001111111 : node1802;
													assign node1802 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1806 = (inp[6]) ? node1816 : node1807;
											assign node1807 = (inp[3]) ? node1809 : 15'b000000011111111;
												assign node1809 = (inp[11]) ? node1811 : 15'b000000011111111;
													assign node1811 = (inp[5]) ? 15'b000000000011111 : node1812;
														assign node1812 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node1816 = (inp[11]) ? node1824 : node1817;
												assign node1817 = (inp[13]) ? node1819 : 15'b000000011111111;
													assign node1819 = (inp[3]) ? 15'b000000000111111 : node1820;
														assign node1820 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node1824 = (inp[1]) ? node1826 : 15'b000000000111111;
													assign node1826 = (inp[5]) ? 15'b000000000011111 : node1827;
														assign node1827 = (inp[3]) ? node1829 : 15'b000000001111111;
															assign node1829 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node1833 = (inp[2]) ? node1953 : node1834;
								assign node1834 = (inp[11]) ? node1898 : node1835;
									assign node1835 = (inp[13]) ? node1873 : node1836;
										assign node1836 = (inp[0]) ? node1852 : node1837;
											assign node1837 = (inp[6]) ? node1845 : node1838;
												assign node1838 = (inp[14]) ? 15'b000001111111111 : node1839;
													assign node1839 = (inp[3]) ? 15'b000011111111111 : node1840;
														assign node1840 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node1845 = (inp[5]) ? node1847 : 15'b000001111111111;
													assign node1847 = (inp[3]) ? 15'b000000011111111 : node1848;
														assign node1848 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1852 = (inp[1]) ? node1858 : node1853;
												assign node1853 = (inp[6]) ? 15'b000000111111111 : node1854;
													assign node1854 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1858 = (inp[5]) ? node1864 : node1859;
													assign node1859 = (inp[3]) ? node1861 : 15'b000000111111111;
														assign node1861 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1864 = (inp[6]) ? node1870 : node1865;
														assign node1865 = (inp[3]) ? 15'b000000011111111 : node1866;
															assign node1866 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node1870 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node1873 = (inp[3]) ? node1887 : node1874;
											assign node1874 = (inp[5]) ? node1882 : node1875;
												assign node1875 = (inp[6]) ? 15'b000001111111111 : node1876;
													assign node1876 = (inp[1]) ? node1878 : 15'b000000111111111;
														assign node1878 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node1882 = (inp[14]) ? 15'b000000011111111 : node1883;
													assign node1883 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1887 = (inp[5]) ? node1893 : node1888;
												assign node1888 = (inp[14]) ? node1890 : 15'b000000011111111;
													assign node1890 = (inp[0]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node1893 = (inp[14]) ? node1895 : 15'b000000001111111;
													assign node1895 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node1898 = (inp[14]) ? node1932 : node1899;
										assign node1899 = (inp[3]) ? node1915 : node1900;
											assign node1900 = (inp[1]) ? node1906 : node1901;
												assign node1901 = (inp[5]) ? 15'b000000011111111 : node1902;
													assign node1902 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1906 = (inp[13]) ? node1912 : node1907;
													assign node1907 = (inp[5]) ? node1909 : 15'b000000111111111;
														assign node1909 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1912 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1915 = (inp[0]) ? node1927 : node1916;
												assign node1916 = (inp[1]) ? node1920 : node1917;
													assign node1917 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node1920 = (inp[6]) ? 15'b000000001111111 : node1921;
														assign node1921 = (inp[5]) ? node1923 : 15'b000000011111111;
															assign node1923 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1927 = (inp[6]) ? node1929 : 15'b000000001111111;
													assign node1929 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
										assign node1932 = (inp[6]) ? node1944 : node1933;
											assign node1933 = (inp[13]) ? node1939 : node1934;
												assign node1934 = (inp[5]) ? 15'b000000011111111 : node1935;
													assign node1935 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1939 = (inp[0]) ? 15'b000000000111111 : node1940;
													assign node1940 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node1944 = (inp[3]) ? node1950 : node1945;
												assign node1945 = (inp[1]) ? 15'b000000000011111 : node1946;
													assign node1946 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node1950 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node1953 = (inp[6]) ? node2029 : node1954;
									assign node1954 = (inp[1]) ? node1988 : node1955;
										assign node1955 = (inp[5]) ? node1969 : node1956;
											assign node1956 = (inp[11]) ? node1962 : node1957;
												assign node1957 = (inp[3]) ? 15'b000000111111111 : node1958;
													assign node1958 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node1962 = (inp[13]) ? 15'b000000011111111 : node1963;
													assign node1963 = (inp[0]) ? node1965 : 15'b000000111111111;
														assign node1965 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node1969 = (inp[11]) ? node1979 : node1970;
												assign node1970 = (inp[14]) ? node1976 : node1971;
													assign node1971 = (inp[3]) ? node1973 : 15'b000000111111111;
														assign node1973 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node1976 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1979 = (inp[3]) ? node1983 : node1980;
													assign node1980 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node1983 = (inp[13]) ? node1985 : 15'b000000001111111;
														assign node1985 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node1988 = (inp[11]) ? node2008 : node1989;
											assign node1989 = (inp[0]) ? node1997 : node1990;
												assign node1990 = (inp[14]) ? node1992 : 15'b000000011111111;
													assign node1992 = (inp[5]) ? node1994 : 15'b000000011111111;
														assign node1994 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node1997 = (inp[3]) ? node2003 : node1998;
													assign node1998 = (inp[5]) ? node2000 : 15'b000000011111111;
														assign node2000 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2003 = (inp[14]) ? node2005 : 15'b000000001111111;
														assign node2005 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2008 = (inp[5]) ? node2018 : node2009;
												assign node2009 = (inp[13]) ? node2015 : node2010;
													assign node2010 = (inp[3]) ? 15'b000000001111111 : node2011;
														assign node2011 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2015 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2018 = (inp[13]) ? node2020 : 15'b000000000111111;
													assign node2020 = (inp[3]) ? node2026 : node2021;
														assign node2021 = (inp[0]) ? node2023 : 15'b000000000111111;
															assign node2023 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
														assign node2026 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node2029 = (inp[5]) ? node2057 : node2030;
										assign node2030 = (inp[14]) ? node2042 : node2031;
											assign node2031 = (inp[0]) ? node2037 : node2032;
												assign node2032 = (inp[13]) ? 15'b000000011111111 : node2033;
													assign node2033 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2037 = (inp[1]) ? node2039 : 15'b000000001111111;
													assign node2039 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2042 = (inp[0]) ? node2050 : node2043;
												assign node2043 = (inp[3]) ? node2045 : 15'b000000001111111;
													assign node2045 = (inp[11]) ? 15'b000000000111111 : node2046;
														assign node2046 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2050 = (inp[3]) ? 15'b000000000111111 : node2051;
													assign node2051 = (inp[11]) ? 15'b000000000111111 : node2052;
														assign node2052 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2057 = (inp[1]) ? node2079 : node2058;
											assign node2058 = (inp[3]) ? node2066 : node2059;
												assign node2059 = (inp[11]) ? node2061 : 15'b000000011111111;
													assign node2061 = (inp[13]) ? 15'b000000000111111 : node2062;
														assign node2062 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2066 = (inp[11]) ? node2072 : node2067;
													assign node2067 = (inp[13]) ? 15'b000000000111111 : node2068;
														assign node2068 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2072 = (inp[13]) ? 15'b000000000011111 : node2073;
														assign node2073 = (inp[14]) ? node2075 : 15'b000000000111111;
															assign node2075 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2079 = (inp[0]) ? node2087 : node2080;
												assign node2080 = (inp[14]) ? node2084 : node2081;
													assign node2081 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2084 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node2087 = (inp[14]) ? node2089 : 15'b000000000011111;
													assign node2089 = (inp[11]) ? node2095 : node2090;
														assign node2090 = (inp[3]) ? node2092 : 15'b000000000011111;
															assign node2092 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
														assign node2095 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
				assign node2098 = (inp[14]) ? node3138 : node2099;
					assign node2099 = (inp[2]) ? node2649 : node2100;
						assign node2100 = (inp[4]) ? node2372 : node2101;
							assign node2101 = (inp[5]) ? node2247 : node2102;
								assign node2102 = (inp[0]) ? node2172 : node2103;
									assign node2103 = (inp[6]) ? node2137 : node2104;
										assign node2104 = (inp[1]) ? node2122 : node2105;
											assign node2105 = (inp[10]) ? node2111 : node2106;
												assign node2106 = (inp[11]) ? node2108 : 15'b000111111111111;
													assign node2108 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node2111 = (inp[3]) ? node2117 : node2112;
													assign node2112 = (inp[11]) ? node2114 : 15'b000111111111111;
														assign node2114 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2117 = (inp[13]) ? node2119 : 15'b000011111111111;
														assign node2119 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2122 = (inp[9]) ? node2130 : node2123;
												assign node2123 = (inp[10]) ? node2127 : node2124;
													assign node2124 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node2127 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2130 = (inp[11]) ? 15'b000001111111111 : node2131;
													assign node2131 = (inp[10]) ? node2133 : 15'b000011111111111;
														assign node2133 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node2137 = (inp[1]) ? node2155 : node2138;
											assign node2138 = (inp[3]) ? node2146 : node2139;
												assign node2139 = (inp[13]) ? node2143 : node2140;
													assign node2140 = (inp[9]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node2143 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2146 = (inp[9]) ? node2150 : node2147;
													assign node2147 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2150 = (inp[10]) ? node2152 : 15'b000001111111111;
														assign node2152 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2155 = (inp[3]) ? node2163 : node2156;
												assign node2156 = (inp[10]) ? 15'b000000111111111 : node2157;
													assign node2157 = (inp[13]) ? 15'b000001111111111 : node2158;
														assign node2158 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2163 = (inp[11]) ? node2169 : node2164;
													assign node2164 = (inp[13]) ? 15'b000000111111111 : node2165;
														assign node2165 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2169 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2172 = (inp[10]) ? node2210 : node2173;
										assign node2173 = (inp[11]) ? node2191 : node2174;
											assign node2174 = (inp[1]) ? node2182 : node2175;
												assign node2175 = (inp[3]) ? 15'b000011111111111 : node2176;
													assign node2176 = (inp[6]) ? node2178 : 15'b000111111111111;
														assign node2178 = (inp[9]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node2182 = (inp[9]) ? node2188 : node2183;
													assign node2183 = (inp[3]) ? node2185 : 15'b000011111111111;
														assign node2185 = (inp[13]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node2188 = (inp[6]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node2191 = (inp[1]) ? node2203 : node2192;
												assign node2192 = (inp[13]) ? node2196 : node2193;
													assign node2193 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2196 = (inp[6]) ? 15'b000000111111111 : node2197;
														assign node2197 = (inp[3]) ? node2199 : 15'b000001111111111;
															assign node2199 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2203 = (inp[13]) ? 15'b000000011111111 : node2204;
													assign node2204 = (inp[9]) ? 15'b000000111111111 : node2205;
														assign node2205 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2210 = (inp[9]) ? node2228 : node2211;
											assign node2211 = (inp[3]) ? node2215 : node2212;
												assign node2212 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2215 = (inp[11]) ? node2223 : node2216;
													assign node2216 = (inp[6]) ? 15'b000000111111111 : node2217;
														assign node2217 = (inp[1]) ? node2219 : 15'b000001111111111;
															assign node2219 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2223 = (inp[6]) ? 15'b000000011111111 : node2224;
														assign node2224 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2228 = (inp[3]) ? node2238 : node2229;
												assign node2229 = (inp[13]) ? node2235 : node2230;
													assign node2230 = (inp[6]) ? node2232 : 15'b000001111111111;
														assign node2232 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2235 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2238 = (inp[11]) ? node2244 : node2239;
													assign node2239 = (inp[13]) ? 15'b000000011111111 : node2240;
														assign node2240 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2244 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2247 = (inp[9]) ? node2315 : node2248;
									assign node2248 = (inp[13]) ? node2286 : node2249;
										assign node2249 = (inp[11]) ? node2269 : node2250;
											assign node2250 = (inp[3]) ? node2254 : node2251;
												assign node2251 = (inp[10]) ? 15'b000011111111111 : 15'b001111111111111;
												assign node2254 = (inp[0]) ? node2264 : node2255;
													assign node2255 = (inp[1]) ? node2259 : node2256;
														assign node2256 = (inp[6]) ? 15'b000011111111111 : 15'b000111111111111;
														assign node2259 = (inp[10]) ? 15'b000001111111111 : node2260;
															assign node2260 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2264 = (inp[1]) ? node2266 : 15'b000001111111111;
														assign node2266 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2269 = (inp[3]) ? node2275 : node2270;
												assign node2270 = (inp[6]) ? 15'b000000111111111 : node2271;
													assign node2271 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2275 = (inp[1]) ? node2283 : node2276;
													assign node2276 = (inp[10]) ? 15'b000000111111111 : node2277;
														assign node2277 = (inp[0]) ? node2279 : 15'b000001111111111;
															assign node2279 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2283 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2286 = (inp[11]) ? node2300 : node2287;
											assign node2287 = (inp[3]) ? 15'b000000111111111 : node2288;
												assign node2288 = (inp[6]) ? node2290 : 15'b000001111111111;
													assign node2290 = (inp[1]) ? node2296 : node2291;
														assign node2291 = (inp[10]) ? node2293 : 15'b000001111111111;
															assign node2293 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node2296 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2300 = (inp[1]) ? node2308 : node2301;
												assign node2301 = (inp[0]) ? node2303 : 15'b000000111111111;
													assign node2303 = (inp[3]) ? node2305 : 15'b000000111111111;
														assign node2305 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2308 = (inp[0]) ? 15'b000000011111111 : node2309;
													assign node2309 = (inp[10]) ? 15'b000000011111111 : node2310;
														assign node2310 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node2315 = (inp[10]) ? node2351 : node2316;
										assign node2316 = (inp[13]) ? node2332 : node2317;
											assign node2317 = (inp[0]) ? node2325 : node2318;
												assign node2318 = (inp[1]) ? node2320 : 15'b000011111111111;
													assign node2320 = (inp[3]) ? 15'b000000111111111 : node2321;
														assign node2321 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2325 = (inp[11]) ? node2329 : node2326;
													assign node2326 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2329 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2332 = (inp[6]) ? node2340 : node2333;
												assign node2333 = (inp[11]) ? node2335 : 15'b000001111111111;
													assign node2335 = (inp[1]) ? 15'b000000111111111 : node2336;
														assign node2336 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2340 = (inp[11]) ? node2344 : node2341;
													assign node2341 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2344 = (inp[3]) ? node2348 : node2345;
														assign node2345 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node2348 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2351 = (inp[11]) ? node2359 : node2352;
											assign node2352 = (inp[6]) ? node2354 : 15'b000000111111111;
												assign node2354 = (inp[13]) ? 15'b000000001111111 : node2355;
													assign node2355 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2359 = (inp[0]) ? node2369 : node2360;
												assign node2360 = (inp[1]) ? node2362 : 15'b000000111111111;
													assign node2362 = (inp[3]) ? node2364 : 15'b000000011111111;
														assign node2364 = (inp[13]) ? 15'b000000001111111 : node2365;
															assign node2365 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2369 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node2372 = (inp[0]) ? node2500 : node2373;
								assign node2373 = (inp[11]) ? node2433 : node2374;
									assign node2374 = (inp[3]) ? node2394 : node2375;
										assign node2375 = (inp[6]) ? node2387 : node2376;
											assign node2376 = (inp[1]) ? node2380 : node2377;
												assign node2377 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node2380 = (inp[9]) ? node2384 : node2381;
													assign node2381 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2384 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2387 = (inp[1]) ? node2389 : 15'b000001111111111;
												assign node2389 = (inp[10]) ? 15'b000000111111111 : node2390;
													assign node2390 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2394 = (inp[1]) ? node2416 : node2395;
											assign node2395 = (inp[13]) ? node2407 : node2396;
												assign node2396 = (inp[5]) ? node2402 : node2397;
													assign node2397 = (inp[6]) ? 15'b000001111111111 : node2398;
														assign node2398 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node2402 = (inp[9]) ? node2404 : 15'b000001111111111;
														assign node2404 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2407 = (inp[10]) ? 15'b000000011111111 : node2408;
													assign node2408 = (inp[5]) ? 15'b000000111111111 : node2409;
														assign node2409 = (inp[6]) ? node2411 : 15'b000001111111111;
															assign node2411 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2416 = (inp[6]) ? node2422 : node2417;
												assign node2417 = (inp[9]) ? node2419 : 15'b000001111111111;
													assign node2419 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2422 = (inp[13]) ? node2426 : node2423;
													assign node2423 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2426 = (inp[5]) ? 15'b000000001111111 : node2427;
														assign node2427 = (inp[9]) ? node2429 : 15'b000000011111111;
															assign node2429 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node2433 = (inp[9]) ? node2465 : node2434;
										assign node2434 = (inp[6]) ? node2452 : node2435;
											assign node2435 = (inp[3]) ? node2445 : node2436;
												assign node2436 = (inp[10]) ? 15'b000001111111111 : node2437;
													assign node2437 = (inp[1]) ? 15'b000001111111111 : node2438;
														assign node2438 = (inp[5]) ? node2440 : 15'b000011111111111;
															assign node2440 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2445 = (inp[13]) ? 15'b000000011111111 : node2446;
													assign node2446 = (inp[5]) ? 15'b000000111111111 : node2447;
														assign node2447 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2452 = (inp[10]) ? node2458 : node2453;
												assign node2453 = (inp[1]) ? node2455 : 15'b000001111111111;
													assign node2455 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2458 = (inp[3]) ? node2462 : node2459;
													assign node2459 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2462 = (inp[1]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node2465 = (inp[10]) ? node2483 : node2466;
											assign node2466 = (inp[3]) ? node2474 : node2467;
												assign node2467 = (inp[13]) ? node2469 : 15'b000000111111111;
													assign node2469 = (inp[6]) ? 15'b000000111111111 : node2470;
														assign node2470 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2474 = (inp[13]) ? node2478 : node2475;
													assign node2475 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2478 = (inp[1]) ? node2480 : 15'b000000011111111;
														assign node2480 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node2483 = (inp[3]) ? node2493 : node2484;
												assign node2484 = (inp[1]) ? node2488 : node2485;
													assign node2485 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2488 = (inp[5]) ? node2490 : 15'b000000011111111;
														assign node2490 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2493 = (inp[5]) ? 15'b000000001111111 : node2494;
													assign node2494 = (inp[6]) ? 15'b000000001111111 : node2495;
														assign node2495 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node2500 = (inp[6]) ? node2574 : node2501;
									assign node2501 = (inp[5]) ? node2533 : node2502;
										assign node2502 = (inp[10]) ? node2520 : node2503;
											assign node2503 = (inp[9]) ? node2511 : node2504;
												assign node2504 = (inp[1]) ? node2506 : 15'b000001111111111;
													assign node2506 = (inp[13]) ? 15'b000001111111111 : node2507;
														assign node2507 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2511 = (inp[11]) ? node2513 : 15'b000001111111111;
													assign node2513 = (inp[1]) ? 15'b000000111111111 : node2514;
														assign node2514 = (inp[13]) ? 15'b000000111111111 : node2515;
															assign node2515 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node2520 = (inp[11]) ? node2528 : node2521;
												assign node2521 = (inp[1]) ? 15'b000000111111111 : node2522;
													assign node2522 = (inp[13]) ? 15'b000000111111111 : node2523;
														assign node2523 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2528 = (inp[1]) ? 15'b000000011111111 : node2529;
													assign node2529 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2533 = (inp[3]) ? node2553 : node2534;
											assign node2534 = (inp[1]) ? node2542 : node2535;
												assign node2535 = (inp[11]) ? 15'b000000111111111 : node2536;
													assign node2536 = (inp[13]) ? node2538 : 15'b000001111111111;
														assign node2538 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2542 = (inp[10]) ? node2550 : node2543;
													assign node2543 = (inp[9]) ? 15'b000000011111111 : node2544;
														assign node2544 = (inp[13]) ? node2546 : 15'b000000111111111;
															assign node2546 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2550 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2553 = (inp[11]) ? node2567 : node2554;
												assign node2554 = (inp[1]) ? node2560 : node2555;
													assign node2555 = (inp[13]) ? 15'b000000011111111 : node2556;
														assign node2556 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2560 = (inp[9]) ? 15'b000000001111111 : node2561;
														assign node2561 = (inp[13]) ? node2563 : 15'b000000011111111;
															assign node2563 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2567 = (inp[10]) ? node2571 : node2568;
													assign node2568 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2571 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2574 = (inp[5]) ? node2614 : node2575;
										assign node2575 = (inp[10]) ? node2593 : node2576;
											assign node2576 = (inp[3]) ? node2584 : node2577;
												assign node2577 = (inp[11]) ? node2581 : node2578;
													assign node2578 = (inp[1]) ? 15'b000001111111111 : 15'b000000111111111;
													assign node2581 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2584 = (inp[13]) ? 15'b000000011111111 : node2585;
													assign node2585 = (inp[9]) ? 15'b000000011111111 : node2586;
														assign node2586 = (inp[11]) ? node2588 : 15'b000000111111111;
															assign node2588 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2593 = (inp[1]) ? node2605 : node2594;
												assign node2594 = (inp[11]) ? node2598 : node2595;
													assign node2595 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2598 = (inp[3]) ? node2600 : 15'b000000011111111;
														assign node2600 = (inp[13]) ? 15'b000000001111111 : node2601;
															assign node2601 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2605 = (inp[9]) ? node2609 : node2606;
													assign node2606 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2609 = (inp[3]) ? node2611 : 15'b000000000111111;
														assign node2611 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node2614 = (inp[10]) ? node2636 : node2615;
											assign node2615 = (inp[1]) ? node2625 : node2616;
												assign node2616 = (inp[13]) ? node2618 : 15'b000000011111111;
													assign node2618 = (inp[9]) ? 15'b000000001111111 : node2619;
														assign node2619 = (inp[3]) ? 15'b000000001111111 : node2620;
															assign node2620 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2625 = (inp[9]) ? node2629 : node2626;
													assign node2626 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2629 = (inp[13]) ? node2631 : 15'b000000001111111;
														assign node2631 = (inp[3]) ? node2633 : 15'b000000000111111;
															assign node2633 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node2636 = (inp[11]) ? node2638 : 15'b000000001111111;
												assign node2638 = (inp[3]) ? node2646 : node2639;
													assign node2639 = (inp[9]) ? node2641 : 15'b000000001111111;
														assign node2641 = (inp[13]) ? 15'b000000000111111 : node2642;
															assign node2642 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2646 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node2649 = (inp[10]) ? node2897 : node2650;
							assign node2650 = (inp[3]) ? node2776 : node2651;
								assign node2651 = (inp[9]) ? node2703 : node2652;
									assign node2652 = (inp[6]) ? node2680 : node2653;
										assign node2653 = (inp[4]) ? node2667 : node2654;
											assign node2654 = (inp[5]) ? node2662 : node2655;
												assign node2655 = (inp[11]) ? node2659 : node2656;
													assign node2656 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node2659 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2662 = (inp[13]) ? 15'b000001111111111 : node2663;
													assign node2663 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node2667 = (inp[11]) ? node2673 : node2668;
												assign node2668 = (inp[13]) ? node2670 : 15'b000011111111111;
													assign node2670 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2673 = (inp[0]) ? 15'b000000111111111 : node2674;
													assign node2674 = (inp[1]) ? 15'b000000111111111 : node2675;
														assign node2675 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node2680 = (inp[0]) ? node2692 : node2681;
											assign node2681 = (inp[11]) ? node2687 : node2682;
												assign node2682 = (inp[5]) ? 15'b000000111111111 : node2683;
													assign node2683 = (inp[13]) ? 15'b000001111111111 : 15'b000111111111111;
												assign node2687 = (inp[13]) ? node2689 : 15'b000000111111111;
													assign node2689 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2692 = (inp[4]) ? node2698 : node2693;
												assign node2693 = (inp[5]) ? node2695 : 15'b000000111111111;
													assign node2695 = (inp[1]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node2698 = (inp[1]) ? 15'b000000011111111 : node2699;
													assign node2699 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node2703 = (inp[13]) ? node2747 : node2704;
										assign node2704 = (inp[11]) ? node2726 : node2705;
											assign node2705 = (inp[6]) ? node2719 : node2706;
												assign node2706 = (inp[4]) ? node2712 : node2707;
													assign node2707 = (inp[1]) ? node2709 : 15'b000001111111111;
														assign node2709 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2712 = (inp[5]) ? 15'b000000111111111 : node2713;
														assign node2713 = (inp[1]) ? node2715 : 15'b000001111111111;
															assign node2715 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node2719 = (inp[4]) ? node2723 : node2720;
													assign node2720 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2723 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2726 = (inp[4]) ? node2736 : node2727;
												assign node2727 = (inp[0]) ? node2733 : node2728;
													assign node2728 = (inp[6]) ? 15'b000000111111111 : node2729;
														assign node2729 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2733 = (inp[6]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node2736 = (inp[1]) ? node2738 : 15'b000000111111111;
													assign node2738 = (inp[6]) ? node2742 : node2739;
														assign node2739 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node2742 = (inp[5]) ? 15'b000000001111111 : node2743;
															assign node2743 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2747 = (inp[0]) ? node2759 : node2748;
											assign node2748 = (inp[5]) ? 15'b000000011111111 : node2749;
												assign node2749 = (inp[6]) ? node2753 : node2750;
													assign node2750 = (inp[4]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node2753 = (inp[1]) ? node2755 : 15'b000000111111111;
														assign node2755 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2759 = (inp[6]) ? node2773 : node2760;
												assign node2760 = (inp[1]) ? node2766 : node2761;
													assign node2761 = (inp[4]) ? 15'b000000011111111 : node2762;
														assign node2762 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2766 = (inp[4]) ? 15'b000000000111111 : node2767;
														assign node2767 = (inp[5]) ? node2769 : 15'b000000011111111;
															assign node2769 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2773 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node2776 = (inp[1]) ? node2836 : node2777;
									assign node2777 = (inp[13]) ? node2807 : node2778;
										assign node2778 = (inp[4]) ? node2792 : node2779;
											assign node2779 = (inp[5]) ? node2787 : node2780;
												assign node2780 = (inp[0]) ? 15'b000000111111111 : node2781;
													assign node2781 = (inp[9]) ? 15'b000001111111111 : node2782;
														assign node2782 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2787 = (inp[6]) ? node2789 : 15'b000000111111111;
													assign node2789 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2792 = (inp[6]) ? node2794 : 15'b000000111111111;
												assign node2794 = (inp[5]) ? node2802 : node2795;
													assign node2795 = (inp[0]) ? node2797 : 15'b000001111111111;
														assign node2797 = (inp[11]) ? 15'b000000011111111 : node2798;
															assign node2798 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2802 = (inp[11]) ? node2804 : 15'b000000011111111;
														assign node2804 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2807 = (inp[11]) ? node2823 : node2808;
											assign node2808 = (inp[9]) ? node2814 : node2809;
												assign node2809 = (inp[5]) ? 15'b000000111111111 : node2810;
													assign node2810 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2814 = (inp[6]) ? node2818 : node2815;
													assign node2815 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2818 = (inp[5]) ? node2820 : 15'b000000011111111;
														assign node2820 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2823 = (inp[5]) ? node2827 : node2824;
												assign node2824 = (inp[9]) ? 15'b000000011111111 : 15'b000000001111111;
												assign node2827 = (inp[9]) ? node2829 : 15'b000000011111111;
													assign node2829 = (inp[4]) ? node2831 : 15'b000000001111111;
														assign node2831 = (inp[0]) ? 15'b000000000111111 : node2832;
															assign node2832 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2836 = (inp[9]) ? node2874 : node2837;
										assign node2837 = (inp[0]) ? node2857 : node2838;
											assign node2838 = (inp[6]) ? node2848 : node2839;
												assign node2839 = (inp[11]) ? node2841 : 15'b000011111111111;
													assign node2841 = (inp[5]) ? node2843 : 15'b000000111111111;
														assign node2843 = (inp[4]) ? 15'b000000011111111 : node2844;
															assign node2844 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2848 = (inp[5]) ? node2852 : node2849;
													assign node2849 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2852 = (inp[13]) ? 15'b000000011111111 : node2853;
														assign node2853 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2857 = (inp[11]) ? node2867 : node2858;
												assign node2858 = (inp[4]) ? node2862 : node2859;
													assign node2859 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2862 = (inp[13]) ? node2864 : 15'b000000011111111;
														assign node2864 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2867 = (inp[13]) ? node2871 : node2868;
													assign node2868 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node2871 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node2874 = (inp[0]) ? node2882 : node2875;
											assign node2875 = (inp[5]) ? node2877 : 15'b000000011111111;
												assign node2877 = (inp[13]) ? 15'b000000000111111 : node2878;
													assign node2878 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2882 = (inp[4]) ? node2890 : node2883;
												assign node2883 = (inp[6]) ? node2885 : 15'b000000011111111;
													assign node2885 = (inp[5]) ? 15'b000000000111111 : node2886;
														assign node2886 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node2890 = (inp[11]) ? node2894 : node2891;
													assign node2891 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node2894 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node2897 = (inp[0]) ? node3017 : node2898;
								assign node2898 = (inp[6]) ? node2954 : node2899;
									assign node2899 = (inp[1]) ? node2921 : node2900;
										assign node2900 = (inp[3]) ? node2914 : node2901;
											assign node2901 = (inp[13]) ? node2907 : node2902;
												assign node2902 = (inp[9]) ? 15'b000001111111111 : node2903;
													assign node2903 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node2907 = (inp[5]) ? node2911 : node2908;
													assign node2908 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2911 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node2914 = (inp[11]) ? node2916 : 15'b000000111111111;
												assign node2916 = (inp[13]) ? 15'b000000011111111 : node2917;
													assign node2917 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node2921 = (inp[9]) ? node2941 : node2922;
											assign node2922 = (inp[4]) ? node2934 : node2923;
												assign node2923 = (inp[5]) ? node2927 : node2924;
													assign node2924 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node2927 = (inp[3]) ? node2929 : 15'b000000111111111;
														assign node2929 = (inp[11]) ? 15'b000000011111111 : node2930;
															assign node2930 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2934 = (inp[5]) ? node2938 : node2935;
													assign node2935 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node2938 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2941 = (inp[11]) ? node2949 : node2942;
												assign node2942 = (inp[3]) ? node2944 : 15'b000000011111111;
													assign node2944 = (inp[13]) ? 15'b000000001111111 : node2945;
														assign node2945 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2949 = (inp[3]) ? node2951 : 15'b000000001111111;
													assign node2951 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node2954 = (inp[13]) ? node2988 : node2955;
										assign node2955 = (inp[4]) ? node2969 : node2956;
											assign node2956 = (inp[5]) ? node2964 : node2957;
												assign node2957 = (inp[3]) ? node2959 : 15'b000001111111111;
													assign node2959 = (inp[9]) ? 15'b000000011111111 : node2960;
														assign node2960 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node2964 = (inp[1]) ? 15'b000000011111111 : node2965;
													assign node2965 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node2969 = (inp[3]) ? node2979 : node2970;
												assign node2970 = (inp[5]) ? 15'b000000111111111 : node2971;
													assign node2971 = (inp[1]) ? node2973 : 15'b000000011111111;
														assign node2973 = (inp[11]) ? node2975 : 15'b000000011111111;
															assign node2975 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node2979 = (inp[11]) ? 15'b000000001111111 : node2980;
													assign node2980 = (inp[9]) ? node2982 : 15'b000000011111111;
														assign node2982 = (inp[1]) ? 15'b000000001111111 : node2983;
															assign node2983 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node2988 = (inp[11]) ? node3008 : node2989;
											assign node2989 = (inp[5]) ? node3001 : node2990;
												assign node2990 = (inp[4]) ? node2992 : 15'b000000011111111;
													assign node2992 = (inp[1]) ? node2998 : node2993;
														assign node2993 = (inp[9]) ? node2995 : 15'b000000011111111;
															assign node2995 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node2998 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3001 = (inp[9]) ? 15'b000000001111111 : node3002;
													assign node3002 = (inp[4]) ? 15'b000000001111111 : node3003;
														assign node3003 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3008 = (inp[3]) ? node3010 : 15'b000000001111111;
												assign node3010 = (inp[1]) ? 15'b000000000011111 : node3011;
													assign node3011 = (inp[4]) ? 15'b000000000111111 : node3012;
														assign node3012 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node3017 = (inp[4]) ? node3067 : node3018;
									assign node3018 = (inp[13]) ? node3040 : node3019;
										assign node3019 = (inp[1]) ? node3027 : node3020;
											assign node3020 = (inp[11]) ? node3024 : node3021;
												assign node3021 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3024 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3027 = (inp[3]) ? 15'b000000001111111 : node3028;
												assign node3028 = (inp[11]) ? node3034 : node3029;
													assign node3029 = (inp[5]) ? 15'b000000011111111 : node3030;
														assign node3030 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3034 = (inp[5]) ? node3036 : 15'b000000011111111;
														assign node3036 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3040 = (inp[1]) ? node3058 : node3041;
											assign node3041 = (inp[6]) ? node3053 : node3042;
												assign node3042 = (inp[3]) ? node3046 : node3043;
													assign node3043 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3046 = (inp[11]) ? node3048 : 15'b000000111111111;
														assign node3048 = (inp[5]) ? 15'b000000001111111 : node3049;
															assign node3049 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3053 = (inp[11]) ? 15'b000000001111111 : node3054;
													assign node3054 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3058 = (inp[6]) ? node3060 : 15'b000000001111111;
												assign node3060 = (inp[3]) ? node3064 : node3061;
													assign node3061 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3064 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3067 = (inp[13]) ? node3101 : node3068;
										assign node3068 = (inp[5]) ? node3084 : node3069;
											assign node3069 = (inp[1]) ? node3075 : node3070;
												assign node3070 = (inp[9]) ? 15'b000000001111111 : node3071;
													assign node3071 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3075 = (inp[11]) ? node3077 : 15'b000000011111111;
													assign node3077 = (inp[3]) ? 15'b000000001111111 : node3078;
														assign node3078 = (inp[9]) ? 15'b000000001111111 : node3079;
															assign node3079 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3084 = (inp[11]) ? node3094 : node3085;
												assign node3085 = (inp[1]) ? node3087 : 15'b000000011111111;
													assign node3087 = (inp[3]) ? 15'b000000000111111 : node3088;
														assign node3088 = (inp[9]) ? 15'b000000001111111 : node3089;
															assign node3089 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3094 = (inp[1]) ? node3098 : node3095;
													assign node3095 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3098 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node3101 = (inp[3]) ? node3127 : node3102;
											assign node3102 = (inp[5]) ? node3110 : node3103;
												assign node3103 = (inp[11]) ? node3107 : node3104;
													assign node3104 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3107 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3110 = (inp[9]) ? node3120 : node3111;
													assign node3111 = (inp[1]) ? node3115 : node3112;
														assign node3112 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
														assign node3115 = (inp[11]) ? node3117 : 15'b000000000111111;
															assign node3117 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3120 = (inp[6]) ? node3122 : 15'b000000000111111;
														assign node3122 = (inp[1]) ? node3124 : 15'b000000000011111;
															assign node3124 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node3127 = (inp[6]) ? node3131 : node3128;
												assign node3128 = (inp[1]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node3131 = (inp[9]) ? node3133 : 15'b000000000011111;
													assign node3133 = (inp[5]) ? node3135 : 15'b000000000011111;
														assign node3135 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node3138 = (inp[9]) ? node3644 : node3139;
						assign node3139 = (inp[1]) ? node3367 : node3140;
							assign node3140 = (inp[11]) ? node3260 : node3141;
								assign node3141 = (inp[3]) ? node3197 : node3142;
									assign node3142 = (inp[5]) ? node3174 : node3143;
										assign node3143 = (inp[0]) ? node3163 : node3144;
											assign node3144 = (inp[2]) ? node3152 : node3145;
												assign node3145 = (inp[4]) ? 15'b000111111111111 : node3146;
													assign node3146 = (inp[10]) ? 15'b000111111111111 : node3147;
														assign node3147 = (inp[13]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node3152 = (inp[10]) ? node3158 : node3153;
													assign node3153 = (inp[13]) ? 15'b000011111111111 : node3154;
														assign node3154 = (inp[6]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node3158 = (inp[4]) ? 15'b000001111111111 : node3159;
														assign node3159 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node3163 = (inp[2]) ? node3169 : node3164;
												assign node3164 = (inp[10]) ? 15'b000001111111111 : node3165;
													assign node3165 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3169 = (inp[6]) ? 15'b000000011111111 : node3170;
													assign node3170 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node3174 = (inp[13]) ? node3184 : node3175;
											assign node3175 = (inp[6]) ? node3181 : node3176;
												assign node3176 = (inp[2]) ? node3178 : 15'b000001111111111;
													assign node3178 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3181 = (inp[2]) ? 15'b000001111111111 : 15'b000000111111111;
											assign node3184 = (inp[6]) ? node3190 : node3185;
												assign node3185 = (inp[0]) ? node3187 : 15'b000000111111111;
													assign node3187 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3190 = (inp[10]) ? node3194 : node3191;
													assign node3191 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3194 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node3197 = (inp[10]) ? node3223 : node3198;
										assign node3198 = (inp[13]) ? node3208 : node3199;
											assign node3199 = (inp[0]) ? node3205 : node3200;
												assign node3200 = (inp[4]) ? 15'b000001111111111 : node3201;
													assign node3201 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3205 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3208 = (inp[5]) ? node3216 : node3209;
												assign node3209 = (inp[6]) ? 15'b000000111111111 : node3210;
													assign node3210 = (inp[4]) ? 15'b000000111111111 : node3211;
														assign node3211 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3216 = (inp[6]) ? 15'b000000011111111 : node3217;
													assign node3217 = (inp[0]) ? node3219 : 15'b000000111111111;
														assign node3219 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3223 = (inp[6]) ? node3247 : node3224;
											assign node3224 = (inp[13]) ? node3236 : node3225;
												assign node3225 = (inp[5]) ? node3231 : node3226;
													assign node3226 = (inp[0]) ? node3228 : 15'b000001111111111;
														assign node3228 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3231 = (inp[2]) ? node3233 : 15'b000000111111111;
														assign node3233 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3236 = (inp[0]) ? node3244 : node3237;
													assign node3237 = (inp[4]) ? node3239 : 15'b000000111111111;
														assign node3239 = (inp[2]) ? 15'b000000011111111 : node3240;
															assign node3240 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3244 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3247 = (inp[5]) ? node3255 : node3248;
												assign node3248 = (inp[2]) ? node3250 : 15'b000000011111111;
													assign node3250 = (inp[4]) ? 15'b000000011111111 : node3251;
														assign node3251 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3255 = (inp[2]) ? node3257 : 15'b000000011111111;
													assign node3257 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node3260 = (inp[4]) ? node3310 : node3261;
									assign node3261 = (inp[3]) ? node3287 : node3262;
										assign node3262 = (inp[5]) ? node3274 : node3263;
											assign node3263 = (inp[10]) ? node3269 : node3264;
												assign node3264 = (inp[13]) ? 15'b000001111111111 : node3265;
													assign node3265 = (inp[6]) ? 15'b000001111111111 : 15'b000111111111111;
												assign node3269 = (inp[2]) ? node3271 : 15'b000000111111111;
													assign node3271 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3274 = (inp[2]) ? 15'b000000011111111 : node3275;
												assign node3275 = (inp[6]) ? node3279 : node3276;
													assign node3276 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3279 = (inp[0]) ? node3281 : 15'b000000111111111;
														assign node3281 = (inp[13]) ? 15'b000000011111111 : node3282;
															assign node3282 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3287 = (inp[5]) ? node3301 : node3288;
											assign node3288 = (inp[6]) ? node3294 : node3289;
												assign node3289 = (inp[10]) ? node3291 : 15'b000000111111111;
													assign node3291 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3294 = (inp[0]) ? node3296 : 15'b000000001111111;
													assign node3296 = (inp[10]) ? 15'b000000011111111 : node3297;
														assign node3297 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3301 = (inp[0]) ? 15'b000000001111111 : node3302;
												assign node3302 = (inp[10]) ? 15'b000000011111111 : node3303;
													assign node3303 = (inp[13]) ? node3305 : 15'b000000111111111;
														assign node3305 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node3310 = (inp[2]) ? node3340 : node3311;
										assign node3311 = (inp[10]) ? node3325 : node3312;
											assign node3312 = (inp[3]) ? node3320 : node3313;
												assign node3313 = (inp[5]) ? node3317 : node3314;
													assign node3314 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3317 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3320 = (inp[13]) ? 15'b000000001111111 : node3321;
													assign node3321 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3325 = (inp[6]) ? node3335 : node3326;
												assign node3326 = (inp[3]) ? node3328 : 15'b000000011111111;
													assign node3328 = (inp[0]) ? node3330 : 15'b000000011111111;
														assign node3330 = (inp[5]) ? 15'b000000001111111 : node3331;
															assign node3331 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3335 = (inp[0]) ? 15'b000000001111111 : node3336;
													assign node3336 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3340 = (inp[0]) ? node3348 : node3341;
											assign node3341 = (inp[13]) ? 15'b000000001111111 : node3342;
												assign node3342 = (inp[5]) ? node3344 : 15'b000000001111111;
													assign node3344 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3348 = (inp[3]) ? node3356 : node3349;
												assign node3349 = (inp[13]) ? 15'b000000000111111 : node3350;
													assign node3350 = (inp[6]) ? 15'b000000001111111 : node3351;
														assign node3351 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3356 = (inp[6]) ? node3362 : node3357;
													assign node3357 = (inp[10]) ? 15'b000000000111111 : node3358;
														assign node3358 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3362 = (inp[13]) ? 15'b000000000011111 : node3363;
														assign node3363 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node3367 = (inp[0]) ? node3511 : node3368;
								assign node3368 = (inp[2]) ? node3450 : node3369;
									assign node3369 = (inp[6]) ? node3407 : node3370;
										assign node3370 = (inp[10]) ? node3384 : node3371;
											assign node3371 = (inp[11]) ? node3377 : node3372;
												assign node3372 = (inp[13]) ? 15'b000000111111111 : node3373;
													assign node3373 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3377 = (inp[3]) ? node3379 : 15'b000000111111111;
													assign node3379 = (inp[4]) ? 15'b000000111111111 : node3380;
														assign node3380 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3384 = (inp[4]) ? node3398 : node3385;
												assign node3385 = (inp[3]) ? node3393 : node3386;
													assign node3386 = (inp[13]) ? node3388 : 15'b000001111111111;
														assign node3388 = (inp[5]) ? 15'b000000011111111 : node3389;
															assign node3389 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3393 = (inp[5]) ? node3395 : 15'b000000111111111;
														assign node3395 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3398 = (inp[3]) ? node3402 : node3399;
													assign node3399 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3402 = (inp[5]) ? node3404 : 15'b000000011111111;
														assign node3404 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3407 = (inp[5]) ? node3427 : node3408;
											assign node3408 = (inp[11]) ? node3420 : node3409;
												assign node3409 = (inp[3]) ? node3413 : node3410;
													assign node3410 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3413 = (inp[4]) ? 15'b000000011111111 : node3414;
														assign node3414 = (inp[13]) ? node3416 : 15'b000000111111111;
															assign node3416 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3420 = (inp[4]) ? node3424 : node3421;
													assign node3421 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node3424 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3427 = (inp[11]) ? node3441 : node3428;
												assign node3428 = (inp[3]) ? node3436 : node3429;
													assign node3429 = (inp[4]) ? node3431 : 15'b000000111111111;
														assign node3431 = (inp[10]) ? 15'b000000011111111 : node3432;
															assign node3432 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3436 = (inp[10]) ? node3438 : 15'b000000011111111;
														assign node3438 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3441 = (inp[13]) ? 15'b000000000111111 : node3442;
													assign node3442 = (inp[3]) ? node3444 : 15'b000000011111111;
														assign node3444 = (inp[10]) ? node3446 : 15'b000000001111111;
															assign node3446 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3450 = (inp[5]) ? node3480 : node3451;
										assign node3451 = (inp[11]) ? node3465 : node3452;
											assign node3452 = (inp[10]) ? node3458 : node3453;
												assign node3453 = (inp[3]) ? node3455 : 15'b000000111111111;
													assign node3455 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3458 = (inp[13]) ? 15'b000000011111111 : node3459;
													assign node3459 = (inp[3]) ? 15'b000000011111111 : node3460;
														assign node3460 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3465 = (inp[10]) ? node3473 : node3466;
												assign node3466 = (inp[3]) ? node3470 : node3467;
													assign node3467 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3470 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3473 = (inp[6]) ? node3477 : node3474;
													assign node3474 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3477 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3480 = (inp[11]) ? node3502 : node3481;
											assign node3481 = (inp[6]) ? node3491 : node3482;
												assign node3482 = (inp[4]) ? node3484 : 15'b000000011111111;
													assign node3484 = (inp[10]) ? node3486 : 15'b000000011111111;
														assign node3486 = (inp[3]) ? 15'b000000001111111 : node3487;
															assign node3487 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3491 = (inp[10]) ? node3497 : node3492;
													assign node3492 = (inp[3]) ? 15'b000000001111111 : node3493;
														assign node3493 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3497 = (inp[13]) ? node3499 : 15'b000000001111111;
														assign node3499 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3502 = (inp[4]) ? node3508 : node3503;
												assign node3503 = (inp[6]) ? 15'b000000001111111 : node3504;
													assign node3504 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3508 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3511 = (inp[3]) ? node3571 : node3512;
									assign node3512 = (inp[2]) ? node3544 : node3513;
										assign node3513 = (inp[11]) ? node3531 : node3514;
											assign node3514 = (inp[13]) ? node3524 : node3515;
												assign node3515 = (inp[10]) ? node3521 : node3516;
													assign node3516 = (inp[4]) ? 15'b000000111111111 : node3517;
														assign node3517 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3521 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3524 = (inp[6]) ? node3526 : 15'b000000011111111;
													assign node3526 = (inp[10]) ? node3528 : 15'b000000011111111;
														assign node3528 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3531 = (inp[5]) ? node3535 : node3532;
												assign node3532 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3535 = (inp[6]) ? 15'b000000001111111 : node3536;
													assign node3536 = (inp[13]) ? 15'b000000001111111 : node3537;
														assign node3537 = (inp[10]) ? node3539 : 15'b000000011111111;
															assign node3539 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3544 = (inp[13]) ? node3558 : node3545;
											assign node3545 = (inp[6]) ? node3549 : node3546;
												assign node3546 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3549 = (inp[10]) ? node3553 : node3550;
													assign node3550 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3553 = (inp[11]) ? node3555 : 15'b000000001111111;
														assign node3555 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3558 = (inp[10]) ? node3564 : node3559;
												assign node3559 = (inp[5]) ? 15'b000000000111111 : node3560;
													assign node3560 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3564 = (inp[4]) ? node3566 : 15'b000000000111111;
													assign node3566 = (inp[5]) ? 15'b000000000011111 : node3567;
														assign node3567 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3571 = (inp[5]) ? node3611 : node3572;
										assign node3572 = (inp[6]) ? node3590 : node3573;
											assign node3573 = (inp[10]) ? node3577 : node3574;
												assign node3574 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3577 = (inp[4]) ? node3583 : node3578;
													assign node3578 = (inp[2]) ? node3580 : 15'b000000011111111;
														assign node3580 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3583 = (inp[2]) ? 15'b000000001111111 : node3584;
														assign node3584 = (inp[11]) ? 15'b000000001111111 : node3585;
															assign node3585 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3590 = (inp[10]) ? node3598 : node3591;
												assign node3591 = (inp[4]) ? node3595 : node3592;
													assign node3592 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3595 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3598 = (inp[13]) ? node3604 : node3599;
													assign node3599 = (inp[2]) ? node3601 : 15'b000000001111111;
														assign node3601 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node3604 = (inp[2]) ? node3608 : node3605;
														assign node3605 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
														assign node3608 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node3611 = (inp[4]) ? node3633 : node3612;
											assign node3612 = (inp[2]) ? node3624 : node3613;
												assign node3613 = (inp[10]) ? node3617 : node3614;
													assign node3614 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3617 = (inp[13]) ? 15'b000000000111111 : node3618;
														assign node3618 = (inp[11]) ? node3620 : 15'b000000001111111;
															assign node3620 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3624 = (inp[13]) ? node3630 : node3625;
													assign node3625 = (inp[10]) ? 15'b000000000111111 : node3626;
														assign node3626 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3630 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node3633 = (inp[6]) ? node3639 : node3634;
												assign node3634 = (inp[11]) ? node3636 : 15'b000000000111111;
													assign node3636 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node3639 = (inp[10]) ? 15'b000000000001111 : node3640;
													assign node3640 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node3644 = (inp[4]) ? node3890 : node3645;
							assign node3645 = (inp[11]) ? node3769 : node3646;
								assign node3646 = (inp[10]) ? node3708 : node3647;
									assign node3647 = (inp[13]) ? node3669 : node3648;
										assign node3648 = (inp[1]) ? node3662 : node3649;
											assign node3649 = (inp[3]) ? node3653 : node3650;
												assign node3650 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node3653 = (inp[5]) ? 15'b000000011111111 : node3654;
													assign node3654 = (inp[6]) ? 15'b000000111111111 : node3655;
														assign node3655 = (inp[0]) ? node3657 : 15'b000001111111111;
															assign node3657 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node3662 = (inp[3]) ? node3664 : 15'b000000111111111;
												assign node3664 = (inp[2]) ? 15'b000000011111111 : node3665;
													assign node3665 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node3669 = (inp[6]) ? node3689 : node3670;
											assign node3670 = (inp[2]) ? node3678 : node3671;
												assign node3671 = (inp[3]) ? 15'b000000111111111 : node3672;
													assign node3672 = (inp[0]) ? node3674 : 15'b000011111111111;
														assign node3674 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node3678 = (inp[3]) ? node3686 : node3679;
													assign node3679 = (inp[1]) ? 15'b000000011111111 : node3680;
														assign node3680 = (inp[0]) ? node3682 : 15'b000000111111111;
															assign node3682 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3686 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3689 = (inp[0]) ? node3701 : node3690;
												assign node3690 = (inp[1]) ? node3696 : node3691;
													assign node3691 = (inp[2]) ? node3693 : 15'b000000111111111;
														assign node3693 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node3696 = (inp[3]) ? node3698 : 15'b000000011111111;
														assign node3698 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3701 = (inp[3]) ? node3703 : 15'b000000001111111;
													assign node3703 = (inp[5]) ? node3705 : 15'b000000001111111;
														assign node3705 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node3708 = (inp[1]) ? node3736 : node3709;
										assign node3709 = (inp[0]) ? node3723 : node3710;
											assign node3710 = (inp[3]) ? node3720 : node3711;
												assign node3711 = (inp[2]) ? node3715 : node3712;
													assign node3712 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3715 = (inp[6]) ? node3717 : 15'b000000111111111;
														assign node3717 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3720 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3723 = (inp[6]) ? node3725 : 15'b000000011111111;
												assign node3725 = (inp[3]) ? node3731 : node3726;
													assign node3726 = (inp[13]) ? node3728 : 15'b000000001111111;
														assign node3728 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3731 = (inp[13]) ? 15'b000000001111111 : node3732;
														assign node3732 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3736 = (inp[2]) ? node3754 : node3737;
											assign node3737 = (inp[3]) ? node3747 : node3738;
												assign node3738 = (inp[5]) ? 15'b000000001111111 : node3739;
													assign node3739 = (inp[13]) ? 15'b000000011111111 : node3740;
														assign node3740 = (inp[0]) ? node3742 : 15'b000000111111111;
															assign node3742 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3747 = (inp[6]) ? node3751 : node3748;
													assign node3748 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3751 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3754 = (inp[0]) ? node3764 : node3755;
												assign node3755 = (inp[6]) ? node3759 : node3756;
													assign node3756 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node3759 = (inp[3]) ? node3761 : 15'b000000001111111;
														assign node3761 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3764 = (inp[13]) ? node3766 : 15'b000000000111111;
													assign node3766 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node3769 = (inp[5]) ? node3839 : node3770;
									assign node3770 = (inp[0]) ? node3800 : node3771;
										assign node3771 = (inp[6]) ? node3787 : node3772;
											assign node3772 = (inp[13]) ? node3782 : node3773;
												assign node3773 = (inp[2]) ? node3777 : node3774;
													assign node3774 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node3777 = (inp[3]) ? node3779 : 15'b000000111111111;
														assign node3779 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3782 = (inp[2]) ? 15'b000000011111111 : node3783;
													assign node3783 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node3787 = (inp[13]) ? node3797 : node3788;
												assign node3788 = (inp[1]) ? node3792 : node3789;
													assign node3789 = (inp[3]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node3792 = (inp[10]) ? 15'b000000001111111 : node3793;
														assign node3793 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node3797 = (inp[1]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node3800 = (inp[13]) ? node3820 : node3801;
											assign node3801 = (inp[3]) ? node3807 : node3802;
												assign node3802 = (inp[1]) ? 15'b000000011111111 : node3803;
													assign node3803 = (inp[6]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node3807 = (inp[1]) ? node3815 : node3808;
													assign node3808 = (inp[2]) ? node3810 : 15'b000000011111111;
														assign node3810 = (inp[10]) ? 15'b000000000111111 : node3811;
															assign node3811 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3815 = (inp[2]) ? node3817 : 15'b000000001111111;
														assign node3817 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3820 = (inp[1]) ? node3830 : node3821;
												assign node3821 = (inp[2]) ? node3823 : 15'b000000001111111;
													assign node3823 = (inp[3]) ? node3825 : 15'b000000001111111;
														assign node3825 = (inp[10]) ? 15'b000000000111111 : node3826;
															assign node3826 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3830 = (inp[10]) ? node3834 : node3831;
													assign node3831 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3834 = (inp[3]) ? 15'b000000000011111 : node3835;
														assign node3835 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3839 = (inp[1]) ? node3861 : node3840;
										assign node3840 = (inp[0]) ? node3848 : node3841;
											assign node3841 = (inp[3]) ? 15'b000000001111111 : node3842;
												assign node3842 = (inp[2]) ? node3844 : 15'b000000111111111;
													assign node3844 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3848 = (inp[13]) ? node3856 : node3849;
												assign node3849 = (inp[3]) ? node3853 : node3850;
													assign node3850 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3853 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3856 = (inp[10]) ? node3858 : 15'b000000000111111;
													assign node3858 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node3861 = (inp[13]) ? node3881 : node3862;
											assign node3862 = (inp[10]) ? node3872 : node3863;
												assign node3863 = (inp[3]) ? node3865 : 15'b000000001111111;
													assign node3865 = (inp[6]) ? 15'b000000000111111 : node3866;
														assign node3866 = (inp[0]) ? node3868 : 15'b000000001111111;
															assign node3868 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3872 = (inp[0]) ? node3878 : node3873;
													assign node3873 = (inp[3]) ? 15'b000000000111111 : node3874;
														assign node3874 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3878 = (inp[6]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node3881 = (inp[6]) ? node3887 : node3882;
												assign node3882 = (inp[0]) ? 15'b000000000111111 : node3883;
													assign node3883 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3887 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node3890 = (inp[2]) ? node4040 : node3891;
								assign node3891 = (inp[11]) ? node3951 : node3892;
									assign node3892 = (inp[13]) ? node3920 : node3893;
										assign node3893 = (inp[10]) ? node3909 : node3894;
											assign node3894 = (inp[3]) ? node3904 : node3895;
												assign node3895 = (inp[5]) ? node3901 : node3896;
													assign node3896 = (inp[0]) ? 15'b000000111111111 : node3897;
														assign node3897 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node3901 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3904 = (inp[6]) ? node3906 : 15'b000000111111111;
													assign node3906 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node3909 = (inp[5]) ? node3915 : node3910;
												assign node3910 = (inp[0]) ? 15'b000000011111111 : node3911;
													assign node3911 = (inp[1]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node3915 = (inp[1]) ? 15'b000000001111111 : node3916;
													assign node3916 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node3920 = (inp[10]) ? node3934 : node3921;
											assign node3921 = (inp[0]) ? node3929 : node3922;
												assign node3922 = (inp[3]) ? node3924 : 15'b000000111111111;
													assign node3924 = (inp[6]) ? 15'b000000001111111 : node3925;
														assign node3925 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3929 = (inp[1]) ? 15'b000000001111111 : node3930;
													assign node3930 = (inp[5]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node3934 = (inp[5]) ? node3942 : node3935;
												assign node3935 = (inp[0]) ? node3939 : node3936;
													assign node3936 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3939 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3942 = (inp[3]) ? node3946 : node3943;
													assign node3943 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node3946 = (inp[0]) ? 15'b000000000001111 : node3947;
														assign node3947 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node3951 = (inp[5]) ? node3989 : node3952;
										assign node3952 = (inp[10]) ? node3972 : node3953;
											assign node3953 = (inp[6]) ? node3963 : node3954;
												assign node3954 = (inp[13]) ? 15'b000000011111111 : node3955;
													assign node3955 = (inp[0]) ? 15'b000000011111111 : node3956;
														assign node3956 = (inp[1]) ? node3958 : 15'b000000111111111;
															assign node3958 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node3963 = (inp[1]) ? node3967 : node3964;
													assign node3964 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node3967 = (inp[0]) ? node3969 : 15'b000000001111111;
														assign node3969 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node3972 = (inp[13]) ? node3984 : node3973;
												assign node3973 = (inp[0]) ? node3979 : node3974;
													assign node3974 = (inp[3]) ? 15'b000000001111111 : node3975;
														assign node3975 = (inp[6]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node3979 = (inp[1]) ? 15'b000000000111111 : node3980;
														assign node3980 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3984 = (inp[6]) ? 15'b000000000111111 : node3985;
													assign node3985 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node3989 = (inp[3]) ? node4017 : node3990;
											assign node3990 = (inp[13]) ? node3998 : node3991;
												assign node3991 = (inp[6]) ? node3993 : 15'b000000001111111;
													assign node3993 = (inp[10]) ? node3995 : 15'b000000001111111;
														assign node3995 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node3998 = (inp[1]) ? node4006 : node3999;
													assign node3999 = (inp[0]) ? node4001 : 15'b000000001111111;
														assign node4001 = (inp[10]) ? 15'b000000000111111 : node4002;
															assign node4002 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4006 = (inp[6]) ? node4012 : node4007;
														assign node4007 = (inp[10]) ? 15'b000000000111111 : node4008;
															assign node4008 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
														assign node4012 = (inp[10]) ? 15'b000000000001111 : node4013;
															assign node4013 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4017 = (inp[0]) ? node4027 : node4018;
												assign node4018 = (inp[6]) ? node4020 : 15'b000000001111111;
													assign node4020 = (inp[1]) ? node4022 : 15'b000000000111111;
														assign node4022 = (inp[13]) ? node4024 : 15'b000000000011111;
															assign node4024 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node4027 = (inp[10]) ? node4029 : 15'b000000000011111;
													assign node4029 = (inp[13]) ? node4035 : node4030;
														assign node4030 = (inp[1]) ? node4032 : 15'b000000000111111;
															assign node4032 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
														assign node4035 = (inp[6]) ? node4037 : 15'b000000000001111;
															assign node4037 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node4040 = (inp[0]) ? node4116 : node4041;
									assign node4041 = (inp[13]) ? node4087 : node4042;
										assign node4042 = (inp[3]) ? node4060 : node4043;
											assign node4043 = (inp[11]) ? node4053 : node4044;
												assign node4044 = (inp[10]) ? node4046 : 15'b000000111111111;
													assign node4046 = (inp[6]) ? 15'b000000011111111 : node4047;
														assign node4047 = (inp[5]) ? 15'b000000011111111 : node4048;
															assign node4048 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4053 = (inp[1]) ? 15'b000000000111111 : node4054;
													assign node4054 = (inp[6]) ? 15'b000000001111111 : node4055;
														assign node4055 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4060 = (inp[6]) ? node4068 : node4061;
												assign node4061 = (inp[10]) ? node4065 : node4062;
													assign node4062 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4065 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4068 = (inp[11]) ? node4080 : node4069;
													assign node4069 = (inp[1]) ? node4075 : node4070;
														assign node4070 = (inp[5]) ? node4072 : 15'b000000001111111;
															assign node4072 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
														assign node4075 = (inp[10]) ? node4077 : 15'b000000000111111;
															assign node4077 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node4080 = (inp[10]) ? node4084 : node4081;
														assign node4081 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
														assign node4084 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node4087 = (inp[11]) ? node4097 : node4088;
											assign node4088 = (inp[5]) ? 15'b000000000111111 : node4089;
												assign node4089 = (inp[1]) ? node4091 : 15'b000000001111111;
													assign node4091 = (inp[3]) ? 15'b000000000111111 : node4092;
														assign node4092 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node4097 = (inp[6]) ? node4105 : node4098;
												assign node4098 = (inp[1]) ? node4100 : 15'b000000001111111;
													assign node4100 = (inp[5]) ? node4102 : 15'b000000000111111;
														assign node4102 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4105 = (inp[5]) ? node4111 : node4106;
													assign node4106 = (inp[1]) ? 15'b000000000011111 : node4107;
														assign node4107 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node4111 = (inp[3]) ? node4113 : 15'b000000000011111;
														assign node4113 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node4116 = (inp[13]) ? node4150 : node4117;
										assign node4117 = (inp[11]) ? node4131 : node4118;
											assign node4118 = (inp[6]) ? node4124 : node4119;
												assign node4119 = (inp[5]) ? 15'b000000000111111 : node4120;
													assign node4120 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4124 = (inp[3]) ? node4126 : 15'b000000000111111;
													assign node4126 = (inp[10]) ? node4128 : 15'b000000000111111;
														assign node4128 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4131 = (inp[3]) ? node4141 : node4132;
												assign node4132 = (inp[5]) ? node4138 : node4133;
													assign node4133 = (inp[1]) ? 15'b000000000111111 : node4134;
														assign node4134 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node4138 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node4141 = (inp[6]) ? node4145 : node4142;
													assign node4142 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node4145 = (inp[5]) ? node4147 : 15'b000000000001111;
														assign node4147 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node4150 = (inp[1]) ? node4166 : node4151;
											assign node4151 = (inp[3]) ? node4159 : node4152;
												assign node4152 = (inp[11]) ? node4154 : 15'b000000000111111;
													assign node4154 = (inp[10]) ? node4156 : 15'b000000000111111;
														assign node4156 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node4159 = (inp[5]) ? node4161 : 15'b000000000011111;
													assign node4161 = (inp[11]) ? node4163 : 15'b000000000011111;
														assign node4163 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node4166 = (inp[11]) ? node4174 : node4167;
												assign node4167 = (inp[5]) ? node4169 : 15'b000000000011111;
													assign node4169 = (inp[10]) ? 15'b000000000000111 : node4170;
														assign node4170 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node4174 = (inp[5]) ? 15'b000000000000111 : node4175;
													assign node4175 = (inp[6]) ? node4177 : 15'b000000000001111;
														assign node4177 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
			assign node4181 = (inp[11]) ? node6219 : node4182;
				assign node4182 = (inp[10]) ? node5222 : node4183;
					assign node4183 = (inp[9]) ? node4711 : node4184;
						assign node4184 = (inp[0]) ? node4438 : node4185;
							assign node4185 = (inp[3]) ? node4321 : node4186;
								assign node4186 = (inp[6]) ? node4260 : node4187;
									assign node4187 = (inp[5]) ? node4231 : node4188;
										assign node4188 = (inp[4]) ? node4206 : node4189;
											assign node4189 = (inp[1]) ? node4195 : node4190;
												assign node4190 = (inp[2]) ? node4192 : 15'b001111111111111;
													assign node4192 = (inp[14]) ? 15'b000111111111111 : 15'b001111111111111;
												assign node4195 = (inp[14]) ? node4203 : node4196;
													assign node4196 = (inp[13]) ? node4200 : node4197;
														assign node4197 = (inp[8]) ? 15'b000111111111111 : 15'b001111111111111;
														assign node4200 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node4203 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node4206 = (inp[13]) ? node4224 : node4207;
												assign node4207 = (inp[14]) ? node4211 : node4208;
													assign node4208 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node4211 = (inp[1]) ? node4219 : node4212;
														assign node4212 = (inp[8]) ? node4216 : node4213;
															assign node4213 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
															assign node4216 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
														assign node4219 = (inp[2]) ? 15'b000001111111111 : node4220;
															assign node4220 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4224 = (inp[8]) ? node4228 : node4225;
													assign node4225 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4228 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node4231 = (inp[1]) ? node4249 : node4232;
											assign node4232 = (inp[4]) ? node4242 : node4233;
												assign node4233 = (inp[2]) ? 15'b000011111111111 : node4234;
													assign node4234 = (inp[8]) ? node4236 : 15'b000111111111111;
														assign node4236 = (inp[13]) ? 15'b000011111111111 : node4237;
															assign node4237 = (inp[14]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node4242 = (inp[8]) ? node4246 : node4243;
													assign node4243 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4246 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4249 = (inp[2]) ? node4255 : node4250;
												assign node4250 = (inp[14]) ? node4252 : 15'b000001111111111;
													assign node4252 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4255 = (inp[13]) ? 15'b000000111111111 : node4256;
													assign node4256 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node4260 = (inp[5]) ? node4290 : node4261;
										assign node4261 = (inp[2]) ? node4273 : node4262;
											assign node4262 = (inp[14]) ? 15'b000001111111111 : node4263;
												assign node4263 = (inp[4]) ? node4267 : node4264;
													assign node4264 = (inp[8]) ? 15'b000011111111111 : 15'b001111111111111;
													assign node4267 = (inp[8]) ? node4269 : 15'b000011111111111;
														assign node4269 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node4273 = (inp[13]) ? node4285 : node4274;
												assign node4274 = (inp[8]) ? node4280 : node4275;
													assign node4275 = (inp[14]) ? 15'b000001111111111 : node4276;
														assign node4276 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node4280 = (inp[14]) ? node4282 : 15'b000001111111111;
														assign node4282 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4285 = (inp[8]) ? 15'b000000111111111 : node4286;
													assign node4286 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node4290 = (inp[1]) ? node4308 : node4291;
											assign node4291 = (inp[13]) ? node4305 : node4292;
												assign node4292 = (inp[8]) ? node4298 : node4293;
													assign node4293 = (inp[4]) ? node4295 : 15'b000011111111111;
														assign node4295 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4298 = (inp[14]) ? node4300 : 15'b000001111111111;
														assign node4300 = (inp[4]) ? 15'b000000111111111 : node4301;
															assign node4301 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4305 = (inp[14]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node4308 = (inp[8]) ? node4312 : node4309;
												assign node4309 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4312 = (inp[4]) ? 15'b000000001111111 : node4313;
													assign node4313 = (inp[2]) ? 15'b000000011111111 : node4314;
														assign node4314 = (inp[14]) ? node4316 : 15'b000000111111111;
															assign node4316 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node4321 = (inp[1]) ? node4385 : node4322;
									assign node4322 = (inp[14]) ? node4352 : node4323;
										assign node4323 = (inp[6]) ? node4339 : node4324;
											assign node4324 = (inp[2]) ? node4330 : node4325;
												assign node4325 = (inp[4]) ? 15'b000011111111111 : node4326;
													assign node4326 = (inp[13]) ? 15'b000011111111111 : 15'b001111111111111;
												assign node4330 = (inp[4]) ? 15'b000000111111111 : node4331;
													assign node4331 = (inp[8]) ? node4333 : 15'b000011111111111;
														assign node4333 = (inp[13]) ? 15'b000001111111111 : node4334;
															assign node4334 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node4339 = (inp[4]) ? node4347 : node4340;
												assign node4340 = (inp[8]) ? 15'b000001111111111 : node4341;
													assign node4341 = (inp[5]) ? 15'b000001111111111 : node4342;
														assign node4342 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4347 = (inp[2]) ? 15'b000000111111111 : node4348;
													assign node4348 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node4352 = (inp[8]) ? node4370 : node4353;
											assign node4353 = (inp[2]) ? node4365 : node4354;
												assign node4354 = (inp[5]) ? node4362 : node4355;
													assign node4355 = (inp[4]) ? 15'b000001111111111 : node4356;
														assign node4356 = (inp[6]) ? node4358 : 15'b000011111111111;
															assign node4358 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4362 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4365 = (inp[4]) ? 15'b000000111111111 : node4366;
													assign node4366 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4370 = (inp[4]) ? node4380 : node4371;
												assign node4371 = (inp[5]) ? node4375 : node4372;
													assign node4372 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4375 = (inp[2]) ? node4377 : 15'b000000111111111;
														assign node4377 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4380 = (inp[6]) ? node4382 : 15'b000000011111111;
													assign node4382 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node4385 = (inp[6]) ? node4415 : node4386;
										assign node4386 = (inp[13]) ? node4402 : node4387;
											assign node4387 = (inp[2]) ? node4395 : node4388;
												assign node4388 = (inp[8]) ? 15'b000001111111111 : node4389;
													assign node4389 = (inp[4]) ? node4391 : 15'b000111111111111;
														assign node4391 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4395 = (inp[8]) ? node4399 : node4396;
													assign node4396 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4399 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4402 = (inp[14]) ? 15'b000000011111111 : node4403;
												assign node4403 = (inp[5]) ? node4407 : node4404;
													assign node4404 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4407 = (inp[4]) ? node4409 : 15'b000001111111111;
														assign node4409 = (inp[8]) ? 15'b000000011111111 : node4410;
															assign node4410 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4415 = (inp[14]) ? node4433 : node4416;
											assign node4416 = (inp[4]) ? node4422 : node4417;
												assign node4417 = (inp[5]) ? node4419 : 15'b000000111111111;
													assign node4419 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node4422 = (inp[8]) ? node4428 : node4423;
													assign node4423 = (inp[5]) ? 15'b000000011111111 : node4424;
														assign node4424 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4428 = (inp[13]) ? node4430 : 15'b000000011111111;
														assign node4430 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4433 = (inp[5]) ? node4435 : 15'b000000011111111;
												assign node4435 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node4438 = (inp[6]) ? node4584 : node4439;
								assign node4439 = (inp[14]) ? node4509 : node4440;
									assign node4440 = (inp[8]) ? node4468 : node4441;
										assign node4441 = (inp[2]) ? node4455 : node4442;
											assign node4442 = (inp[4]) ? node4450 : node4443;
												assign node4443 = (inp[13]) ? node4445 : 15'b000011111111111;
													assign node4445 = (inp[1]) ? node4447 : 15'b000011111111111;
														assign node4447 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4450 = (inp[5]) ? 15'b000001111111111 : node4451;
													assign node4451 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node4455 = (inp[13]) ? node4461 : node4456;
												assign node4456 = (inp[3]) ? node4458 : 15'b000001111111111;
													assign node4458 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4461 = (inp[4]) ? 15'b000000111111111 : node4462;
													assign node4462 = (inp[1]) ? node4464 : 15'b000001111111111;
														assign node4464 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node4468 = (inp[1]) ? node4490 : node4469;
											assign node4469 = (inp[2]) ? node4479 : node4470;
												assign node4470 = (inp[4]) ? node4476 : node4471;
													assign node4471 = (inp[5]) ? 15'b000001111111111 : node4472;
														assign node4472 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4476 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4479 = (inp[4]) ? node4483 : node4480;
													assign node4480 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4483 = (inp[3]) ? node4485 : 15'b000000111111111;
														assign node4485 = (inp[13]) ? 15'b000000011111111 : node4486;
															assign node4486 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4490 = (inp[5]) ? node4498 : node4491;
												assign node4491 = (inp[13]) ? node4495 : node4492;
													assign node4492 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4495 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4498 = (inp[4]) ? node4502 : node4499;
													assign node4499 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4502 = (inp[13]) ? node4504 : 15'b000000111111111;
														assign node4504 = (inp[3]) ? node4506 : 15'b000000001111111;
															assign node4506 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4509 = (inp[4]) ? node4547 : node4510;
										assign node4510 = (inp[3]) ? node4526 : node4511;
											assign node4511 = (inp[13]) ? node4513 : 15'b000001111111111;
												assign node4513 = (inp[1]) ? 15'b000000111111111 : node4514;
													assign node4514 = (inp[2]) ? node4520 : node4515;
														assign node4515 = (inp[8]) ? node4517 : 15'b000001111111111;
															assign node4517 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node4520 = (inp[8]) ? 15'b000000111111111 : node4521;
															assign node4521 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4526 = (inp[8]) ? node4534 : node4527;
												assign node4527 = (inp[1]) ? node4529 : 15'b000001111111111;
													assign node4529 = (inp[13]) ? node4531 : 15'b000000111111111;
														assign node4531 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4534 = (inp[13]) ? node4542 : node4535;
													assign node4535 = (inp[2]) ? 15'b000000011111111 : node4536;
														assign node4536 = (inp[1]) ? node4538 : 15'b000000111111111;
															assign node4538 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4542 = (inp[2]) ? node4544 : 15'b000000011111111;
														assign node4544 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node4547 = (inp[1]) ? node4563 : node4548;
											assign node4548 = (inp[8]) ? node4558 : node4549;
												assign node4549 = (inp[2]) ? node4551 : 15'b000000111111111;
													assign node4551 = (inp[13]) ? node4553 : 15'b000000111111111;
														assign node4553 = (inp[5]) ? 15'b000000011111111 : node4554;
															assign node4554 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4558 = (inp[5]) ? 15'b000000011111111 : node4559;
													assign node4559 = (inp[13]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node4563 = (inp[5]) ? node4575 : node4564;
												assign node4564 = (inp[13]) ? node4572 : node4565;
													assign node4565 = (inp[3]) ? 15'b000000011111111 : node4566;
														assign node4566 = (inp[8]) ? node4568 : 15'b000000111111111;
															assign node4568 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4572 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4575 = (inp[2]) ? node4581 : node4576;
													assign node4576 = (inp[3]) ? 15'b000000001111111 : node4577;
														assign node4577 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4581 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node4584 = (inp[13]) ? node4656 : node4585;
									assign node4585 = (inp[8]) ? node4625 : node4586;
										assign node4586 = (inp[1]) ? node4602 : node4587;
											assign node4587 = (inp[2]) ? node4595 : node4588;
												assign node4588 = (inp[3]) ? node4590 : 15'b000011111111111;
													assign node4590 = (inp[5]) ? node4592 : 15'b000001111111111;
														assign node4592 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4595 = (inp[14]) ? node4597 : 15'b000001111111111;
													assign node4597 = (inp[3]) ? node4599 : 15'b000000111111111;
														assign node4599 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4602 = (inp[5]) ? node4612 : node4603;
												assign node4603 = (inp[3]) ? node4609 : node4604;
													assign node4604 = (inp[4]) ? 15'b000000111111111 : node4605;
														assign node4605 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node4609 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4612 = (inp[4]) ? node4620 : node4613;
													assign node4613 = (inp[2]) ? node4615 : 15'b000000111111111;
														assign node4615 = (inp[14]) ? 15'b000000011111111 : node4616;
															assign node4616 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4620 = (inp[14]) ? node4622 : 15'b000000011111111;
														assign node4622 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4625 = (inp[4]) ? node4647 : node4626;
											assign node4626 = (inp[3]) ? node4632 : node4627;
												assign node4627 = (inp[5]) ? node4629 : 15'b000000111111111;
													assign node4629 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4632 = (inp[2]) ? node4642 : node4633;
													assign node4633 = (inp[1]) ? node4639 : node4634;
														assign node4634 = (inp[14]) ? node4636 : 15'b000000111111111;
															assign node4636 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node4639 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4642 = (inp[14]) ? node4644 : 15'b000000011111111;
														assign node4644 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4647 = (inp[1]) ? node4651 : node4648;
												assign node4648 = (inp[3]) ? 15'b000000001111111 : 15'b000001111111111;
												assign node4651 = (inp[2]) ? node4653 : 15'b000000001111111;
													assign node4653 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4656 = (inp[5]) ? node4688 : node4657;
										assign node4657 = (inp[1]) ? node4681 : node4658;
											assign node4658 = (inp[8]) ? node4670 : node4659;
												assign node4659 = (inp[2]) ? node4663 : node4660;
													assign node4660 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4663 = (inp[4]) ? node4665 : 15'b000000111111111;
														assign node4665 = (inp[3]) ? 15'b000000011111111 : node4666;
															assign node4666 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4670 = (inp[14]) ? node4678 : node4671;
													assign node4671 = (inp[2]) ? node4675 : node4672;
														assign node4672 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node4675 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4678 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4681 = (inp[4]) ? 15'b000000001111111 : node4682;
												assign node4682 = (inp[14]) ? node4684 : 15'b000000011111111;
													assign node4684 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4688 = (inp[2]) ? node4700 : node4689;
											assign node4689 = (inp[14]) ? node4693 : node4690;
												assign node4690 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4693 = (inp[3]) ? 15'b000000001111111 : node4694;
													assign node4694 = (inp[4]) ? node4696 : 15'b000000111111111;
														assign node4696 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4700 = (inp[4]) ? node4704 : node4701;
												assign node4701 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4704 = (inp[8]) ? 15'b000000000011111 : node4705;
													assign node4705 = (inp[1]) ? node4707 : 15'b000000001111111;
														assign node4707 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node4711 = (inp[5]) ? node4967 : node4712;
							assign node4712 = (inp[3]) ? node4838 : node4713;
								assign node4713 = (inp[2]) ? node4781 : node4714;
									assign node4714 = (inp[6]) ? node4750 : node4715;
										assign node4715 = (inp[4]) ? node4735 : node4716;
											assign node4716 = (inp[8]) ? node4728 : node4717;
												assign node4717 = (inp[14]) ? node4723 : node4718;
													assign node4718 = (inp[0]) ? 15'b000011111111111 : node4719;
														assign node4719 = (inp[1]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node4723 = (inp[13]) ? node4725 : 15'b000011111111111;
														assign node4725 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node4728 = (inp[14]) ? 15'b000000111111111 : node4729;
													assign node4729 = (inp[0]) ? 15'b000001111111111 : node4730;
														assign node4730 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node4735 = (inp[1]) ? node4741 : node4736;
												assign node4736 = (inp[0]) ? 15'b000001111111111 : node4737;
													assign node4737 = (inp[8]) ? 15'b000001111111111 : 15'b000111111111111;
												assign node4741 = (inp[8]) ? 15'b000000111111111 : node4742;
													assign node4742 = (inp[13]) ? 15'b000000111111111 : node4743;
														assign node4743 = (inp[0]) ? node4745 : 15'b000001111111111;
															assign node4745 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node4750 = (inp[13]) ? node4766 : node4751;
											assign node4751 = (inp[4]) ? node4759 : node4752;
												assign node4752 = (inp[0]) ? 15'b000001111111111 : node4753;
													assign node4753 = (inp[1]) ? 15'b000011111111111 : node4754;
														assign node4754 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node4759 = (inp[8]) ? node4763 : node4760;
													assign node4760 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4763 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4766 = (inp[1]) ? node4776 : node4767;
												assign node4767 = (inp[8]) ? node4771 : node4768;
													assign node4768 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4771 = (inp[4]) ? node4773 : 15'b000000111111111;
														assign node4773 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4776 = (inp[8]) ? 15'b000000011111111 : node4777;
													assign node4777 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node4781 = (inp[6]) ? node4803 : node4782;
										assign node4782 = (inp[1]) ? node4794 : node4783;
											assign node4783 = (inp[13]) ? node4789 : node4784;
												assign node4784 = (inp[14]) ? node4786 : 15'b000001111111111;
													assign node4786 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4789 = (inp[4]) ? node4791 : 15'b000001111111111;
													assign node4791 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4794 = (inp[0]) ? node4796 : 15'b000000111111111;
												assign node4796 = (inp[14]) ? node4800 : node4797;
													assign node4797 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4800 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4803 = (inp[4]) ? node4825 : node4804;
											assign node4804 = (inp[14]) ? node4816 : node4805;
												assign node4805 = (inp[13]) ? node4813 : node4806;
													assign node4806 = (inp[1]) ? node4808 : 15'b000001111111111;
														assign node4808 = (inp[0]) ? 15'b000000111111111 : node4809;
															assign node4809 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4813 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4816 = (inp[8]) ? node4822 : node4817;
													assign node4817 = (inp[1]) ? 15'b000000011111111 : node4818;
														assign node4818 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4822 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4825 = (inp[13]) ? node4831 : node4826;
												assign node4826 = (inp[14]) ? node4828 : 15'b000000011111111;
													assign node4828 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4831 = (inp[8]) ? 15'b000000001111111 : node4832;
													assign node4832 = (inp[0]) ? 15'b000000011111111 : node4833;
														assign node4833 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
								assign node4838 = (inp[4]) ? node4896 : node4839;
									assign node4839 = (inp[6]) ? node4877 : node4840;
										assign node4840 = (inp[1]) ? node4858 : node4841;
											assign node4841 = (inp[13]) ? node4849 : node4842;
												assign node4842 = (inp[14]) ? node4844 : 15'b000001111111111;
													assign node4844 = (inp[0]) ? node4846 : 15'b000001111111111;
														assign node4846 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4849 = (inp[14]) ? node4853 : node4850;
													assign node4850 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4853 = (inp[8]) ? 15'b000000001111111 : node4854;
														assign node4854 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node4858 = (inp[8]) ? node4866 : node4859;
												assign node4859 = (inp[14]) ? node4861 : 15'b000011111111111;
													assign node4861 = (inp[0]) ? 15'b000000111111111 : node4862;
														assign node4862 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4866 = (inp[14]) ? node4874 : node4867;
													assign node4867 = (inp[13]) ? node4869 : 15'b000000111111111;
														assign node4869 = (inp[2]) ? 15'b000000011111111 : node4870;
															assign node4870 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4874 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4877 = (inp[14]) ? node4889 : node4878;
											assign node4878 = (inp[2]) ? node4884 : node4879;
												assign node4879 = (inp[0]) ? node4881 : 15'b000000111111111;
													assign node4881 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4884 = (inp[0]) ? node4886 : 15'b000000011111111;
													assign node4886 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node4889 = (inp[8]) ? node4891 : 15'b000000011111111;
												assign node4891 = (inp[2]) ? node4893 : 15'b000000011111111;
													assign node4893 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node4896 = (inp[14]) ? node4926 : node4897;
										assign node4897 = (inp[13]) ? node4913 : node4898;
											assign node4898 = (inp[0]) ? node4906 : node4899;
												assign node4899 = (inp[6]) ? node4903 : node4900;
													assign node4900 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node4903 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4906 = (inp[1]) ? node4910 : node4907;
													assign node4907 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node4910 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node4913 = (inp[6]) ? node4921 : node4914;
												assign node4914 = (inp[8]) ? node4916 : 15'b000000011111111;
													assign node4916 = (inp[1]) ? node4918 : 15'b000000011111111;
														assign node4918 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node4921 = (inp[1]) ? node4923 : 15'b000000001111111;
													assign node4923 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node4926 = (inp[2]) ? node4954 : node4927;
											assign node4927 = (inp[13]) ? node4935 : node4928;
												assign node4928 = (inp[6]) ? node4930 : 15'b000000111111111;
													assign node4930 = (inp[1]) ? 15'b000000011111111 : node4931;
														assign node4931 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node4935 = (inp[1]) ? node4945 : node4936;
													assign node4936 = (inp[6]) ? 15'b000000001111111 : node4937;
														assign node4937 = (inp[0]) ? node4941 : node4938;
															assign node4938 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
															assign node4941 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node4945 = (inp[0]) ? node4947 : 15'b000000001111111;
														assign node4947 = (inp[8]) ? node4951 : node4948;
															assign node4948 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
															assign node4951 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node4954 = (inp[6]) ? node4960 : node4955;
												assign node4955 = (inp[1]) ? node4957 : 15'b000000001111111;
													assign node4957 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node4960 = (inp[13]) ? 15'b000000000011111 : node4961;
													assign node4961 = (inp[0]) ? node4963 : 15'b000000000111111;
														assign node4963 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node4967 = (inp[1]) ? node5085 : node4968;
								assign node4968 = (inp[0]) ? node5024 : node4969;
									assign node4969 = (inp[14]) ? node4999 : node4970;
										assign node4970 = (inp[6]) ? node4988 : node4971;
											assign node4971 = (inp[2]) ? node4979 : node4972;
												assign node4972 = (inp[8]) ? node4974 : 15'b000011111111111;
													assign node4974 = (inp[4]) ? node4976 : 15'b000001111111111;
														assign node4976 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node4979 = (inp[3]) ? 15'b000000111111111 : node4980;
													assign node4980 = (inp[8]) ? node4982 : 15'b000001111111111;
														assign node4982 = (inp[13]) ? 15'b000000111111111 : node4983;
															assign node4983 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node4988 = (inp[13]) ? node4990 : 15'b000000111111111;
												assign node4990 = (inp[3]) ? 15'b000000011111111 : node4991;
													assign node4991 = (inp[8]) ? node4993 : 15'b000001111111111;
														assign node4993 = (inp[2]) ? 15'b000000011111111 : node4994;
															assign node4994 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node4999 = (inp[8]) ? node5009 : node5000;
											assign node5000 = (inp[4]) ? node5004 : node5001;
												assign node5001 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5004 = (inp[2]) ? 15'b000000001111111 : node5005;
													assign node5005 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5009 = (inp[4]) ? node5017 : node5010;
												assign node5010 = (inp[13]) ? node5012 : 15'b000000001111111;
													assign node5012 = (inp[6]) ? node5014 : 15'b000000011111111;
														assign node5014 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5017 = (inp[3]) ? node5019 : 15'b000000001111111;
													assign node5019 = (inp[6]) ? 15'b000000000111111 : node5020;
														assign node5020 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5024 = (inp[8]) ? node5052 : node5025;
										assign node5025 = (inp[6]) ? node5039 : node5026;
											assign node5026 = (inp[2]) ? node5032 : node5027;
												assign node5027 = (inp[4]) ? node5029 : 15'b000000111111111;
													assign node5029 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5032 = (inp[4]) ? node5034 : 15'b000000011111111;
													assign node5034 = (inp[13]) ? 15'b000000011111111 : node5035;
														assign node5035 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5039 = (inp[13]) ? node5047 : node5040;
												assign node5040 = (inp[2]) ? node5042 : 15'b000000011111111;
													assign node5042 = (inp[4]) ? node5044 : 15'b000000011111111;
														assign node5044 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5047 = (inp[14]) ? 15'b000000001111111 : node5048;
													assign node5048 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5052 = (inp[2]) ? node5074 : node5053;
											assign node5053 = (inp[13]) ? node5065 : node5054;
												assign node5054 = (inp[3]) ? node5062 : node5055;
													assign node5055 = (inp[14]) ? 15'b000000011111111 : node5056;
														assign node5056 = (inp[4]) ? 15'b000000111111111 : node5057;
															assign node5057 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5062 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node5065 = (inp[6]) ? node5069 : node5066;
													assign node5066 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5069 = (inp[14]) ? 15'b000000000111111 : node5070;
														assign node5070 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5074 = (inp[3]) ? node5078 : node5075;
												assign node5075 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node5078 = (inp[6]) ? node5080 : 15'b000000000011111;
													assign node5080 = (inp[13]) ? 15'b000000000111111 : node5081;
														assign node5081 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node5085 = (inp[6]) ? node5147 : node5086;
									assign node5086 = (inp[2]) ? node5110 : node5087;
										assign node5087 = (inp[3]) ? node5095 : node5088;
											assign node5088 = (inp[8]) ? node5092 : node5089;
												assign node5089 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5092 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5095 = (inp[0]) ? node5103 : node5096;
												assign node5096 = (inp[4]) ? node5098 : 15'b000000111111111;
													assign node5098 = (inp[14]) ? node5100 : 15'b000000011111111;
														assign node5100 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5103 = (inp[8]) ? 15'b000000000111111 : node5104;
													assign node5104 = (inp[4]) ? 15'b000000001111111 : node5105;
														assign node5105 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5110 = (inp[4]) ? node5132 : node5111;
											assign node5111 = (inp[8]) ? node5121 : node5112;
												assign node5112 = (inp[3]) ? node5118 : node5113;
													assign node5113 = (inp[14]) ? 15'b000000011111111 : node5114;
														assign node5114 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5118 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5121 = (inp[0]) ? node5125 : node5122;
													assign node5122 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5125 = (inp[13]) ? node5127 : 15'b000000001111111;
														assign node5127 = (inp[3]) ? 15'b000000000111111 : node5128;
															assign node5128 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5132 = (inp[14]) ? node5142 : node5133;
												assign node5133 = (inp[13]) ? node5139 : node5134;
													assign node5134 = (inp[0]) ? node5136 : 15'b000000001111111;
														assign node5136 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5139 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5142 = (inp[13]) ? 15'b000000000111111 : node5143;
													assign node5143 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node5147 = (inp[4]) ? node5187 : node5148;
										assign node5148 = (inp[8]) ? node5168 : node5149;
											assign node5149 = (inp[14]) ? node5155 : node5150;
												assign node5150 = (inp[13]) ? 15'b000000111111111 : node5151;
													assign node5151 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5155 = (inp[3]) ? node5165 : node5156;
													assign node5156 = (inp[0]) ? node5162 : node5157;
														assign node5157 = (inp[13]) ? 15'b000000011111111 : node5158;
															assign node5158 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node5162 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5165 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node5168 = (inp[14]) ? node5176 : node5169;
												assign node5169 = (inp[13]) ? node5173 : node5170;
													assign node5170 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5173 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5176 = (inp[13]) ? node5182 : node5177;
													assign node5177 = (inp[0]) ? 15'b000000000111111 : node5178;
														assign node5178 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5182 = (inp[2]) ? 15'b000000000011111 : node5183;
														assign node5183 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5187 = (inp[14]) ? node5201 : node5188;
											assign node5188 = (inp[0]) ? node5194 : node5189;
												assign node5189 = (inp[2]) ? node5191 : 15'b000000001111111;
													assign node5191 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5194 = (inp[13]) ? node5196 : 15'b000000001111111;
													assign node5196 = (inp[3]) ? 15'b000000000011111 : node5197;
														assign node5197 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5201 = (inp[0]) ? node5211 : node5202;
												assign node5202 = (inp[8]) ? 15'b000000000011111 : node5203;
													assign node5203 = (inp[13]) ? node5205 : 15'b000000000111111;
														assign node5205 = (inp[3]) ? node5207 : 15'b000000000111111;
															assign node5207 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5211 = (inp[13]) ? node5215 : node5212;
													assign node5212 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node5215 = (inp[8]) ? 15'b000000000001111 : node5216;
														assign node5216 = (inp[2]) ? node5218 : 15'b000000000011111;
															assign node5218 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node5222 = (inp[3]) ? node5740 : node5223;
						assign node5223 = (inp[0]) ? node5477 : node5224;
							assign node5224 = (inp[8]) ? node5350 : node5225;
								assign node5225 = (inp[13]) ? node5301 : node5226;
									assign node5226 = (inp[14]) ? node5264 : node5227;
										assign node5227 = (inp[2]) ? node5247 : node5228;
											assign node5228 = (inp[4]) ? node5240 : node5229;
												assign node5229 = (inp[6]) ? node5235 : node5230;
													assign node5230 = (inp[9]) ? 15'b000011111111111 : node5231;
														assign node5231 = (inp[5]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node5235 = (inp[1]) ? node5237 : 15'b000011111111111;
														assign node5237 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5240 = (inp[6]) ? node5244 : node5241;
													assign node5241 = (inp[1]) ? 15'b000011111111111 : 15'b000001111111111;
													assign node5244 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5247 = (inp[1]) ? node5249 : 15'b000001111111111;
												assign node5249 = (inp[6]) ? node5259 : node5250;
													assign node5250 = (inp[5]) ? node5254 : node5251;
														assign node5251 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
														assign node5254 = (inp[4]) ? 15'b000000111111111 : node5255;
															assign node5255 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5259 = (inp[5]) ? node5261 : 15'b000000111111111;
														assign node5261 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5264 = (inp[6]) ? node5286 : node5265;
											assign node5265 = (inp[2]) ? node5271 : node5266;
												assign node5266 = (inp[9]) ? 15'b000001111111111 : node5267;
													assign node5267 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5271 = (inp[1]) ? node5279 : node5272;
													assign node5272 = (inp[5]) ? node5274 : 15'b000001111111111;
														assign node5274 = (inp[4]) ? 15'b000000111111111 : node5275;
															assign node5275 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5279 = (inp[4]) ? node5281 : 15'b000000111111111;
														assign node5281 = (inp[5]) ? 15'b000000011111111 : node5282;
															assign node5282 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5286 = (inp[1]) ? node5294 : node5287;
												assign node5287 = (inp[2]) ? node5291 : node5288;
													assign node5288 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5291 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5294 = (inp[4]) ? node5298 : node5295;
													assign node5295 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5298 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node5301 = (inp[1]) ? node5325 : node5302;
										assign node5302 = (inp[6]) ? node5314 : node5303;
											assign node5303 = (inp[9]) ? node5309 : node5304;
												assign node5304 = (inp[2]) ? node5306 : 15'b000011111111111;
													assign node5306 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5309 = (inp[5]) ? node5311 : 15'b000000111111111;
													assign node5311 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5314 = (inp[9]) ? node5320 : node5315;
												assign node5315 = (inp[5]) ? node5317 : 15'b000001111111111;
													assign node5317 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5320 = (inp[14]) ? 15'b000000011111111 : node5321;
													assign node5321 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5325 = (inp[6]) ? node5339 : node5326;
											assign node5326 = (inp[5]) ? node5334 : node5327;
												assign node5327 = (inp[9]) ? node5331 : node5328;
													assign node5328 = (inp[4]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node5331 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5334 = (inp[4]) ? 15'b000000011111111 : node5335;
													assign node5335 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5339 = (inp[5]) ? node5343 : node5340;
												assign node5340 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5343 = (inp[2]) ? 15'b000000000111111 : node5344;
													assign node5344 = (inp[4]) ? node5346 : 15'b000000011111111;
														assign node5346 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node5350 = (inp[2]) ? node5422 : node5351;
									assign node5351 = (inp[6]) ? node5387 : node5352;
										assign node5352 = (inp[1]) ? node5368 : node5353;
											assign node5353 = (inp[14]) ? node5363 : node5354;
												assign node5354 = (inp[9]) ? 15'b000001111111111 : node5355;
													assign node5355 = (inp[5]) ? 15'b000001111111111 : node5356;
														assign node5356 = (inp[13]) ? node5358 : 15'b000011111111111;
															assign node5358 = (inp[4]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5363 = (inp[4]) ? 15'b000000011111111 : node5364;
													assign node5364 = (inp[13]) ? 15'b000000111111111 : 15'b000011111111111;
											assign node5368 = (inp[9]) ? node5378 : node5369;
												assign node5369 = (inp[13]) ? node5373 : node5370;
													assign node5370 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5373 = (inp[14]) ? node5375 : 15'b000000111111111;
														assign node5375 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5378 = (inp[13]) ? 15'b000000001111111 : node5379;
													assign node5379 = (inp[4]) ? 15'b000000011111111 : node5380;
														assign node5380 = (inp[14]) ? node5382 : 15'b000000111111111;
															assign node5382 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node5387 = (inp[13]) ? node5411 : node5388;
											assign node5388 = (inp[4]) ? node5400 : node5389;
												assign node5389 = (inp[9]) ? node5397 : node5390;
													assign node5390 = (inp[1]) ? 15'b000000111111111 : node5391;
														assign node5391 = (inp[14]) ? 15'b000001111111111 : node5392;
															assign node5392 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node5397 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5400 = (inp[5]) ? node5408 : node5401;
													assign node5401 = (inp[9]) ? 15'b000000011111111 : node5402;
														assign node5402 = (inp[14]) ? node5404 : 15'b000000111111111;
															assign node5404 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5408 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5411 = (inp[4]) ? node5417 : node5412;
												assign node5412 = (inp[5]) ? node5414 : 15'b000000011111111;
													assign node5414 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5417 = (inp[14]) ? 15'b000000000111111 : node5418;
													assign node5418 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node5422 = (inp[5]) ? node5444 : node5423;
										assign node5423 = (inp[14]) ? node5435 : node5424;
											assign node5424 = (inp[1]) ? node5428 : node5425;
												assign node5425 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5428 = (inp[6]) ? 15'b000000011111111 : node5429;
													assign node5429 = (inp[13]) ? 15'b000000011111111 : node5430;
														assign node5430 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5435 = (inp[1]) ? node5441 : node5436;
												assign node5436 = (inp[6]) ? 15'b000000011111111 : node5437;
													assign node5437 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5441 = (inp[4]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node5444 = (inp[1]) ? node5462 : node5445;
											assign node5445 = (inp[4]) ? node5453 : node5446;
												assign node5446 = (inp[9]) ? node5450 : node5447;
													assign node5447 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5450 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5453 = (inp[9]) ? node5459 : node5454;
													assign node5454 = (inp[13]) ? 15'b000000001111111 : node5455;
														assign node5455 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5459 = (inp[14]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node5462 = (inp[6]) ? node5470 : node5463;
												assign node5463 = (inp[4]) ? node5465 : 15'b000000001111111;
													assign node5465 = (inp[14]) ? node5467 : 15'b000000001111111;
														assign node5467 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5470 = (inp[14]) ? node5472 : 15'b000000000111111;
													assign node5472 = (inp[4]) ? 15'b000000000001111 : node5473;
														assign node5473 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node5477 = (inp[5]) ? node5603 : node5478;
								assign node5478 = (inp[1]) ? node5542 : node5479;
									assign node5479 = (inp[14]) ? node5513 : node5480;
										assign node5480 = (inp[8]) ? node5498 : node5481;
											assign node5481 = (inp[4]) ? node5491 : node5482;
												assign node5482 = (inp[9]) ? node5488 : node5483;
													assign node5483 = (inp[2]) ? node5485 : 15'b000001111111111;
														assign node5485 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5488 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5491 = (inp[13]) ? node5493 : 15'b000000111111111;
													assign node5493 = (inp[6]) ? 15'b000000111111111 : node5494;
														assign node5494 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5498 = (inp[13]) ? node5510 : node5499;
												assign node5499 = (inp[6]) ? node5507 : node5500;
													assign node5500 = (inp[2]) ? 15'b000000111111111 : node5501;
														assign node5501 = (inp[9]) ? node5503 : 15'b000001111111111;
															assign node5503 = (inp[4]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5507 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5510 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5513 = (inp[4]) ? node5525 : node5514;
											assign node5514 = (inp[13]) ? node5520 : node5515;
												assign node5515 = (inp[8]) ? node5517 : 15'b000000111111111;
													assign node5517 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node5520 = (inp[2]) ? 15'b000000011111111 : node5521;
													assign node5521 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5525 = (inp[8]) ? 15'b000000001111111 : node5526;
												assign node5526 = (inp[2]) ? node5534 : node5527;
													assign node5527 = (inp[9]) ? node5529 : 15'b000000111111111;
														assign node5529 = (inp[6]) ? 15'b000000011111111 : node5530;
															assign node5530 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5534 = (inp[13]) ? node5536 : 15'b000000011111111;
														assign node5536 = (inp[6]) ? 15'b000000001111111 : node5537;
															assign node5537 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node5542 = (inp[9]) ? node5570 : node5543;
										assign node5543 = (inp[13]) ? node5551 : node5544;
											assign node5544 = (inp[8]) ? node5548 : node5545;
												assign node5545 = (inp[2]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node5548 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5551 = (inp[2]) ? node5559 : node5552;
												assign node5552 = (inp[4]) ? 15'b000000011111111 : node5553;
													assign node5553 = (inp[8]) ? node5555 : 15'b000000111111111;
														assign node5555 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5559 = (inp[14]) ? node5567 : node5560;
													assign node5560 = (inp[8]) ? node5562 : 15'b000000011111111;
														assign node5562 = (inp[6]) ? 15'b000000001111111 : node5563;
															assign node5563 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5567 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5570 = (inp[6]) ? node5586 : node5571;
											assign node5571 = (inp[13]) ? node5581 : node5572;
												assign node5572 = (inp[14]) ? node5578 : node5573;
													assign node5573 = (inp[4]) ? 15'b000000011111111 : node5574;
														assign node5574 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5578 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5581 = (inp[2]) ? 15'b000000001111111 : node5582;
													assign node5582 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5586 = (inp[2]) ? node5596 : node5587;
												assign node5587 = (inp[8]) ? 15'b000000001111111 : node5588;
													assign node5588 = (inp[4]) ? 15'b000000001111111 : node5589;
														assign node5589 = (inp[14]) ? node5591 : 15'b000000011111111;
															assign node5591 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5596 = (inp[4]) ? node5600 : node5597;
													assign node5597 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5600 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node5603 = (inp[8]) ? node5673 : node5604;
									assign node5604 = (inp[13]) ? node5638 : node5605;
										assign node5605 = (inp[14]) ? node5623 : node5606;
											assign node5606 = (inp[6]) ? node5618 : node5607;
												assign node5607 = (inp[4]) ? node5615 : node5608;
													assign node5608 = (inp[1]) ? node5610 : 15'b000001111111111;
														assign node5610 = (inp[9]) ? 15'b000000111111111 : node5611;
															assign node5611 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5615 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5618 = (inp[2]) ? 15'b000000001111111 : node5619;
													assign node5619 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5623 = (inp[4]) ? node5633 : node5624;
												assign node5624 = (inp[6]) ? node5630 : node5625;
													assign node5625 = (inp[9]) ? 15'b000000011111111 : node5626;
														assign node5626 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5630 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5633 = (inp[6]) ? 15'b000000000111111 : node5634;
													assign node5634 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node5638 = (inp[4]) ? node5658 : node5639;
											assign node5639 = (inp[2]) ? node5647 : node5640;
												assign node5640 = (inp[9]) ? 15'b000000011111111 : node5641;
													assign node5641 = (inp[1]) ? 15'b000000011111111 : node5642;
														assign node5642 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5647 = (inp[6]) ? node5651 : node5648;
													assign node5648 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5651 = (inp[14]) ? 15'b000000000011111 : node5652;
														assign node5652 = (inp[1]) ? node5654 : 15'b000000001111111;
															assign node5654 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5658 = (inp[14]) ? node5664 : node5659;
												assign node5659 = (inp[6]) ? 15'b000000000111111 : node5660;
													assign node5660 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5664 = (inp[6]) ? node5666 : 15'b000000000111111;
													assign node5666 = (inp[2]) ? node5670 : node5667;
														assign node5667 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
														assign node5670 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node5673 = (inp[2]) ? node5709 : node5674;
										assign node5674 = (inp[14]) ? node5692 : node5675;
											assign node5675 = (inp[1]) ? node5685 : node5676;
												assign node5676 = (inp[4]) ? node5680 : node5677;
													assign node5677 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5680 = (inp[13]) ? node5682 : 15'b000000011111111;
														assign node5682 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5685 = (inp[9]) ? node5689 : node5686;
													assign node5686 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5689 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5692 = (inp[4]) ? node5698 : node5693;
												assign node5693 = (inp[9]) ? node5695 : 15'b000000011111111;
													assign node5695 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5698 = (inp[1]) ? node5704 : node5699;
													assign node5699 = (inp[13]) ? 15'b000000000111111 : node5700;
														assign node5700 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5704 = (inp[9]) ? node5706 : 15'b000000000111111;
														assign node5706 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node5709 = (inp[1]) ? node5723 : node5710;
											assign node5710 = (inp[14]) ? node5718 : node5711;
												assign node5711 = (inp[13]) ? node5713 : 15'b000000001111111;
													assign node5713 = (inp[9]) ? node5715 : 15'b000000001111111;
														assign node5715 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5718 = (inp[13]) ? node5720 : 15'b000000000111111;
													assign node5720 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node5723 = (inp[9]) ? node5729 : node5724;
												assign node5724 = (inp[4]) ? node5726 : 15'b000000000111111;
													assign node5726 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5729 = (inp[13]) ? node5733 : node5730;
													assign node5730 = (inp[14]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node5733 = (inp[4]) ? 15'b000000000001111 : node5734;
														assign node5734 = (inp[14]) ? node5736 : 15'b000000000011111;
															assign node5736 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node5740 = (inp[5]) ? node5990 : node5741;
							assign node5741 = (inp[13]) ? node5851 : node5742;
								assign node5742 = (inp[6]) ? node5784 : node5743;
									assign node5743 = (inp[2]) ? node5761 : node5744;
										assign node5744 = (inp[0]) ? node5754 : node5745;
											assign node5745 = (inp[4]) ? node5751 : node5746;
												assign node5746 = (inp[8]) ? 15'b000001111111111 : node5747;
													assign node5747 = (inp[9]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node5751 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node5754 = (inp[1]) ? 15'b000000001111111 : node5755;
												assign node5755 = (inp[14]) ? 15'b000000111111111 : node5756;
													assign node5756 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node5761 = (inp[0]) ? node5773 : node5762;
											assign node5762 = (inp[8]) ? node5768 : node5763;
												assign node5763 = (inp[4]) ? 15'b000000111111111 : node5764;
													assign node5764 = (inp[14]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node5768 = (inp[1]) ? 15'b000000001111111 : node5769;
													assign node5769 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node5773 = (inp[9]) ? node5779 : node5774;
												assign node5774 = (inp[8]) ? node5776 : 15'b000000011111111;
													assign node5776 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5779 = (inp[1]) ? 15'b000000000111111 : node5780;
													assign node5780 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node5784 = (inp[8]) ? node5824 : node5785;
										assign node5785 = (inp[9]) ? node5805 : node5786;
											assign node5786 = (inp[0]) ? node5800 : node5787;
												assign node5787 = (inp[2]) ? node5793 : node5788;
													assign node5788 = (inp[4]) ? node5790 : 15'b000011111111111;
														assign node5790 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node5793 = (inp[4]) ? 15'b000000011111111 : node5794;
														assign node5794 = (inp[1]) ? 15'b000000111111111 : node5795;
															assign node5795 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node5800 = (inp[2]) ? node5802 : 15'b000000011111111;
													assign node5802 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5805 = (inp[4]) ? node5815 : node5806;
												assign node5806 = (inp[0]) ? 15'b000000011111111 : node5807;
													assign node5807 = (inp[14]) ? node5809 : 15'b000000011111111;
														assign node5809 = (inp[1]) ? node5811 : 15'b000000011111111;
															assign node5811 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5815 = (inp[0]) ? node5819 : node5816;
													assign node5816 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5819 = (inp[2]) ? node5821 : 15'b000000001111111;
														assign node5821 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5824 = (inp[1]) ? node5838 : node5825;
											assign node5825 = (inp[14]) ? node5829 : node5826;
												assign node5826 = (inp[9]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node5829 = (inp[4]) ? node5833 : node5830;
													assign node5830 = (inp[2]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node5833 = (inp[9]) ? node5835 : 15'b000000001111111;
														assign node5835 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5838 = (inp[2]) ? node5840 : 15'b000000001111111;
												assign node5840 = (inp[4]) ? node5846 : node5841;
													assign node5841 = (inp[0]) ? node5843 : 15'b000000000111111;
														assign node5843 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node5846 = (inp[9]) ? node5848 : 15'b000000000111111;
														assign node5848 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node5851 = (inp[14]) ? node5921 : node5852;
									assign node5852 = (inp[4]) ? node5892 : node5853;
										assign node5853 = (inp[0]) ? node5871 : node5854;
											assign node5854 = (inp[6]) ? node5862 : node5855;
												assign node5855 = (inp[9]) ? node5857 : 15'b000000111111111;
													assign node5857 = (inp[2]) ? 15'b000000011111111 : node5858;
														assign node5858 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5862 = (inp[2]) ? node5868 : node5863;
													assign node5863 = (inp[9]) ? 15'b000000011111111 : node5864;
														assign node5864 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node5868 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5871 = (inp[9]) ? node5879 : node5872;
												assign node5872 = (inp[1]) ? node5874 : 15'b000000011111111;
													assign node5874 = (inp[8]) ? node5876 : 15'b000000011111111;
														assign node5876 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5879 = (inp[2]) ? node5887 : node5880;
													assign node5880 = (inp[8]) ? node5882 : 15'b000000011111111;
														assign node5882 = (inp[6]) ? 15'b000000001111111 : node5883;
															assign node5883 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5887 = (inp[1]) ? node5889 : 15'b000000001111111;
														assign node5889 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node5892 = (inp[8]) ? node5906 : node5893;
											assign node5893 = (inp[6]) ? node5901 : node5894;
												assign node5894 = (inp[1]) ? node5898 : node5895;
													assign node5895 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node5898 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node5901 = (inp[2]) ? 15'b000000001111111 : node5902;
													assign node5902 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node5906 = (inp[2]) ? node5912 : node5907;
												assign node5907 = (inp[0]) ? node5909 : 15'b000000001111111;
													assign node5909 = (inp[9]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node5912 = (inp[0]) ? node5918 : node5913;
													assign node5913 = (inp[1]) ? 15'b000000000111111 : node5914;
														assign node5914 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5918 = (inp[6]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node5921 = (inp[2]) ? node5957 : node5922;
										assign node5922 = (inp[4]) ? node5938 : node5923;
											assign node5923 = (inp[6]) ? node5929 : node5924;
												assign node5924 = (inp[0]) ? 15'b000000001111111 : node5925;
													assign node5925 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node5929 = (inp[9]) ? node5933 : node5930;
													assign node5930 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5933 = (inp[1]) ? node5935 : 15'b000000001111111;
														assign node5935 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node5938 = (inp[1]) ? node5948 : node5939;
												assign node5939 = (inp[6]) ? node5945 : node5940;
													assign node5940 = (inp[0]) ? node5942 : 15'b000000111111111;
														assign node5942 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5945 = (inp[9]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node5948 = (inp[6]) ? node5954 : node5949;
													assign node5949 = (inp[8]) ? 15'b000000000111111 : node5950;
														assign node5950 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5954 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node5957 = (inp[6]) ? node5971 : node5958;
											assign node5958 = (inp[4]) ? node5966 : node5959;
												assign node5959 = (inp[1]) ? node5963 : node5960;
													assign node5960 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node5963 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node5966 = (inp[8]) ? 15'b000000000111111 : node5967;
													assign node5967 = (inp[1]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node5971 = (inp[8]) ? node5985 : node5972;
												assign node5972 = (inp[4]) ? node5980 : node5973;
													assign node5973 = (inp[1]) ? 15'b000000000111111 : node5974;
														assign node5974 = (inp[9]) ? node5976 : 15'b000000001111111;
															assign node5976 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node5980 = (inp[9]) ? node5982 : 15'b000000000111111;
														assign node5982 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node5985 = (inp[9]) ? 15'b000000000011111 : node5986;
													assign node5986 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node5990 = (inp[8]) ? node6104 : node5991;
								assign node5991 = (inp[14]) ? node6039 : node5992;
									assign node5992 = (inp[9]) ? node6012 : node5993;
										assign node5993 = (inp[2]) ? node6003 : node5994;
											assign node5994 = (inp[6]) ? node6000 : node5995;
												assign node5995 = (inp[1]) ? node5997 : 15'b000001111111111;
													assign node5997 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6000 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6003 = (inp[6]) ? node6007 : node6004;
												assign node6004 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6007 = (inp[0]) ? 15'b000000001111111 : node6008;
													assign node6008 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node6012 = (inp[1]) ? node6030 : node6013;
											assign node6013 = (inp[13]) ? node6021 : node6014;
												assign node6014 = (inp[0]) ? node6018 : node6015;
													assign node6015 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6018 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6021 = (inp[6]) ? node6027 : node6022;
													assign node6022 = (inp[2]) ? 15'b000000001111111 : node6023;
														assign node6023 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6027 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6030 = (inp[0]) ? node6032 : 15'b000000001111111;
												assign node6032 = (inp[6]) ? node6036 : node6033;
													assign node6033 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6036 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node6039 = (inp[6]) ? node6083 : node6040;
										assign node6040 = (inp[1]) ? node6064 : node6041;
											assign node6041 = (inp[0]) ? node6051 : node6042;
												assign node6042 = (inp[9]) ? node6046 : node6043;
													assign node6043 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6046 = (inp[4]) ? node6048 : 15'b000000011111111;
														assign node6048 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6051 = (inp[2]) ? node6059 : node6052;
													assign node6052 = (inp[4]) ? node6054 : 15'b000000011111111;
														assign node6054 = (inp[13]) ? 15'b000000001111111 : node6055;
															assign node6055 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6059 = (inp[9]) ? node6061 : 15'b000000001111111;
														assign node6061 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6064 = (inp[2]) ? node6072 : node6065;
												assign node6065 = (inp[13]) ? node6069 : node6066;
													assign node6066 = (inp[0]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node6069 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6072 = (inp[13]) ? node6078 : node6073;
													assign node6073 = (inp[4]) ? 15'b000000000111111 : node6074;
														assign node6074 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6078 = (inp[4]) ? 15'b000000000011111 : node6079;
														assign node6079 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6083 = (inp[0]) ? node6091 : node6084;
											assign node6084 = (inp[4]) ? node6086 : 15'b000000001111111;
												assign node6086 = (inp[13]) ? 15'b000000000111111 : node6087;
													assign node6087 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6091 = (inp[1]) ? node6099 : node6092;
												assign node6092 = (inp[9]) ? 15'b000000000011111 : node6093;
													assign node6093 = (inp[4]) ? node6095 : 15'b000000001111111;
														assign node6095 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6099 = (inp[2]) ? node6101 : 15'b000000000011111;
													assign node6101 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node6104 = (inp[2]) ? node6154 : node6105;
									assign node6105 = (inp[14]) ? node6129 : node6106;
										assign node6106 = (inp[1]) ? node6118 : node6107;
											assign node6107 = (inp[13]) ? node6111 : node6108;
												assign node6108 = (inp[6]) ? 15'b000000001111111 : 15'b000001111111111;
												assign node6111 = (inp[9]) ? node6115 : node6112;
													assign node6112 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6115 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6118 = (inp[6]) ? node6124 : node6119;
												assign node6119 = (inp[9]) ? node6121 : 15'b000000001111111;
													assign node6121 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6124 = (inp[9]) ? node6126 : 15'b000000000111111;
													assign node6126 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6129 = (inp[6]) ? node6143 : node6130;
											assign node6130 = (inp[9]) ? node6134 : node6131;
												assign node6131 = (inp[0]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node6134 = (inp[13]) ? node6140 : node6135;
													assign node6135 = (inp[1]) ? 15'b000000000111111 : node6136;
														assign node6136 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6140 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node6143 = (inp[13]) ? node6149 : node6144;
												assign node6144 = (inp[0]) ? node6146 : 15'b000000000111111;
													assign node6146 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6149 = (inp[4]) ? node6151 : 15'b000000000011111;
													assign node6151 = (inp[9]) ? 15'b000000000000111 : 15'b000000000011111;
									assign node6154 = (inp[9]) ? node6186 : node6155;
										assign node6155 = (inp[6]) ? node6167 : node6156;
											assign node6156 = (inp[13]) ? node6162 : node6157;
												assign node6157 = (inp[14]) ? node6159 : 15'b000000001111111;
													assign node6159 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6162 = (inp[4]) ? 15'b000000000111111 : node6163;
													assign node6163 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node6167 = (inp[4]) ? node6177 : node6168;
												assign node6168 = (inp[1]) ? node6170 : 15'b000000001111111;
													assign node6170 = (inp[13]) ? 15'b000000000011111 : node6171;
														assign node6171 = (inp[0]) ? node6173 : 15'b000000000111111;
															assign node6173 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6177 = (inp[0]) ? node6181 : node6178;
													assign node6178 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node6181 = (inp[13]) ? node6183 : 15'b000000000011111;
														assign node6183 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node6186 = (inp[6]) ? node6200 : node6187;
											assign node6187 = (inp[4]) ? 15'b000000000011111 : node6188;
												assign node6188 = (inp[1]) ? node6194 : node6189;
													assign node6189 = (inp[0]) ? 15'b000000000111111 : node6190;
														assign node6190 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6194 = (inp[14]) ? node6196 : 15'b000000000111111;
														assign node6196 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node6200 = (inp[0]) ? node6210 : node6201;
												assign node6201 = (inp[14]) ? node6207 : node6202;
													assign node6202 = (inp[4]) ? 15'b000000000011111 : node6203;
														assign node6203 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node6207 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node6210 = (inp[14]) ? node6214 : node6211;
													assign node6211 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node6214 = (inp[1]) ? node6216 : 15'b000000000001111;
														assign node6216 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
				assign node6219 = (inp[14]) ? node7233 : node6220;
					assign node6220 = (inp[2]) ? node6708 : node6221;
						assign node6221 = (inp[13]) ? node6447 : node6222;
							assign node6222 = (inp[4]) ? node6326 : node6223;
								assign node6223 = (inp[6]) ? node6273 : node6224;
									assign node6224 = (inp[1]) ? node6248 : node6225;
										assign node6225 = (inp[8]) ? node6237 : node6226;
											assign node6226 = (inp[5]) ? node6228 : 15'b000011111111111;
												assign node6228 = (inp[9]) ? node6234 : node6229;
													assign node6229 = (inp[10]) ? 15'b000001111111111 : node6230;
														assign node6230 = (inp[3]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node6234 = (inp[0]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node6237 = (inp[9]) ? node6243 : node6238;
												assign node6238 = (inp[5]) ? 15'b000001111111111 : node6239;
													assign node6239 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node6243 = (inp[10]) ? node6245 : 15'b000000111111111;
													assign node6245 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node6248 = (inp[0]) ? node6260 : node6249;
											assign node6249 = (inp[3]) ? node6253 : node6250;
												assign node6250 = (inp[8]) ? 15'b000001111111111 : 15'b000111111111111;
												assign node6253 = (inp[9]) ? node6257 : node6254;
													assign node6254 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6257 = (inp[10]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node6260 = (inp[3]) ? node6262 : 15'b000000111111111;
												assign node6262 = (inp[8]) ? node6270 : node6263;
													assign node6263 = (inp[9]) ? 15'b000000011111111 : node6264;
														assign node6264 = (inp[5]) ? node6266 : 15'b000000111111111;
															assign node6266 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6270 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node6273 = (inp[5]) ? node6295 : node6274;
										assign node6274 = (inp[10]) ? node6282 : node6275;
											assign node6275 = (inp[0]) ? node6277 : 15'b000001111111111;
												assign node6277 = (inp[8]) ? 15'b000000111111111 : node6278;
													assign node6278 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6282 = (inp[8]) ? node6286 : node6283;
												assign node6283 = (inp[3]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node6286 = (inp[9]) ? 15'b000000011111111 : node6287;
													assign node6287 = (inp[1]) ? node6289 : 15'b000000111111111;
														assign node6289 = (inp[3]) ? 15'b000000011111111 : node6290;
															assign node6290 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node6295 = (inp[3]) ? node6311 : node6296;
											assign node6296 = (inp[8]) ? node6302 : node6297;
												assign node6297 = (inp[10]) ? 15'b000000111111111 : node6298;
													assign node6298 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6302 = (inp[0]) ? node6306 : node6303;
													assign node6303 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6306 = (inp[9]) ? node6308 : 15'b000000011111111;
														assign node6308 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6311 = (inp[0]) ? node6319 : node6312;
												assign node6312 = (inp[9]) ? node6314 : 15'b000000011111111;
													assign node6314 = (inp[10]) ? node6316 : 15'b000000011111111;
														assign node6316 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6319 = (inp[1]) ? 15'b000000001111111 : node6320;
													assign node6320 = (inp[10]) ? node6322 : 15'b000000011111111;
														assign node6322 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node6326 = (inp[9]) ? node6402 : node6327;
									assign node6327 = (inp[5]) ? node6375 : node6328;
										assign node6328 = (inp[10]) ? node6356 : node6329;
											assign node6329 = (inp[0]) ? node6343 : node6330;
												assign node6330 = (inp[1]) ? node6336 : node6331;
													assign node6331 = (inp[6]) ? node6333 : 15'b000011111111111;
														assign node6333 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6336 = (inp[3]) ? 15'b000000111111111 : node6337;
														assign node6337 = (inp[6]) ? node6339 : 15'b000001111111111;
															assign node6339 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6343 = (inp[3]) ? node6353 : node6344;
													assign node6344 = (inp[1]) ? node6350 : node6345;
														assign node6345 = (inp[6]) ? node6347 : 15'b000001111111111;
															assign node6347 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node6350 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6353 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6356 = (inp[6]) ? node6366 : node6357;
												assign node6357 = (inp[1]) ? node6361 : node6358;
													assign node6358 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6361 = (inp[0]) ? node6363 : 15'b000000111111111;
														assign node6363 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6366 = (inp[3]) ? node6368 : 15'b000000111111111;
													assign node6368 = (inp[0]) ? 15'b000000001111111 : node6369;
														assign node6369 = (inp[8]) ? node6371 : 15'b000000011111111;
															assign node6371 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6375 = (inp[1]) ? node6389 : node6376;
											assign node6376 = (inp[0]) ? node6384 : node6377;
												assign node6377 = (inp[6]) ? node6381 : node6378;
													assign node6378 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6381 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6384 = (inp[8]) ? node6386 : 15'b000000111111111;
													assign node6386 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6389 = (inp[0]) ? node6395 : node6390;
												assign node6390 = (inp[10]) ? 15'b000000001111111 : node6391;
													assign node6391 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6395 = (inp[10]) ? node6397 : 15'b000000001111111;
													assign node6397 = (inp[3]) ? 15'b000000000111111 : node6398;
														assign node6398 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node6402 = (inp[3]) ? node6420 : node6403;
										assign node6403 = (inp[6]) ? node6411 : node6404;
											assign node6404 = (inp[10]) ? node6406 : 15'b000000111111111;
												assign node6406 = (inp[1]) ? node6408 : 15'b000000111111111;
													assign node6408 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6411 = (inp[10]) ? node6413 : 15'b000000011111111;
												assign node6413 = (inp[5]) ? 15'b000000001111111 : node6414;
													assign node6414 = (inp[0]) ? 15'b000000001111111 : node6415;
														assign node6415 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6420 = (inp[10]) ? node6432 : node6421;
											assign node6421 = (inp[1]) ? node6427 : node6422;
												assign node6422 = (inp[6]) ? node6424 : 15'b000000011111111;
													assign node6424 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6427 = (inp[0]) ? 15'b000000001111111 : node6428;
													assign node6428 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6432 = (inp[0]) ? node6442 : node6433;
												assign node6433 = (inp[8]) ? node6435 : 15'b000000111111111;
													assign node6435 = (inp[6]) ? node6437 : 15'b000000001111111;
														assign node6437 = (inp[1]) ? 15'b000000000111111 : node6438;
															assign node6438 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6442 = (inp[8]) ? 15'b000000000111111 : node6443;
													assign node6443 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node6447 = (inp[10]) ? node6593 : node6448;
								assign node6448 = (inp[9]) ? node6516 : node6449;
									assign node6449 = (inp[4]) ? node6487 : node6450;
										assign node6450 = (inp[0]) ? node6472 : node6451;
											assign node6451 = (inp[3]) ? node6467 : node6452;
												assign node6452 = (inp[6]) ? node6456 : node6453;
													assign node6453 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node6456 = (inp[5]) ? node6462 : node6457;
														assign node6457 = (inp[8]) ? node6459 : 15'b000001111111111;
															assign node6459 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node6462 = (inp[8]) ? 15'b000000111111111 : node6463;
															assign node6463 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6467 = (inp[5]) ? 15'b000000111111111 : node6468;
													assign node6468 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node6472 = (inp[6]) ? node6482 : node6473;
												assign node6473 = (inp[8]) ? node6479 : node6474;
													assign node6474 = (inp[3]) ? 15'b000000111111111 : node6475;
														assign node6475 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6479 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6482 = (inp[1]) ? node6484 : 15'b000000111111111;
													assign node6484 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6487 = (inp[3]) ? node6501 : node6488;
											assign node6488 = (inp[1]) ? node6496 : node6489;
												assign node6489 = (inp[8]) ? node6493 : node6490;
													assign node6490 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6493 = (inp[0]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node6496 = (inp[6]) ? node6498 : 15'b000000011111111;
													assign node6498 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6501 = (inp[1]) ? node6511 : node6502;
												assign node6502 = (inp[6]) ? node6506 : node6503;
													assign node6503 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6506 = (inp[0]) ? 15'b000000000111111 : node6507;
														assign node6507 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6511 = (inp[5]) ? 15'b000000001111111 : node6512;
													assign node6512 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node6516 = (inp[0]) ? node6564 : node6517;
										assign node6517 = (inp[3]) ? node6539 : node6518;
											assign node6518 = (inp[1]) ? node6526 : node6519;
												assign node6519 = (inp[5]) ? 15'b000000111111111 : node6520;
													assign node6520 = (inp[8]) ? node6522 : 15'b000011111111111;
														assign node6522 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6526 = (inp[5]) ? node6532 : node6527;
													assign node6527 = (inp[8]) ? node6529 : 15'b000000111111111;
														assign node6529 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6532 = (inp[8]) ? node6534 : 15'b000000011111111;
														assign node6534 = (inp[4]) ? 15'b000000001111111 : node6535;
															assign node6535 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6539 = (inp[5]) ? node6551 : node6540;
												assign node6540 = (inp[8]) ? node6546 : node6541;
													assign node6541 = (inp[1]) ? node6543 : 15'b000000111111111;
														assign node6543 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6546 = (inp[4]) ? node6548 : 15'b000000011111111;
														assign node6548 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6551 = (inp[8]) ? node6559 : node6552;
													assign node6552 = (inp[4]) ? 15'b000000001111111 : node6553;
														assign node6553 = (inp[6]) ? node6555 : 15'b000000011111111;
															assign node6555 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6559 = (inp[6]) ? node6561 : 15'b000000001111111;
														assign node6561 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node6564 = (inp[1]) ? node6578 : node6565;
											assign node6565 = (inp[3]) ? node6569 : node6566;
												assign node6566 = (inp[8]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node6569 = (inp[5]) ? 15'b000000001111111 : node6570;
													assign node6570 = (inp[6]) ? 15'b000000001111111 : node6571;
														assign node6571 = (inp[8]) ? node6573 : 15'b000000011111111;
															assign node6573 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6578 = (inp[5]) ? node6590 : node6579;
												assign node6579 = (inp[6]) ? node6585 : node6580;
													assign node6580 = (inp[3]) ? 15'b000000001111111 : node6581;
														assign node6581 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6585 = (inp[3]) ? 15'b000000000111111 : node6586;
														assign node6586 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6590 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node6593 = (inp[0]) ? node6663 : node6594;
									assign node6594 = (inp[9]) ? node6632 : node6595;
										assign node6595 = (inp[1]) ? node6611 : node6596;
											assign node6596 = (inp[8]) ? node6602 : node6597;
												assign node6597 = (inp[6]) ? node6599 : 15'b000001111111111;
													assign node6599 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node6602 = (inp[6]) ? node6608 : node6603;
													assign node6603 = (inp[5]) ? 15'b000000011111111 : node6604;
														assign node6604 = (inp[4]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6608 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6611 = (inp[8]) ? node6623 : node6612;
												assign node6612 = (inp[3]) ? node6614 : 15'b000000011111111;
													assign node6614 = (inp[4]) ? node6620 : node6615;
														assign node6615 = (inp[5]) ? node6617 : 15'b000000011111111;
															assign node6617 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node6620 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6623 = (inp[5]) ? node6627 : node6624;
													assign node6624 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node6627 = (inp[6]) ? node6629 : 15'b000000001111111;
														assign node6629 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6632 = (inp[3]) ? node6650 : node6633;
											assign node6633 = (inp[4]) ? node6641 : node6634;
												assign node6634 = (inp[6]) ? 15'b000000001111111 : node6635;
													assign node6635 = (inp[5]) ? node6637 : 15'b000000011111111;
														assign node6637 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6641 = (inp[8]) ? node6647 : node6642;
													assign node6642 = (inp[5]) ? 15'b000000001111111 : node6643;
														assign node6643 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6647 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6650 = (inp[4]) ? node6652 : 15'b000000001111111;
												assign node6652 = (inp[5]) ? 15'b000000000011111 : node6653;
													assign node6653 = (inp[8]) ? node6657 : node6654;
														assign node6654 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node6657 = (inp[6]) ? node6659 : 15'b000000000111111;
															assign node6659 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node6663 = (inp[5]) ? node6683 : node6664;
										assign node6664 = (inp[4]) ? node6678 : node6665;
											assign node6665 = (inp[3]) ? node6673 : node6666;
												assign node6666 = (inp[8]) ? node6670 : node6667;
													assign node6667 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6670 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6673 = (inp[8]) ? 15'b000000000111111 : node6674;
													assign node6674 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6678 = (inp[9]) ? 15'b000000000001111 : node6679;
												assign node6679 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6683 = (inp[8]) ? node6695 : node6684;
											assign node6684 = (inp[3]) ? node6690 : node6685;
												assign node6685 = (inp[1]) ? 15'b000000000111111 : node6686;
													assign node6686 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6690 = (inp[6]) ? node6692 : 15'b000000000111111;
													assign node6692 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node6695 = (inp[1]) ? node6703 : node6696;
												assign node6696 = (inp[4]) ? node6700 : node6697;
													assign node6697 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6700 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6703 = (inp[4]) ? 15'b000000000001111 : node6704;
													assign node6704 = (inp[3]) ? 15'b000000000001111 : 15'b000000000111111;
						assign node6708 = (inp[4]) ? node6974 : node6709;
							assign node6709 = (inp[13]) ? node6823 : node6710;
								assign node6710 = (inp[3]) ? node6774 : node6711;
									assign node6711 = (inp[9]) ? node6741 : node6712;
										assign node6712 = (inp[6]) ? node6734 : node6713;
											assign node6713 = (inp[0]) ? node6723 : node6714;
												assign node6714 = (inp[10]) ? node6720 : node6715;
													assign node6715 = (inp[1]) ? node6717 : 15'b000011111111111;
														assign node6717 = (inp[5]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node6720 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6723 = (inp[1]) ? node6731 : node6724;
													assign node6724 = (inp[5]) ? 15'b000000111111111 : node6725;
														assign node6725 = (inp[8]) ? node6727 : 15'b000001111111111;
															assign node6727 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6731 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6734 = (inp[8]) ? 15'b000000011111111 : node6735;
												assign node6735 = (inp[0]) ? node6737 : 15'b000001111111111;
													assign node6737 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node6741 = (inp[1]) ? node6763 : node6742;
											assign node6742 = (inp[10]) ? node6754 : node6743;
												assign node6743 = (inp[8]) ? node6749 : node6744;
													assign node6744 = (inp[5]) ? node6746 : 15'b000001111111111;
														assign node6746 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6749 = (inp[6]) ? node6751 : 15'b000000111111111;
														assign node6751 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6754 = (inp[0]) ? 15'b000000011111111 : node6755;
													assign node6755 = (inp[6]) ? node6757 : 15'b000000111111111;
														assign node6757 = (inp[5]) ? 15'b000000011111111 : node6758;
															assign node6758 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6763 = (inp[10]) ? node6769 : node6764;
												assign node6764 = (inp[5]) ? node6766 : 15'b000000011111111;
													assign node6766 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6769 = (inp[0]) ? 15'b000000001111111 : node6770;
													assign node6770 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node6774 = (inp[5]) ? node6796 : node6775;
										assign node6775 = (inp[1]) ? node6789 : node6776;
											assign node6776 = (inp[10]) ? node6784 : node6777;
												assign node6777 = (inp[0]) ? 15'b000000111111111 : node6778;
													assign node6778 = (inp[6]) ? node6780 : 15'b000001111111111;
														assign node6780 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6784 = (inp[0]) ? 15'b000000001111111 : node6785;
													assign node6785 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6789 = (inp[0]) ? 15'b000000001111111 : node6790;
												assign node6790 = (inp[9]) ? node6792 : 15'b000000011111111;
													assign node6792 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node6796 = (inp[0]) ? node6810 : node6797;
											assign node6797 = (inp[6]) ? node6805 : node6798;
												assign node6798 = (inp[1]) ? node6802 : node6799;
													assign node6799 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6802 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6805 = (inp[10]) ? node6807 : 15'b000000001111111;
													assign node6807 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6810 = (inp[8]) ? node6812 : 15'b000000001111111;
												assign node6812 = (inp[1]) ? node6816 : node6813;
													assign node6813 = (inp[9]) ? 15'b000000001111111 : 15'b000000000111111;
													assign node6816 = (inp[10]) ? 15'b000000000011111 : node6817;
														assign node6817 = (inp[9]) ? node6819 : 15'b000000000111111;
															assign node6819 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node6823 = (inp[10]) ? node6897 : node6824;
									assign node6824 = (inp[0]) ? node6862 : node6825;
										assign node6825 = (inp[8]) ? node6841 : node6826;
											assign node6826 = (inp[3]) ? node6836 : node6827;
												assign node6827 = (inp[5]) ? node6831 : node6828;
													assign node6828 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node6831 = (inp[9]) ? 15'b000000011111111 : node6832;
														assign node6832 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node6836 = (inp[1]) ? 15'b000000011111111 : node6837;
													assign node6837 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node6841 = (inp[9]) ? node6855 : node6842;
												assign node6842 = (inp[3]) ? node6850 : node6843;
													assign node6843 = (inp[1]) ? node6845 : 15'b000000011111111;
														assign node6845 = (inp[5]) ? node6847 : 15'b000000011111111;
															assign node6847 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6850 = (inp[1]) ? 15'b000000011111111 : node6851;
														assign node6851 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6855 = (inp[6]) ? node6857 : 15'b000000011111111;
													assign node6857 = (inp[1]) ? node6859 : 15'b000000001111111;
														assign node6859 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node6862 = (inp[9]) ? node6880 : node6863;
											assign node6863 = (inp[1]) ? node6871 : node6864;
												assign node6864 = (inp[3]) ? node6866 : 15'b000000011111111;
													assign node6866 = (inp[5]) ? 15'b000000001111111 : node6867;
														assign node6867 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6871 = (inp[6]) ? node6877 : node6872;
													assign node6872 = (inp[8]) ? 15'b000000001111111 : node6873;
														assign node6873 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6877 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6880 = (inp[3]) ? node6892 : node6881;
												assign node6881 = (inp[1]) ? node6885 : node6882;
													assign node6882 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6885 = (inp[8]) ? 15'b000000000111111 : node6886;
														assign node6886 = (inp[6]) ? node6888 : 15'b000000001111111;
															assign node6888 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6892 = (inp[1]) ? 15'b000000000011111 : node6893;
													assign node6893 = (inp[6]) ? 15'b000000000111111 : 15'b000000011111111;
									assign node6897 = (inp[1]) ? node6939 : node6898;
										assign node6898 = (inp[8]) ? node6918 : node6899;
											assign node6899 = (inp[3]) ? node6911 : node6900;
												assign node6900 = (inp[6]) ? node6908 : node6901;
													assign node6901 = (inp[9]) ? 15'b000000011111111 : node6902;
														assign node6902 = (inp[5]) ? node6904 : 15'b000000111111111;
															assign node6904 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6908 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node6911 = (inp[5]) ? node6915 : node6912;
													assign node6912 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6915 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node6918 = (inp[5]) ? node6928 : node6919;
												assign node6919 = (inp[0]) ? node6925 : node6920;
													assign node6920 = (inp[9]) ? 15'b000000001111111 : node6921;
														assign node6921 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6925 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6928 = (inp[3]) ? node6934 : node6929;
													assign node6929 = (inp[0]) ? 15'b000000000111111 : node6930;
														assign node6930 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6934 = (inp[6]) ? node6936 : 15'b000000000111111;
														assign node6936 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node6939 = (inp[8]) ? node6965 : node6940;
											assign node6940 = (inp[3]) ? node6952 : node6941;
												assign node6941 = (inp[6]) ? node6945 : node6942;
													assign node6942 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node6945 = (inp[0]) ? 15'b000000000011111 : node6946;
														assign node6946 = (inp[5]) ? node6948 : 15'b000000001111111;
															assign node6948 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node6952 = (inp[9]) ? node6958 : node6953;
													assign node6953 = (inp[5]) ? 15'b000000000111111 : node6954;
														assign node6954 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node6958 = (inp[0]) ? 15'b000000000001111 : node6959;
														assign node6959 = (inp[5]) ? node6961 : 15'b000000000111111;
															assign node6961 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node6965 = (inp[5]) ? node6971 : node6966;
												assign node6966 = (inp[3]) ? node6968 : 15'b000000000111111;
													assign node6968 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node6971 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node6974 = (inp[10]) ? node7108 : node6975;
								assign node6975 = (inp[6]) ? node7051 : node6976;
									assign node6976 = (inp[5]) ? node7018 : node6977;
										assign node6977 = (inp[0]) ? node6997 : node6978;
											assign node6978 = (inp[13]) ? node6988 : node6979;
												assign node6979 = (inp[3]) ? node6981 : 15'b000001111111111;
													assign node6981 = (inp[9]) ? node6983 : 15'b000000111111111;
														assign node6983 = (inp[1]) ? 15'b000000011111111 : node6984;
															assign node6984 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node6988 = (inp[3]) ? node6994 : node6989;
													assign node6989 = (inp[1]) ? 15'b000000011111111 : node6990;
														assign node6990 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node6994 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node6997 = (inp[9]) ? node7007 : node6998;
												assign node6998 = (inp[1]) ? node7002 : node6999;
													assign node6999 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7002 = (inp[8]) ? node7004 : 15'b000000011111111;
														assign node7004 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7007 = (inp[3]) ? node7015 : node7008;
													assign node7008 = (inp[13]) ? 15'b000000001111111 : node7009;
														assign node7009 = (inp[8]) ? node7011 : 15'b000000011111111;
															assign node7011 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7015 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7018 = (inp[0]) ? node7034 : node7019;
											assign node7019 = (inp[9]) ? node7027 : node7020;
												assign node7020 = (inp[8]) ? node7022 : 15'b000000111111111;
													assign node7022 = (inp[3]) ? node7024 : 15'b000000011111111;
														assign node7024 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7027 = (inp[3]) ? 15'b000000000111111 : node7028;
													assign node7028 = (inp[13]) ? 15'b000000001111111 : node7029;
														assign node7029 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7034 = (inp[1]) ? node7042 : node7035;
												assign node7035 = (inp[8]) ? node7039 : node7036;
													assign node7036 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7039 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7042 = (inp[3]) ? node7046 : node7043;
													assign node7043 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7046 = (inp[9]) ? node7048 : 15'b000000000111111;
														assign node7048 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node7051 = (inp[8]) ? node7083 : node7052;
										assign node7052 = (inp[1]) ? node7066 : node7053;
											assign node7053 = (inp[13]) ? node7059 : node7054;
												assign node7054 = (inp[0]) ? 15'b000000011111111 : node7055;
													assign node7055 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7059 = (inp[5]) ? node7063 : node7060;
													assign node7060 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7063 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7066 = (inp[13]) ? node7072 : node7067;
												assign node7067 = (inp[5]) ? node7069 : 15'b000000001111111;
													assign node7069 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7072 = (inp[0]) ? node7080 : node7073;
													assign node7073 = (inp[3]) ? node7075 : 15'b000000011111111;
														assign node7075 = (inp[9]) ? 15'b000000000111111 : node7076;
															assign node7076 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7080 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7083 = (inp[9]) ? node7093 : node7084;
											assign node7084 = (inp[5]) ? node7088 : node7085;
												assign node7085 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node7088 = (inp[13]) ? 15'b000000000111111 : node7089;
													assign node7089 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7093 = (inp[3]) ? node7099 : node7094;
												assign node7094 = (inp[13]) ? node7096 : 15'b000000000111111;
													assign node7096 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7099 = (inp[0]) ? node7101 : 15'b000000000111111;
													assign node7101 = (inp[5]) ? node7103 : 15'b000000000011111;
														assign node7103 = (inp[13]) ? 15'b000000000001111 : node7104;
															assign node7104 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node7108 = (inp[8]) ? node7168 : node7109;
									assign node7109 = (inp[1]) ? node7137 : node7110;
										assign node7110 = (inp[6]) ? node7124 : node7111;
											assign node7111 = (inp[5]) ? node7117 : node7112;
												assign node7112 = (inp[3]) ? 15'b000000001111111 : node7113;
													assign node7113 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7117 = (inp[13]) ? node7121 : node7118;
													assign node7118 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7121 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7124 = (inp[0]) ? node7130 : node7125;
												assign node7125 = (inp[13]) ? node7127 : 15'b000000011111111;
													assign node7127 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7130 = (inp[9]) ? 15'b000000000011111 : node7131;
													assign node7131 = (inp[13]) ? 15'b000000000111111 : node7132;
														assign node7132 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7137 = (inp[5]) ? node7157 : node7138;
											assign node7138 = (inp[13]) ? node7146 : node7139;
												assign node7139 = (inp[3]) ? 15'b000000001111111 : node7140;
													assign node7140 = (inp[0]) ? node7142 : 15'b000000011111111;
														assign node7142 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7146 = (inp[9]) ? node7154 : node7147;
													assign node7147 = (inp[3]) ? 15'b000000000111111 : node7148;
														assign node7148 = (inp[0]) ? node7150 : 15'b000000001111111;
															assign node7150 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7154 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7157 = (inp[13]) ? 15'b000000000011111 : node7158;
												assign node7158 = (inp[3]) ? node7160 : 15'b000000000111111;
													assign node7160 = (inp[0]) ? node7164 : node7161;
														assign node7161 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
														assign node7164 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7168 = (inp[13]) ? node7202 : node7169;
										assign node7169 = (inp[6]) ? node7187 : node7170;
											assign node7170 = (inp[3]) ? node7176 : node7171;
												assign node7171 = (inp[5]) ? 15'b000000001111111 : node7172;
													assign node7172 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7176 = (inp[1]) ? node7184 : node7177;
													assign node7177 = (inp[0]) ? 15'b000000000111111 : node7178;
														assign node7178 = (inp[5]) ? node7180 : 15'b000000011111111;
															assign node7180 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7184 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7187 = (inp[1]) ? node7197 : node7188;
												assign node7188 = (inp[9]) ? node7192 : node7189;
													assign node7189 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7192 = (inp[3]) ? node7194 : 15'b000000000111111;
														assign node7194 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7197 = (inp[5]) ? 15'b000000000011111 : node7198;
													assign node7198 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7202 = (inp[3]) ? node7218 : node7203;
											assign node7203 = (inp[0]) ? node7211 : node7204;
												assign node7204 = (inp[9]) ? node7206 : 15'b000000000111111;
													assign node7206 = (inp[1]) ? node7208 : 15'b000000000111111;
														assign node7208 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7211 = (inp[5]) ? node7215 : node7212;
													assign node7212 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7215 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7218 = (inp[0]) ? node7226 : node7219;
												assign node7219 = (inp[9]) ? node7221 : 15'b000000000011111;
													assign node7221 = (inp[1]) ? node7223 : 15'b000000000011111;
														assign node7223 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7226 = (inp[1]) ? node7230 : node7227;
													assign node7227 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node7230 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
					assign node7233 = (inp[9]) ? node7739 : node7234;
						assign node7234 = (inp[6]) ? node7482 : node7235;
							assign node7235 = (inp[0]) ? node7363 : node7236;
								assign node7236 = (inp[2]) ? node7304 : node7237;
									assign node7237 = (inp[4]) ? node7277 : node7238;
										assign node7238 = (inp[8]) ? node7258 : node7239;
											assign node7239 = (inp[3]) ? node7251 : node7240;
												assign node7240 = (inp[10]) ? node7246 : node7241;
													assign node7241 = (inp[1]) ? node7243 : 15'b000011111111111;
														assign node7243 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node7246 = (inp[5]) ? 15'b000001111111111 : node7247;
														assign node7247 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node7251 = (inp[13]) ? node7253 : 15'b000011111111111;
													assign node7253 = (inp[5]) ? node7255 : 15'b000000111111111;
														assign node7255 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7258 = (inp[1]) ? node7268 : node7259;
												assign node7259 = (inp[13]) ? 15'b000000111111111 : node7260;
													assign node7260 = (inp[3]) ? node7262 : 15'b000001111111111;
														assign node7262 = (inp[10]) ? 15'b000000111111111 : node7263;
															assign node7263 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7268 = (inp[3]) ? 15'b000000001111111 : node7269;
													assign node7269 = (inp[13]) ? 15'b000000011111111 : node7270;
														assign node7270 = (inp[10]) ? node7272 : 15'b000001111111111;
															assign node7272 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node7277 = (inp[13]) ? node7299 : node7278;
											assign node7278 = (inp[8]) ? node7284 : node7279;
												assign node7279 = (inp[10]) ? node7281 : 15'b000000111111111;
													assign node7281 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7284 = (inp[1]) ? node7292 : node7285;
													assign node7285 = (inp[3]) ? 15'b000000011111111 : node7286;
														assign node7286 = (inp[5]) ? node7288 : 15'b000000111111111;
															assign node7288 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7292 = (inp[3]) ? 15'b000000001111111 : node7293;
														assign node7293 = (inp[5]) ? node7295 : 15'b000000011111111;
															assign node7295 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7299 = (inp[10]) ? 15'b000000000111111 : node7300;
												assign node7300 = (inp[3]) ? 15'b000000011111111 : 15'b000000001111111;
									assign node7304 = (inp[10]) ? node7344 : node7305;
										assign node7305 = (inp[5]) ? node7319 : node7306;
											assign node7306 = (inp[4]) ? node7310 : node7307;
												assign node7307 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7310 = (inp[1]) ? 15'b000000011111111 : node7311;
													assign node7311 = (inp[13]) ? node7313 : 15'b000000111111111;
														assign node7313 = (inp[3]) ? 15'b000000011111111 : node7314;
															assign node7314 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7319 = (inp[13]) ? node7333 : node7320;
												assign node7320 = (inp[8]) ? node7326 : node7321;
													assign node7321 = (inp[3]) ? node7323 : 15'b000000111111111;
														assign node7323 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7326 = (inp[4]) ? 15'b000000001111111 : node7327;
														assign node7327 = (inp[1]) ? 15'b000000011111111 : node7328;
															assign node7328 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7333 = (inp[3]) ? node7337 : node7334;
													assign node7334 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7337 = (inp[4]) ? node7339 : 15'b000000001111111;
														assign node7339 = (inp[1]) ? node7341 : 15'b000000000111111;
															assign node7341 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7344 = (inp[8]) ? node7360 : node7345;
											assign node7345 = (inp[1]) ? node7347 : 15'b000000011111111;
												assign node7347 = (inp[3]) ? node7353 : node7348;
													assign node7348 = (inp[13]) ? node7350 : 15'b000000011111111;
														assign node7350 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7353 = (inp[5]) ? 15'b000000000111111 : node7354;
														assign node7354 = (inp[4]) ? 15'b000000001111111 : node7355;
															assign node7355 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7360 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node7363 = (inp[5]) ? node7427 : node7364;
									assign node7364 = (inp[4]) ? node7400 : node7365;
										assign node7365 = (inp[1]) ? node7387 : node7366;
											assign node7366 = (inp[8]) ? node7376 : node7367;
												assign node7367 = (inp[2]) ? node7373 : node7368;
													assign node7368 = (inp[3]) ? 15'b000000111111111 : node7369;
														assign node7369 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node7373 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7376 = (inp[3]) ? node7382 : node7377;
													assign node7377 = (inp[13]) ? node7379 : 15'b000000111111111;
														assign node7379 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7382 = (inp[2]) ? node7384 : 15'b000000011111111;
														assign node7384 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7387 = (inp[10]) ? node7395 : node7388;
												assign node7388 = (inp[2]) ? node7392 : node7389;
													assign node7389 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7392 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7395 = (inp[13]) ? 15'b000000000111111 : node7396;
													assign node7396 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node7400 = (inp[8]) ? node7416 : node7401;
											assign node7401 = (inp[10]) ? node7411 : node7402;
												assign node7402 = (inp[1]) ? 15'b000000001111111 : node7403;
													assign node7403 = (inp[13]) ? node7405 : 15'b000000111111111;
														assign node7405 = (inp[3]) ? node7407 : 15'b000000011111111;
															assign node7407 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7411 = (inp[13]) ? node7413 : 15'b000000011111111;
													assign node7413 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7416 = (inp[2]) ? node7422 : node7417;
												assign node7417 = (inp[10]) ? node7419 : 15'b000000001111111;
													assign node7419 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node7422 = (inp[13]) ? node7424 : 15'b000000000111111;
													assign node7424 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7427 = (inp[8]) ? node7455 : node7428;
										assign node7428 = (inp[1]) ? node7438 : node7429;
											assign node7429 = (inp[10]) ? node7431 : 15'b000000011111111;
												assign node7431 = (inp[3]) ? node7435 : node7432;
													assign node7432 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7435 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7438 = (inp[13]) ? node7448 : node7439;
												assign node7439 = (inp[2]) ? node7441 : 15'b000000011111111;
													assign node7441 = (inp[3]) ? node7443 : 15'b000000001111111;
														assign node7443 = (inp[10]) ? 15'b000000000111111 : node7444;
															assign node7444 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7448 = (inp[4]) ? 15'b000000000111111 : node7449;
													assign node7449 = (inp[3]) ? 15'b000000000111111 : node7450;
														assign node7450 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7455 = (inp[2]) ? node7469 : node7456;
											assign node7456 = (inp[4]) ? node7466 : node7457;
												assign node7457 = (inp[10]) ? node7461 : node7458;
													assign node7458 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7461 = (inp[1]) ? 15'b000000000111111 : node7462;
														assign node7462 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7466 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7469 = (inp[3]) ? node7477 : node7470;
												assign node7470 = (inp[13]) ? node7472 : 15'b000000000111111;
													assign node7472 = (inp[10]) ? node7474 : 15'b000000000111111;
														assign node7474 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7477 = (inp[1]) ? node7479 : 15'b000000000011111;
													assign node7479 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node7482 = (inp[1]) ? node7608 : node7483;
								assign node7483 = (inp[13]) ? node7551 : node7484;
									assign node7484 = (inp[8]) ? node7528 : node7485;
										assign node7485 = (inp[4]) ? node7501 : node7486;
											assign node7486 = (inp[2]) ? node7492 : node7487;
												assign node7487 = (inp[10]) ? 15'b000000111111111 : node7488;
													assign node7488 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7492 = (inp[0]) ? node7494 : 15'b000000111111111;
													assign node7494 = (inp[10]) ? 15'b000000011111111 : node7495;
														assign node7495 = (inp[5]) ? 15'b000000011111111 : node7496;
															assign node7496 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node7501 = (inp[0]) ? node7517 : node7502;
												assign node7502 = (inp[3]) ? node7510 : node7503;
													assign node7503 = (inp[5]) ? 15'b000000011111111 : node7504;
														assign node7504 = (inp[10]) ? node7506 : 15'b000000111111111;
															assign node7506 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7510 = (inp[5]) ? 15'b000000001111111 : node7511;
														assign node7511 = (inp[10]) ? node7513 : 15'b000000011111111;
															assign node7513 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7517 = (inp[10]) ? node7521 : node7518;
													assign node7518 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7521 = (inp[3]) ? node7523 : 15'b000000001111111;
														assign node7523 = (inp[5]) ? node7525 : 15'b000000000111111;
															assign node7525 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7528 = (inp[10]) ? node7544 : node7529;
											assign node7529 = (inp[0]) ? node7535 : node7530;
												assign node7530 = (inp[4]) ? node7532 : 15'b000000111111111;
													assign node7532 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7535 = (inp[2]) ? node7539 : node7536;
													assign node7536 = (inp[5]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node7539 = (inp[4]) ? 15'b000000000111111 : node7540;
														assign node7540 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7544 = (inp[5]) ? 15'b000000000111111 : node7545;
												assign node7545 = (inp[4]) ? node7547 : 15'b000000001111111;
													assign node7547 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node7551 = (inp[4]) ? node7581 : node7552;
										assign node7552 = (inp[8]) ? node7572 : node7553;
											assign node7553 = (inp[10]) ? node7559 : node7554;
												assign node7554 = (inp[3]) ? node7556 : 15'b000000011111111;
													assign node7556 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7559 = (inp[0]) ? node7565 : node7560;
													assign node7560 = (inp[3]) ? 15'b000000001111111 : node7561;
														assign node7561 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7565 = (inp[5]) ? 15'b000000000111111 : node7566;
														assign node7566 = (inp[2]) ? node7568 : 15'b000000001111111;
															assign node7568 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7572 = (inp[5]) ? node7574 : 15'b000000001111111;
												assign node7574 = (inp[2]) ? 15'b000000000011111 : node7575;
													assign node7575 = (inp[3]) ? 15'b000000000111111 : node7576;
														assign node7576 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7581 = (inp[3]) ? node7597 : node7582;
											assign node7582 = (inp[0]) ? 15'b000000000111111 : node7583;
												assign node7583 = (inp[2]) ? node7589 : node7584;
													assign node7584 = (inp[10]) ? node7586 : 15'b000000011111111;
														assign node7586 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7589 = (inp[5]) ? node7591 : 15'b000000001111111;
														assign node7591 = (inp[10]) ? node7593 : 15'b000000000111111;
															assign node7593 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7597 = (inp[10]) ? node7603 : node7598;
												assign node7598 = (inp[0]) ? 15'b000000000011111 : node7599;
													assign node7599 = (inp[8]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node7603 = (inp[0]) ? node7605 : 15'b000000000011111;
													assign node7605 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node7608 = (inp[0]) ? node7682 : node7609;
									assign node7609 = (inp[8]) ? node7645 : node7610;
										assign node7610 = (inp[13]) ? node7624 : node7611;
											assign node7611 = (inp[5]) ? node7617 : node7612;
												assign node7612 = (inp[4]) ? node7614 : 15'b000000011111111;
													assign node7614 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7617 = (inp[2]) ? node7619 : 15'b000000001111111;
													assign node7619 = (inp[3]) ? 15'b000000001111111 : node7620;
														assign node7620 = (inp[4]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7624 = (inp[5]) ? node7638 : node7625;
												assign node7625 = (inp[3]) ? 15'b000000000111111 : node7626;
													assign node7626 = (inp[2]) ? node7632 : node7627;
														assign node7627 = (inp[4]) ? 15'b000000011111111 : node7628;
															assign node7628 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node7632 = (inp[4]) ? node7634 : 15'b000000001111111;
															assign node7634 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7638 = (inp[2]) ? node7642 : node7639;
													assign node7639 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7642 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7645 = (inp[4]) ? node7665 : node7646;
											assign node7646 = (inp[10]) ? node7650 : node7647;
												assign node7647 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7650 = (inp[13]) ? node7660 : node7651;
													assign node7651 = (inp[3]) ? node7653 : 15'b000000001111111;
														assign node7653 = (inp[5]) ? node7657 : node7654;
															assign node7654 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
															assign node7657 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7660 = (inp[2]) ? 15'b000000000011111 : node7661;
														assign node7661 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7665 = (inp[5]) ? node7669 : node7666;
												assign node7666 = (inp[3]) ? 15'b000000000111111 : 15'b000000000011111;
												assign node7669 = (inp[2]) ? node7677 : node7670;
													assign node7670 = (inp[10]) ? 15'b000000000011111 : node7671;
														assign node7671 = (inp[13]) ? node7673 : 15'b000000000111111;
															assign node7673 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7677 = (inp[13]) ? node7679 : 15'b000000000011111;
														assign node7679 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7682 = (inp[2]) ? node7706 : node7683;
										assign node7683 = (inp[4]) ? node7691 : node7684;
											assign node7684 = (inp[10]) ? 15'b000000000111111 : node7685;
												assign node7685 = (inp[13]) ? 15'b000000001111111 : node7686;
													assign node7686 = (inp[5]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node7691 = (inp[5]) ? node7701 : node7692;
												assign node7692 = (inp[3]) ? node7698 : node7693;
													assign node7693 = (inp[8]) ? node7695 : 15'b000000001111111;
														assign node7695 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7698 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7701 = (inp[3]) ? 15'b000000000011111 : node7702;
													assign node7702 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7706 = (inp[5]) ? node7726 : node7707;
											assign node7707 = (inp[3]) ? node7719 : node7708;
												assign node7708 = (inp[13]) ? node7712 : node7709;
													assign node7709 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7712 = (inp[10]) ? 15'b000000000011111 : node7713;
														assign node7713 = (inp[4]) ? node7715 : 15'b000000000111111;
															assign node7715 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7719 = (inp[13]) ? 15'b000000000001111 : node7720;
													assign node7720 = (inp[4]) ? node7722 : 15'b000000000011111;
														assign node7722 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7726 = (inp[4]) ? node7728 : 15'b000000000011111;
												assign node7728 = (inp[8]) ? node7734 : node7729;
													assign node7729 = (inp[3]) ? 15'b000000000001111 : node7730;
														assign node7730 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node7734 = (inp[10]) ? 15'b000000000000111 : node7735;
														assign node7735 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node7739 = (inp[8]) ? node7981 : node7740;
							assign node7740 = (inp[6]) ? node7854 : node7741;
								assign node7741 = (inp[4]) ? node7797 : node7742;
									assign node7742 = (inp[10]) ? node7772 : node7743;
										assign node7743 = (inp[0]) ? node7757 : node7744;
											assign node7744 = (inp[3]) ? node7752 : node7745;
												assign node7745 = (inp[1]) ? 15'b000000111111111 : node7746;
													assign node7746 = (inp[5]) ? node7748 : 15'b000000111111111;
														assign node7748 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7752 = (inp[2]) ? node7754 : 15'b000000011111111;
													assign node7754 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node7757 = (inp[2]) ? node7769 : node7758;
												assign node7758 = (inp[5]) ? node7764 : node7759;
													assign node7759 = (inp[13]) ? node7761 : 15'b000000111111111;
														assign node7761 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7764 = (inp[13]) ? node7766 : 15'b000000011111111;
														assign node7766 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7769 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node7772 = (inp[5]) ? node7786 : node7773;
											assign node7773 = (inp[13]) ? node7779 : node7774;
												assign node7774 = (inp[3]) ? 15'b000000011111111 : node7775;
													assign node7775 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node7779 = (inp[1]) ? node7783 : node7780;
													assign node7780 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node7783 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7786 = (inp[1]) ? node7790 : node7787;
												assign node7787 = (inp[0]) ? 15'b000000011111111 : 15'b000000001111111;
												assign node7790 = (inp[13]) ? node7792 : 15'b000000000111111;
													assign node7792 = (inp[0]) ? node7794 : 15'b000000000111111;
														assign node7794 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7797 = (inp[2]) ? node7829 : node7798;
										assign node7798 = (inp[13]) ? node7816 : node7799;
											assign node7799 = (inp[1]) ? node7809 : node7800;
												assign node7800 = (inp[0]) ? node7802 : 15'b000000111111111;
													assign node7802 = (inp[5]) ? node7804 : 15'b000000011111111;
														assign node7804 = (inp[10]) ? 15'b000000001111111 : node7805;
															assign node7805 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7809 = (inp[3]) ? 15'b000000001111111 : node7810;
													assign node7810 = (inp[5]) ? 15'b000000001111111 : node7811;
														assign node7811 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7816 = (inp[1]) ? node7818 : 15'b000000001111111;
												assign node7818 = (inp[10]) ? node7826 : node7819;
													assign node7819 = (inp[3]) ? node7821 : 15'b000000001111111;
														assign node7821 = (inp[0]) ? 15'b000000000111111 : node7822;
															assign node7822 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7826 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7829 = (inp[0]) ? node7839 : node7830;
											assign node7830 = (inp[10]) ? node7834 : node7831;
												assign node7831 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7834 = (inp[5]) ? 15'b000000000111111 : node7835;
													assign node7835 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7839 = (inp[13]) ? node7849 : node7840;
												assign node7840 = (inp[1]) ? node7844 : node7841;
													assign node7841 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7844 = (inp[10]) ? node7846 : 15'b000000000111111;
														assign node7846 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7849 = (inp[5]) ? 15'b000000000011111 : node7850;
													assign node7850 = (inp[1]) ? 15'b000000000011111 : 15'b000000001111111;
								assign node7854 = (inp[5]) ? node7912 : node7855;
									assign node7855 = (inp[13]) ? node7891 : node7856;
										assign node7856 = (inp[3]) ? node7870 : node7857;
											assign node7857 = (inp[4]) ? node7865 : node7858;
												assign node7858 = (inp[10]) ? node7862 : node7859;
													assign node7859 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node7862 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7865 = (inp[0]) ? 15'b000000000111111 : node7866;
													assign node7866 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node7870 = (inp[1]) ? node7878 : node7871;
												assign node7871 = (inp[10]) ? 15'b000000001111111 : node7872;
													assign node7872 = (inp[2]) ? node7874 : 15'b000000001111111;
														assign node7874 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node7878 = (inp[2]) ? node7886 : node7879;
													assign node7879 = (inp[10]) ? node7881 : 15'b000000001111111;
														assign node7881 = (inp[0]) ? 15'b000000000111111 : node7882;
															assign node7882 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7886 = (inp[0]) ? 15'b000000000011111 : node7887;
														assign node7887 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node7891 = (inp[1]) ? node7899 : node7892;
											assign node7892 = (inp[0]) ? 15'b000000000111111 : node7893;
												assign node7893 = (inp[4]) ? node7895 : 15'b000000001111111;
													assign node7895 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node7899 = (inp[0]) ? node7907 : node7900;
												assign node7900 = (inp[4]) ? node7904 : node7901;
													assign node7901 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7904 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7907 = (inp[4]) ? 15'b000000000011111 : node7908;
													assign node7908 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node7912 = (inp[1]) ? node7946 : node7913;
										assign node7913 = (inp[0]) ? node7929 : node7914;
											assign node7914 = (inp[10]) ? node7920 : node7915;
												assign node7915 = (inp[3]) ? 15'b000000001111111 : node7916;
													assign node7916 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node7920 = (inp[13]) ? node7926 : node7921;
													assign node7921 = (inp[2]) ? node7923 : 15'b000000001111111;
														assign node7923 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7926 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node7929 = (inp[4]) ? node7935 : node7930;
												assign node7930 = (inp[2]) ? node7932 : 15'b000000000111111;
													assign node7932 = (inp[10]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node7935 = (inp[10]) ? node7943 : node7936;
													assign node7936 = (inp[3]) ? 15'b000000000011111 : node7937;
														assign node7937 = (inp[13]) ? node7939 : 15'b000000000111111;
															assign node7939 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node7943 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node7946 = (inp[2]) ? node7960 : node7947;
											assign node7947 = (inp[0]) ? node7955 : node7948;
												assign node7948 = (inp[4]) ? node7952 : node7949;
													assign node7949 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node7952 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node7955 = (inp[13]) ? node7957 : 15'b000000000011111;
													assign node7957 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node7960 = (inp[10]) ? node7970 : node7961;
												assign node7961 = (inp[13]) ? node7963 : 15'b000000000011111;
													assign node7963 = (inp[0]) ? 15'b000000000001111 : node7964;
														assign node7964 = (inp[3]) ? node7966 : 15'b000000000011111;
															assign node7966 = (inp[4]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node7970 = (inp[4]) ? node7978 : node7971;
													assign node7971 = (inp[3]) ? node7973 : 15'b000000000011111;
														assign node7973 = (inp[0]) ? 15'b000000000001111 : node7974;
															assign node7974 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node7978 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node7981 = (inp[3]) ? node8085 : node7982;
								assign node7982 = (inp[13]) ? node8030 : node7983;
									assign node7983 = (inp[2]) ? node8007 : node7984;
										assign node7984 = (inp[5]) ? node7998 : node7985;
											assign node7985 = (inp[0]) ? node7993 : node7986;
												assign node7986 = (inp[1]) ? 15'b000000011111111 : node7987;
													assign node7987 = (inp[4]) ? 15'b000000011111111 : node7988;
														assign node7988 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node7993 = (inp[10]) ? 15'b000000000111111 : node7994;
													assign node7994 = (inp[4]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node7998 = (inp[4]) ? node8004 : node7999;
												assign node7999 = (inp[6]) ? 15'b000000001111111 : node8000;
													assign node8000 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8004 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8007 = (inp[4]) ? node8021 : node8008;
											assign node8008 = (inp[0]) ? node8010 : 15'b000000001111111;
												assign node8010 = (inp[5]) ? node8018 : node8011;
													assign node8011 = (inp[1]) ? 15'b000000000111111 : node8012;
														assign node8012 = (inp[6]) ? node8014 : 15'b000000001111111;
															assign node8014 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8018 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node8021 = (inp[1]) ? node8023 : 15'b000000000111111;
												assign node8023 = (inp[10]) ? node8027 : node8024;
													assign node8024 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node8027 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node8030 = (inp[1]) ? node8064 : node8031;
										assign node8031 = (inp[6]) ? node8043 : node8032;
											assign node8032 = (inp[4]) ? node8034 : 15'b000000001111111;
												assign node8034 = (inp[0]) ? 15'b000000000111111 : node8035;
													assign node8035 = (inp[5]) ? node8037 : 15'b000000001111111;
														assign node8037 = (inp[10]) ? 15'b000000000111111 : node8038;
															assign node8038 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8043 = (inp[0]) ? node8055 : node8044;
												assign node8044 = (inp[2]) ? node8048 : node8045;
													assign node8045 = (inp[4]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8048 = (inp[10]) ? node8050 : 15'b000000000111111;
														assign node8050 = (inp[4]) ? 15'b000000000011111 : node8051;
															assign node8051 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8055 = (inp[5]) ? node8059 : node8056;
													assign node8056 = (inp[4]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node8059 = (inp[4]) ? node8061 : 15'b000000000011111;
														assign node8061 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node8064 = (inp[10]) ? node8076 : node8065;
											assign node8065 = (inp[4]) ? node8071 : node8066;
												assign node8066 = (inp[2]) ? node8068 : 15'b000000000111111;
													assign node8068 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8071 = (inp[6]) ? node8073 : 15'b000000000011111;
													assign node8073 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node8076 = (inp[0]) ? 15'b000000000001111 : node8077;
												assign node8077 = (inp[4]) ? node8079 : 15'b000000000011111;
													assign node8079 = (inp[6]) ? node8081 : 15'b000000000011111;
														assign node8081 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node8085 = (inp[4]) ? node8163 : node8086;
									assign node8086 = (inp[2]) ? node8122 : node8087;
										assign node8087 = (inp[0]) ? node8105 : node8088;
											assign node8088 = (inp[5]) ? node8094 : node8089;
												assign node8089 = (inp[10]) ? 15'b000000001111111 : node8090;
													assign node8090 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8094 = (inp[10]) ? node8100 : node8095;
													assign node8095 = (inp[1]) ? node8097 : 15'b000000011111111;
														assign node8097 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node8100 = (inp[6]) ? node8102 : 15'b000000000111111;
														assign node8102 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node8105 = (inp[6]) ? node8111 : node8106;
												assign node8106 = (inp[5]) ? 15'b000000000011111 : node8107;
													assign node8107 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8111 = (inp[1]) ? node8117 : node8112;
													assign node8112 = (inp[5]) ? node8114 : 15'b000000000111111;
														assign node8114 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node8117 = (inp[13]) ? node8119 : 15'b000000000011111;
														assign node8119 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node8122 = (inp[10]) ? node8138 : node8123;
											assign node8123 = (inp[1]) ? node8129 : node8124;
												assign node8124 = (inp[0]) ? 15'b000000000111111 : node8125;
													assign node8125 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8129 = (inp[0]) ? node8135 : node8130;
													assign node8130 = (inp[13]) ? 15'b000000000011111 : node8131;
														assign node8131 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node8135 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node8138 = (inp[6]) ? node8148 : node8139;
												assign node8139 = (inp[0]) ? node8143 : node8140;
													assign node8140 = (inp[1]) ? 15'b000000000111111 : 15'b000000000011111;
													assign node8143 = (inp[13]) ? node8145 : 15'b000000000011111;
														assign node8145 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node8148 = (inp[5]) ? node8156 : node8149;
													assign node8149 = (inp[0]) ? node8151 : 15'b000000000001111;
														assign node8151 = (inp[1]) ? node8153 : 15'b000000000001111;
															assign node8153 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node8156 = (inp[1]) ? 15'b000000000001111 : node8157;
														assign node8157 = (inp[13]) ? 15'b000000000001111 : node8158;
															assign node8158 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node8163 = (inp[0]) ? node8191 : node8164;
										assign node8164 = (inp[1]) ? node8178 : node8165;
											assign node8165 = (inp[6]) ? node8173 : node8166;
												assign node8166 = (inp[2]) ? node8168 : 15'b000000001111111;
													assign node8168 = (inp[13]) ? node8170 : 15'b000000000111111;
														assign node8170 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node8173 = (inp[10]) ? 15'b000000000011111 : node8174;
													assign node8174 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node8178 = (inp[2]) ? node8184 : node8179;
												assign node8179 = (inp[6]) ? node8181 : 15'b000000000011111;
													assign node8181 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node8184 = (inp[6]) ? 15'b000000000000011 : node8185;
													assign node8185 = (inp[13]) ? 15'b000000000001111 : node8186;
														assign node8186 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node8191 = (inp[13]) ? node8211 : node8192;
											assign node8192 = (inp[1]) ? node8202 : node8193;
												assign node8193 = (inp[6]) ? node8199 : node8194;
													assign node8194 = (inp[10]) ? 15'b000000000011111 : node8195;
														assign node8195 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node8199 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node8202 = (inp[2]) ? node8208 : node8203;
													assign node8203 = (inp[10]) ? 15'b000000000001111 : node8204;
														assign node8204 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node8208 = (inp[6]) ? 15'b000000000000011 : 15'b000000000001111;
											assign node8211 = (inp[10]) ? node8223 : node8212;
												assign node8212 = (inp[6]) ? node8216 : node8213;
													assign node8213 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node8216 = (inp[5]) ? node8218 : 15'b000000000001111;
														assign node8218 = (inp[2]) ? 15'b000000000000111 : node8219;
															assign node8219 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node8223 = (inp[6]) ? node8231 : node8224;
													assign node8224 = (inp[5]) ? node8226 : 15'b000000000001111;
														assign node8226 = (inp[2]) ? 15'b000000000000111 : node8227;
															assign node8227 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node8231 = (inp[5]) ? node8233 : 15'b000000000000111;
														assign node8233 = (inp[1]) ? node8235 : 15'b000000000000011;
															assign node8235 = (inp[2]) ? 15'b000000000000001 : 15'b000000000000011;
		assign node8238 = (inp[4]) ? node12518 : node8239;
			assign node8239 = (inp[9]) ? node10419 : node8240;
				assign node8240 = (inp[3]) ? node9344 : node8241;
					assign node8241 = (inp[11]) ? node8789 : node8242;
						assign node8242 = (inp[1]) ? node8528 : node8243;
							assign node8243 = (inp[0]) ? node8381 : node8244;
								assign node8244 = (inp[5]) ? node8314 : node8245;
									assign node8245 = (inp[10]) ? node8281 : node8246;
										assign node8246 = (inp[13]) ? node8266 : node8247;
											assign node8247 = (inp[2]) ? node8255 : node8248;
												assign node8248 = (inp[14]) ? node8252 : node8249;
													assign node8249 = (inp[12]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node8252 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node8255 = (inp[8]) ? node8259 : node8256;
													assign node8256 = (inp[12]) ? 15'b000011111111111 : 15'b001111111111111;
													assign node8259 = (inp[12]) ? 15'b000011111111111 : node8260;
														assign node8260 = (inp[14]) ? 15'b000011111111111 : node8261;
															assign node8261 = (inp[6]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node8266 = (inp[6]) ? node8276 : node8267;
												assign node8267 = (inp[14]) ? node8273 : node8268;
													assign node8268 = (inp[8]) ? 15'b000011111111111 : node8269;
														assign node8269 = (inp[2]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node8273 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8276 = (inp[8]) ? node8278 : 15'b000001111111111;
													assign node8278 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node8281 = (inp[8]) ? node8301 : node8282;
											assign node8282 = (inp[2]) ? node8292 : node8283;
												assign node8283 = (inp[6]) ? 15'b000011111111111 : node8284;
													assign node8284 = (inp[13]) ? node8286 : 15'b000111111111111;
														assign node8286 = (inp[12]) ? 15'b000011111111111 : node8287;
															assign node8287 = (inp[14]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node8292 = (inp[14]) ? node8296 : node8293;
													assign node8293 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8296 = (inp[6]) ? node8298 : 15'b000001111111111;
														assign node8298 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8301 = (inp[12]) ? node8303 : 15'b000001111111111;
												assign node8303 = (inp[2]) ? 15'b000000111111111 : node8304;
													assign node8304 = (inp[6]) ? node8308 : node8305;
														assign node8305 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
														assign node8308 = (inp[13]) ? 15'b000000111111111 : node8309;
															assign node8309 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
									assign node8314 = (inp[10]) ? node8350 : node8315;
										assign node8315 = (inp[13]) ? node8331 : node8316;
											assign node8316 = (inp[14]) ? node8326 : node8317;
												assign node8317 = (inp[12]) ? node8321 : node8318;
													assign node8318 = (inp[6]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node8321 = (inp[8]) ? node8323 : 15'b000011111111111;
														assign node8323 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8326 = (inp[8]) ? 15'b000001111111111 : node8327;
													assign node8327 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node8331 = (inp[8]) ? node8341 : node8332;
												assign node8332 = (inp[12]) ? node8338 : node8333;
													assign node8333 = (inp[14]) ? node8335 : 15'b000011111111111;
														assign node8335 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8338 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8341 = (inp[12]) ? node8347 : node8342;
													assign node8342 = (inp[14]) ? 15'b000000111111111 : node8343;
														assign node8343 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8347 = (inp[2]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node8350 = (inp[14]) ? node8362 : node8351;
											assign node8351 = (inp[6]) ? node8355 : node8352;
												assign node8352 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8355 = (inp[13]) ? node8359 : node8356;
													assign node8356 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8359 = (inp[2]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node8362 = (inp[2]) ? node8368 : node8363;
												assign node8363 = (inp[13]) ? node8365 : 15'b000001111111111;
													assign node8365 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8368 = (inp[8]) ? node8376 : node8369;
													assign node8369 = (inp[6]) ? node8371 : 15'b000000111111111;
														assign node8371 = (inp[13]) ? node8373 : 15'b000000011111111;
															assign node8373 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8376 = (inp[13]) ? 15'b000000001111111 : node8377;
														assign node8377 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
								assign node8381 = (inp[10]) ? node8453 : node8382;
									assign node8382 = (inp[14]) ? node8418 : node8383;
										assign node8383 = (inp[2]) ? node8399 : node8384;
											assign node8384 = (inp[12]) ? node8392 : node8385;
												assign node8385 = (inp[6]) ? node8387 : 15'b000111111111111;
													assign node8387 = (inp[8]) ? node8389 : 15'b000011111111111;
														assign node8389 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8392 = (inp[13]) ? node8396 : node8393;
													assign node8393 = (inp[6]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8396 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8399 = (inp[12]) ? node8407 : node8400;
												assign node8400 = (inp[6]) ? node8404 : node8401;
													assign node8401 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8404 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8407 = (inp[8]) ? node8415 : node8408;
													assign node8408 = (inp[6]) ? node8410 : 15'b000001111111111;
														assign node8410 = (inp[5]) ? 15'b000000111111111 : node8411;
															assign node8411 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8415 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node8418 = (inp[8]) ? node8438 : node8419;
											assign node8419 = (inp[5]) ? node8427 : node8420;
												assign node8420 = (inp[6]) ? node8424 : node8421;
													assign node8421 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8424 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8427 = (inp[2]) ? node8435 : node8428;
													assign node8428 = (inp[12]) ? node8430 : 15'b000001111111111;
														assign node8430 = (inp[6]) ? 15'b000000111111111 : node8431;
															assign node8431 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8435 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8438 = (inp[12]) ? node8448 : node8439;
												assign node8439 = (inp[6]) ? node8445 : node8440;
													assign node8440 = (inp[13]) ? 15'b000000111111111 : node8441;
														assign node8441 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8445 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node8448 = (inp[5]) ? 15'b000000011111111 : node8449;
													assign node8449 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node8453 = (inp[6]) ? node8493 : node8454;
										assign node8454 = (inp[14]) ? node8474 : node8455;
											assign node8455 = (inp[12]) ? node8467 : node8456;
												assign node8456 = (inp[2]) ? node8460 : node8457;
													assign node8457 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8460 = (inp[8]) ? 15'b000000111111111 : node8461;
														assign node8461 = (inp[13]) ? node8463 : 15'b000001111111111;
															assign node8463 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8467 = (inp[8]) ? 15'b000000011111111 : node8468;
													assign node8468 = (inp[5]) ? 15'b000000111111111 : node8469;
														assign node8469 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8474 = (inp[2]) ? node8482 : node8475;
												assign node8475 = (inp[12]) ? node8477 : 15'b000000111111111;
													assign node8477 = (inp[13]) ? node8479 : 15'b000000111111111;
														assign node8479 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8482 = (inp[5]) ? node8490 : node8483;
													assign node8483 = (inp[8]) ? 15'b000000011111111 : node8484;
														assign node8484 = (inp[12]) ? node8486 : 15'b000000111111111;
															assign node8486 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8490 = (inp[8]) ? 15'b000000011111111 : 15'b000000001111111;
										assign node8493 = (inp[8]) ? node8513 : node8494;
											assign node8494 = (inp[14]) ? node8508 : node8495;
												assign node8495 = (inp[5]) ? node8501 : node8496;
													assign node8496 = (inp[13]) ? 15'b000000111111111 : node8497;
														assign node8497 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8501 = (inp[12]) ? node8503 : 15'b000000111111111;
														assign node8503 = (inp[13]) ? 15'b000000011111111 : node8504;
															assign node8504 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8508 = (inp[13]) ? 15'b000000011111111 : node8509;
													assign node8509 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8513 = (inp[2]) ? node8517 : node8514;
												assign node8514 = (inp[13]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node8517 = (inp[12]) ? 15'b000000001111111 : node8518;
													assign node8518 = (inp[14]) ? node8522 : node8519;
														assign node8519 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node8522 = (inp[5]) ? 15'b000000001111111 : node8523;
															assign node8523 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
							assign node8528 = (inp[2]) ? node8672 : node8529;
								assign node8529 = (inp[8]) ? node8597 : node8530;
									assign node8530 = (inp[10]) ? node8572 : node8531;
										assign node8531 = (inp[6]) ? node8553 : node8532;
											assign node8532 = (inp[12]) ? node8548 : node8533;
												assign node8533 = (inp[13]) ? node8539 : node8534;
													assign node8534 = (inp[14]) ? 15'b000011111111111 : node8535;
														assign node8535 = (inp[5]) ? 15'b000111111111111 : 15'b001111111111111;
													assign node8539 = (inp[5]) ? node8543 : node8540;
														assign node8540 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
														assign node8543 = (inp[0]) ? 15'b000001111111111 : node8544;
															assign node8544 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8548 = (inp[13]) ? 15'b000001111111111 : node8549;
													assign node8549 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node8553 = (inp[5]) ? node8561 : node8554;
												assign node8554 = (inp[14]) ? node8556 : 15'b000011111111111;
													assign node8556 = (inp[0]) ? 15'b000000111111111 : node8557;
														assign node8557 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8561 = (inp[13]) ? node8567 : node8562;
													assign node8562 = (inp[12]) ? node8564 : 15'b000001111111111;
														assign node8564 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8567 = (inp[12]) ? 15'b000000011111111 : node8568;
														assign node8568 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node8572 = (inp[0]) ? node8584 : node8573;
											assign node8573 = (inp[14]) ? node8579 : node8574;
												assign node8574 = (inp[6]) ? node8576 : 15'b000011111111111;
													assign node8576 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8579 = (inp[6]) ? node8581 : 15'b000000111111111;
													assign node8581 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8584 = (inp[5]) ? node8592 : node8585;
												assign node8585 = (inp[12]) ? node8589 : node8586;
													assign node8586 = (inp[13]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node8589 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8592 = (inp[14]) ? 15'b000000001111111 : node8593;
													assign node8593 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
									assign node8597 = (inp[13]) ? node8637 : node8598;
										assign node8598 = (inp[5]) ? node8612 : node8599;
											assign node8599 = (inp[0]) ? node8601 : 15'b000011111111111;
												assign node8601 = (inp[14]) ? node8609 : node8602;
													assign node8602 = (inp[6]) ? node8604 : 15'b000001111111111;
														assign node8604 = (inp[12]) ? 15'b000000111111111 : node8605;
															assign node8605 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8609 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8612 = (inp[6]) ? node8626 : node8613;
												assign node8613 = (inp[14]) ? node8617 : node8614;
													assign node8614 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8617 = (inp[10]) ? 15'b000000011111111 : node8618;
														assign node8618 = (inp[12]) ? node8622 : node8619;
															assign node8619 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
															assign node8622 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8626 = (inp[14]) ? node8632 : node8627;
													assign node8627 = (inp[0]) ? node8629 : 15'b000000111111111;
														assign node8629 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8632 = (inp[10]) ? node8634 : 15'b000000011111111;
														assign node8634 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8637 = (inp[6]) ? node8653 : node8638;
											assign node8638 = (inp[5]) ? node8642 : node8639;
												assign node8639 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8642 = (inp[0]) ? node8648 : node8643;
													assign node8643 = (inp[10]) ? 15'b000000011111111 : node8644;
														assign node8644 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8648 = (inp[12]) ? 15'b000000001111111 : node8649;
														assign node8649 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8653 = (inp[12]) ? node8665 : node8654;
												assign node8654 = (inp[14]) ? node8660 : node8655;
													assign node8655 = (inp[5]) ? 15'b000000011111111 : node8656;
														assign node8656 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8660 = (inp[10]) ? 15'b000000001111111 : node8661;
														assign node8661 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8665 = (inp[14]) ? 15'b000000001111111 : node8666;
													assign node8666 = (inp[5]) ? node8668 : 15'b000000001111111;
														assign node8668 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node8672 = (inp[12]) ? node8734 : node8673;
									assign node8673 = (inp[10]) ? node8699 : node8674;
										assign node8674 = (inp[5]) ? node8688 : node8675;
											assign node8675 = (inp[6]) ? node8683 : node8676;
												assign node8676 = (inp[13]) ? node8678 : 15'b000011111111111;
													assign node8678 = (inp[14]) ? node8680 : 15'b000001111111111;
														assign node8680 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8683 = (inp[14]) ? node8685 : 15'b000000111111111;
													assign node8685 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node8688 = (inp[13]) ? node8696 : node8689;
												assign node8689 = (inp[0]) ? node8691 : 15'b000000111111111;
													assign node8691 = (inp[8]) ? node8693 : 15'b000000111111111;
														assign node8693 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8696 = (inp[0]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node8699 = (inp[6]) ? node8721 : node8700;
											assign node8700 = (inp[13]) ? node8710 : node8701;
												assign node8701 = (inp[14]) ? node8705 : node8702;
													assign node8702 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8705 = (inp[5]) ? node8707 : 15'b000000111111111;
														assign node8707 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8710 = (inp[5]) ? node8714 : node8711;
													assign node8711 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8714 = (inp[14]) ? 15'b000000001111111 : node8715;
														assign node8715 = (inp[8]) ? node8717 : 15'b000000011111111;
															assign node8717 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8721 = (inp[14]) ? node8729 : node8722;
												assign node8722 = (inp[0]) ? node8726 : node8723;
													assign node8723 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8726 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8729 = (inp[0]) ? 15'b000000001111111 : node8730;
													assign node8730 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node8734 = (inp[13]) ? node8762 : node8735;
										assign node8735 = (inp[0]) ? node8747 : node8736;
											assign node8736 = (inp[6]) ? node8742 : node8737;
												assign node8737 = (inp[14]) ? node8739 : 15'b000000111111111;
													assign node8739 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8742 = (inp[14]) ? 15'b000000011111111 : node8743;
													assign node8743 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8747 = (inp[5]) ? node8753 : node8748;
												assign node8748 = (inp[14]) ? node8750 : 15'b000000111111111;
													assign node8750 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8753 = (inp[14]) ? node8757 : node8754;
													assign node8754 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8757 = (inp[8]) ? node8759 : 15'b000000001111111;
														assign node8759 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8762 = (inp[14]) ? node8776 : node8763;
											assign node8763 = (inp[8]) ? node8769 : node8764;
												assign node8764 = (inp[10]) ? 15'b000000001111111 : node8765;
													assign node8765 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8769 = (inp[6]) ? node8773 : node8770;
													assign node8770 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8773 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node8776 = (inp[0]) ? node8782 : node8777;
												assign node8777 = (inp[6]) ? node8779 : 15'b000000001111111;
													assign node8779 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node8782 = (inp[6]) ? 15'b000000000011111 : node8783;
													assign node8783 = (inp[10]) ? node8785 : 15'b000000001111111;
														assign node8785 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
						assign node8789 = (inp[5]) ? node9077 : node8790;
							assign node8790 = (inp[13]) ? node8930 : node8791;
								assign node8791 = (inp[0]) ? node8857 : node8792;
									assign node8792 = (inp[1]) ? node8832 : node8793;
										assign node8793 = (inp[8]) ? node8817 : node8794;
											assign node8794 = (inp[12]) ? node8810 : node8795;
												assign node8795 = (inp[6]) ? node8807 : node8796;
													assign node8796 = (inp[10]) ? node8802 : node8797;
														assign node8797 = (inp[2]) ? node8799 : 15'b000111111111111;
															assign node8799 = (inp[14]) ? 15'b000011111111111 : 15'b000111111111111;
														assign node8802 = (inp[2]) ? node8804 : 15'b000011111111111;
															assign node8804 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8807 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node8810 = (inp[10]) ? node8814 : node8811;
													assign node8811 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8814 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8817 = (inp[14]) ? node8823 : node8818;
												assign node8818 = (inp[12]) ? node8820 : 15'b000001111111111;
													assign node8820 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8823 = (inp[10]) ? node8829 : node8824;
													assign node8824 = (inp[12]) ? node8826 : 15'b000001111111111;
														assign node8826 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8829 = (inp[6]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node8832 = (inp[10]) ? node8842 : node8833;
											assign node8833 = (inp[2]) ? node8839 : node8834;
												assign node8834 = (inp[14]) ? 15'b000001111111111 : node8835;
													assign node8835 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8839 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8842 = (inp[6]) ? node8852 : node8843;
												assign node8843 = (inp[12]) ? 15'b000000111111111 : node8844;
													assign node8844 = (inp[8]) ? 15'b000000111111111 : node8845;
														assign node8845 = (inp[2]) ? node8847 : 15'b000001111111111;
															assign node8847 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8852 = (inp[14]) ? 15'b000000011111111 : node8853;
													assign node8853 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node8857 = (inp[14]) ? node8891 : node8858;
										assign node8858 = (inp[12]) ? node8880 : node8859;
											assign node8859 = (inp[6]) ? node8873 : node8860;
												assign node8860 = (inp[10]) ? node8866 : node8861;
													assign node8861 = (inp[1]) ? 15'b000001111111111 : node8862;
														assign node8862 = (inp[2]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node8866 = (inp[2]) ? 15'b000000111111111 : node8867;
														assign node8867 = (inp[8]) ? node8869 : 15'b000001111111111;
															assign node8869 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8873 = (inp[2]) ? node8877 : node8874;
													assign node8874 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node8877 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8880 = (inp[2]) ? node8888 : node8881;
												assign node8881 = (inp[10]) ? node8883 : 15'b000000111111111;
													assign node8883 = (inp[8]) ? node8885 : 15'b000000111111111;
														assign node8885 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8888 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node8891 = (inp[10]) ? node8911 : node8892;
											assign node8892 = (inp[6]) ? node8898 : node8893;
												assign node8893 = (inp[12]) ? 15'b000000111111111 : node8894;
													assign node8894 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node8898 = (inp[12]) ? node8906 : node8899;
													assign node8899 = (inp[1]) ? node8901 : 15'b000000111111111;
														assign node8901 = (inp[8]) ? 15'b000000011111111 : node8902;
															assign node8902 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8906 = (inp[2]) ? 15'b000000001111111 : node8907;
														assign node8907 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node8911 = (inp[2]) ? node8925 : node8912;
												assign node8912 = (inp[8]) ? node8916 : node8913;
													assign node8913 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node8916 = (inp[1]) ? node8920 : node8917;
														assign node8917 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node8920 = (inp[12]) ? 15'b000000001111111 : node8921;
															assign node8921 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node8925 = (inp[1]) ? 15'b000000001111111 : node8926;
													assign node8926 = (inp[6]) ? 15'b000000000111111 : 15'b000000011111111;
								assign node8930 = (inp[2]) ? node8994 : node8931;
									assign node8931 = (inp[8]) ? node8967 : node8932;
										assign node8932 = (inp[14]) ? node8948 : node8933;
											assign node8933 = (inp[0]) ? node8939 : node8934;
												assign node8934 = (inp[10]) ? node8936 : 15'b000001111111111;
													assign node8936 = (inp[1]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node8939 = (inp[6]) ? 15'b000000111111111 : node8940;
													assign node8940 = (inp[10]) ? node8942 : 15'b000001111111111;
														assign node8942 = (inp[12]) ? 15'b000000111111111 : node8943;
															assign node8943 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node8948 = (inp[0]) ? node8958 : node8949;
												assign node8949 = (inp[12]) ? node8955 : node8950;
													assign node8950 = (inp[6]) ? 15'b000001111111111 : node8951;
														assign node8951 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node8955 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8958 = (inp[12]) ? node8962 : node8959;
													assign node8959 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node8962 = (inp[1]) ? node8964 : 15'b000000001111111;
														assign node8964 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node8967 = (inp[1]) ? node8983 : node8968;
											assign node8968 = (inp[12]) ? node8976 : node8969;
												assign node8969 = (inp[0]) ? node8971 : 15'b000000111111111;
													assign node8971 = (inp[10]) ? node8973 : 15'b000000111111111;
														assign node8973 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8976 = (inp[6]) ? 15'b000000011111111 : node8977;
													assign node8977 = (inp[14]) ? node8979 : 15'b000000111111111;
														assign node8979 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node8983 = (inp[6]) ? node8989 : node8984;
												assign node8984 = (inp[14]) ? 15'b000000011111111 : node8985;
													assign node8985 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node8989 = (inp[10]) ? 15'b000000000111111 : node8990;
													assign node8990 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node8994 = (inp[14]) ? node9032 : node8995;
										assign node8995 = (inp[0]) ? node9017 : node8996;
											assign node8996 = (inp[8]) ? node9010 : node8997;
												assign node8997 = (inp[1]) ? node9003 : node8998;
													assign node8998 = (inp[10]) ? 15'b000000111111111 : node8999;
														assign node8999 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9003 = (inp[6]) ? node9005 : 15'b000001111111111;
														assign node9005 = (inp[10]) ? 15'b000000011111111 : node9006;
															assign node9006 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9010 = (inp[10]) ? node9014 : node9011;
													assign node9011 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9014 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9017 = (inp[8]) ? node9025 : node9018;
												assign node9018 = (inp[6]) ? 15'b000000011111111 : node9019;
													assign node9019 = (inp[10]) ? 15'b000000011111111 : node9020;
														assign node9020 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9025 = (inp[6]) ? node9029 : node9026;
													assign node9026 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9029 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9032 = (inp[10]) ? node9054 : node9033;
											assign node9033 = (inp[1]) ? node9049 : node9034;
												assign node9034 = (inp[6]) ? node9042 : node9035;
													assign node9035 = (inp[0]) ? node9037 : 15'b000000111111111;
														assign node9037 = (inp[8]) ? 15'b000000011111111 : node9038;
															assign node9038 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9042 = (inp[0]) ? 15'b000000001111111 : node9043;
														assign node9043 = (inp[8]) ? node9045 : 15'b000000011111111;
															assign node9045 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9049 = (inp[8]) ? node9051 : 15'b000000011111111;
													assign node9051 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9054 = (inp[0]) ? node9066 : node9055;
												assign node9055 = (inp[1]) ? node9061 : node9056;
													assign node9056 = (inp[12]) ? node9058 : 15'b000000011111111;
														assign node9058 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9061 = (inp[12]) ? 15'b000000000111111 : node9062;
														assign node9062 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9066 = (inp[12]) ? node9072 : node9067;
													assign node9067 = (inp[1]) ? 15'b000000000111111 : node9068;
														assign node9068 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9072 = (inp[8]) ? node9074 : 15'b000000000111111;
														assign node9074 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node9077 = (inp[14]) ? node9219 : node9078;
								assign node9078 = (inp[6]) ? node9148 : node9079;
									assign node9079 = (inp[12]) ? node9113 : node9080;
										assign node9080 = (inp[10]) ? node9100 : node9081;
											assign node9081 = (inp[8]) ? node9089 : node9082;
												assign node9082 = (inp[13]) ? node9086 : node9083;
													assign node9083 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node9086 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9089 = (inp[2]) ? node9091 : 15'b000001111111111;
													assign node9091 = (inp[0]) ? node9097 : node9092;
														assign node9092 = (inp[13]) ? 15'b000000111111111 : node9093;
															assign node9093 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node9097 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9100 = (inp[13]) ? node9108 : node9101;
												assign node9101 = (inp[8]) ? node9105 : node9102;
													assign node9102 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9105 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9108 = (inp[8]) ? 15'b000000011111111 : node9109;
													assign node9109 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node9113 = (inp[2]) ? node9135 : node9114;
											assign node9114 = (inp[13]) ? node9122 : node9115;
												assign node9115 = (inp[8]) ? node9119 : node9116;
													assign node9116 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9119 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9122 = (inp[10]) ? node9128 : node9123;
													assign node9123 = (inp[8]) ? node9125 : 15'b000000111111111;
														assign node9125 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9128 = (inp[0]) ? node9130 : 15'b000000011111111;
														assign node9130 = (inp[8]) ? 15'b000000001111111 : node9131;
															assign node9131 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9135 = (inp[1]) ? node9143 : node9136;
												assign node9136 = (inp[8]) ? node9138 : 15'b000000011111111;
													assign node9138 = (inp[0]) ? node9140 : 15'b000000011111111;
														assign node9140 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9143 = (inp[0]) ? 15'b000000001111111 : node9144;
													assign node9144 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node9148 = (inp[13]) ? node9182 : node9149;
										assign node9149 = (inp[1]) ? node9169 : node9150;
											assign node9150 = (inp[12]) ? node9158 : node9151;
												assign node9151 = (inp[0]) ? node9155 : node9152;
													assign node9152 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9155 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9158 = (inp[8]) ? node9162 : node9159;
													assign node9159 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9162 = (inp[2]) ? 15'b000000001111111 : node9163;
														assign node9163 = (inp[0]) ? node9165 : 15'b000000011111111;
															assign node9165 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9169 = (inp[0]) ? node9177 : node9170;
												assign node9170 = (inp[2]) ? node9174 : node9171;
													assign node9171 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9174 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9177 = (inp[2]) ? node9179 : 15'b000000001111111;
													assign node9179 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9182 = (inp[2]) ? node9198 : node9183;
											assign node9183 = (inp[1]) ? node9195 : node9184;
												assign node9184 = (inp[8]) ? node9188 : node9185;
													assign node9185 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9188 = (inp[12]) ? 15'b000000001111111 : node9189;
														assign node9189 = (inp[0]) ? node9191 : 15'b000000111111111;
															assign node9191 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9195 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9198 = (inp[8]) ? node9210 : node9199;
												assign node9199 = (inp[10]) ? node9203 : node9200;
													assign node9200 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9203 = (inp[12]) ? 15'b000000000111111 : node9204;
														assign node9204 = (inp[0]) ? node9206 : 15'b000000001111111;
															assign node9206 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9210 = (inp[12]) ? node9216 : node9211;
													assign node9211 = (inp[1]) ? 15'b000000000111111 : node9212;
														assign node9212 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9216 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node9219 = (inp[10]) ? node9271 : node9220;
									assign node9220 = (inp[13]) ? node9242 : node9221;
										assign node9221 = (inp[0]) ? node9231 : node9222;
											assign node9222 = (inp[6]) ? node9226 : node9223;
												assign node9223 = (inp[2]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node9226 = (inp[8]) ? 15'b000000011111111 : node9227;
													assign node9227 = (inp[1]) ? 15'b000000011111111 : 15'b000001111111111;
											assign node9231 = (inp[6]) ? node9233 : 15'b000000011111111;
												assign node9233 = (inp[12]) ? node9239 : node9234;
													assign node9234 = (inp[8]) ? node9236 : 15'b000000011111111;
														assign node9236 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9239 = (inp[1]) ? 15'b000000001111111 : 15'b000000000111111;
										assign node9242 = (inp[2]) ? node9258 : node9243;
											assign node9243 = (inp[0]) ? node9253 : node9244;
												assign node9244 = (inp[6]) ? node9250 : node9245;
													assign node9245 = (inp[8]) ? 15'b000000011111111 : node9246;
														assign node9246 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9250 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9253 = (inp[6]) ? 15'b000000000111111 : node9254;
													assign node9254 = (inp[1]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node9258 = (inp[8]) ? node9266 : node9259;
												assign node9259 = (inp[1]) ? node9263 : node9260;
													assign node9260 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9263 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9266 = (inp[1]) ? node9268 : 15'b000000000111111;
													assign node9268 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node9271 = (inp[8]) ? node9297 : node9272;
										assign node9272 = (inp[13]) ? node9286 : node9273;
											assign node9273 = (inp[12]) ? node9279 : node9274;
												assign node9274 = (inp[1]) ? node9276 : 15'b000000111111111;
													assign node9276 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9279 = (inp[0]) ? 15'b000000001111111 : node9280;
													assign node9280 = (inp[1]) ? 15'b000000001111111 : node9281;
														assign node9281 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9286 = (inp[2]) ? node9292 : node9287;
												assign node9287 = (inp[0]) ? node9289 : 15'b000000001111111;
													assign node9289 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9292 = (inp[6]) ? node9294 : 15'b000000000111111;
													assign node9294 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9297 = (inp[12]) ? node9319 : node9298;
											assign node9298 = (inp[0]) ? node9304 : node9299;
												assign node9299 = (inp[13]) ? node9301 : 15'b000000001111111;
													assign node9301 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9304 = (inp[13]) ? node9310 : node9305;
													assign node9305 = (inp[6]) ? node9307 : 15'b000000001111111;
														assign node9307 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9310 = (inp[1]) ? node9316 : node9311;
														assign node9311 = (inp[2]) ? 15'b000000000111111 : node9312;
															assign node9312 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
														assign node9316 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9319 = (inp[1]) ? node9329 : node9320;
												assign node9320 = (inp[6]) ? node9326 : node9321;
													assign node9321 = (inp[2]) ? 15'b000000000111111 : node9322;
														assign node9322 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9326 = (inp[13]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node9329 = (inp[6]) ? node9339 : node9330;
													assign node9330 = (inp[0]) ? node9334 : node9331;
														assign node9331 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
														assign node9334 = (inp[13]) ? node9336 : 15'b000000000011111;
															assign node9336 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node9339 = (inp[13]) ? 15'b000000000001111 : node9340;
														assign node9340 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
					assign node9344 = (inp[1]) ? node9870 : node9345;
						assign node9345 = (inp[12]) ? node9597 : node9346;
							assign node9346 = (inp[11]) ? node9486 : node9347;
								assign node9347 = (inp[2]) ? node9421 : node9348;
									assign node9348 = (inp[5]) ? node9384 : node9349;
										assign node9349 = (inp[6]) ? node9367 : node9350;
											assign node9350 = (inp[13]) ? node9358 : node9351;
												assign node9351 = (inp[8]) ? node9353 : 15'b000111111111111;
													assign node9353 = (inp[10]) ? 15'b000011111111111 : node9354;
														assign node9354 = (inp[0]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node9358 = (inp[0]) ? 15'b000001111111111 : node9359;
													assign node9359 = (inp[10]) ? 15'b000011111111111 : node9360;
														assign node9360 = (inp[14]) ? 15'b000011111111111 : node9361;
															assign node9361 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
											assign node9367 = (inp[0]) ? node9379 : node9368;
												assign node9368 = (inp[13]) ? 15'b000001111111111 : node9369;
													assign node9369 = (inp[14]) ? node9373 : node9370;
														assign node9370 = (inp[8]) ? 15'b000011111111111 : 15'b000111111111111;
														assign node9373 = (inp[8]) ? 15'b000001111111111 : node9374;
															assign node9374 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node9379 = (inp[10]) ? 15'b000000011111111 : node9380;
													assign node9380 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node9384 = (inp[8]) ? node9406 : node9385;
											assign node9385 = (inp[10]) ? node9397 : node9386;
												assign node9386 = (inp[14]) ? node9390 : node9387;
													assign node9387 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node9390 = (inp[0]) ? node9392 : 15'b000011111111111;
														assign node9392 = (inp[13]) ? 15'b000000111111111 : node9393;
															assign node9393 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9397 = (inp[0]) ? node9401 : node9398;
													assign node9398 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9401 = (inp[6]) ? node9403 : 15'b000000111111111;
														assign node9403 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9406 = (inp[6]) ? node9414 : node9407;
												assign node9407 = (inp[10]) ? 15'b000000011111111 : node9408;
													assign node9408 = (inp[0]) ? 15'b000000111111111 : node9409;
														assign node9409 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9414 = (inp[14]) ? 15'b000000001111111 : node9415;
													assign node9415 = (inp[13]) ? 15'b000000011111111 : node9416;
														assign node9416 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node9421 = (inp[0]) ? node9457 : node9422;
										assign node9422 = (inp[13]) ? node9442 : node9423;
											assign node9423 = (inp[14]) ? node9431 : node9424;
												assign node9424 = (inp[8]) ? node9426 : 15'b000001111111111;
													assign node9426 = (inp[5]) ? node9428 : 15'b000001111111111;
														assign node9428 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9431 = (inp[5]) ? node9435 : node9432;
													assign node9432 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9435 = (inp[6]) ? node9437 : 15'b000000111111111;
														assign node9437 = (inp[10]) ? 15'b000000011111111 : node9438;
															assign node9438 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9442 = (inp[8]) ? node9450 : node9443;
												assign node9443 = (inp[6]) ? 15'b000000111111111 : node9444;
													assign node9444 = (inp[5]) ? 15'b000000111111111 : node9445;
														assign node9445 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9450 = (inp[14]) ? node9454 : node9451;
													assign node9451 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9454 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node9457 = (inp[6]) ? node9471 : node9458;
											assign node9458 = (inp[10]) ? node9464 : node9459;
												assign node9459 = (inp[8]) ? 15'b000000111111111 : node9460;
													assign node9460 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9464 = (inp[8]) ? 15'b000000000111111 : node9465;
													assign node9465 = (inp[13]) ? 15'b000000011111111 : node9466;
														assign node9466 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9471 = (inp[5]) ? node9477 : node9472;
												assign node9472 = (inp[8]) ? node9474 : 15'b000000011111111;
													assign node9474 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node9477 = (inp[10]) ? node9481 : node9478;
													assign node9478 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9481 = (inp[14]) ? node9483 : 15'b000000001111111;
														assign node9483 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node9486 = (inp[14]) ? node9534 : node9487;
									assign node9487 = (inp[6]) ? node9517 : node9488;
										assign node9488 = (inp[13]) ? node9506 : node9489;
											assign node9489 = (inp[10]) ? node9499 : node9490;
												assign node9490 = (inp[8]) ? 15'b000001111111111 : node9491;
													assign node9491 = (inp[0]) ? 15'b000001111111111 : node9492;
														assign node9492 = (inp[2]) ? node9494 : 15'b000011111111111;
															assign node9494 = (inp[5]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node9499 = (inp[5]) ? node9501 : 15'b000001111111111;
													assign node9501 = (inp[2]) ? 15'b000000011111111 : node9502;
														assign node9502 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node9506 = (inp[0]) ? node9508 : 15'b000000111111111;
												assign node9508 = (inp[2]) ? node9510 : 15'b000001111111111;
													assign node9510 = (inp[8]) ? 15'b000000011111111 : node9511;
														assign node9511 = (inp[5]) ? 15'b000000011111111 : node9512;
															assign node9512 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node9517 = (inp[10]) ? node9525 : node9518;
											assign node9518 = (inp[5]) ? 15'b000000011111111 : node9519;
												assign node9519 = (inp[8]) ? 15'b000000011111111 : node9520;
													assign node9520 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node9525 = (inp[0]) ? node9527 : 15'b000000011111111;
												assign node9527 = (inp[8]) ? 15'b000000001111111 : node9528;
													assign node9528 = (inp[2]) ? node9530 : 15'b000000001111111;
														assign node9530 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node9534 = (inp[13]) ? node9572 : node9535;
										assign node9535 = (inp[6]) ? node9549 : node9536;
											assign node9536 = (inp[0]) ? node9546 : node9537;
												assign node9537 = (inp[2]) ? node9539 : 15'b000001111111111;
													assign node9539 = (inp[10]) ? node9541 : 15'b000000111111111;
														assign node9541 = (inp[8]) ? 15'b000000011111111 : node9542;
															assign node9542 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9546 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9549 = (inp[2]) ? node9559 : node9550;
												assign node9550 = (inp[0]) ? node9556 : node9551;
													assign node9551 = (inp[10]) ? 15'b000000011111111 : node9552;
														assign node9552 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9556 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9559 = (inp[5]) ? node9565 : node9560;
													assign node9560 = (inp[10]) ? 15'b000000001111111 : node9561;
														assign node9561 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9565 = (inp[8]) ? node9567 : 15'b000000001111111;
														assign node9567 = (inp[10]) ? 15'b000000000111111 : node9568;
															assign node9568 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9572 = (inp[2]) ? node9580 : node9573;
											assign node9573 = (inp[0]) ? 15'b000000001111111 : node9574;
												assign node9574 = (inp[5]) ? node9576 : 15'b000000111111111;
													assign node9576 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9580 = (inp[10]) ? node9590 : node9581;
												assign node9581 = (inp[8]) ? node9587 : node9582;
													assign node9582 = (inp[0]) ? 15'b000000001111111 : node9583;
														assign node9583 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9587 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node9590 = (inp[6]) ? node9592 : 15'b000000000111111;
													assign node9592 = (inp[5]) ? node9594 : 15'b000000000111111;
														assign node9594 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node9597 = (inp[13]) ? node9731 : node9598;
								assign node9598 = (inp[5]) ? node9670 : node9599;
									assign node9599 = (inp[8]) ? node9639 : node9600;
										assign node9600 = (inp[0]) ? node9622 : node9601;
											assign node9601 = (inp[6]) ? node9615 : node9602;
												assign node9602 = (inp[14]) ? node9610 : node9603;
													assign node9603 = (inp[10]) ? node9605 : 15'b000111111111111;
														assign node9605 = (inp[2]) ? 15'b000001111111111 : node9606;
															assign node9606 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node9610 = (inp[10]) ? node9612 : 15'b000001111111111;
														assign node9612 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9615 = (inp[14]) ? node9619 : node9616;
													assign node9616 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9619 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9622 = (inp[14]) ? node9632 : node9623;
												assign node9623 = (inp[10]) ? node9627 : node9624;
													assign node9624 = (inp[2]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node9627 = (inp[6]) ? node9629 : 15'b000000111111111;
														assign node9629 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9632 = (inp[10]) ? 15'b000000011111111 : node9633;
													assign node9633 = (inp[6]) ? 15'b000000011111111 : node9634;
														assign node9634 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node9639 = (inp[14]) ? node9655 : node9640;
											assign node9640 = (inp[6]) ? node9648 : node9641;
												assign node9641 = (inp[2]) ? node9643 : 15'b000000111111111;
													assign node9643 = (inp[11]) ? node9645 : 15'b000000111111111;
														assign node9645 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9648 = (inp[11]) ? 15'b000000001111111 : node9649;
													assign node9649 = (inp[10]) ? 15'b000000011111111 : node9650;
														assign node9650 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9655 = (inp[10]) ? node9661 : node9656;
												assign node9656 = (inp[11]) ? node9658 : 15'b000000111111111;
													assign node9658 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9661 = (inp[2]) ? node9667 : node9662;
													assign node9662 = (inp[6]) ? 15'b000000001111111 : node9663;
														assign node9663 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9667 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node9670 = (inp[0]) ? node9700 : node9671;
										assign node9671 = (inp[14]) ? node9687 : node9672;
											assign node9672 = (inp[11]) ? node9682 : node9673;
												assign node9673 = (inp[6]) ? node9679 : node9674;
													assign node9674 = (inp[10]) ? node9676 : 15'b000001111111111;
														assign node9676 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9679 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9682 = (inp[8]) ? 15'b000000011111111 : node9683;
													assign node9683 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node9687 = (inp[2]) ? node9693 : node9688;
												assign node9688 = (inp[10]) ? node9690 : 15'b000000111111111;
													assign node9690 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9693 = (inp[11]) ? node9695 : 15'b000000001111111;
													assign node9695 = (inp[6]) ? node9697 : 15'b000000001111111;
														assign node9697 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9700 = (inp[11]) ? node9716 : node9701;
											assign node9701 = (inp[8]) ? node9713 : node9702;
												assign node9702 = (inp[14]) ? node9708 : node9703;
													assign node9703 = (inp[6]) ? 15'b000000011111111 : node9704;
														assign node9704 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9708 = (inp[10]) ? 15'b000000001111111 : node9709;
														assign node9709 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9713 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node9716 = (inp[6]) ? node9726 : node9717;
												assign node9717 = (inp[10]) ? node9721 : node9718;
													assign node9718 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9721 = (inp[8]) ? 15'b000000000111111 : node9722;
														assign node9722 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9726 = (inp[10]) ? node9728 : 15'b000000000111111;
													assign node9728 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node9731 = (inp[8]) ? node9793 : node9732;
									assign node9732 = (inp[10]) ? node9768 : node9733;
										assign node9733 = (inp[14]) ? node9751 : node9734;
											assign node9734 = (inp[2]) ? node9742 : node9735;
												assign node9735 = (inp[5]) ? 15'b000000111111111 : node9736;
													assign node9736 = (inp[11]) ? 15'b000001111111111 : node9737;
														assign node9737 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node9742 = (inp[11]) ? node9746 : node9743;
													assign node9743 = (inp[5]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node9746 = (inp[6]) ? node9748 : 15'b000000011111111;
														assign node9748 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9751 = (inp[2]) ? node9761 : node9752;
												assign node9752 = (inp[0]) ? node9756 : node9753;
													assign node9753 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9756 = (inp[11]) ? node9758 : 15'b000000011111111;
														assign node9758 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9761 = (inp[11]) ? 15'b000000001111111 : node9762;
													assign node9762 = (inp[6]) ? 15'b000000001111111 : node9763;
														assign node9763 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node9768 = (inp[0]) ? node9776 : node9769;
											assign node9769 = (inp[5]) ? node9771 : 15'b000000011111111;
												assign node9771 = (inp[14]) ? 15'b000000001111111 : node9772;
													assign node9772 = (inp[11]) ? 15'b000000011111111 : 15'b000000001111111;
											assign node9776 = (inp[2]) ? node9786 : node9777;
												assign node9777 = (inp[6]) ? node9781 : node9778;
													assign node9778 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9781 = (inp[5]) ? 15'b000000000111111 : node9782;
														assign node9782 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9786 = (inp[6]) ? node9788 : 15'b000000000111111;
													assign node9788 = (inp[11]) ? 15'b000000000011111 : node9789;
														assign node9789 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node9793 = (inp[14]) ? node9835 : node9794;
										assign node9794 = (inp[11]) ? node9822 : node9795;
											assign node9795 = (inp[5]) ? node9811 : node9796;
												assign node9796 = (inp[10]) ? node9800 : node9797;
													assign node9797 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9800 = (inp[0]) ? node9806 : node9801;
														assign node9801 = (inp[6]) ? node9803 : 15'b000000011111111;
															assign node9803 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node9806 = (inp[6]) ? node9808 : 15'b000000001111111;
															assign node9808 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9811 = (inp[6]) ? node9815 : node9812;
													assign node9812 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9815 = (inp[10]) ? node9817 : 15'b000000001111111;
														assign node9817 = (inp[0]) ? 15'b000000000111111 : node9818;
															assign node9818 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node9822 = (inp[0]) ? node9830 : node9823;
												assign node9823 = (inp[2]) ? node9825 : 15'b000000011111111;
													assign node9825 = (inp[6]) ? node9827 : 15'b000000001111111;
														assign node9827 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9830 = (inp[10]) ? node9832 : 15'b000000000111111;
													assign node9832 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node9835 = (inp[0]) ? node9853 : node9836;
											assign node9836 = (inp[11]) ? node9842 : node9837;
												assign node9837 = (inp[5]) ? node9839 : 15'b000000011111111;
													assign node9839 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node9842 = (inp[2]) ? node9848 : node9843;
													assign node9843 = (inp[10]) ? 15'b000000000111111 : node9844;
														assign node9844 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9848 = (inp[6]) ? 15'b000000000011111 : node9849;
														assign node9849 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node9853 = (inp[6]) ? node9859 : node9854;
												assign node9854 = (inp[2]) ? 15'b000000000111111 : node9855;
													assign node9855 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node9859 = (inp[11]) ? node9863 : node9860;
													assign node9860 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node9863 = (inp[10]) ? node9865 : 15'b000000000011111;
														assign node9865 = (inp[5]) ? node9867 : 15'b000000000001111;
															assign node9867 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node9870 = (inp[6]) ? node10154 : node9871;
							assign node9871 = (inp[5]) ? node10031 : node9872;
								assign node9872 = (inp[0]) ? node9964 : node9873;
									assign node9873 = (inp[14]) ? node9911 : node9874;
										assign node9874 = (inp[13]) ? node9894 : node9875;
											assign node9875 = (inp[2]) ? node9887 : node9876;
												assign node9876 = (inp[10]) ? node9882 : node9877;
													assign node9877 = (inp[8]) ? 15'b000001111111111 : node9878;
														assign node9878 = (inp[12]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node9882 = (inp[11]) ? node9884 : 15'b000001111111111;
														assign node9884 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node9887 = (inp[10]) ? node9891 : node9888;
													assign node9888 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node9891 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9894 = (inp[8]) ? node9904 : node9895;
												assign node9895 = (inp[2]) ? node9901 : node9896;
													assign node9896 = (inp[11]) ? 15'b000000111111111 : node9897;
														assign node9897 = (inp[12]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node9901 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9904 = (inp[12]) ? 15'b000000011111111 : node9905;
													assign node9905 = (inp[10]) ? 15'b000000011111111 : node9906;
														assign node9906 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node9911 = (inp[12]) ? node9941 : node9912;
											assign node9912 = (inp[10]) ? node9926 : node9913;
												assign node9913 = (inp[2]) ? node9917 : node9914;
													assign node9914 = (inp[8]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node9917 = (inp[8]) ? 15'b000000011111111 : node9918;
														assign node9918 = (inp[13]) ? node9922 : node9919;
															assign node9919 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
															assign node9922 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9926 = (inp[2]) ? node9938 : node9927;
													assign node9927 = (inp[11]) ? node9933 : node9928;
														assign node9928 = (inp[8]) ? node9930 : 15'b000000111111111;
															assign node9930 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node9933 = (inp[8]) ? 15'b000000011111111 : node9934;
															assign node9934 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9938 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node9941 = (inp[11]) ? node9951 : node9942;
												assign node9942 = (inp[10]) ? node9944 : 15'b000000111111111;
													assign node9944 = (inp[2]) ? 15'b000000001111111 : node9945;
														assign node9945 = (inp[8]) ? node9947 : 15'b000000011111111;
															assign node9947 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9951 = (inp[13]) ? node9961 : node9952;
													assign node9952 = (inp[8]) ? node9958 : node9953;
														assign node9953 = (inp[2]) ? node9955 : 15'b000000011111111;
															assign node9955 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node9958 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node9961 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node9964 = (inp[11]) ? node9998 : node9965;
										assign node9965 = (inp[12]) ? node9973 : node9966;
											assign node9966 = (inp[14]) ? node9970 : node9967;
												assign node9967 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node9970 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node9973 = (inp[14]) ? node9987 : node9974;
												assign node9974 = (inp[10]) ? node9980 : node9975;
													assign node9975 = (inp[13]) ? 15'b000000011111111 : node9976;
														assign node9976 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node9980 = (inp[2]) ? node9982 : 15'b000000011111111;
														assign node9982 = (inp[8]) ? 15'b000000001111111 : node9983;
															assign node9983 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node9987 = (inp[13]) ? node9995 : node9988;
													assign node9988 = (inp[8]) ? node9990 : 15'b000000011111111;
														assign node9990 = (inp[2]) ? 15'b000000001111111 : node9991;
															assign node9991 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node9995 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node9998 = (inp[13]) ? node10012 : node9999;
											assign node9999 = (inp[2]) ? 15'b000000001111111 : node10000;
												assign node10000 = (inp[8]) ? node10006 : node10001;
													assign node10001 = (inp[12]) ? 15'b000000011111111 : node10002;
														assign node10002 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10006 = (inp[12]) ? 15'b000000001111111 : node10007;
														assign node10007 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10012 = (inp[10]) ? node10016 : node10013;
												assign node10013 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node10016 = (inp[14]) ? node10024 : node10017;
													assign node10017 = (inp[12]) ? 15'b000000000111111 : node10018;
														assign node10018 = (inp[2]) ? node10020 : 15'b000000001111111;
															assign node10020 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10024 = (inp[12]) ? 15'b000000000011111 : node10025;
														assign node10025 = (inp[8]) ? 15'b000000000011111 : node10026;
															assign node10026 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node10031 = (inp[14]) ? node10091 : node10032;
									assign node10032 = (inp[0]) ? node10058 : node10033;
										assign node10033 = (inp[8]) ? node10047 : node10034;
											assign node10034 = (inp[12]) ? node10042 : node10035;
												assign node10035 = (inp[2]) ? node10039 : node10036;
													assign node10036 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10039 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10042 = (inp[13]) ? 15'b000000011111111 : node10043;
													assign node10043 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10047 = (inp[13]) ? node10051 : node10048;
												assign node10048 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10051 = (inp[11]) ? 15'b000000000111111 : node10052;
													assign node10052 = (inp[2]) ? node10054 : 15'b000000001111111;
														assign node10054 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10058 = (inp[2]) ? node10072 : node10059;
											assign node10059 = (inp[12]) ? node10065 : node10060;
												assign node10060 = (inp[13]) ? node10062 : 15'b000000011111111;
													assign node10062 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10065 = (inp[13]) ? node10067 : 15'b000000001111111;
													assign node10067 = (inp[10]) ? 15'b000000001111111 : node10068;
														assign node10068 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10072 = (inp[12]) ? node10084 : node10073;
												assign node10073 = (inp[8]) ? node10081 : node10074;
													assign node10074 = (inp[13]) ? 15'b000000001111111 : node10075;
														assign node10075 = (inp[10]) ? node10077 : 15'b000000011111111;
															assign node10077 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10081 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10084 = (inp[11]) ? 15'b000000000011111 : node10085;
													assign node10085 = (inp[8]) ? 15'b000000000111111 : node10086;
														assign node10086 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node10091 = (inp[11]) ? node10113 : node10092;
										assign node10092 = (inp[10]) ? node10106 : node10093;
											assign node10093 = (inp[8]) ? node10101 : node10094;
												assign node10094 = (inp[13]) ? 15'b000000011111111 : node10095;
													assign node10095 = (inp[0]) ? 15'b000000011111111 : node10096;
														assign node10096 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10101 = (inp[12]) ? 15'b000000000111111 : node10102;
													assign node10102 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10106 = (inp[0]) ? node10108 : 15'b000000001111111;
												assign node10108 = (inp[12]) ? node10110 : 15'b000000000111111;
													assign node10110 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node10113 = (inp[8]) ? node10131 : node10114;
											assign node10114 = (inp[13]) ? node10122 : node10115;
												assign node10115 = (inp[12]) ? node10119 : node10116;
													assign node10116 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10119 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10122 = (inp[12]) ? node10128 : node10123;
													assign node10123 = (inp[10]) ? 15'b000000000111111 : node10124;
														assign node10124 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10128 = (inp[2]) ? 15'b000000000111111 : 15'b000000000011111;
											assign node10131 = (inp[0]) ? node10143 : node10132;
												assign node10132 = (inp[2]) ? node10136 : node10133;
													assign node10133 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10136 = (inp[13]) ? node10138 : 15'b000000000111111;
														assign node10138 = (inp[12]) ? node10140 : 15'b000000000111111;
															assign node10140 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10143 = (inp[10]) ? node10151 : node10144;
													assign node10144 = (inp[13]) ? node10146 : 15'b000000000111111;
														assign node10146 = (inp[2]) ? 15'b000000000011111 : node10147;
															assign node10147 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10151 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node10154 = (inp[12]) ? node10286 : node10155;
								assign node10155 = (inp[14]) ? node10221 : node10156;
									assign node10156 = (inp[8]) ? node10188 : node10157;
										assign node10157 = (inp[2]) ? node10169 : node10158;
											assign node10158 = (inp[0]) ? 15'b000000011111111 : node10159;
												assign node10159 = (inp[10]) ? node10161 : 15'b000000111111111;
													assign node10161 = (inp[5]) ? 15'b000000011111111 : node10162;
														assign node10162 = (inp[11]) ? node10164 : 15'b000000111111111;
															assign node10164 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10169 = (inp[10]) ? node10181 : node10170;
												assign node10170 = (inp[13]) ? node10178 : node10171;
													assign node10171 = (inp[11]) ? node10173 : 15'b000000111111111;
														assign node10173 = (inp[5]) ? 15'b000000011111111 : node10174;
															assign node10174 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10178 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10181 = (inp[11]) ? node10185 : node10182;
													assign node10182 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10185 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10188 = (inp[5]) ? node10204 : node10189;
											assign node10189 = (inp[11]) ? node10199 : node10190;
												assign node10190 = (inp[0]) ? 15'b000000001111111 : node10191;
													assign node10191 = (inp[10]) ? node10193 : 15'b000000111111111;
														assign node10193 = (inp[2]) ? 15'b000000011111111 : node10194;
															assign node10194 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10199 = (inp[10]) ? 15'b000000001111111 : node10200;
													assign node10200 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10204 = (inp[2]) ? node10214 : node10205;
												assign node10205 = (inp[13]) ? node10207 : 15'b000000011111111;
													assign node10207 = (inp[11]) ? node10209 : 15'b000000001111111;
														assign node10209 = (inp[10]) ? 15'b000000000111111 : node10210;
															assign node10210 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10214 = (inp[10]) ? node10216 : 15'b000000001111111;
													assign node10216 = (inp[11]) ? 15'b000000000011111 : node10217;
														assign node10217 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node10221 = (inp[10]) ? node10255 : node10222;
										assign node10222 = (inp[13]) ? node10242 : node10223;
											assign node10223 = (inp[8]) ? node10233 : node10224;
												assign node10224 = (inp[11]) ? node10226 : 15'b000000011111111;
													assign node10226 = (inp[2]) ? 15'b000000001111111 : node10227;
														assign node10227 = (inp[0]) ? 15'b000000001111111 : node10228;
															assign node10228 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10233 = (inp[5]) ? node10237 : node10234;
													assign node10234 = (inp[0]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node10237 = (inp[0]) ? node10239 : 15'b000000001111111;
														assign node10239 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10242 = (inp[5]) ? node10248 : node10243;
												assign node10243 = (inp[11]) ? node10245 : 15'b000000001111111;
													assign node10245 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10248 = (inp[2]) ? 15'b000000000111111 : node10249;
													assign node10249 = (inp[11]) ? node10251 : 15'b000000011111111;
														assign node10251 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10255 = (inp[8]) ? node10271 : node10256;
											assign node10256 = (inp[2]) ? node10266 : node10257;
												assign node10257 = (inp[5]) ? node10259 : 15'b000000001111111;
													assign node10259 = (inp[13]) ? node10261 : 15'b000000001111111;
														assign node10261 = (inp[11]) ? 15'b000000000111111 : node10262;
															assign node10262 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10266 = (inp[5]) ? 15'b000000000111111 : node10267;
													assign node10267 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10271 = (inp[13]) ? node10279 : node10272;
												assign node10272 = (inp[0]) ? node10276 : node10273;
													assign node10273 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10276 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10279 = (inp[0]) ? 15'b000000000001111 : node10280;
													assign node10280 = (inp[2]) ? node10282 : 15'b000000000111111;
														assign node10282 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node10286 = (inp[10]) ? node10348 : node10287;
									assign node10287 = (inp[2]) ? node10323 : node10288;
										assign node10288 = (inp[14]) ? node10306 : node10289;
											assign node10289 = (inp[5]) ? node10295 : node10290;
												assign node10290 = (inp[0]) ? 15'b000000011111111 : node10291;
													assign node10291 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10295 = (inp[0]) ? node10301 : node10296;
													assign node10296 = (inp[13]) ? node10298 : 15'b000000011111111;
														assign node10298 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10301 = (inp[13]) ? 15'b000000000111111 : node10302;
														assign node10302 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10306 = (inp[0]) ? node10314 : node10307;
												assign node10307 = (inp[5]) ? node10311 : node10308;
													assign node10308 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10311 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10314 = (inp[13]) ? node10320 : node10315;
													assign node10315 = (inp[5]) ? node10317 : 15'b000000001111111;
														assign node10317 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10320 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node10323 = (inp[5]) ? node10335 : node10324;
											assign node10324 = (inp[11]) ? node10330 : node10325;
												assign node10325 = (inp[14]) ? 15'b000000001111111 : node10326;
													assign node10326 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10330 = (inp[0]) ? node10332 : 15'b000000001111111;
													assign node10332 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10335 = (inp[11]) ? node10343 : node10336;
												assign node10336 = (inp[8]) ? 15'b000000000011111 : node10337;
													assign node10337 = (inp[0]) ? node10339 : 15'b000000000111111;
														assign node10339 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10343 = (inp[0]) ? node10345 : 15'b000000000011111;
													assign node10345 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node10348 = (inp[8]) ? node10374 : node10349;
										assign node10349 = (inp[2]) ? node10361 : node10350;
											assign node10350 = (inp[13]) ? node10356 : node10351;
												assign node10351 = (inp[14]) ? 15'b000000001111111 : node10352;
													assign node10352 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10356 = (inp[0]) ? 15'b000000000111111 : node10357;
													assign node10357 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10361 = (inp[13]) ? node10365 : node10362;
												assign node10362 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10365 = (inp[0]) ? node10371 : node10366;
													assign node10366 = (inp[14]) ? 15'b000000000011111 : node10367;
														assign node10367 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10371 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node10374 = (inp[14]) ? node10394 : node10375;
											assign node10375 = (inp[0]) ? node10387 : node10376;
												assign node10376 = (inp[5]) ? node10384 : node10377;
													assign node10377 = (inp[11]) ? node10379 : 15'b000000001111111;
														assign node10379 = (inp[2]) ? 15'b000000000111111 : node10380;
															assign node10380 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10384 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10387 = (inp[13]) ? node10391 : node10388;
													assign node10388 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10391 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node10394 = (inp[5]) ? node10408 : node10395;
												assign node10395 = (inp[2]) ? node10401 : node10396;
													assign node10396 = (inp[11]) ? 15'b000000000011111 : node10397;
														assign node10397 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10401 = (inp[0]) ? node10403 : 15'b000000000011111;
														assign node10403 = (inp[13]) ? 15'b000000000001111 : node10404;
															assign node10404 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node10408 = (inp[0]) ? node10412 : node10409;
													assign node10409 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node10412 = (inp[13]) ? node10414 : 15'b000000000011111;
														assign node10414 = (inp[2]) ? 15'b000000000000111 : node10415;
															assign node10415 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
				assign node10419 = (inp[10]) ? node11465 : node10420;
					assign node10420 = (inp[13]) ? node10974 : node10421;
						assign node10421 = (inp[11]) ? node10699 : node10422;
							assign node10422 = (inp[2]) ? node10564 : node10423;
								assign node10423 = (inp[3]) ? node10493 : node10424;
									assign node10424 = (inp[6]) ? node10464 : node10425;
										assign node10425 = (inp[0]) ? node10443 : node10426;
											assign node10426 = (inp[14]) ? node10438 : node10427;
												assign node10427 = (inp[8]) ? node10435 : node10428;
													assign node10428 = (inp[1]) ? node10430 : 15'b000111111111111;
														assign node10430 = (inp[12]) ? 15'b000011111111111 : node10431;
															assign node10431 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node10435 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node10438 = (inp[8]) ? node10440 : 15'b000001111111111;
													assign node10440 = (inp[12]) ? 15'b000000111111111 : 15'b000011111111111;
											assign node10443 = (inp[12]) ? node10449 : node10444;
												assign node10444 = (inp[8]) ? 15'b000001111111111 : node10445;
													assign node10445 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node10449 = (inp[1]) ? node10457 : node10450;
													assign node10450 = (inp[8]) ? node10452 : 15'b000001111111111;
														assign node10452 = (inp[14]) ? 15'b000000111111111 : node10453;
															assign node10453 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10457 = (inp[8]) ? 15'b000000011111111 : node10458;
														assign node10458 = (inp[5]) ? 15'b000000111111111 : node10459;
															assign node10459 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
										assign node10464 = (inp[12]) ? node10480 : node10465;
											assign node10465 = (inp[1]) ? node10475 : node10466;
												assign node10466 = (inp[5]) ? node10470 : node10467;
													assign node10467 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node10470 = (inp[0]) ? 15'b000000011111111 : node10471;
														assign node10471 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10475 = (inp[5]) ? node10477 : 15'b000000111111111;
													assign node10477 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10480 = (inp[14]) ? node10488 : node10481;
												assign node10481 = (inp[5]) ? node10485 : node10482;
													assign node10482 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10485 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10488 = (inp[5]) ? node10490 : 15'b000000011111111;
													assign node10490 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node10493 = (inp[0]) ? node10537 : node10494;
										assign node10494 = (inp[1]) ? node10518 : node10495;
											assign node10495 = (inp[14]) ? node10507 : node10496;
												assign node10496 = (inp[6]) ? node10504 : node10497;
													assign node10497 = (inp[12]) ? 15'b000001111111111 : node10498;
														assign node10498 = (inp[5]) ? node10500 : 15'b000011111111111;
															assign node10500 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node10504 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10507 = (inp[12]) ? node10509 : 15'b000001111111111;
													assign node10509 = (inp[8]) ? node10513 : node10510;
														assign node10510 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node10513 = (inp[6]) ? 15'b000000011111111 : node10514;
															assign node10514 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10518 = (inp[12]) ? node10526 : node10519;
												assign node10519 = (inp[5]) ? node10523 : node10520;
													assign node10520 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10523 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node10526 = (inp[5]) ? 15'b000000001111111 : node10527;
													assign node10527 = (inp[8]) ? node10531 : node10528;
														assign node10528 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node10531 = (inp[6]) ? node10533 : 15'b000000011111111;
															assign node10533 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node10537 = (inp[5]) ? node10551 : node10538;
											assign node10538 = (inp[6]) ? node10544 : node10539;
												assign node10539 = (inp[14]) ? node10541 : 15'b000000111111111;
													assign node10541 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10544 = (inp[14]) ? node10546 : 15'b000000001111111;
													assign node10546 = (inp[8]) ? 15'b000000011111111 : node10547;
														assign node10547 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10551 = (inp[12]) ? node10553 : 15'b000000011111111;
												assign node10553 = (inp[14]) ? node10561 : node10554;
													assign node10554 = (inp[8]) ? node10556 : 15'b000000011111111;
														assign node10556 = (inp[6]) ? 15'b000000001111111 : node10557;
															assign node10557 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10561 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node10564 = (inp[8]) ? node10640 : node10565;
									assign node10565 = (inp[1]) ? node10593 : node10566;
										assign node10566 = (inp[6]) ? node10582 : node10567;
											assign node10567 = (inp[12]) ? node10573 : node10568;
												assign node10568 = (inp[5]) ? node10570 : 15'b000001111111111;
													assign node10570 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10573 = (inp[3]) ? node10577 : node10574;
													assign node10574 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10577 = (inp[0]) ? node10579 : 15'b000000111111111;
														assign node10579 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10582 = (inp[5]) ? node10586 : node10583;
												assign node10583 = (inp[14]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node10586 = (inp[12]) ? 15'b000000011111111 : node10587;
													assign node10587 = (inp[14]) ? node10589 : 15'b000000111111111;
														assign node10589 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node10593 = (inp[5]) ? node10613 : node10594;
											assign node10594 = (inp[12]) ? node10602 : node10595;
												assign node10595 = (inp[6]) ? node10599 : node10596;
													assign node10596 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10599 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10602 = (inp[14]) ? node10604 : 15'b000000111111111;
													assign node10604 = (inp[6]) ? node10610 : node10605;
														assign node10605 = (inp[3]) ? 15'b000000011111111 : node10606;
															assign node10606 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node10610 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10613 = (inp[0]) ? node10627 : node10614;
												assign node10614 = (inp[3]) ? node10622 : node10615;
													assign node10615 = (inp[6]) ? node10619 : node10616;
														assign node10616 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node10619 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10622 = (inp[6]) ? node10624 : 15'b000000011111111;
														assign node10624 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10627 = (inp[3]) ? node10635 : node10628;
													assign node10628 = (inp[12]) ? node10630 : 15'b000000011111111;
														assign node10630 = (inp[14]) ? 15'b000000001111111 : node10631;
															assign node10631 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10635 = (inp[6]) ? 15'b000000000011111 : node10636;
														assign node10636 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node10640 = (inp[3]) ? node10672 : node10641;
										assign node10641 = (inp[5]) ? node10655 : node10642;
											assign node10642 = (inp[12]) ? node10648 : node10643;
												assign node10643 = (inp[1]) ? 15'b000000111111111 : node10644;
													assign node10644 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10648 = (inp[6]) ? node10652 : node10649;
													assign node10649 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10652 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10655 = (inp[12]) ? node10667 : node10656;
												assign node10656 = (inp[14]) ? node10662 : node10657;
													assign node10657 = (inp[0]) ? 15'b000000011111111 : node10658;
														assign node10658 = (inp[1]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node10662 = (inp[1]) ? node10664 : 15'b000000011111111;
														assign node10664 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10667 = (inp[0]) ? node10669 : 15'b000000001111111;
													assign node10669 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node10672 = (inp[12]) ? node10686 : node10673;
											assign node10673 = (inp[1]) ? node10679 : node10674;
												assign node10674 = (inp[6]) ? node10676 : 15'b000000011111111;
													assign node10676 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10679 = (inp[14]) ? node10681 : 15'b000000011111111;
													assign node10681 = (inp[5]) ? node10683 : 15'b000000001111111;
														assign node10683 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10686 = (inp[14]) ? node10694 : node10687;
												assign node10687 = (inp[1]) ? node10689 : 15'b000000001111111;
													assign node10689 = (inp[6]) ? node10691 : 15'b000000001111111;
														assign node10691 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10694 = (inp[0]) ? node10696 : 15'b000000001111111;
													assign node10696 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node10699 = (inp[2]) ? node10833 : node10700;
								assign node10700 = (inp[5]) ? node10766 : node10701;
									assign node10701 = (inp[6]) ? node10731 : node10702;
										assign node10702 = (inp[0]) ? node10714 : node10703;
											assign node10703 = (inp[1]) ? node10709 : node10704;
												assign node10704 = (inp[8]) ? 15'b000001111111111 : node10705;
													assign node10705 = (inp[3]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node10709 = (inp[12]) ? 15'b000000111111111 : node10710;
													assign node10710 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node10714 = (inp[1]) ? node10728 : node10715;
												assign node10715 = (inp[8]) ? node10723 : node10716;
													assign node10716 = (inp[12]) ? 15'b000000111111111 : node10717;
														assign node10717 = (inp[3]) ? node10719 : 15'b000001111111111;
															assign node10719 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10723 = (inp[14]) ? 15'b000000011111111 : node10724;
														assign node10724 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10728 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node10731 = (inp[8]) ? node10743 : node10732;
											assign node10732 = (inp[3]) ? node10738 : node10733;
												assign node10733 = (inp[14]) ? node10735 : 15'b000001111111111;
													assign node10735 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10738 = (inp[1]) ? 15'b000000011111111 : node10739;
													assign node10739 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10743 = (inp[12]) ? node10759 : node10744;
												assign node10744 = (inp[0]) ? node10750 : node10745;
													assign node10745 = (inp[3]) ? 15'b000000011111111 : node10746;
														assign node10746 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10750 = (inp[14]) ? node10754 : node10751;
														assign node10751 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node10754 = (inp[1]) ? 15'b000000001111111 : node10755;
															assign node10755 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10759 = (inp[3]) ? 15'b000000000111111 : node10760;
													assign node10760 = (inp[14]) ? node10762 : 15'b000000011111111;
														assign node10762 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node10766 = (inp[12]) ? node10798 : node10767;
										assign node10767 = (inp[0]) ? node10783 : node10768;
											assign node10768 = (inp[3]) ? node10778 : node10769;
												assign node10769 = (inp[1]) ? node10775 : node10770;
													assign node10770 = (inp[6]) ? 15'b000000111111111 : node10771;
														assign node10771 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10775 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10778 = (inp[1]) ? 15'b000000011111111 : node10779;
													assign node10779 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10783 = (inp[1]) ? node10793 : node10784;
												assign node10784 = (inp[14]) ? node10788 : node10785;
													assign node10785 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10788 = (inp[6]) ? node10790 : 15'b000000011111111;
														assign node10790 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10793 = (inp[6]) ? 15'b000000000011111 : node10794;
													assign node10794 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node10798 = (inp[14]) ? node10814 : node10799;
											assign node10799 = (inp[8]) ? node10809 : node10800;
												assign node10800 = (inp[3]) ? node10802 : 15'b000000111111111;
													assign node10802 = (inp[1]) ? node10804 : 15'b000000011111111;
														assign node10804 = (inp[0]) ? 15'b000000001111111 : node10805;
															assign node10805 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10809 = (inp[0]) ? 15'b000000001111111 : node10810;
													assign node10810 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node10814 = (inp[3]) ? node10826 : node10815;
												assign node10815 = (inp[8]) ? node10821 : node10816;
													assign node10816 = (inp[6]) ? 15'b000000001111111 : node10817;
														assign node10817 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10821 = (inp[1]) ? node10823 : 15'b000000001111111;
														assign node10823 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10826 = (inp[1]) ? node10830 : node10827;
													assign node10827 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node10830 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node10833 = (inp[1]) ? node10895 : node10834;
									assign node10834 = (inp[0]) ? node10860 : node10835;
										assign node10835 = (inp[8]) ? node10845 : node10836;
											assign node10836 = (inp[12]) ? 15'b000000011111111 : node10837;
												assign node10837 = (inp[14]) ? node10841 : node10838;
													assign node10838 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10841 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10845 = (inp[3]) ? node10853 : node10846;
												assign node10846 = (inp[5]) ? 15'b000000001111111 : node10847;
													assign node10847 = (inp[12]) ? node10849 : 15'b000000111111111;
														assign node10849 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node10853 = (inp[6]) ? 15'b000000001111111 : node10854;
													assign node10854 = (inp[5]) ? 15'b000000001111111 : node10855;
														assign node10855 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node10860 = (inp[3]) ? node10882 : node10861;
											assign node10861 = (inp[6]) ? node10871 : node10862;
												assign node10862 = (inp[5]) ? node10866 : node10863;
													assign node10863 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10866 = (inp[12]) ? 15'b000000001111111 : node10867;
														assign node10867 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10871 = (inp[14]) ? node10877 : node10872;
													assign node10872 = (inp[12]) ? 15'b000000001111111 : node10873;
														assign node10873 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10877 = (inp[5]) ? node10879 : 15'b000000001111111;
														assign node10879 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node10882 = (inp[12]) ? node10888 : node10883;
												assign node10883 = (inp[14]) ? node10885 : 15'b000000001111111;
													assign node10885 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10888 = (inp[5]) ? node10890 : 15'b000000001111111;
													assign node10890 = (inp[14]) ? node10892 : 15'b000000000011111;
														assign node10892 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node10895 = (inp[6]) ? node10937 : node10896;
										assign node10896 = (inp[3]) ? node10918 : node10897;
											assign node10897 = (inp[14]) ? node10905 : node10898;
												assign node10898 = (inp[8]) ? node10902 : node10899;
													assign node10899 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node10902 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node10905 = (inp[0]) ? node10913 : node10906;
													assign node10906 = (inp[8]) ? 15'b000000001111111 : node10907;
														assign node10907 = (inp[12]) ? node10909 : 15'b000000011111111;
															assign node10909 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10913 = (inp[8]) ? 15'b000000000111111 : node10914;
														assign node10914 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10918 = (inp[5]) ? node10932 : node10919;
												assign node10919 = (inp[0]) ? node10921 : 15'b000000001111111;
													assign node10921 = (inp[14]) ? node10927 : node10922;
														assign node10922 = (inp[8]) ? node10924 : 15'b000000001111111;
															assign node10924 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
														assign node10927 = (inp[8]) ? 15'b000000000111111 : node10928;
															assign node10928 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10932 = (inp[12]) ? node10934 : 15'b000000000111111;
													assign node10934 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node10937 = (inp[5]) ? node10957 : node10938;
											assign node10938 = (inp[0]) ? node10948 : node10939;
												assign node10939 = (inp[3]) ? node10945 : node10940;
													assign node10940 = (inp[8]) ? 15'b000000001111111 : node10941;
														assign node10941 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node10945 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node10948 = (inp[8]) ? node10952 : node10949;
													assign node10949 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node10952 = (inp[3]) ? 15'b000000000111111 : node10953;
														assign node10953 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node10957 = (inp[8]) ? node10967 : node10958;
												assign node10958 = (inp[0]) ? node10960 : 15'b000000000111111;
													assign node10960 = (inp[12]) ? node10962 : 15'b000000000111111;
														assign node10962 = (inp[3]) ? 15'b000000000011111 : node10963;
															assign node10963 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node10967 = (inp[14]) ? node10971 : node10968;
													assign node10968 = (inp[12]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node10971 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node10974 = (inp[8]) ? node11202 : node10975;
							assign node10975 = (inp[5]) ? node11093 : node10976;
								assign node10976 = (inp[3]) ? node11034 : node10977;
									assign node10977 = (inp[6]) ? node11005 : node10978;
										assign node10978 = (inp[1]) ? node10998 : node10979;
											assign node10979 = (inp[2]) ? node10987 : node10980;
												assign node10980 = (inp[0]) ? node10984 : node10981;
													assign node10981 = (inp[11]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node10984 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node10987 = (inp[14]) ? node10995 : node10988;
													assign node10988 = (inp[0]) ? 15'b000000111111111 : node10989;
														assign node10989 = (inp[11]) ? node10991 : 15'b000001111111111;
															assign node10991 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node10995 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node10998 = (inp[12]) ? 15'b000000011111111 : node10999;
												assign node10999 = (inp[0]) ? node11001 : 15'b000000111111111;
													assign node11001 = (inp[2]) ? 15'b000000001111111 : 15'b000000111111111;
										assign node11005 = (inp[0]) ? node11023 : node11006;
											assign node11006 = (inp[14]) ? node11016 : node11007;
												assign node11007 = (inp[11]) ? node11013 : node11008;
													assign node11008 = (inp[1]) ? 15'b000000111111111 : node11009;
														assign node11009 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11013 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11016 = (inp[12]) ? node11018 : 15'b000000011111111;
													assign node11018 = (inp[11]) ? node11020 : 15'b000000011111111;
														assign node11020 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11023 = (inp[2]) ? node11029 : node11024;
												assign node11024 = (inp[14]) ? node11026 : 15'b000000011111111;
													assign node11026 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11029 = (inp[11]) ? 15'b000000000111111 : node11030;
													assign node11030 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node11034 = (inp[12]) ? node11062 : node11035;
										assign node11035 = (inp[2]) ? node11041 : node11036;
											assign node11036 = (inp[0]) ? 15'b000000011111111 : node11037;
												assign node11037 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node11041 = (inp[11]) ? node11053 : node11042;
												assign node11042 = (inp[6]) ? node11050 : node11043;
													assign node11043 = (inp[14]) ? 15'b000000011111111 : node11044;
														assign node11044 = (inp[1]) ? node11046 : 15'b000000111111111;
															assign node11046 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11050 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11053 = (inp[0]) ? 15'b000000001111111 : node11054;
													assign node11054 = (inp[1]) ? node11056 : 15'b000000011111111;
														assign node11056 = (inp[6]) ? 15'b000000001111111 : node11057;
															assign node11057 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node11062 = (inp[2]) ? node11074 : node11063;
											assign node11063 = (inp[11]) ? node11071 : node11064;
												assign node11064 = (inp[6]) ? node11066 : 15'b000000111111111;
													assign node11066 = (inp[14]) ? 15'b000000011111111 : node11067;
														assign node11067 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11071 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11074 = (inp[1]) ? node11082 : node11075;
												assign node11075 = (inp[14]) ? node11079 : node11076;
													assign node11076 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11079 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11082 = (inp[0]) ? node11088 : node11083;
													assign node11083 = (inp[11]) ? 15'b000000000111111 : node11084;
														assign node11084 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11088 = (inp[14]) ? node11090 : 15'b000000000111111;
														assign node11090 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node11093 = (inp[2]) ? node11149 : node11094;
									assign node11094 = (inp[0]) ? node11122 : node11095;
										assign node11095 = (inp[3]) ? node11109 : node11096;
											assign node11096 = (inp[12]) ? node11104 : node11097;
												assign node11097 = (inp[6]) ? node11099 : 15'b000000111111111;
													assign node11099 = (inp[14]) ? 15'b000000111111111 : node11100;
														assign node11100 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node11104 = (inp[1]) ? node11106 : 15'b000000011111111;
													assign node11106 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11109 = (inp[14]) ? node11117 : node11110;
												assign node11110 = (inp[6]) ? node11112 : 15'b000000011111111;
													assign node11112 = (inp[11]) ? node11114 : 15'b000000011111111;
														assign node11114 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11117 = (inp[11]) ? node11119 : 15'b000000001111111;
													assign node11119 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node11122 = (inp[11]) ? node11138 : node11123;
											assign node11123 = (inp[1]) ? node11127 : node11124;
												assign node11124 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11127 = (inp[6]) ? node11135 : node11128;
													assign node11128 = (inp[3]) ? 15'b000000001111111 : node11129;
														assign node11129 = (inp[14]) ? node11131 : 15'b000000011111111;
															assign node11131 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11135 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11138 = (inp[12]) ? node11144 : node11139;
												assign node11139 = (inp[1]) ? node11141 : 15'b000000001111111;
													assign node11141 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11144 = (inp[14]) ? node11146 : 15'b000000000111111;
													assign node11146 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node11149 = (inp[14]) ? node11175 : node11150;
										assign node11150 = (inp[3]) ? node11160 : node11151;
											assign node11151 = (inp[12]) ? node11157 : node11152;
												assign node11152 = (inp[0]) ? 15'b000000011111111 : node11153;
													assign node11153 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11157 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11160 = (inp[11]) ? node11166 : node11161;
												assign node11161 = (inp[6]) ? node11163 : 15'b000000011111111;
													assign node11163 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11166 = (inp[0]) ? node11170 : node11167;
													assign node11167 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11170 = (inp[6]) ? node11172 : 15'b000000000111111;
														assign node11172 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11175 = (inp[1]) ? node11185 : node11176;
											assign node11176 = (inp[6]) ? 15'b000000000111111 : node11177;
												assign node11177 = (inp[12]) ? node11179 : 15'b000000001111111;
													assign node11179 = (inp[0]) ? node11181 : 15'b000000001111111;
														assign node11181 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11185 = (inp[3]) ? node11193 : node11186;
												assign node11186 = (inp[6]) ? node11190 : node11187;
													assign node11187 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11190 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11193 = (inp[12]) ? node11197 : node11194;
													assign node11194 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11197 = (inp[11]) ? node11199 : 15'b000000000011111;
														assign node11199 = (inp[6]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node11202 = (inp[11]) ? node11350 : node11203;
								assign node11203 = (inp[5]) ? node11273 : node11204;
									assign node11204 = (inp[2]) ? node11238 : node11205;
										assign node11205 = (inp[3]) ? node11219 : node11206;
											assign node11206 = (inp[1]) ? 15'b000000011111111 : node11207;
												assign node11207 = (inp[0]) ? node11211 : node11208;
													assign node11208 = (inp[14]) ? 15'b000001111111111 : 15'b000000111111111;
													assign node11211 = (inp[6]) ? 15'b000000011111111 : node11212;
														assign node11212 = (inp[14]) ? node11214 : 15'b000000111111111;
															assign node11214 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node11219 = (inp[14]) ? node11229 : node11220;
												assign node11220 = (inp[1]) ? node11224 : node11221;
													assign node11221 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11224 = (inp[6]) ? 15'b000000000111111 : node11225;
														assign node11225 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11229 = (inp[6]) ? 15'b000000001111111 : node11230;
													assign node11230 = (inp[12]) ? node11232 : 15'b000000011111111;
														assign node11232 = (inp[1]) ? 15'b000000001111111 : node11233;
															assign node11233 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node11238 = (inp[1]) ? node11250 : node11239;
											assign node11239 = (inp[0]) ? node11241 : 15'b000000011111111;
												assign node11241 = (inp[3]) ? 15'b000000000111111 : node11242;
													assign node11242 = (inp[12]) ? 15'b000000001111111 : node11243;
														assign node11243 = (inp[6]) ? node11245 : 15'b000000011111111;
															assign node11245 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11250 = (inp[14]) ? node11264 : node11251;
												assign node11251 = (inp[12]) ? node11257 : node11252;
													assign node11252 = (inp[3]) ? 15'b000000001111111 : node11253;
														assign node11253 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11257 = (inp[3]) ? 15'b000000000011111 : node11258;
														assign node11258 = (inp[0]) ? node11260 : 15'b000000001111111;
															assign node11260 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11264 = (inp[3]) ? node11268 : node11265;
													assign node11265 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11268 = (inp[6]) ? node11270 : 15'b000000000111111;
														assign node11270 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node11273 = (inp[14]) ? node11319 : node11274;
										assign node11274 = (inp[12]) ? node11294 : node11275;
											assign node11275 = (inp[6]) ? node11285 : node11276;
												assign node11276 = (inp[0]) ? 15'b000000011111111 : node11277;
													assign node11277 = (inp[3]) ? 15'b000000111111111 : node11278;
														assign node11278 = (inp[1]) ? 15'b000000111111111 : node11279;
															assign node11279 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node11285 = (inp[3]) ? node11291 : node11286;
													assign node11286 = (inp[1]) ? 15'b000000001111111 : node11287;
														assign node11287 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11291 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11294 = (inp[0]) ? node11308 : node11295;
												assign node11295 = (inp[1]) ? node11303 : node11296;
													assign node11296 = (inp[6]) ? node11298 : 15'b000000011111111;
														assign node11298 = (inp[2]) ? node11300 : 15'b000000001111111;
															assign node11300 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11303 = (inp[6]) ? 15'b000000000111111 : node11304;
														assign node11304 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11308 = (inp[1]) ? node11314 : node11309;
													assign node11309 = (inp[2]) ? 15'b000000000111111 : node11310;
														assign node11310 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11314 = (inp[2]) ? node11316 : 15'b000000000111111;
														assign node11316 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11319 = (inp[6]) ? node11337 : node11320;
											assign node11320 = (inp[0]) ? node11326 : node11321;
												assign node11321 = (inp[1]) ? node11323 : 15'b000000001111111;
													assign node11323 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11326 = (inp[2]) ? node11332 : node11327;
													assign node11327 = (inp[12]) ? 15'b000000000111111 : node11328;
														assign node11328 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11332 = (inp[1]) ? 15'b000000000011111 : node11333;
														assign node11333 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node11337 = (inp[0]) ? node11343 : node11338;
												assign node11338 = (inp[1]) ? node11340 : 15'b000000000111111;
													assign node11340 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11343 = (inp[2]) ? node11347 : node11344;
													assign node11344 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11347 = (inp[1]) ? 15'b000000000000111 : 15'b000000000011111;
								assign node11350 = (inp[6]) ? node11408 : node11351;
									assign node11351 = (inp[14]) ? node11383 : node11352;
										assign node11352 = (inp[0]) ? node11366 : node11353;
											assign node11353 = (inp[2]) ? node11359 : node11354;
												assign node11354 = (inp[1]) ? node11356 : 15'b000000011111111;
													assign node11356 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11359 = (inp[12]) ? node11363 : node11360;
													assign node11360 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11363 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11366 = (inp[5]) ? node11376 : node11367;
												assign node11367 = (inp[3]) ? 15'b000000000111111 : node11368;
													assign node11368 = (inp[1]) ? node11370 : 15'b000000011111111;
														assign node11370 = (inp[12]) ? 15'b000000001111111 : node11371;
															assign node11371 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11376 = (inp[1]) ? node11378 : 15'b000000000111111;
													assign node11378 = (inp[3]) ? 15'b000000000001111 : node11379;
														assign node11379 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11383 = (inp[3]) ? node11391 : node11384;
											assign node11384 = (inp[0]) ? 15'b000000000111111 : node11385;
												assign node11385 = (inp[1]) ? 15'b000000000111111 : node11386;
													assign node11386 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11391 = (inp[12]) ? node11401 : node11392;
												assign node11392 = (inp[5]) ? node11394 : 15'b000000000111111;
													assign node11394 = (inp[0]) ? 15'b000000000011111 : node11395;
														assign node11395 = (inp[2]) ? node11397 : 15'b000000000111111;
															assign node11397 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11401 = (inp[2]) ? node11405 : node11402;
													assign node11402 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11405 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node11408 = (inp[1]) ? node11426 : node11409;
										assign node11409 = (inp[2]) ? node11421 : node11410;
											assign node11410 = (inp[12]) ? node11416 : node11411;
												assign node11411 = (inp[3]) ? node11413 : 15'b000000011111111;
													assign node11413 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11416 = (inp[14]) ? 15'b000000000011111 : node11417;
													assign node11417 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11421 = (inp[12]) ? 15'b000000000011111 : node11422;
												assign node11422 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11426 = (inp[0]) ? node11448 : node11427;
											assign node11427 = (inp[3]) ? node11441 : node11428;
												assign node11428 = (inp[12]) ? node11436 : node11429;
													assign node11429 = (inp[5]) ? node11431 : 15'b000000001111111;
														assign node11431 = (inp[14]) ? node11433 : 15'b000000000111111;
															assign node11433 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11436 = (inp[2]) ? 15'b000000000011111 : node11437;
														assign node11437 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11441 = (inp[14]) ? node11445 : node11442;
													assign node11442 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11445 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node11448 = (inp[2]) ? node11456 : node11449;
												assign node11449 = (inp[12]) ? node11453 : node11450;
													assign node11450 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11453 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node11456 = (inp[3]) ? node11462 : node11457;
													assign node11457 = (inp[12]) ? 15'b000000000001111 : node11458;
														assign node11458 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node11462 = (inp[14]) ? 15'b000000000000011 : 15'b000000000001111;
					assign node11465 = (inp[8]) ? node12007 : node11466;
						assign node11466 = (inp[6]) ? node11732 : node11467;
							assign node11467 = (inp[0]) ? node11599 : node11468;
								assign node11468 = (inp[11]) ? node11532 : node11469;
									assign node11469 = (inp[12]) ? node11505 : node11470;
										assign node11470 = (inp[3]) ? node11484 : node11471;
											assign node11471 = (inp[5]) ? node11479 : node11472;
												assign node11472 = (inp[14]) ? 15'b000001111111111 : node11473;
													assign node11473 = (inp[2]) ? 15'b000001111111111 : node11474;
														assign node11474 = (inp[13]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node11479 = (inp[14]) ? 15'b000000111111111 : node11480;
													assign node11480 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node11484 = (inp[13]) ? node11500 : node11485;
												assign node11485 = (inp[1]) ? node11497 : node11486;
													assign node11486 = (inp[14]) ? node11492 : node11487;
														assign node11487 = (inp[2]) ? node11489 : 15'b000001111111111;
															assign node11489 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node11492 = (inp[2]) ? 15'b000000111111111 : node11493;
															assign node11493 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11497 = (inp[14]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node11500 = (inp[14]) ? 15'b000000011111111 : node11501;
													assign node11501 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node11505 = (inp[5]) ? node11521 : node11506;
											assign node11506 = (inp[2]) ? node11512 : node11507;
												assign node11507 = (inp[3]) ? 15'b000000111111111 : node11508;
													assign node11508 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node11512 = (inp[13]) ? 15'b000000001111111 : node11513;
													assign node11513 = (inp[14]) ? node11515 : 15'b000000111111111;
														assign node11515 = (inp[3]) ? 15'b000000011111111 : node11516;
															assign node11516 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node11521 = (inp[3]) ? node11527 : node11522;
												assign node11522 = (inp[13]) ? 15'b000000001111111 : node11523;
													assign node11523 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11527 = (inp[1]) ? node11529 : 15'b000000001111111;
													assign node11529 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node11532 = (inp[1]) ? node11572 : node11533;
										assign node11533 = (inp[12]) ? node11553 : node11534;
											assign node11534 = (inp[5]) ? node11544 : node11535;
												assign node11535 = (inp[14]) ? 15'b000000111111111 : node11536;
													assign node11536 = (inp[3]) ? node11538 : 15'b000011111111111;
														assign node11538 = (inp[13]) ? 15'b000000111111111 : node11539;
															assign node11539 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node11544 = (inp[13]) ? node11546 : 15'b000000111111111;
													assign node11546 = (inp[14]) ? 15'b000000001111111 : node11547;
														assign node11547 = (inp[2]) ? node11549 : 15'b000000011111111;
															assign node11549 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11553 = (inp[2]) ? node11565 : node11554;
												assign node11554 = (inp[3]) ? node11558 : node11555;
													assign node11555 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11558 = (inp[5]) ? node11560 : 15'b000000011111111;
														assign node11560 = (inp[14]) ? 15'b000000001111111 : node11561;
															assign node11561 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11565 = (inp[3]) ? 15'b000000000111111 : node11566;
													assign node11566 = (inp[5]) ? 15'b000000001111111 : node11567;
														assign node11567 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node11572 = (inp[14]) ? node11580 : node11573;
											assign node11573 = (inp[13]) ? node11575 : 15'b000000011111111;
												assign node11575 = (inp[2]) ? 15'b000000001111111 : node11576;
													assign node11576 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11580 = (inp[5]) ? node11588 : node11581;
												assign node11581 = (inp[2]) ? 15'b000000001111111 : node11582;
													assign node11582 = (inp[13]) ? node11584 : 15'b000000001111111;
														assign node11584 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11588 = (inp[2]) ? node11594 : node11589;
													assign node11589 = (inp[3]) ? node11591 : 15'b000000001111111;
														assign node11591 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11594 = (inp[12]) ? node11596 : 15'b000000000111111;
														assign node11596 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node11599 = (inp[11]) ? node11675 : node11600;
									assign node11600 = (inp[1]) ? node11646 : node11601;
										assign node11601 = (inp[2]) ? node11623 : node11602;
											assign node11602 = (inp[5]) ? node11612 : node11603;
												assign node11603 = (inp[14]) ? node11609 : node11604;
													assign node11604 = (inp[13]) ? node11606 : 15'b000001111111111;
														assign node11606 = (inp[12]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node11609 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11612 = (inp[13]) ? node11616 : node11613;
													assign node11613 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11616 = (inp[14]) ? node11618 : 15'b000000011111111;
														assign node11618 = (inp[3]) ? 15'b000000001111111 : node11619;
															assign node11619 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11623 = (inp[3]) ? node11631 : node11624;
												assign node11624 = (inp[14]) ? node11626 : 15'b000000011111111;
													assign node11626 = (inp[13]) ? node11628 : 15'b000000011111111;
														assign node11628 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11631 = (inp[13]) ? node11643 : node11632;
													assign node11632 = (inp[12]) ? node11638 : node11633;
														assign node11633 = (inp[5]) ? node11635 : 15'b000000011111111;
															assign node11635 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node11638 = (inp[14]) ? 15'b000000001111111 : node11639;
															assign node11639 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11643 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node11646 = (inp[5]) ? node11664 : node11647;
											assign node11647 = (inp[14]) ? node11653 : node11648;
												assign node11648 = (inp[2]) ? 15'b000000011111111 : node11649;
													assign node11649 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node11653 = (inp[2]) ? node11657 : node11654;
													assign node11654 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11657 = (inp[3]) ? 15'b000000000111111 : node11658;
														assign node11658 = (inp[12]) ? node11660 : 15'b000000001111111;
															assign node11660 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11664 = (inp[14]) ? node11672 : node11665;
												assign node11665 = (inp[12]) ? node11669 : node11666;
													assign node11666 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11669 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11672 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node11675 = (inp[13]) ? node11703 : node11676;
										assign node11676 = (inp[14]) ? node11694 : node11677;
											assign node11677 = (inp[3]) ? node11687 : node11678;
												assign node11678 = (inp[5]) ? node11684 : node11679;
													assign node11679 = (inp[2]) ? 15'b000000011111111 : node11680;
														assign node11680 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11684 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11687 = (inp[1]) ? node11691 : node11688;
													assign node11688 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11691 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11694 = (inp[12]) ? node11700 : node11695;
												assign node11695 = (inp[2]) ? node11697 : 15'b000000011111111;
													assign node11697 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11700 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11703 = (inp[2]) ? node11719 : node11704;
											assign node11704 = (inp[5]) ? node11714 : node11705;
												assign node11705 = (inp[14]) ? node11711 : node11706;
													assign node11706 = (inp[3]) ? 15'b000000001111111 : node11707;
														assign node11707 = (inp[12]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11711 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11714 = (inp[3]) ? node11716 : 15'b000000000111111;
													assign node11716 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node11719 = (inp[3]) ? node11727 : node11720;
												assign node11720 = (inp[14]) ? 15'b000000000011111 : node11721;
													assign node11721 = (inp[12]) ? node11723 : 15'b000000000111111;
														assign node11723 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11727 = (inp[14]) ? node11729 : 15'b000000000011111;
													assign node11729 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node11732 = (inp[1]) ? node11872 : node11733;
								assign node11733 = (inp[0]) ? node11797 : node11734;
									assign node11734 = (inp[12]) ? node11764 : node11735;
										assign node11735 = (inp[13]) ? node11747 : node11736;
											assign node11736 = (inp[5]) ? node11738 : 15'b000000111111111;
												assign node11738 = (inp[2]) ? node11742 : node11739;
													assign node11739 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11742 = (inp[11]) ? node11744 : 15'b000000011111111;
														assign node11744 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11747 = (inp[11]) ? node11757 : node11748;
												assign node11748 = (inp[3]) ? node11750 : 15'b000000011111111;
													assign node11750 = (inp[14]) ? 15'b000000001111111 : node11751;
														assign node11751 = (inp[2]) ? node11753 : 15'b000000011111111;
															assign node11753 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11757 = (inp[5]) ? 15'b000000001111111 : node11758;
													assign node11758 = (inp[14]) ? 15'b000000001111111 : node11759;
														assign node11759 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node11764 = (inp[5]) ? node11778 : node11765;
											assign node11765 = (inp[3]) ? node11773 : node11766;
												assign node11766 = (inp[13]) ? node11770 : node11767;
													assign node11767 = (inp[14]) ? 15'b000000011111111 : 15'b000001111111111;
													assign node11770 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11773 = (inp[11]) ? 15'b000000000111111 : node11774;
													assign node11774 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node11778 = (inp[14]) ? node11786 : node11779;
												assign node11779 = (inp[2]) ? node11781 : 15'b000000111111111;
													assign node11781 = (inp[11]) ? node11783 : 15'b000000001111111;
														assign node11783 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11786 = (inp[11]) ? node11794 : node11787;
													assign node11787 = (inp[13]) ? node11789 : 15'b000000001111111;
														assign node11789 = (inp[2]) ? 15'b000000000111111 : node11790;
															assign node11790 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11794 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node11797 = (inp[2]) ? node11831 : node11798;
										assign node11798 = (inp[5]) ? node11814 : node11799;
											assign node11799 = (inp[13]) ? node11805 : node11800;
												assign node11800 = (inp[11]) ? 15'b000000011111111 : node11801;
													assign node11801 = (inp[12]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node11805 = (inp[11]) ? node11809 : node11806;
													assign node11806 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11809 = (inp[14]) ? node11811 : 15'b000000001111111;
														assign node11811 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11814 = (inp[11]) ? node11826 : node11815;
												assign node11815 = (inp[14]) ? node11819 : node11816;
													assign node11816 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11819 = (inp[3]) ? node11821 : 15'b000000001111111;
														assign node11821 = (inp[13]) ? 15'b000000000111111 : node11822;
															assign node11822 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11826 = (inp[12]) ? node11828 : 15'b000000001111111;
													assign node11828 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11831 = (inp[14]) ? node11855 : node11832;
											assign node11832 = (inp[3]) ? node11842 : node11833;
												assign node11833 = (inp[13]) ? node11837 : node11834;
													assign node11834 = (inp[11]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node11837 = (inp[11]) ? node11839 : 15'b000000001111111;
														assign node11839 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11842 = (inp[12]) ? node11848 : node11843;
													assign node11843 = (inp[11]) ? node11845 : 15'b000000001111111;
														assign node11845 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11848 = (inp[13]) ? node11850 : 15'b000000000111111;
														assign node11850 = (inp[11]) ? 15'b000000000011111 : node11851;
															assign node11851 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node11855 = (inp[5]) ? node11865 : node11856;
												assign node11856 = (inp[13]) ? node11860 : node11857;
													assign node11857 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11860 = (inp[3]) ? node11862 : 15'b000000000111111;
														assign node11862 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11865 = (inp[13]) ? node11869 : node11866;
													assign node11866 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node11869 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node11872 = (inp[2]) ? node11946 : node11873;
									assign node11873 = (inp[11]) ? node11915 : node11874;
										assign node11874 = (inp[0]) ? node11896 : node11875;
											assign node11875 = (inp[14]) ? node11885 : node11876;
												assign node11876 = (inp[3]) ? node11882 : node11877;
													assign node11877 = (inp[13]) ? 15'b000000011111111 : node11878;
														assign node11878 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11882 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11885 = (inp[12]) ? node11893 : node11886;
													assign node11886 = (inp[13]) ? node11888 : 15'b000000011111111;
														assign node11888 = (inp[3]) ? 15'b000000001111111 : node11889;
															assign node11889 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node11893 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11896 = (inp[3]) ? node11906 : node11897;
												assign node11897 = (inp[12]) ? node11901 : node11898;
													assign node11898 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node11901 = (inp[5]) ? node11903 : 15'b000000001111111;
														assign node11903 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11906 = (inp[5]) ? node11910 : node11907;
													assign node11907 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11910 = (inp[14]) ? node11912 : 15'b000000000111111;
														assign node11912 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node11915 = (inp[14]) ? node11929 : node11916;
											assign node11916 = (inp[5]) ? node11918 : 15'b000000001111111;
												assign node11918 = (inp[0]) ? node11924 : node11919;
													assign node11919 = (inp[12]) ? node11921 : 15'b000000001111111;
														assign node11921 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11924 = (inp[12]) ? 15'b000000000011111 : node11925;
														assign node11925 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node11929 = (inp[3]) ? node11941 : node11930;
												assign node11930 = (inp[5]) ? node11936 : node11931;
													assign node11931 = (inp[0]) ? 15'b000000000111111 : node11932;
														assign node11932 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11936 = (inp[13]) ? 15'b000000000011111 : node11937;
														assign node11937 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node11941 = (inp[5]) ? 15'b000000000001111 : node11942;
													assign node11942 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node11946 = (inp[13]) ? node11980 : node11947;
										assign node11947 = (inp[5]) ? node11963 : node11948;
											assign node11948 = (inp[14]) ? node11956 : node11949;
												assign node11949 = (inp[11]) ? 15'b000000000111111 : node11950;
													assign node11950 = (inp[3]) ? 15'b000000001111111 : node11951;
														assign node11951 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node11956 = (inp[12]) ? node11960 : node11957;
													assign node11957 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11960 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node11963 = (inp[0]) ? node11975 : node11964;
												assign node11964 = (inp[3]) ? node11968 : node11965;
													assign node11965 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node11968 = (inp[14]) ? 15'b000000000011111 : node11969;
														assign node11969 = (inp[11]) ? node11971 : 15'b000000000111111;
															assign node11971 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11975 = (inp[14]) ? 15'b000000000001111 : node11976;
													assign node11976 = (inp[12]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node11980 = (inp[3]) ? node11992 : node11981;
											assign node11981 = (inp[5]) ? node11989 : node11982;
												assign node11982 = (inp[0]) ? node11984 : 15'b000000000111111;
													assign node11984 = (inp[14]) ? node11986 : 15'b000000000111111;
														assign node11986 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node11989 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node11992 = (inp[11]) ? node11998 : node11993;
												assign node11993 = (inp[0]) ? node11995 : 15'b000000000111111;
													assign node11995 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node11998 = (inp[12]) ? node12002 : node11999;
													assign node11999 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node12002 = (inp[14]) ? node12004 : 15'b000000000001111;
														assign node12004 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node12007 = (inp[5]) ? node12263 : node12008;
							assign node12008 = (inp[6]) ? node12134 : node12009;
								assign node12009 = (inp[0]) ? node12063 : node12010;
									assign node12010 = (inp[3]) ? node12044 : node12011;
										assign node12011 = (inp[12]) ? node12023 : node12012;
											assign node12012 = (inp[13]) ? node12014 : 15'b000000111111111;
												assign node12014 = (inp[14]) ? 15'b000000011111111 : node12015;
													assign node12015 = (inp[2]) ? node12017 : 15'b000000111111111;
														assign node12017 = (inp[1]) ? 15'b000000011111111 : node12018;
															assign node12018 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node12023 = (inp[14]) ? node12035 : node12024;
												assign node12024 = (inp[11]) ? node12032 : node12025;
													assign node12025 = (inp[13]) ? 15'b000000011111111 : node12026;
														assign node12026 = (inp[2]) ? 15'b000000111111111 : node12027;
															assign node12027 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12032 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12035 = (inp[11]) ? node12037 : 15'b000000001111111;
													assign node12037 = (inp[13]) ? node12039 : 15'b000000001111111;
														assign node12039 = (inp[1]) ? node12041 : 15'b000000000111111;
															assign node12041 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node12044 = (inp[12]) ? node12052 : node12045;
											assign node12045 = (inp[13]) ? 15'b000000001111111 : node12046;
												assign node12046 = (inp[1]) ? 15'b000000000111111 : node12047;
													assign node12047 = (inp[14]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node12052 = (inp[14]) ? node12058 : node12053;
												assign node12053 = (inp[1]) ? node12055 : 15'b000000011111111;
													assign node12055 = (inp[13]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node12058 = (inp[2]) ? node12060 : 15'b000000000111111;
													assign node12060 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node12063 = (inp[1]) ? node12105 : node12064;
										assign node12064 = (inp[11]) ? node12082 : node12065;
											assign node12065 = (inp[14]) ? node12075 : node12066;
												assign node12066 = (inp[12]) ? node12072 : node12067;
													assign node12067 = (inp[2]) ? node12069 : 15'b000000111111111;
														assign node12069 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12072 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12075 = (inp[2]) ? 15'b000000000111111 : node12076;
													assign node12076 = (inp[13]) ? 15'b000000001111111 : node12077;
														assign node12077 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12082 = (inp[12]) ? node12094 : node12083;
												assign node12083 = (inp[3]) ? node12091 : node12084;
													assign node12084 = (inp[13]) ? node12086 : 15'b000000001111111;
														assign node12086 = (inp[2]) ? node12088 : 15'b000000001111111;
															assign node12088 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12091 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12094 = (inp[3]) ? node12102 : node12095;
													assign node12095 = (inp[2]) ? 15'b000000000111111 : node12096;
														assign node12096 = (inp[14]) ? node12098 : 15'b000000001111111;
															assign node12098 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12102 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node12105 = (inp[14]) ? node12119 : node12106;
											assign node12106 = (inp[2]) ? node12108 : 15'b000000001111111;
												assign node12108 = (inp[13]) ? node12112 : node12109;
													assign node12109 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12112 = (inp[11]) ? 15'b000000000011111 : node12113;
														assign node12113 = (inp[3]) ? 15'b000000000111111 : node12114;
															assign node12114 = (inp[12]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12119 = (inp[12]) ? node12129 : node12120;
												assign node12120 = (inp[2]) ? node12126 : node12121;
													assign node12121 = (inp[3]) ? 15'b000000000111111 : node12122;
														assign node12122 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12126 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12129 = (inp[2]) ? node12131 : 15'b000000000011111;
													assign node12131 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node12134 = (inp[13]) ? node12194 : node12135;
									assign node12135 = (inp[3]) ? node12167 : node12136;
										assign node12136 = (inp[0]) ? node12154 : node12137;
											assign node12137 = (inp[11]) ? node12145 : node12138;
												assign node12138 = (inp[1]) ? node12142 : node12139;
													assign node12139 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12142 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12145 = (inp[14]) ? node12149 : node12146;
													assign node12146 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12149 = (inp[1]) ? node12151 : 15'b000000001111111;
														assign node12151 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12154 = (inp[11]) ? node12162 : node12155;
												assign node12155 = (inp[1]) ? 15'b000000000111111 : node12156;
													assign node12156 = (inp[14]) ? 15'b000000001111111 : node12157;
														assign node12157 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12162 = (inp[1]) ? node12164 : 15'b000000000111111;
													assign node12164 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node12167 = (inp[2]) ? node12177 : node12168;
											assign node12168 = (inp[11]) ? node12172 : node12169;
												assign node12169 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12172 = (inp[1]) ? 15'b000000000111111 : node12173;
													assign node12173 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node12177 = (inp[12]) ? node12185 : node12178;
												assign node12178 = (inp[1]) ? node12182 : node12179;
													assign node12179 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12182 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12185 = (inp[0]) ? 15'b000000000001111 : node12186;
													assign node12186 = (inp[14]) ? node12188 : 15'b000000000111111;
														assign node12188 = (inp[1]) ? 15'b000000000011111 : node12189;
															assign node12189 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node12194 = (inp[12]) ? node12226 : node12195;
										assign node12195 = (inp[2]) ? node12215 : node12196;
											assign node12196 = (inp[0]) ? node12208 : node12197;
												assign node12197 = (inp[3]) ? node12203 : node12198;
													assign node12198 = (inp[11]) ? node12200 : 15'b000000011111111;
														assign node12200 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12203 = (inp[14]) ? node12205 : 15'b000000001111111;
														assign node12205 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12208 = (inp[11]) ? node12212 : node12209;
													assign node12209 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12212 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12215 = (inp[11]) ? node12221 : node12216;
												assign node12216 = (inp[0]) ? node12218 : 15'b000000000111111;
													assign node12218 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12221 = (inp[0]) ? 15'b000000000011111 : node12222;
													assign node12222 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node12226 = (inp[11]) ? node12246 : node12227;
											assign node12227 = (inp[2]) ? node12235 : node12228;
												assign node12228 = (inp[3]) ? node12232 : node12229;
													assign node12229 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12232 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12235 = (inp[1]) ? node12241 : node12236;
													assign node12236 = (inp[0]) ? 15'b000000000011111 : node12237;
														assign node12237 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node12241 = (inp[14]) ? 15'b000000000001111 : node12242;
														assign node12242 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node12246 = (inp[3]) ? node12256 : node12247;
												assign node12247 = (inp[2]) ? node12249 : 15'b000000000011111;
													assign node12249 = (inp[1]) ? node12251 : 15'b000000000011111;
														assign node12251 = (inp[0]) ? 15'b000000000001111 : node12252;
															assign node12252 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node12256 = (inp[0]) ? node12258 : 15'b000000000001111;
													assign node12258 = (inp[2]) ? node12260 : 15'b000000000001111;
														assign node12260 = (inp[14]) ? 15'b000000000000011 : 15'b000000000000111;
							assign node12263 = (inp[0]) ? node12389 : node12264;
								assign node12264 = (inp[1]) ? node12334 : node12265;
									assign node12265 = (inp[2]) ? node12291 : node12266;
										assign node12266 = (inp[14]) ? node12282 : node12267;
											assign node12267 = (inp[13]) ? node12279 : node12268;
												assign node12268 = (inp[6]) ? node12274 : node12269;
													assign node12269 = (inp[11]) ? 15'b000000111111111 : node12270;
														assign node12270 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12274 = (inp[3]) ? node12276 : 15'b000000011111111;
														assign node12276 = (inp[12]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12279 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12282 = (inp[3]) ? node12286 : node12283;
												assign node12283 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node12286 = (inp[11]) ? 15'b000000000111111 : node12287;
													assign node12287 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node12291 = (inp[14]) ? node12315 : node12292;
											assign node12292 = (inp[3]) ? node12304 : node12293;
												assign node12293 = (inp[11]) ? node12301 : node12294;
													assign node12294 = (inp[12]) ? 15'b000000001111111 : node12295;
														assign node12295 = (inp[6]) ? 15'b000000011111111 : node12296;
															assign node12296 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12301 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12304 = (inp[11]) ? node12312 : node12305;
													assign node12305 = (inp[12]) ? node12307 : 15'b000000001111111;
														assign node12307 = (inp[6]) ? 15'b000000000111111 : node12308;
															assign node12308 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12312 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12315 = (inp[11]) ? node12327 : node12316;
												assign node12316 = (inp[12]) ? node12320 : node12317;
													assign node12317 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12320 = (inp[3]) ? node12322 : 15'b000000000111111;
														assign node12322 = (inp[13]) ? 15'b000000000011111 : node12323;
															assign node12323 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12327 = (inp[3]) ? node12331 : node12328;
													assign node12328 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node12331 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node12334 = (inp[14]) ? node12364 : node12335;
										assign node12335 = (inp[2]) ? node12349 : node12336;
											assign node12336 = (inp[13]) ? node12342 : node12337;
												assign node12337 = (inp[11]) ? node12339 : 15'b000000001111111;
													assign node12339 = (inp[6]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node12342 = (inp[11]) ? node12346 : node12343;
													assign node12343 = (inp[3]) ? 15'b000000001111111 : 15'b000000000111111;
													assign node12346 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12349 = (inp[6]) ? node12351 : 15'b000000000111111;
												assign node12351 = (inp[12]) ? node12361 : node12352;
													assign node12352 = (inp[13]) ? node12354 : 15'b000000000111111;
														assign node12354 = (inp[11]) ? node12358 : node12355;
															assign node12355 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
															assign node12358 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node12361 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node12364 = (inp[6]) ? node12376 : node12365;
											assign node12365 = (inp[13]) ? node12373 : node12366;
												assign node12366 = (inp[2]) ? node12368 : 15'b000000011111111;
													assign node12368 = (inp[12]) ? node12370 : 15'b000000000111111;
														assign node12370 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12373 = (inp[3]) ? 15'b000000000011111 : 15'b000000000001111;
											assign node12376 = (inp[12]) ? node12380 : node12377;
												assign node12377 = (inp[13]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node12380 = (inp[3]) ? node12382 : 15'b000000000001111;
													assign node12382 = (inp[13]) ? node12386 : node12383;
														assign node12383 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
														assign node12386 = (inp[11]) ? 15'b000000000000011 : 15'b000000000000111;
								assign node12389 = (inp[13]) ? node12453 : node12390;
									assign node12390 = (inp[11]) ? node12428 : node12391;
										assign node12391 = (inp[12]) ? node12411 : node12392;
											assign node12392 = (inp[14]) ? node12400 : node12393;
												assign node12393 = (inp[2]) ? 15'b000000000111111 : node12394;
													assign node12394 = (inp[3]) ? 15'b000000001111111 : node12395;
														assign node12395 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12400 = (inp[3]) ? node12404 : node12401;
													assign node12401 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12404 = (inp[2]) ? node12408 : node12405;
														assign node12405 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
														assign node12408 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node12411 = (inp[2]) ? node12421 : node12412;
												assign node12412 = (inp[6]) ? node12414 : 15'b000000000111111;
													assign node12414 = (inp[14]) ? node12416 : 15'b000000000111111;
														assign node12416 = (inp[1]) ? 15'b000000000011111 : node12417;
															assign node12417 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12421 = (inp[14]) ? node12425 : node12422;
													assign node12422 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node12425 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node12428 = (inp[1]) ? node12446 : node12429;
											assign node12429 = (inp[12]) ? node12439 : node12430;
												assign node12430 = (inp[14]) ? node12432 : 15'b000000000111111;
													assign node12432 = (inp[6]) ? 15'b000000000011111 : node12433;
														assign node12433 = (inp[3]) ? node12435 : 15'b000000000111111;
															assign node12435 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12439 = (inp[2]) ? node12443 : node12440;
													assign node12440 = (inp[14]) ? 15'b000000000111111 : 15'b000000000011111;
													assign node12443 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node12446 = (inp[3]) ? node12448 : 15'b000000000011111;
												assign node12448 = (inp[14]) ? 15'b000000000000111 : node12449;
													assign node12449 = (inp[12]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node12453 = (inp[12]) ? node12479 : node12454;
										assign node12454 = (inp[11]) ? node12462 : node12455;
											assign node12455 = (inp[3]) ? node12459 : node12456;
												assign node12456 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12459 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node12462 = (inp[1]) ? node12468 : node12463;
												assign node12463 = (inp[14]) ? 15'b000000000011111 : node12464;
													assign node12464 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12468 = (inp[3]) ? node12472 : node12469;
													assign node12469 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node12472 = (inp[2]) ? node12474 : 15'b000000000001111;
														assign node12474 = (inp[14]) ? node12476 : 15'b000000000000111;
															assign node12476 = (inp[6]) ? 15'b000000000000011 : 15'b000000000000111;
										assign node12479 = (inp[6]) ? node12501 : node12480;
											assign node12480 = (inp[3]) ? node12492 : node12481;
												assign node12481 = (inp[14]) ? node12485 : node12482;
													assign node12482 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node12485 = (inp[2]) ? node12487 : 15'b000000000011111;
														assign node12487 = (inp[1]) ? node12489 : 15'b000000000001111;
															assign node12489 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node12492 = (inp[14]) ? 15'b000000000000111 : node12493;
													assign node12493 = (inp[11]) ? node12495 : 15'b000000000011111;
														assign node12495 = (inp[2]) ? node12497 : 15'b000000000001111;
															assign node12497 = (inp[1]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node12501 = (inp[14]) ? node12505 : node12502;
												assign node12502 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node12505 = (inp[1]) ? node12511 : node12506;
													assign node12506 = (inp[2]) ? 15'b000000000000111 : node12507;
														assign node12507 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node12511 = (inp[11]) ? 15'b000000000000011 : node12512;
														assign node12512 = (inp[3]) ? node12514 : 15'b000000000000111;
															assign node12514 = (inp[2]) ? 15'b000000000000011 : 15'b000000000000111;
			assign node12518 = (inp[12]) ? node14602 : node12519;
				assign node12519 = (inp[9]) ? node13539 : node12520;
					assign node12520 = (inp[8]) ? node13024 : node12521;
						assign node12521 = (inp[6]) ? node12775 : node12522;
							assign node12522 = (inp[3]) ? node12654 : node12523;
								assign node12523 = (inp[2]) ? node12581 : node12524;
									assign node12524 = (inp[14]) ? node12556 : node12525;
										assign node12525 = (inp[5]) ? node12549 : node12526;
											assign node12526 = (inp[0]) ? node12538 : node12527;
												assign node12527 = (inp[11]) ? node12535 : node12528;
													assign node12528 = (inp[13]) ? node12532 : node12529;
														assign node12529 = (inp[10]) ? 15'b000111111111111 : 15'b001111111111111;
														assign node12532 = (inp[10]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node12535 = (inp[10]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node12538 = (inp[13]) ? node12546 : node12539;
													assign node12539 = (inp[10]) ? node12541 : 15'b000011111111111;
														assign node12541 = (inp[11]) ? 15'b000001111111111 : node12542;
															assign node12542 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node12546 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node12549 = (inp[10]) ? 15'b000000111111111 : node12550;
												assign node12550 = (inp[11]) ? 15'b000000111111111 : node12551;
													assign node12551 = (inp[1]) ? 15'b000001111111111 : 15'b000011111111111;
										assign node12556 = (inp[5]) ? node12572 : node12557;
											assign node12557 = (inp[13]) ? node12563 : node12558;
												assign node12558 = (inp[10]) ? 15'b000001111111111 : node12559;
													assign node12559 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
												assign node12563 = (inp[11]) ? node12569 : node12564;
													assign node12564 = (inp[10]) ? 15'b000000111111111 : node12565;
														assign node12565 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12569 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node12572 = (inp[1]) ? 15'b000000011111111 : node12573;
												assign node12573 = (inp[10]) ? node12577 : node12574;
													assign node12574 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12577 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
									assign node12581 = (inp[10]) ? node12617 : node12582;
										assign node12582 = (inp[14]) ? node12606 : node12583;
											assign node12583 = (inp[11]) ? node12595 : node12584;
												assign node12584 = (inp[1]) ? node12592 : node12585;
													assign node12585 = (inp[0]) ? 15'b000001111111111 : node12586;
														assign node12586 = (inp[13]) ? 15'b000011111111111 : node12587;
															assign node12587 = (inp[5]) ? 15'b000011111111111 : 15'b000111111111111;
													assign node12592 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node12595 = (inp[5]) ? node12603 : node12596;
													assign node12596 = (inp[13]) ? 15'b000000111111111 : node12597;
														assign node12597 = (inp[0]) ? node12599 : 15'b000001111111111;
															assign node12599 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12603 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node12606 = (inp[13]) ? node12612 : node12607;
												assign node12607 = (inp[5]) ? node12609 : 15'b000001111111111;
													assign node12609 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12612 = (inp[11]) ? node12614 : 15'b000000011111111;
													assign node12614 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node12617 = (inp[5]) ? node12637 : node12618;
											assign node12618 = (inp[13]) ? node12630 : node12619;
												assign node12619 = (inp[1]) ? node12623 : node12620;
													assign node12620 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12623 = (inp[11]) ? node12625 : 15'b000000111111111;
														assign node12625 = (inp[0]) ? 15'b000000011111111 : node12626;
															assign node12626 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12630 = (inp[0]) ? node12634 : node12631;
													assign node12631 = (inp[1]) ? 15'b000000111111111 : 15'b000000011111111;
													assign node12634 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12637 = (inp[0]) ? node12649 : node12638;
												assign node12638 = (inp[1]) ? node12644 : node12639;
													assign node12639 = (inp[14]) ? node12641 : 15'b000000111111111;
														assign node12641 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12644 = (inp[14]) ? node12646 : 15'b000000011111111;
														assign node12646 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12649 = (inp[11]) ? 15'b000000001111111 : node12650;
													assign node12650 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node12654 = (inp[0]) ? node12712 : node12655;
									assign node12655 = (inp[11]) ? node12691 : node12656;
										assign node12656 = (inp[2]) ? node12680 : node12657;
											assign node12657 = (inp[10]) ? node12667 : node12658;
												assign node12658 = (inp[5]) ? node12664 : node12659;
													assign node12659 = (inp[1]) ? node12661 : 15'b000011111111111;
														assign node12661 = (inp[13]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node12664 = (inp[14]) ? 15'b000001111111111 : 15'b000000111111111;
												assign node12667 = (inp[1]) ? node12673 : node12668;
													assign node12668 = (inp[14]) ? node12670 : 15'b000001111111111;
														assign node12670 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12673 = (inp[5]) ? 15'b000000011111111 : node12674;
														assign node12674 = (inp[14]) ? 15'b000000111111111 : node12675;
															assign node12675 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node12680 = (inp[13]) ? node12682 : 15'b000000111111111;
												assign node12682 = (inp[5]) ? node12688 : node12683;
													assign node12683 = (inp[10]) ? node12685 : 15'b000000111111111;
														assign node12685 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12688 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node12691 = (inp[10]) ? node12701 : node12692;
											assign node12692 = (inp[2]) ? node12696 : node12693;
												assign node12693 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node12696 = (inp[1]) ? 15'b000000001111111 : node12697;
													assign node12697 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node12701 = (inp[2]) ? node12707 : node12702;
												assign node12702 = (inp[5]) ? node12704 : 15'b000000011111111;
													assign node12704 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12707 = (inp[1]) ? 15'b000000001111111 : node12708;
													assign node12708 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node12712 = (inp[5]) ? node12750 : node12713;
										assign node12713 = (inp[2]) ? node12733 : node12714;
											assign node12714 = (inp[1]) ? node12728 : node12715;
												assign node12715 = (inp[13]) ? node12723 : node12716;
													assign node12716 = (inp[14]) ? 15'b000000111111111 : node12717;
														assign node12717 = (inp[10]) ? node12719 : 15'b000001111111111;
															assign node12719 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12723 = (inp[11]) ? node12725 : 15'b000000111111111;
														assign node12725 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12728 = (inp[10]) ? 15'b000000001111111 : node12729;
													assign node12729 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node12733 = (inp[14]) ? node12741 : node12734;
												assign node12734 = (inp[13]) ? 15'b000000011111111 : node12735;
													assign node12735 = (inp[10]) ? node12737 : 15'b000000011111111;
														assign node12737 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12741 = (inp[10]) ? 15'b000000000111111 : node12742;
													assign node12742 = (inp[13]) ? 15'b000000001111111 : node12743;
														assign node12743 = (inp[1]) ? node12745 : 15'b000000011111111;
															assign node12745 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node12750 = (inp[13]) ? node12762 : node12751;
											assign node12751 = (inp[2]) ? node12755 : node12752;
												assign node12752 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12755 = (inp[11]) ? 15'b000000001111111 : node12756;
													assign node12756 = (inp[14]) ? 15'b000000001111111 : node12757;
														assign node12757 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12762 = (inp[10]) ? node12766 : node12763;
												assign node12763 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12766 = (inp[14]) ? 15'b000000000111111 : node12767;
													assign node12767 = (inp[2]) ? 15'b000000000111111 : node12768;
														assign node12768 = (inp[11]) ? node12770 : 15'b000000001111111;
															assign node12770 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
							assign node12775 = (inp[1]) ? node12881 : node12776;
								assign node12776 = (inp[10]) ? node12834 : node12777;
									assign node12777 = (inp[13]) ? node12797 : node12778;
										assign node12778 = (inp[3]) ? node12788 : node12779;
											assign node12779 = (inp[5]) ? 15'b000001111111111 : node12780;
												assign node12780 = (inp[0]) ? node12782 : 15'b000011111111111;
													assign node12782 = (inp[11]) ? 15'b000001111111111 : node12783;
														assign node12783 = (inp[14]) ? 15'b000001111111111 : 15'b000011111111111;
											assign node12788 = (inp[14]) ? node12792 : node12789;
												assign node12789 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12792 = (inp[11]) ? 15'b000000011111111 : node12793;
													assign node12793 = (inp[5]) ? 15'b000000111111111 : 15'b000000011111111;
										assign node12797 = (inp[14]) ? node12821 : node12798;
											assign node12798 = (inp[2]) ? node12810 : node12799;
												assign node12799 = (inp[3]) ? node12807 : node12800;
													assign node12800 = (inp[11]) ? 15'b000000111111111 : node12801;
														assign node12801 = (inp[0]) ? node12803 : 15'b000001111111111;
															assign node12803 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node12807 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node12810 = (inp[0]) ? 15'b000000011111111 : node12811;
													assign node12811 = (inp[3]) ? node12813 : 15'b000000111111111;
														assign node12813 = (inp[5]) ? node12817 : node12814;
															assign node12814 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
															assign node12817 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12821 = (inp[5]) ? node12825 : node12822;
												assign node12822 = (inp[2]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node12825 = (inp[11]) ? 15'b000000001111111 : node12826;
													assign node12826 = (inp[2]) ? 15'b000000001111111 : node12827;
														assign node12827 = (inp[0]) ? node12829 : 15'b000000011111111;
															assign node12829 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node12834 = (inp[5]) ? node12856 : node12835;
										assign node12835 = (inp[3]) ? node12849 : node12836;
											assign node12836 = (inp[2]) ? node12842 : node12837;
												assign node12837 = (inp[11]) ? 15'b000000111111111 : node12838;
													assign node12838 = (inp[0]) ? 15'b000000111111111 : 15'b000011111111111;
												assign node12842 = (inp[14]) ? node12846 : node12843;
													assign node12843 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12846 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12849 = (inp[0]) ? 15'b000000001111111 : node12850;
												assign node12850 = (inp[2]) ? 15'b000000000111111 : node12851;
													assign node12851 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node12856 = (inp[13]) ? node12872 : node12857;
											assign node12857 = (inp[2]) ? node12865 : node12858;
												assign node12858 = (inp[14]) ? 15'b000000011111111 : node12859;
													assign node12859 = (inp[3]) ? node12861 : 15'b000000011111111;
														assign node12861 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12865 = (inp[0]) ? 15'b000000000111111 : node12866;
													assign node12866 = (inp[11]) ? node12868 : 15'b000000011111111;
														assign node12868 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12872 = (inp[14]) ? node12876 : node12873;
												assign node12873 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12876 = (inp[0]) ? 15'b000000000011111 : node12877;
													assign node12877 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
								assign node12881 = (inp[11]) ? node12951 : node12882;
									assign node12882 = (inp[14]) ? node12914 : node12883;
										assign node12883 = (inp[0]) ? node12901 : node12884;
											assign node12884 = (inp[5]) ? node12886 : 15'b000001111111111;
												assign node12886 = (inp[10]) ? node12896 : node12887;
													assign node12887 = (inp[3]) ? node12893 : node12888;
														assign node12888 = (inp[2]) ? 15'b000000111111111 : node12889;
															assign node12889 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node12893 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12896 = (inp[2]) ? 15'b000000011111111 : node12897;
														assign node12897 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node12901 = (inp[10]) ? node12907 : node12902;
												assign node12902 = (inp[13]) ? node12904 : 15'b000000011111111;
													assign node12904 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12907 = (inp[2]) ? 15'b000000001111111 : node12908;
													assign node12908 = (inp[5]) ? node12910 : 15'b000000011111111;
														assign node12910 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node12914 = (inp[5]) ? node12932 : node12915;
											assign node12915 = (inp[13]) ? 15'b000000001111111 : node12916;
												assign node12916 = (inp[10]) ? node12924 : node12917;
													assign node12917 = (inp[3]) ? node12919 : 15'b000000111111111;
														assign node12919 = (inp[2]) ? node12921 : 15'b000000011111111;
															assign node12921 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12924 = (inp[3]) ? 15'b000000001111111 : node12925;
														assign node12925 = (inp[0]) ? node12927 : 15'b000000011111111;
															assign node12927 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node12932 = (inp[10]) ? node12944 : node12933;
												assign node12933 = (inp[13]) ? node12939 : node12934;
													assign node12934 = (inp[3]) ? 15'b000000001111111 : node12935;
														assign node12935 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12939 = (inp[2]) ? node12941 : 15'b000000001111111;
														assign node12941 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node12944 = (inp[0]) ? node12948 : node12945;
													assign node12945 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node12948 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node12951 = (inp[14]) ? node12985 : node12952;
										assign node12952 = (inp[10]) ? node12972 : node12953;
											assign node12953 = (inp[5]) ? node12963 : node12954;
												assign node12954 = (inp[3]) ? node12960 : node12955;
													assign node12955 = (inp[0]) ? 15'b000000011111111 : node12956;
														assign node12956 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node12960 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12963 = (inp[2]) ? node12969 : node12964;
													assign node12964 = (inp[0]) ? node12966 : 15'b000000011111111;
														assign node12966 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12969 = (inp[0]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node12972 = (inp[13]) ? node12982 : node12973;
												assign node12973 = (inp[5]) ? 15'b000000000111111 : node12974;
													assign node12974 = (inp[0]) ? node12976 : 15'b000000011111111;
														assign node12976 = (inp[2]) ? 15'b000000001111111 : node12977;
															assign node12977 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node12982 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node12985 = (inp[13]) ? node13003 : node12986;
											assign node12986 = (inp[3]) ? node12998 : node12987;
												assign node12987 = (inp[10]) ? node12993 : node12988;
													assign node12988 = (inp[0]) ? node12990 : 15'b000000011111111;
														assign node12990 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node12993 = (inp[5]) ? node12995 : 15'b000000001111111;
														assign node12995 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node12998 = (inp[2]) ? node13000 : 15'b000000000111111;
													assign node13000 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13003 = (inp[2]) ? node13013 : node13004;
												assign node13004 = (inp[0]) ? node13010 : node13005;
													assign node13005 = (inp[10]) ? 15'b000000000111111 : node13006;
														assign node13006 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13010 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13013 = (inp[5]) ? node13019 : node13014;
													assign node13014 = (inp[3]) ? 15'b000000000011111 : node13015;
														assign node13015 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13019 = (inp[10]) ? node13021 : 15'b000000000011111;
														assign node13021 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
						assign node13024 = (inp[10]) ? node13272 : node13025;
							assign node13025 = (inp[0]) ? node13151 : node13026;
								assign node13026 = (inp[6]) ? node13094 : node13027;
									assign node13027 = (inp[3]) ? node13055 : node13028;
										assign node13028 = (inp[2]) ? node13038 : node13029;
											assign node13029 = (inp[1]) ? node13035 : node13030;
												assign node13030 = (inp[5]) ? 15'b000001111111111 : node13031;
													assign node13031 = (inp[11]) ? 15'b000011111111111 : 15'b000111111111111;
												assign node13035 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node13038 = (inp[13]) ? node13050 : node13039;
												assign node13039 = (inp[1]) ? node13047 : node13040;
													assign node13040 = (inp[14]) ? 15'b000000111111111 : node13041;
														assign node13041 = (inp[5]) ? node13043 : 15'b000001111111111;
															assign node13043 = (inp[11]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13047 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13050 = (inp[11]) ? 15'b000000011111111 : node13051;
													assign node13051 = (inp[5]) ? 15'b000000011111111 : 15'b000001111111111;
										assign node13055 = (inp[11]) ? node13079 : node13056;
											assign node13056 = (inp[13]) ? node13070 : node13057;
												assign node13057 = (inp[5]) ? node13065 : node13058;
													assign node13058 = (inp[1]) ? node13060 : 15'b000001111111111;
														assign node13060 = (inp[14]) ? 15'b000000111111111 : node13061;
															assign node13061 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13065 = (inp[14]) ? node13067 : 15'b000000111111111;
														assign node13067 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13070 = (inp[2]) ? node13076 : node13071;
													assign node13071 = (inp[14]) ? node13073 : 15'b000000111111111;
														assign node13073 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13076 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13079 = (inp[13]) ? node13089 : node13080;
												assign node13080 = (inp[1]) ? node13086 : node13081;
													assign node13081 = (inp[14]) ? 15'b000000011111111 : node13082;
														assign node13082 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13086 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13089 = (inp[5]) ? 15'b000000001111111 : node13090;
													assign node13090 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
									assign node13094 = (inp[1]) ? node13118 : node13095;
										assign node13095 = (inp[11]) ? node13107 : node13096;
											assign node13096 = (inp[2]) ? node13100 : node13097;
												assign node13097 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node13100 = (inp[3]) ? node13102 : 15'b000000111111111;
													assign node13102 = (inp[5]) ? 15'b000000001111111 : node13103;
														assign node13103 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node13107 = (inp[2]) ? node13113 : node13108;
												assign node13108 = (inp[5]) ? 15'b000000011111111 : node13109;
													assign node13109 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13113 = (inp[14]) ? node13115 : 15'b000000001111111;
													assign node13115 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node13118 = (inp[2]) ? node13134 : node13119;
											assign node13119 = (inp[13]) ? node13125 : node13120;
												assign node13120 = (inp[14]) ? node13122 : 15'b000000011111111;
													assign node13122 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13125 = (inp[11]) ? node13129 : node13126;
													assign node13126 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13129 = (inp[3]) ? 15'b000000000111111 : node13130;
														assign node13130 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13134 = (inp[11]) ? node13140 : node13135;
												assign node13135 = (inp[13]) ? node13137 : 15'b000000111111111;
													assign node13137 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13140 = (inp[13]) ? node13146 : node13141;
													assign node13141 = (inp[3]) ? 15'b000000000111111 : node13142;
														assign node13142 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13146 = (inp[14]) ? node13148 : 15'b000000000011111;
														assign node13148 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node13151 = (inp[3]) ? node13207 : node13152;
									assign node13152 = (inp[2]) ? node13182 : node13153;
										assign node13153 = (inp[5]) ? node13173 : node13154;
											assign node13154 = (inp[13]) ? node13166 : node13155;
												assign node13155 = (inp[11]) ? node13163 : node13156;
													assign node13156 = (inp[14]) ? 15'b000000111111111 : node13157;
														assign node13157 = (inp[6]) ? node13159 : 15'b000001111111111;
															assign node13159 = (inp[1]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13163 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13166 = (inp[1]) ? node13170 : node13167;
													assign node13167 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13170 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13173 = (inp[6]) ? node13175 : 15'b000000011111111;
												assign node13175 = (inp[13]) ? node13179 : node13176;
													assign node13176 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13179 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node13182 = (inp[11]) ? node13202 : node13183;
											assign node13183 = (inp[13]) ? node13193 : node13184;
												assign node13184 = (inp[5]) ? node13186 : 15'b000000011111111;
													assign node13186 = (inp[14]) ? node13188 : 15'b000000011111111;
														assign node13188 = (inp[1]) ? 15'b000000001111111 : node13189;
															assign node13189 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13193 = (inp[6]) ? node13199 : node13194;
													assign node13194 = (inp[5]) ? 15'b000000001111111 : node13195;
														assign node13195 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13199 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13202 = (inp[5]) ? node13204 : 15'b000000001111111;
												assign node13204 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node13207 = (inp[2]) ? node13239 : node13208;
										assign node13208 = (inp[1]) ? node13222 : node13209;
											assign node13209 = (inp[11]) ? node13215 : node13210;
												assign node13210 = (inp[13]) ? 15'b000000011111111 : node13211;
													assign node13211 = (inp[14]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node13215 = (inp[14]) ? 15'b000000000111111 : node13216;
													assign node13216 = (inp[5]) ? node13218 : 15'b000000011111111;
														assign node13218 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13222 = (inp[6]) ? node13232 : node13223;
												assign node13223 = (inp[5]) ? node13227 : node13224;
													assign node13224 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13227 = (inp[14]) ? node13229 : 15'b000000001111111;
														assign node13229 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13232 = (inp[5]) ? node13236 : node13233;
													assign node13233 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13236 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node13239 = (inp[11]) ? node13259 : node13240;
											assign node13240 = (inp[14]) ? node13252 : node13241;
												assign node13241 = (inp[5]) ? node13245 : node13242;
													assign node13242 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13245 = (inp[1]) ? node13247 : 15'b000000001111111;
														assign node13247 = (inp[13]) ? 15'b000000000111111 : node13248;
															assign node13248 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13252 = (inp[1]) ? node13256 : node13253;
													assign node13253 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13256 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node13259 = (inp[13]) ? node13267 : node13260;
												assign node13260 = (inp[1]) ? node13262 : 15'b000000000111111;
													assign node13262 = (inp[6]) ? node13264 : 15'b000000000111111;
														assign node13264 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node13267 = (inp[6]) ? node13269 : 15'b000000000011111;
													assign node13269 = (inp[1]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node13272 = (inp[14]) ? node13400 : node13273;
								assign node13273 = (inp[2]) ? node13341 : node13274;
									assign node13274 = (inp[11]) ? node13316 : node13275;
										assign node13275 = (inp[3]) ? node13301 : node13276;
											assign node13276 = (inp[6]) ? node13286 : node13277;
												assign node13277 = (inp[1]) ? node13283 : node13278;
													assign node13278 = (inp[0]) ? node13280 : 15'b000001111111111;
														assign node13280 = (inp[5]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13283 = (inp[13]) ? 15'b000000111111111 : 15'b000000011111111;
												assign node13286 = (inp[5]) ? node13294 : node13287;
													assign node13287 = (inp[0]) ? 15'b000000011111111 : node13288;
														assign node13288 = (inp[13]) ? node13290 : 15'b000000111111111;
															assign node13290 = (inp[1]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13294 = (inp[13]) ? node13296 : 15'b000000011111111;
														assign node13296 = (inp[0]) ? 15'b000000001111111 : node13297;
															assign node13297 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13301 = (inp[1]) ? node13313 : node13302;
												assign node13302 = (inp[13]) ? node13310 : node13303;
													assign node13303 = (inp[5]) ? 15'b000000011111111 : node13304;
														assign node13304 = (inp[6]) ? node13306 : 15'b000000111111111;
															assign node13306 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13310 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13313 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node13316 = (inp[0]) ? node13332 : node13317;
											assign node13317 = (inp[1]) ? 15'b000000001111111 : node13318;
												assign node13318 = (inp[6]) ? node13322 : node13319;
													assign node13319 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13322 = (inp[5]) ? node13328 : node13323;
														assign node13323 = (inp[3]) ? node13325 : 15'b000000011111111;
															assign node13325 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node13328 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13332 = (inp[3]) ? node13338 : node13333;
												assign node13333 = (inp[6]) ? node13335 : 15'b000000001111111;
													assign node13335 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13338 = (inp[5]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node13341 = (inp[0]) ? node13363 : node13342;
										assign node13342 = (inp[3]) ? node13354 : node13343;
											assign node13343 = (inp[6]) ? node13349 : node13344;
												assign node13344 = (inp[11]) ? 15'b000000011111111 : node13345;
													assign node13345 = (inp[5]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node13349 = (inp[5]) ? 15'b000000000111111 : node13350;
													assign node13350 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13354 = (inp[5]) ? node13356 : 15'b000000001111111;
												assign node13356 = (inp[6]) ? node13360 : node13357;
													assign node13357 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13360 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node13363 = (inp[1]) ? node13385 : node13364;
											assign node13364 = (inp[13]) ? node13376 : node13365;
												assign node13365 = (inp[5]) ? node13369 : node13366;
													assign node13366 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node13369 = (inp[11]) ? 15'b000000000111111 : node13370;
														assign node13370 = (inp[6]) ? node13372 : 15'b000000001111111;
															assign node13372 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13376 = (inp[11]) ? node13380 : node13377;
													assign node13377 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13380 = (inp[6]) ? node13382 : 15'b000000000111111;
														assign node13382 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13385 = (inp[3]) ? node13393 : node13386;
												assign node13386 = (inp[11]) ? node13390 : node13387;
													assign node13387 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13390 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13393 = (inp[6]) ? node13397 : node13394;
													assign node13394 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node13397 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node13400 = (inp[1]) ? node13466 : node13401;
									assign node13401 = (inp[6]) ? node13425 : node13402;
										assign node13402 = (inp[2]) ? node13418 : node13403;
											assign node13403 = (inp[13]) ? node13409 : node13404;
												assign node13404 = (inp[5]) ? 15'b000000011111111 : node13405;
													assign node13405 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13409 = (inp[11]) ? node13413 : node13410;
													assign node13410 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13413 = (inp[5]) ? node13415 : 15'b000000000111111;
														assign node13415 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13418 = (inp[11]) ? 15'b000000000111111 : node13419;
												assign node13419 = (inp[0]) ? node13421 : 15'b000000001111111;
													assign node13421 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node13425 = (inp[3]) ? node13443 : node13426;
											assign node13426 = (inp[0]) ? node13438 : node13427;
												assign node13427 = (inp[11]) ? node13431 : node13428;
													assign node13428 = (inp[5]) ? 15'b000000011111111 : 15'b000000001111111;
													assign node13431 = (inp[13]) ? 15'b000000000111111 : node13432;
														assign node13432 = (inp[5]) ? node13434 : 15'b000000001111111;
															assign node13434 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13438 = (inp[11]) ? node13440 : 15'b000000000111111;
													assign node13440 = (inp[2]) ? 15'b000000000001111 : 15'b000000001111111;
											assign node13443 = (inp[13]) ? node13459 : node13444;
												assign node13444 = (inp[0]) ? node13452 : node13445;
													assign node13445 = (inp[5]) ? 15'b000000000111111 : node13446;
														assign node13446 = (inp[2]) ? node13448 : 15'b000000001111111;
															assign node13448 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13452 = (inp[11]) ? node13454 : 15'b000000000111111;
														assign node13454 = (inp[5]) ? node13456 : 15'b000000000011111;
															assign node13456 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node13459 = (inp[11]) ? node13463 : node13460;
													assign node13460 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13463 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node13466 = (inp[3]) ? node13506 : node13467;
										assign node13467 = (inp[5]) ? node13495 : node13468;
											assign node13468 = (inp[0]) ? node13476 : node13469;
												assign node13469 = (inp[11]) ? node13473 : node13470;
													assign node13470 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13473 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13476 = (inp[6]) ? node13488 : node13477;
													assign node13477 = (inp[13]) ? node13483 : node13478;
														assign node13478 = (inp[11]) ? node13480 : 15'b000000001111111;
															assign node13480 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
														assign node13483 = (inp[2]) ? node13485 : 15'b000000000111111;
															assign node13485 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13488 = (inp[2]) ? node13490 : 15'b000000000111111;
														assign node13490 = (inp[13]) ? 15'b000000000011111 : node13491;
															assign node13491 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13495 = (inp[6]) ? 15'b000000000011111 : node13496;
												assign node13496 = (inp[11]) ? 15'b000000000011111 : node13497;
													assign node13497 = (inp[2]) ? node13499 : 15'b000000000111111;
														assign node13499 = (inp[0]) ? node13501 : 15'b000000000111111;
															assign node13501 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node13506 = (inp[11]) ? node13516 : node13507;
											assign node13507 = (inp[2]) ? node13509 : 15'b000000000111111;
												assign node13509 = (inp[6]) ? 15'b000000000011111 : node13510;
													assign node13510 = (inp[0]) ? 15'b000000000011111 : node13511;
														assign node13511 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13516 = (inp[6]) ? node13526 : node13517;
												assign node13517 = (inp[5]) ? node13523 : node13518;
													assign node13518 = (inp[2]) ? 15'b000000000011111 : node13519;
														assign node13519 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13523 = (inp[13]) ? 15'b000000000000111 : 15'b000000000011111;
												assign node13526 = (inp[5]) ? node13528 : 15'b000000000001111;
													assign node13528 = (inp[2]) ? node13534 : node13529;
														assign node13529 = (inp[0]) ? node13531 : 15'b000000000001111;
															assign node13531 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
														assign node13534 = (inp[0]) ? node13536 : 15'b000000000000111;
															assign node13536 = (inp[13]) ? 15'b000000000000011 : 15'b000000000000111;
					assign node13539 = (inp[11]) ? node14067 : node13540;
						assign node13540 = (inp[3]) ? node13812 : node13541;
							assign node13541 = (inp[1]) ? node13677 : node13542;
								assign node13542 = (inp[0]) ? node13618 : node13543;
									assign node13543 = (inp[13]) ? node13581 : node13544;
										assign node13544 = (inp[2]) ? node13562 : node13545;
											assign node13545 = (inp[6]) ? node13555 : node13546;
												assign node13546 = (inp[10]) ? node13552 : node13547;
													assign node13547 = (inp[5]) ? 15'b000001111111111 : node13548;
														assign node13548 = (inp[8]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node13552 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node13555 = (inp[14]) ? 15'b000000111111111 : node13556;
													assign node13556 = (inp[10]) ? node13558 : 15'b000001111111111;
														assign node13558 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
											assign node13562 = (inp[8]) ? node13570 : node13563;
												assign node13563 = (inp[10]) ? node13567 : node13564;
													assign node13564 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13567 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13570 = (inp[6]) ? node13578 : node13571;
													assign node13571 = (inp[14]) ? node13573 : 15'b000000111111111;
														assign node13573 = (inp[5]) ? 15'b000000011111111 : node13574;
															assign node13574 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13578 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node13581 = (inp[14]) ? node13599 : node13582;
											assign node13582 = (inp[10]) ? node13594 : node13583;
												assign node13583 = (inp[8]) ? node13585 : 15'b000001111111111;
													assign node13585 = (inp[2]) ? node13589 : node13586;
														assign node13586 = (inp[6]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node13589 = (inp[5]) ? 15'b000000011111111 : node13590;
															assign node13590 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13594 = (inp[2]) ? node13596 : 15'b000000011111111;
													assign node13596 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13599 = (inp[8]) ? node13609 : node13600;
												assign node13600 = (inp[5]) ? node13606 : node13601;
													assign node13601 = (inp[2]) ? 15'b000000011111111 : node13602;
														assign node13602 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13606 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13609 = (inp[2]) ? node13611 : 15'b000000011111111;
													assign node13611 = (inp[10]) ? 15'b000000000111111 : node13612;
														assign node13612 = (inp[5]) ? node13614 : 15'b000000001111111;
															assign node13614 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node13618 = (inp[2]) ? node13646 : node13619;
										assign node13619 = (inp[13]) ? node13635 : node13620;
											assign node13620 = (inp[5]) ? node13628 : node13621;
												assign node13621 = (inp[6]) ? 15'b000000111111111 : node13622;
													assign node13622 = (inp[8]) ? node13624 : 15'b000001111111111;
														assign node13624 = (inp[10]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node13628 = (inp[10]) ? 15'b000000001111111 : node13629;
													assign node13629 = (inp[14]) ? 15'b000000011111111 : node13630;
														assign node13630 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node13635 = (inp[5]) ? node13643 : node13636;
												assign node13636 = (inp[14]) ? node13638 : 15'b000000011111111;
													assign node13638 = (inp[8]) ? 15'b000000001111111 : node13639;
														assign node13639 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13643 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node13646 = (inp[10]) ? node13666 : node13647;
											assign node13647 = (inp[14]) ? node13651 : node13648;
												assign node13648 = (inp[5]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13651 = (inp[8]) ? node13657 : node13652;
													assign node13652 = (inp[13]) ? node13654 : 15'b000000011111111;
														assign node13654 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13657 = (inp[5]) ? node13663 : node13658;
														assign node13658 = (inp[6]) ? 15'b000000001111111 : node13659;
															assign node13659 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node13663 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13666 = (inp[8]) ? node13670 : node13667;
												assign node13667 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13670 = (inp[5]) ? 15'b000000000011111 : node13671;
													assign node13671 = (inp[13]) ? node13673 : 15'b000000000111111;
														assign node13673 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node13677 = (inp[10]) ? node13745 : node13678;
									assign node13678 = (inp[2]) ? node13714 : node13679;
										assign node13679 = (inp[0]) ? node13695 : node13680;
											assign node13680 = (inp[5]) ? node13688 : node13681;
												assign node13681 = (inp[13]) ? node13685 : node13682;
													assign node13682 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13685 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13688 = (inp[8]) ? 15'b000000011111111 : node13689;
													assign node13689 = (inp[6]) ? node13691 : 15'b000000111111111;
														assign node13691 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node13695 = (inp[8]) ? node13705 : node13696;
												assign node13696 = (inp[6]) ? node13702 : node13697;
													assign node13697 = (inp[14]) ? 15'b000000011111111 : node13698;
														assign node13698 = (inp[13]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13702 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13705 = (inp[5]) ? node13711 : node13706;
													assign node13706 = (inp[6]) ? node13708 : 15'b000000001111111;
														assign node13708 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13711 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node13714 = (inp[6]) ? node13736 : node13715;
											assign node13715 = (inp[13]) ? node13727 : node13716;
												assign node13716 = (inp[5]) ? node13724 : node13717;
													assign node13717 = (inp[14]) ? 15'b000000011111111 : node13718;
														assign node13718 = (inp[8]) ? 15'b000000111111111 : node13719;
															assign node13719 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node13724 = (inp[8]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node13727 = (inp[14]) ? 15'b000000000111111 : node13728;
													assign node13728 = (inp[8]) ? node13730 : 15'b000000001111111;
														assign node13730 = (inp[5]) ? node13732 : 15'b000000001111111;
															assign node13732 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13736 = (inp[14]) ? node13742 : node13737;
												assign node13737 = (inp[8]) ? 15'b000000000011111 : node13738;
													assign node13738 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13742 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node13745 = (inp[0]) ? node13783 : node13746;
										assign node13746 = (inp[6]) ? node13764 : node13747;
											assign node13747 = (inp[13]) ? node13755 : node13748;
												assign node13748 = (inp[5]) ? 15'b000000011111111 : node13749;
													assign node13749 = (inp[14]) ? node13751 : 15'b000000011111111;
														assign node13751 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13755 = (inp[5]) ? node13761 : node13756;
													assign node13756 = (inp[8]) ? 15'b000000001111111 : node13757;
														assign node13757 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13761 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13764 = (inp[8]) ? node13772 : node13765;
												assign node13765 = (inp[5]) ? 15'b000000000111111 : node13766;
													assign node13766 = (inp[14]) ? 15'b000000001111111 : node13767;
														assign node13767 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13772 = (inp[2]) ? node13776 : node13773;
													assign node13773 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13776 = (inp[13]) ? node13778 : 15'b000000000111111;
														assign node13778 = (inp[5]) ? node13780 : 15'b000000000011111;
															assign node13780 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node13783 = (inp[8]) ? node13797 : node13784;
											assign node13784 = (inp[2]) ? node13790 : node13785;
												assign node13785 = (inp[6]) ? node13787 : 15'b000000011111111;
													assign node13787 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13790 = (inp[14]) ? node13794 : node13791;
													assign node13791 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13794 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13797 = (inp[5]) ? node13807 : node13798;
												assign node13798 = (inp[13]) ? node13800 : 15'b000000000111111;
													assign node13800 = (inp[2]) ? 15'b000000000011111 : node13801;
														assign node13801 = (inp[6]) ? node13803 : 15'b000000000111111;
															assign node13803 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node13807 = (inp[6]) ? 15'b000000000011111 : node13808;
													assign node13808 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node13812 = (inp[14]) ? node13944 : node13813;
								assign node13813 = (inp[2]) ? node13871 : node13814;
									assign node13814 = (inp[8]) ? node13844 : node13815;
										assign node13815 = (inp[5]) ? node13833 : node13816;
											assign node13816 = (inp[1]) ? node13822 : node13817;
												assign node13817 = (inp[6]) ? node13819 : 15'b000000111111111;
													assign node13819 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13822 = (inp[13]) ? node13830 : node13823;
													assign node13823 = (inp[0]) ? 15'b000000011111111 : node13824;
														assign node13824 = (inp[6]) ? node13826 : 15'b000000111111111;
															assign node13826 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13830 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13833 = (inp[6]) ? node13835 : 15'b000000011111111;
												assign node13835 = (inp[13]) ? 15'b000000001111111 : node13836;
													assign node13836 = (inp[0]) ? 15'b000000001111111 : node13837;
														assign node13837 = (inp[1]) ? 15'b000000011111111 : node13838;
															assign node13838 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
										assign node13844 = (inp[13]) ? node13860 : node13845;
											assign node13845 = (inp[5]) ? node13855 : node13846;
												assign node13846 = (inp[0]) ? node13850 : node13847;
													assign node13847 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13850 = (inp[10]) ? node13852 : 15'b000000011111111;
														assign node13852 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13855 = (inp[1]) ? 15'b000000000111111 : node13856;
													assign node13856 = (inp[10]) ? 15'b000000001111111 : 15'b000000111111111;
											assign node13860 = (inp[5]) ? node13866 : node13861;
												assign node13861 = (inp[6]) ? 15'b000000000111111 : node13862;
													assign node13862 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13866 = (inp[10]) ? node13868 : 15'b000000000111111;
													assign node13868 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node13871 = (inp[10]) ? node13911 : node13872;
										assign node13872 = (inp[5]) ? node13888 : node13873;
											assign node13873 = (inp[0]) ? node13883 : node13874;
												assign node13874 = (inp[1]) ? node13880 : node13875;
													assign node13875 = (inp[8]) ? 15'b000000011111111 : node13876;
														assign node13876 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13880 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13883 = (inp[6]) ? 15'b000000001111111 : node13884;
													assign node13884 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node13888 = (inp[13]) ? node13898 : node13889;
												assign node13889 = (inp[0]) ? node13895 : node13890;
													assign node13890 = (inp[1]) ? 15'b000000001111111 : node13891;
														assign node13891 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13895 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13898 = (inp[8]) ? node13906 : node13899;
													assign node13899 = (inp[0]) ? 15'b000000000111111 : node13900;
														assign node13900 = (inp[6]) ? node13902 : 15'b000000001111111;
															assign node13902 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13906 = (inp[6]) ? node13908 : 15'b000000000111111;
														assign node13908 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node13911 = (inp[5]) ? node13929 : node13912;
											assign node13912 = (inp[13]) ? node13922 : node13913;
												assign node13913 = (inp[0]) ? node13919 : node13914;
													assign node13914 = (inp[8]) ? 15'b000000001111111 : node13915;
														assign node13915 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13919 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13922 = (inp[1]) ? node13926 : node13923;
													assign node13923 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node13926 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node13929 = (inp[6]) ? node13935 : node13930;
												assign node13930 = (inp[8]) ? 15'b000000000111111 : node13931;
													assign node13931 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13935 = (inp[0]) ? 15'b000000000001111 : node13936;
													assign node13936 = (inp[8]) ? 15'b000000000011111 : node13937;
														assign node13937 = (inp[1]) ? node13939 : 15'b000000000111111;
															assign node13939 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
								assign node13944 = (inp[6]) ? node14018 : node13945;
									assign node13945 = (inp[0]) ? node13981 : node13946;
										assign node13946 = (inp[8]) ? node13964 : node13947;
											assign node13947 = (inp[1]) ? node13955 : node13948;
												assign node13948 = (inp[2]) ? node13952 : node13949;
													assign node13949 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node13952 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node13955 = (inp[10]) ? node13961 : node13956;
													assign node13956 = (inp[2]) ? node13958 : 15'b000000011111111;
														assign node13958 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13961 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13964 = (inp[5]) ? node13974 : node13965;
												assign node13965 = (inp[10]) ? node13971 : node13966;
													assign node13966 = (inp[13]) ? 15'b000000001111111 : node13967;
														assign node13967 = (inp[1]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13971 = (inp[1]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node13974 = (inp[2]) ? node13978 : node13975;
													assign node13975 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node13978 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node13981 = (inp[13]) ? node13997 : node13982;
											assign node13982 = (inp[5]) ? node13988 : node13983;
												assign node13983 = (inp[10]) ? 15'b000000001111111 : node13984;
													assign node13984 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node13988 = (inp[10]) ? node13992 : node13989;
													assign node13989 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node13992 = (inp[1]) ? 15'b000000000111111 : node13993;
														assign node13993 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node13997 = (inp[10]) ? node14007 : node13998;
												assign node13998 = (inp[1]) ? 15'b000000000011111 : node13999;
													assign node13999 = (inp[5]) ? node14001 : 15'b000000001111111;
														assign node14001 = (inp[8]) ? node14003 : 15'b000000000111111;
															assign node14003 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14007 = (inp[5]) ? node14011 : node14008;
													assign node14008 = (inp[1]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14011 = (inp[1]) ? 15'b000000000001111 : node14012;
														assign node14012 = (inp[2]) ? node14014 : 15'b000000000011111;
															assign node14014 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node14018 = (inp[1]) ? node14036 : node14019;
										assign node14019 = (inp[5]) ? node14023 : node14020;
											assign node14020 = (inp[10]) ? 15'b000000000111111 : 15'b000000011111111;
											assign node14023 = (inp[13]) ? node14029 : node14024;
												assign node14024 = (inp[2]) ? node14026 : 15'b000000000111111;
													assign node14026 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14029 = (inp[10]) ? 15'b000000000001111 : node14030;
													assign node14030 = (inp[2]) ? 15'b000000000011111 : node14031;
														assign node14031 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node14036 = (inp[8]) ? node14050 : node14037;
											assign node14037 = (inp[2]) ? node14043 : node14038;
												assign node14038 = (inp[10]) ? node14040 : 15'b000000000111111;
													assign node14040 = (inp[13]) ? 15'b000000000001111 : 15'b000000000111111;
												assign node14043 = (inp[5]) ? node14047 : node14044;
													assign node14044 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14047 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node14050 = (inp[2]) ? node14060 : node14051;
												assign node14051 = (inp[13]) ? node14055 : node14052;
													assign node14052 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14055 = (inp[0]) ? node14057 : 15'b000000000011111;
														assign node14057 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node14060 = (inp[13]) ? node14064 : node14061;
													assign node14061 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node14064 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node14067 = (inp[1]) ? node14337 : node14068;
							assign node14068 = (inp[8]) ? node14200 : node14069;
								assign node14069 = (inp[6]) ? node14117 : node14070;
									assign node14070 = (inp[13]) ? node14092 : node14071;
										assign node14071 = (inp[2]) ? node14081 : node14072;
											assign node14072 = (inp[14]) ? node14076 : node14073;
												assign node14073 = (inp[5]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node14076 = (inp[0]) ? node14078 : 15'b000000111111111;
													assign node14078 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node14081 = (inp[14]) ? 15'b000000001111111 : node14082;
												assign node14082 = (inp[5]) ? node14086 : node14083;
													assign node14083 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14086 = (inp[0]) ? 15'b000000001111111 : node14087;
														assign node14087 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node14092 = (inp[3]) ? node14106 : node14093;
											assign node14093 = (inp[14]) ? node14099 : node14094;
												assign node14094 = (inp[10]) ? node14096 : 15'b000000011111111;
													assign node14096 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14099 = (inp[0]) ? node14101 : 15'b000000011111111;
													assign node14101 = (inp[10]) ? node14103 : 15'b000000001111111;
														assign node14103 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14106 = (inp[2]) ? node14112 : node14107;
												assign node14107 = (inp[5]) ? 15'b000000011111111 : node14108;
													assign node14108 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14112 = (inp[14]) ? node14114 : 15'b000000000111111;
													assign node14114 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node14117 = (inp[0]) ? node14153 : node14118;
										assign node14118 = (inp[10]) ? node14132 : node14119;
											assign node14119 = (inp[13]) ? node14125 : node14120;
												assign node14120 = (inp[3]) ? 15'b000000011111111 : node14121;
													assign node14121 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14125 = (inp[14]) ? node14129 : node14126;
													assign node14126 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14129 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14132 = (inp[5]) ? node14138 : node14133;
												assign node14133 = (inp[2]) ? 15'b000000000111111 : node14134;
													assign node14134 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14138 = (inp[13]) ? node14144 : node14139;
													assign node14139 = (inp[2]) ? node14141 : 15'b000000001111111;
														assign node14141 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14144 = (inp[3]) ? node14150 : node14145;
														assign node14145 = (inp[14]) ? 15'b000000000111111 : node14146;
															assign node14146 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
														assign node14150 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node14153 = (inp[13]) ? node14181 : node14154;
											assign node14154 = (inp[3]) ? node14170 : node14155;
												assign node14155 = (inp[2]) ? node14163 : node14156;
													assign node14156 = (inp[5]) ? node14158 : 15'b000000011111111;
														assign node14158 = (inp[14]) ? 15'b000000000111111 : node14159;
															assign node14159 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14163 = (inp[14]) ? 15'b000000000111111 : node14164;
														assign node14164 = (inp[5]) ? node14166 : 15'b000000001111111;
															assign node14166 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14170 = (inp[10]) ? node14174 : node14171;
													assign node14171 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14174 = (inp[14]) ? 15'b000000000011111 : node14175;
														assign node14175 = (inp[5]) ? node14177 : 15'b000000000111111;
															assign node14177 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14181 = (inp[14]) ? node14191 : node14182;
												assign node14182 = (inp[3]) ? node14186 : node14183;
													assign node14183 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14186 = (inp[2]) ? 15'b000000000111111 : node14187;
														assign node14187 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14191 = (inp[3]) ? node14197 : node14192;
													assign node14192 = (inp[10]) ? 15'b000000000011111 : node14193;
														assign node14193 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14197 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node14200 = (inp[10]) ? node14280 : node14201;
									assign node14201 = (inp[0]) ? node14237 : node14202;
										assign node14202 = (inp[5]) ? node14222 : node14203;
											assign node14203 = (inp[13]) ? node14215 : node14204;
												assign node14204 = (inp[6]) ? 15'b000000011111111 : node14205;
													assign node14205 = (inp[2]) ? node14211 : node14206;
														assign node14206 = (inp[3]) ? 15'b000000111111111 : node14207;
															assign node14207 = (inp[14]) ? 15'b000000111111111 : 15'b000001111111111;
														assign node14211 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14215 = (inp[2]) ? node14217 : 15'b000000011111111;
													assign node14217 = (inp[14]) ? node14219 : 15'b000000001111111;
														assign node14219 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14222 = (inp[6]) ? node14228 : node14223;
												assign node14223 = (inp[13]) ? 15'b000000001111111 : node14224;
													assign node14224 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14228 = (inp[14]) ? node14234 : node14229;
													assign node14229 = (inp[13]) ? 15'b000000000111111 : node14230;
														assign node14230 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14234 = (inp[13]) ? 15'b000000000111111 : 15'b000000000011111;
										assign node14237 = (inp[14]) ? node14261 : node14238;
											assign node14238 = (inp[3]) ? node14252 : node14239;
												assign node14239 = (inp[6]) ? node14245 : node14240;
													assign node14240 = (inp[5]) ? 15'b000000001111111 : node14241;
														assign node14241 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14245 = (inp[2]) ? node14247 : 15'b000000001111111;
														assign node14247 = (inp[13]) ? 15'b000000000111111 : node14248;
															assign node14248 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14252 = (inp[2]) ? node14258 : node14253;
													assign node14253 = (inp[13]) ? 15'b000000000111111 : node14254;
														assign node14254 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14258 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14261 = (inp[6]) ? node14269 : node14262;
												assign node14262 = (inp[13]) ? node14266 : node14263;
													assign node14263 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14266 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14269 = (inp[2]) ? node14275 : node14270;
													assign node14270 = (inp[5]) ? node14272 : 15'b000000000111111;
														assign node14272 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node14275 = (inp[3]) ? node14277 : 15'b000000000011111;
														assign node14277 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node14280 = (inp[2]) ? node14304 : node14281;
										assign node14281 = (inp[5]) ? node14289 : node14282;
											assign node14282 = (inp[13]) ? 15'b000000000111111 : node14283;
												assign node14283 = (inp[0]) ? node14285 : 15'b000000011111111;
													assign node14285 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14289 = (inp[0]) ? node14297 : node14290;
												assign node14290 = (inp[3]) ? node14294 : node14291;
													assign node14291 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14294 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14297 = (inp[13]) ? node14301 : node14298;
													assign node14298 = (inp[3]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node14301 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node14304 = (inp[0]) ? node14318 : node14305;
											assign node14305 = (inp[6]) ? node14313 : node14306;
												assign node14306 = (inp[14]) ? node14310 : node14307;
													assign node14307 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14310 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14313 = (inp[3]) ? 15'b000000000011111 : node14314;
													assign node14314 = (inp[5]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14318 = (inp[5]) ? node14328 : node14319;
												assign node14319 = (inp[13]) ? node14323 : node14320;
													assign node14320 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14323 = (inp[6]) ? node14325 : 15'b000000000011111;
														assign node14325 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node14328 = (inp[13]) ? node14332 : node14329;
													assign node14329 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node14332 = (inp[14]) ? node14334 : 15'b000000000001111;
														assign node14334 = (inp[3]) ? 15'b000000000000011 : 15'b000000000000111;
							assign node14337 = (inp[8]) ? node14463 : node14338;
								assign node14338 = (inp[3]) ? node14390 : node14339;
									assign node14339 = (inp[10]) ? node14369 : node14340;
										assign node14340 = (inp[13]) ? node14356 : node14341;
											assign node14341 = (inp[14]) ? node14347 : node14342;
												assign node14342 = (inp[2]) ? 15'b000000011111111 : node14343;
													assign node14343 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14347 = (inp[0]) ? node14353 : node14348;
													assign node14348 = (inp[5]) ? 15'b000000001111111 : node14349;
														assign node14349 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14353 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14356 = (inp[2]) ? node14362 : node14357;
												assign node14357 = (inp[6]) ? node14359 : 15'b000000001111111;
													assign node14359 = (inp[5]) ? 15'b000000001111111 : 15'b000000000111111;
												assign node14362 = (inp[14]) ? 15'b000000000111111 : node14363;
													assign node14363 = (inp[6]) ? 15'b000000000111111 : node14364;
														assign node14364 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node14369 = (inp[6]) ? node14379 : node14370;
											assign node14370 = (inp[2]) ? node14372 : 15'b000000001111111;
												assign node14372 = (inp[14]) ? 15'b000000000011111 : node14373;
													assign node14373 = (inp[0]) ? 15'b000000000111111 : node14374;
														assign node14374 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14379 = (inp[13]) ? node14385 : node14380;
												assign node14380 = (inp[5]) ? node14382 : 15'b000000000111111;
													assign node14382 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14385 = (inp[2]) ? 15'b000000000011111 : node14386;
													assign node14386 = (inp[5]) ? 15'b000000000011111 : 15'b000000001111111;
									assign node14390 = (inp[14]) ? node14424 : node14391;
										assign node14391 = (inp[13]) ? node14411 : node14392;
											assign node14392 = (inp[2]) ? node14404 : node14393;
												assign node14393 = (inp[10]) ? node14397 : node14394;
													assign node14394 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14397 = (inp[0]) ? node14399 : 15'b000000001111111;
														assign node14399 = (inp[5]) ? 15'b000000000111111 : node14400;
															assign node14400 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14404 = (inp[10]) ? 15'b000000000001111 : node14405;
													assign node14405 = (inp[0]) ? 15'b000000000111111 : node14406;
														assign node14406 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14411 = (inp[0]) ? node14421 : node14412;
												assign node14412 = (inp[5]) ? node14418 : node14413;
													assign node14413 = (inp[6]) ? 15'b000000000111111 : node14414;
														assign node14414 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14418 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14421 = (inp[5]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node14424 = (inp[6]) ? node14448 : node14425;
											assign node14425 = (inp[0]) ? node14435 : node14426;
												assign node14426 = (inp[2]) ? node14430 : node14427;
													assign node14427 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14430 = (inp[10]) ? node14432 : 15'b000000000111111;
														assign node14432 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14435 = (inp[13]) ? node14439 : node14436;
													assign node14436 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14439 = (inp[5]) ? node14443 : node14440;
														assign node14440 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
														assign node14443 = (inp[10]) ? 15'b000000000001111 : node14444;
															assign node14444 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node14448 = (inp[2]) ? node14450 : 15'b000000000011111;
												assign node14450 = (inp[13]) ? node14456 : node14451;
													assign node14451 = (inp[0]) ? 15'b000000000001111 : node14452;
														assign node14452 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node14456 = (inp[5]) ? 15'b000000000000111 : node14457;
														assign node14457 = (inp[0]) ? node14459 : 15'b000000000001111;
															assign node14459 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node14463 = (inp[5]) ? node14541 : node14464;
									assign node14464 = (inp[14]) ? node14506 : node14465;
										assign node14465 = (inp[0]) ? node14485 : node14466;
											assign node14466 = (inp[10]) ? node14476 : node14467;
												assign node14467 = (inp[6]) ? 15'b000000000111111 : node14468;
													assign node14468 = (inp[13]) ? 15'b000000001111111 : node14469;
														assign node14469 = (inp[3]) ? node14471 : 15'b000000011111111;
															assign node14471 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14476 = (inp[3]) ? 15'b000000000011111 : node14477;
													assign node14477 = (inp[2]) ? 15'b000000000111111 : node14478;
														assign node14478 = (inp[6]) ? node14480 : 15'b000000001111111;
															assign node14480 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14485 = (inp[10]) ? node14499 : node14486;
												assign node14486 = (inp[6]) ? node14490 : node14487;
													assign node14487 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14490 = (inp[3]) ? 15'b000000000011111 : node14491;
														assign node14491 = (inp[2]) ? node14495 : node14492;
															assign node14492 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
															assign node14495 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14499 = (inp[13]) ? 15'b000000000011111 : node14500;
													assign node14500 = (inp[3]) ? 15'b000000000011111 : node14501;
														assign node14501 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node14506 = (inp[10]) ? node14526 : node14507;
											assign node14507 = (inp[0]) ? node14515 : node14508;
												assign node14508 = (inp[6]) ? node14510 : 15'b000000001111111;
													assign node14510 = (inp[2]) ? node14512 : 15'b000000000111111;
														assign node14512 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14515 = (inp[2]) ? node14523 : node14516;
													assign node14516 = (inp[13]) ? 15'b000000000011111 : node14517;
														assign node14517 = (inp[3]) ? node14519 : 15'b000000000111111;
															assign node14519 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14523 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node14526 = (inp[0]) ? node14534 : node14527;
												assign node14527 = (inp[13]) ? node14531 : node14528;
													assign node14528 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14531 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node14534 = (inp[2]) ? node14536 : 15'b000000000001111;
													assign node14536 = (inp[13]) ? 15'b000000000000111 : node14537;
														assign node14537 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node14541 = (inp[10]) ? node14565 : node14542;
										assign node14542 = (inp[2]) ? node14550 : node14543;
											assign node14543 = (inp[14]) ? node14545 : 15'b000000000111111;
												assign node14545 = (inp[6]) ? node14547 : 15'b000000000111111;
													assign node14547 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node14550 = (inp[6]) ? node14552 : 15'b000000000011111;
												assign node14552 = (inp[14]) ? 15'b000000000000111 : node14553;
													assign node14553 = (inp[0]) ? node14559 : node14554;
														assign node14554 = (inp[13]) ? node14556 : 15'b000000000011111;
															assign node14556 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
														assign node14559 = (inp[3]) ? node14561 : 15'b000000000001111;
															assign node14561 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node14565 = (inp[6]) ? node14591 : node14566;
											assign node14566 = (inp[0]) ? node14576 : node14567;
												assign node14567 = (inp[3]) ? node14569 : 15'b000000000011111;
													assign node14569 = (inp[2]) ? node14571 : 15'b000000000011111;
														assign node14571 = (inp[13]) ? 15'b000000000001111 : node14572;
															assign node14572 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node14576 = (inp[3]) ? node14584 : node14577;
													assign node14577 = (inp[14]) ? 15'b000000000001111 : node14578;
														assign node14578 = (inp[13]) ? node14580 : 15'b000000000111111;
															assign node14580 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node14584 = (inp[2]) ? 15'b000000000000111 : node14585;
														assign node14585 = (inp[13]) ? node14587 : 15'b000000000001111;
															assign node14587 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node14591 = (inp[14]) ? node14593 : 15'b000000000001111;
												assign node14593 = (inp[0]) ? node14595 : 15'b000000000000111;
													assign node14595 = (inp[13]) ? node14597 : 15'b000000000000111;
														assign node14597 = (inp[2]) ? 15'b000000000000011 : node14598;
															assign node14598 = (inp[3]) ? 15'b000000000000011 : 15'b000000000000111;
				assign node14602 = (inp[1]) ? node15690 : node14603;
					assign node14603 = (inp[5]) ? node15145 : node14604;
						assign node14604 = (inp[13]) ? node14850 : node14605;
							assign node14605 = (inp[14]) ? node14735 : node14606;
								assign node14606 = (inp[11]) ? node14684 : node14607;
									assign node14607 = (inp[6]) ? node14653 : node14608;
										assign node14608 = (inp[9]) ? node14630 : node14609;
											assign node14609 = (inp[2]) ? node14619 : node14610;
												assign node14610 = (inp[10]) ? node14616 : node14611;
													assign node14611 = (inp[3]) ? 15'b000001111111111 : node14612;
														assign node14612 = (inp[0]) ? 15'b000001111111111 : 15'b000011111111111;
													assign node14616 = (inp[0]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node14619 = (inp[8]) ? node14627 : node14620;
													assign node14620 = (inp[0]) ? 15'b000000111111111 : node14621;
														assign node14621 = (inp[10]) ? node14623 : 15'b000001111111111;
															assign node14623 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node14627 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node14630 = (inp[10]) ? node14640 : node14631;
												assign node14631 = (inp[8]) ? node14635 : node14632;
													assign node14632 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node14635 = (inp[0]) ? node14637 : 15'b000000111111111;
														assign node14637 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14640 = (inp[0]) ? node14648 : node14641;
													assign node14641 = (inp[2]) ? 15'b000000011111111 : node14642;
														assign node14642 = (inp[8]) ? node14644 : 15'b000000111111111;
															assign node14644 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14648 = (inp[8]) ? node14650 : 15'b000000011111111;
														assign node14650 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node14653 = (inp[8]) ? node14669 : node14654;
											assign node14654 = (inp[10]) ? node14660 : node14655;
												assign node14655 = (inp[0]) ? 15'b000000011111111 : node14656;
													assign node14656 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node14660 = (inp[3]) ? 15'b000000011111111 : node14661;
													assign node14661 = (inp[2]) ? node14663 : 15'b000000111111111;
														assign node14663 = (inp[9]) ? 15'b000000011111111 : node14664;
															assign node14664 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node14669 = (inp[0]) ? node14677 : node14670;
												assign node14670 = (inp[2]) ? 15'b000000011111111 : node14671;
													assign node14671 = (inp[3]) ? 15'b000000011111111 : node14672;
														assign node14672 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14677 = (inp[10]) ? node14681 : node14678;
													assign node14678 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14681 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node14684 = (inp[2]) ? node14720 : node14685;
										assign node14685 = (inp[10]) ? node14701 : node14686;
											assign node14686 = (inp[6]) ? node14694 : node14687;
												assign node14687 = (inp[0]) ? node14691 : node14688;
													assign node14688 = (inp[3]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node14691 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14694 = (inp[8]) ? node14696 : 15'b000000111111111;
													assign node14696 = (inp[9]) ? node14698 : 15'b000000011111111;
														assign node14698 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node14701 = (inp[9]) ? node14715 : node14702;
												assign node14702 = (inp[8]) ? node14708 : node14703;
													assign node14703 = (inp[3]) ? 15'b000000011111111 : node14704;
														assign node14704 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14708 = (inp[6]) ? 15'b000000001111111 : node14709;
														assign node14709 = (inp[0]) ? node14711 : 15'b000000011111111;
															assign node14711 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14715 = (inp[3]) ? node14717 : 15'b000000001111111;
													assign node14717 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node14720 = (inp[0]) ? node14728 : node14721;
											assign node14721 = (inp[9]) ? 15'b000000001111111 : node14722;
												assign node14722 = (inp[8]) ? node14724 : 15'b000000011111111;
													assign node14724 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node14728 = (inp[3]) ? node14732 : node14729;
												assign node14729 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14732 = (inp[9]) ? 15'b000000000111111 : 15'b000000000011111;
								assign node14735 = (inp[8]) ? node14785 : node14736;
									assign node14736 = (inp[3]) ? node14762 : node14737;
										assign node14737 = (inp[9]) ? node14751 : node14738;
											assign node14738 = (inp[2]) ? node14746 : node14739;
												assign node14739 = (inp[10]) ? node14743 : node14740;
													assign node14740 = (inp[11]) ? 15'b000000111111111 : 15'b000011111111111;
													assign node14743 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14746 = (inp[6]) ? 15'b000000011111111 : node14747;
													assign node14747 = (inp[0]) ? 15'b000000111111111 : 15'b000000011111111;
											assign node14751 = (inp[11]) ? node14755 : node14752;
												assign node14752 = (inp[10]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14755 = (inp[6]) ? node14759 : node14756;
													assign node14756 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14759 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node14762 = (inp[2]) ? node14774 : node14763;
											assign node14763 = (inp[9]) ? 15'b000000000111111 : node14764;
												assign node14764 = (inp[0]) ? node14768 : node14765;
													assign node14765 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14768 = (inp[6]) ? node14770 : 15'b000000011111111;
														assign node14770 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node14774 = (inp[11]) ? node14776 : 15'b000000001111111;
												assign node14776 = (inp[10]) ? node14782 : node14777;
													assign node14777 = (inp[9]) ? node14779 : 15'b000000001111111;
														assign node14779 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
													assign node14782 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node14785 = (inp[9]) ? node14817 : node14786;
										assign node14786 = (inp[11]) ? node14798 : node14787;
											assign node14787 = (inp[0]) ? node14793 : node14788;
												assign node14788 = (inp[10]) ? 15'b000000011111111 : node14789;
													assign node14789 = (inp[2]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14793 = (inp[10]) ? node14795 : 15'b000000011111111;
													assign node14795 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node14798 = (inp[0]) ? node14808 : node14799;
												assign node14799 = (inp[2]) ? node14805 : node14800;
													assign node14800 = (inp[10]) ? 15'b000000001111111 : node14801;
														assign node14801 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14805 = (inp[3]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node14808 = (inp[10]) ? node14814 : node14809;
													assign node14809 = (inp[3]) ? 15'b000000000111111 : node14810;
														assign node14810 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14814 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node14817 = (inp[3]) ? node14835 : node14818;
											assign node14818 = (inp[10]) ? node14826 : node14819;
												assign node14819 = (inp[0]) ? node14821 : 15'b000000011111111;
													assign node14821 = (inp[11]) ? 15'b000000000111111 : node14822;
														assign node14822 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14826 = (inp[0]) ? node14832 : node14827;
													assign node14827 = (inp[2]) ? 15'b000000000111111 : node14828;
														assign node14828 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14832 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14835 = (inp[0]) ? node14847 : node14836;
												assign node14836 = (inp[10]) ? node14840 : node14837;
													assign node14837 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14840 = (inp[6]) ? 15'b000000000011111 : node14841;
														assign node14841 = (inp[11]) ? node14843 : 15'b000000000111111;
															assign node14843 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14847 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
							assign node14850 = (inp[0]) ? node15000 : node14851;
								assign node14851 = (inp[3]) ? node14925 : node14852;
									assign node14852 = (inp[8]) ? node14890 : node14853;
										assign node14853 = (inp[14]) ? node14871 : node14854;
											assign node14854 = (inp[10]) ? node14864 : node14855;
												assign node14855 = (inp[6]) ? node14861 : node14856;
													assign node14856 = (inp[2]) ? node14858 : 15'b000001111111111;
														assign node14858 = (inp[9]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node14861 = (inp[9]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14864 = (inp[2]) ? node14866 : 15'b000000111111111;
													assign node14866 = (inp[9]) ? node14868 : 15'b000000011111111;
														assign node14868 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node14871 = (inp[6]) ? node14885 : node14872;
												assign node14872 = (inp[9]) ? node14878 : node14873;
													assign node14873 = (inp[2]) ? node14875 : 15'b000000111111111;
														assign node14875 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14878 = (inp[2]) ? node14880 : 15'b000000011111111;
														assign node14880 = (inp[11]) ? 15'b000000001111111 : node14881;
															assign node14881 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node14885 = (inp[10]) ? 15'b000000001111111 : node14886;
													assign node14886 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
										assign node14890 = (inp[14]) ? node14914 : node14891;
											assign node14891 = (inp[9]) ? node14903 : node14892;
												assign node14892 = (inp[2]) ? node14898 : node14893;
													assign node14893 = (inp[11]) ? node14895 : 15'b000000111111111;
														assign node14895 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node14898 = (inp[6]) ? 15'b000000011111111 : node14899;
														assign node14899 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node14903 = (inp[11]) ? node14907 : node14904;
													assign node14904 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14907 = (inp[2]) ? node14909 : 15'b000000001111111;
														assign node14909 = (inp[10]) ? 15'b000000000111111 : node14910;
															assign node14910 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14914 = (inp[11]) ? node14918 : node14915;
												assign node14915 = (inp[2]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node14918 = (inp[6]) ? 15'b000000000011111 : node14919;
													assign node14919 = (inp[10]) ? node14921 : 15'b000000000111111;
														assign node14921 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node14925 = (inp[9]) ? node14953 : node14926;
										assign node14926 = (inp[6]) ? node14942 : node14927;
											assign node14927 = (inp[8]) ? node14933 : node14928;
												assign node14928 = (inp[11]) ? 15'b000000011111111 : node14929;
													assign node14929 = (inp[2]) ? 15'b000000011111111 : 15'b000001111111111;
												assign node14933 = (inp[11]) ? node14937 : node14934;
													assign node14934 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14937 = (inp[2]) ? node14939 : 15'b000000001111111;
														assign node14939 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node14942 = (inp[8]) ? node14948 : node14943;
												assign node14943 = (inp[10]) ? node14945 : 15'b000000001111111;
													assign node14945 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14948 = (inp[11]) ? 15'b000000000111111 : node14949;
													assign node14949 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node14953 = (inp[8]) ? node14979 : node14954;
											assign node14954 = (inp[10]) ? node14970 : node14955;
												assign node14955 = (inp[11]) ? node14963 : node14956;
													assign node14956 = (inp[14]) ? 15'b000000001111111 : node14957;
														assign node14957 = (inp[6]) ? node14959 : 15'b000000011111111;
															assign node14959 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node14963 = (inp[6]) ? 15'b000000000011111 : node14964;
														assign node14964 = (inp[14]) ? node14966 : 15'b000000001111111;
															assign node14966 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node14970 = (inp[14]) ? node14974 : node14971;
													assign node14971 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node14974 = (inp[11]) ? 15'b000000000011111 : node14975;
														assign node14975 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node14979 = (inp[11]) ? node14993 : node14980;
												assign node14980 = (inp[14]) ? node14988 : node14981;
													assign node14981 = (inp[10]) ? node14983 : 15'b000000000111111;
														assign node14983 = (inp[6]) ? node14985 : 15'b000000000111111;
															assign node14985 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14988 = (inp[2]) ? 15'b000000000011111 : node14989;
														assign node14989 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node14993 = (inp[6]) ? node14997 : node14994;
													assign node14994 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node14997 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node15000 = (inp[10]) ? node15072 : node15001;
									assign node15001 = (inp[14]) ? node15033 : node15002;
										assign node15002 = (inp[8]) ? node15020 : node15003;
											assign node15003 = (inp[2]) ? node15009 : node15004;
												assign node15004 = (inp[6]) ? 15'b000000011111111 : node15005;
													assign node15005 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node15009 = (inp[6]) ? node15017 : node15010;
													assign node15010 = (inp[3]) ? 15'b000000001111111 : node15011;
														assign node15011 = (inp[9]) ? node15013 : 15'b000000011111111;
															assign node15013 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15017 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15020 = (inp[6]) ? node15028 : node15021;
												assign node15021 = (inp[2]) ? node15023 : 15'b000000001111111;
													assign node15023 = (inp[11]) ? node15025 : 15'b000000001111111;
														assign node15025 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15028 = (inp[3]) ? 15'b000000000001111 : node15029;
													assign node15029 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node15033 = (inp[2]) ? node15057 : node15034;
											assign node15034 = (inp[9]) ? node15050 : node15035;
												assign node15035 = (inp[6]) ? node15045 : node15036;
													assign node15036 = (inp[8]) ? node15040 : node15037;
														assign node15037 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node15040 = (inp[11]) ? node15042 : 15'b000000001111111;
															assign node15042 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15045 = (inp[11]) ? 15'b000000000111111 : node15046;
														assign node15046 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15050 = (inp[6]) ? node15052 : 15'b000000000111111;
													assign node15052 = (inp[8]) ? 15'b000000000111111 : node15053;
														assign node15053 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15057 = (inp[9]) ? node15067 : node15058;
												assign node15058 = (inp[3]) ? node15062 : node15059;
													assign node15059 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15062 = (inp[8]) ? 15'b000000000011111 : node15063;
														assign node15063 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
												assign node15067 = (inp[11]) ? 15'b000000000001111 : node15068;
													assign node15068 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node15072 = (inp[2]) ? node15106 : node15073;
										assign node15073 = (inp[11]) ? node15091 : node15074;
											assign node15074 = (inp[9]) ? node15078 : node15075;
												assign node15075 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15078 = (inp[3]) ? node15086 : node15079;
													assign node15079 = (inp[14]) ? 15'b000000000111111 : node15080;
														assign node15080 = (inp[6]) ? node15082 : 15'b000000001111111;
															assign node15082 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15086 = (inp[6]) ? node15088 : 15'b000000000111111;
														assign node15088 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node15091 = (inp[14]) ? node15097 : node15092;
												assign node15092 = (inp[6]) ? 15'b000000000111111 : node15093;
													assign node15093 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15097 = (inp[6]) ? node15101 : node15098;
													assign node15098 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15101 = (inp[8]) ? node15103 : 15'b000000000011111;
														assign node15103 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node15106 = (inp[9]) ? node15122 : node15107;
											assign node15107 = (inp[11]) ? node15113 : node15108;
												assign node15108 = (inp[14]) ? node15110 : 15'b000000000111111;
													assign node15110 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15113 = (inp[3]) ? node15117 : node15114;
													assign node15114 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15117 = (inp[6]) ? node15119 : 15'b000000000011111;
														assign node15119 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15122 = (inp[14]) ? node15132 : node15123;
												assign node15123 = (inp[11]) ? node15129 : node15124;
													assign node15124 = (inp[3]) ? 15'b000000000011111 : node15125;
														assign node15125 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15129 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15132 = (inp[3]) ? node15138 : node15133;
													assign node15133 = (inp[8]) ? node15135 : 15'b000000000011111;
														assign node15135 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15138 = (inp[8]) ? node15140 : 15'b000000000001111;
														assign node15140 = (inp[6]) ? 15'b000000000000111 : node15141;
															assign node15141 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
						assign node15145 = (inp[10]) ? node15429 : node15146;
							assign node15146 = (inp[3]) ? node15280 : node15147;
								assign node15147 = (inp[13]) ? node15225 : node15148;
									assign node15148 = (inp[0]) ? node15176 : node15149;
										assign node15149 = (inp[2]) ? node15157 : node15150;
											assign node15150 = (inp[9]) ? node15152 : 15'b000001111111111;
												assign node15152 = (inp[6]) ? 15'b000000011111111 : node15153;
													assign node15153 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node15157 = (inp[11]) ? node15171 : node15158;
												assign node15158 = (inp[14]) ? node15166 : node15159;
													assign node15159 = (inp[9]) ? node15161 : 15'b000000111111111;
														assign node15161 = (inp[6]) ? node15163 : 15'b000000011111111;
															assign node15163 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15166 = (inp[6]) ? node15168 : 15'b000000011111111;
														assign node15168 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15171 = (inp[6]) ? 15'b000000001111111 : node15172;
													assign node15172 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node15176 = (inp[6]) ? node15206 : node15177;
											assign node15177 = (inp[2]) ? node15197 : node15178;
												assign node15178 = (inp[11]) ? node15190 : node15179;
													assign node15179 = (inp[8]) ? node15185 : node15180;
														assign node15180 = (inp[9]) ? node15182 : 15'b000000111111111;
															assign node15182 = (inp[14]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node15185 = (inp[9]) ? node15187 : 15'b000000011111111;
															assign node15187 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15190 = (inp[9]) ? node15192 : 15'b000000011111111;
														assign node15192 = (inp[8]) ? 15'b000000001111111 : node15193;
															assign node15193 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15197 = (inp[9]) ? node15201 : node15198;
													assign node15198 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15201 = (inp[11]) ? 15'b000000000111111 : node15202;
														assign node15202 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15206 = (inp[9]) ? node15218 : node15207;
												assign node15207 = (inp[8]) ? node15215 : node15208;
													assign node15208 = (inp[14]) ? 15'b000000001111111 : node15209;
														assign node15209 = (inp[11]) ? node15211 : 15'b000000011111111;
															assign node15211 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15215 = (inp[11]) ? 15'b000000000111111 : 15'b000000011111111;
												assign node15218 = (inp[8]) ? 15'b000000000111111 : node15219;
													assign node15219 = (inp[14]) ? 15'b000000000111111 : node15220;
														assign node15220 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node15225 = (inp[2]) ? node15251 : node15226;
										assign node15226 = (inp[14]) ? node15238 : node15227;
											assign node15227 = (inp[11]) ? node15233 : node15228;
												assign node15228 = (inp[0]) ? 15'b000000011111111 : node15229;
													assign node15229 = (inp[8]) ? 15'b000000111111111 : 15'b000001111111111;
												assign node15233 = (inp[0]) ? 15'b000000001111111 : node15234;
													assign node15234 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node15238 = (inp[6]) ? node15246 : node15239;
												assign node15239 = (inp[9]) ? node15243 : node15240;
													assign node15240 = (inp[0]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node15243 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15246 = (inp[8]) ? 15'b000000000111111 : node15247;
													assign node15247 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node15251 = (inp[6]) ? node15269 : node15252;
											assign node15252 = (inp[0]) ? node15258 : node15253;
												assign node15253 = (inp[11]) ? 15'b000000001111111 : node15254;
													assign node15254 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15258 = (inp[11]) ? node15264 : node15259;
													assign node15259 = (inp[9]) ? node15261 : 15'b000000001111111;
														assign node15261 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15264 = (inp[14]) ? 15'b000000000011111 : node15265;
														assign node15265 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node15269 = (inp[14]) ? node15277 : node15270;
												assign node15270 = (inp[11]) ? node15274 : node15271;
													assign node15271 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15274 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15277 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node15280 = (inp[9]) ? node15352 : node15281;
									assign node15281 = (inp[6]) ? node15317 : node15282;
										assign node15282 = (inp[11]) ? node15296 : node15283;
											assign node15283 = (inp[14]) ? node15289 : node15284;
												assign node15284 = (inp[0]) ? 15'b000000011111111 : node15285;
													assign node15285 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node15289 = (inp[2]) ? 15'b000000001111111 : node15290;
													assign node15290 = (inp[13]) ? 15'b000000001111111 : node15291;
														assign node15291 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node15296 = (inp[0]) ? node15312 : node15297;
												assign node15297 = (inp[2]) ? node15307 : node15298;
													assign node15298 = (inp[8]) ? node15304 : node15299;
														assign node15299 = (inp[14]) ? 15'b000000011111111 : node15300;
															assign node15300 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
														assign node15304 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15307 = (inp[13]) ? 15'b000000000111111 : node15308;
														assign node15308 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15312 = (inp[2]) ? node15314 : 15'b000000000111111;
													assign node15314 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node15317 = (inp[2]) ? node15333 : node15318;
											assign node15318 = (inp[8]) ? node15328 : node15319;
												assign node15319 = (inp[14]) ? node15325 : node15320;
													assign node15320 = (inp[13]) ? 15'b000000001111111 : node15321;
														assign node15321 = (inp[0]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15325 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15328 = (inp[11]) ? 15'b000000000111111 : node15329;
													assign node15329 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15333 = (inp[8]) ? node15341 : node15334;
												assign node15334 = (inp[0]) ? node15338 : node15335;
													assign node15335 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15338 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15341 = (inp[0]) ? node15349 : node15342;
													assign node15342 = (inp[14]) ? node15344 : 15'b000000000111111;
														assign node15344 = (inp[13]) ? 15'b000000000011111 : node15345;
															assign node15345 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15349 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node15352 = (inp[6]) ? node15390 : node15353;
										assign node15353 = (inp[0]) ? node15371 : node15354;
											assign node15354 = (inp[2]) ? node15362 : node15355;
												assign node15355 = (inp[14]) ? node15357 : 15'b000000001111111;
													assign node15357 = (inp[13]) ? node15359 : 15'b000000001111111;
														assign node15359 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15362 = (inp[14]) ? node15368 : node15363;
													assign node15363 = (inp[8]) ? 15'b000000000111111 : node15364;
														assign node15364 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15368 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node15371 = (inp[14]) ? node15381 : node15372;
												assign node15372 = (inp[8]) ? node15378 : node15373;
													assign node15373 = (inp[11]) ? 15'b000000000111111 : node15374;
														assign node15374 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15378 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15381 = (inp[2]) ? node15387 : node15382;
													assign node15382 = (inp[11]) ? 15'b000000000011111 : node15383;
														assign node15383 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15387 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node15390 = (inp[8]) ? node15404 : node15391;
											assign node15391 = (inp[2]) ? node15399 : node15392;
												assign node15392 = (inp[0]) ? node15396 : node15393;
													assign node15393 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15396 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15399 = (inp[13]) ? 15'b000000000011111 : node15400;
													assign node15400 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node15404 = (inp[2]) ? node15412 : node15405;
												assign node15405 = (inp[0]) ? node15409 : node15406;
													assign node15406 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15409 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15412 = (inp[13]) ? node15420 : node15413;
													assign node15413 = (inp[14]) ? 15'b000000000001111 : node15414;
														assign node15414 = (inp[11]) ? node15416 : 15'b000000000011111;
															assign node15416 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15420 = (inp[0]) ? node15424 : node15421;
														assign node15421 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
														assign node15424 = (inp[14]) ? node15426 : 15'b000000000000111;
															assign node15426 = (inp[11]) ? 15'b000000000000011 : 15'b000000000000111;
							assign node15429 = (inp[9]) ? node15577 : node15430;
								assign node15430 = (inp[2]) ? node15504 : node15431;
									assign node15431 = (inp[14]) ? node15469 : node15432;
										assign node15432 = (inp[13]) ? node15444 : node15433;
											assign node15433 = (inp[8]) ? node15435 : 15'b000000011111111;
												assign node15435 = (inp[11]) ? 15'b000000001111111 : node15436;
													assign node15436 = (inp[0]) ? node15438 : 15'b000000011111111;
														assign node15438 = (inp[3]) ? 15'b000000001111111 : node15439;
															assign node15439 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node15444 = (inp[11]) ? node15460 : node15445;
												assign node15445 = (inp[0]) ? node15451 : node15446;
													assign node15446 = (inp[6]) ? 15'b000000001111111 : node15447;
														assign node15447 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node15451 = (inp[3]) ? node15455 : node15452;
														assign node15452 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node15455 = (inp[6]) ? 15'b000000000111111 : node15456;
															assign node15456 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15460 = (inp[6]) ? node15466 : node15461;
													assign node15461 = (inp[3]) ? 15'b000000000111111 : node15462;
														assign node15462 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15466 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node15469 = (inp[0]) ? node15485 : node15470;
											assign node15470 = (inp[8]) ? node15478 : node15471;
												assign node15471 = (inp[13]) ? 15'b000000001111111 : node15472;
													assign node15472 = (inp[6]) ? 15'b000000001111111 : node15473;
														assign node15473 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15478 = (inp[13]) ? node15482 : node15479;
													assign node15479 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15482 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node15485 = (inp[11]) ? node15495 : node15486;
												assign node15486 = (inp[13]) ? node15492 : node15487;
													assign node15487 = (inp[3]) ? 15'b000000000111111 : node15488;
														assign node15488 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15492 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15495 = (inp[6]) ? node15499 : node15496;
													assign node15496 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15499 = (inp[8]) ? 15'b000000000000111 : node15500;
														assign node15500 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
									assign node15504 = (inp[13]) ? node15542 : node15505;
										assign node15505 = (inp[11]) ? node15517 : node15506;
											assign node15506 = (inp[0]) ? node15512 : node15507;
												assign node15507 = (inp[3]) ? 15'b000000000111111 : node15508;
													assign node15508 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15512 = (inp[8]) ? 15'b000000000111111 : node15513;
													assign node15513 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15517 = (inp[8]) ? node15529 : node15518;
												assign node15518 = (inp[3]) ? node15522 : node15519;
													assign node15519 = (inp[0]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15522 = (inp[14]) ? node15524 : 15'b000000000111111;
														assign node15524 = (inp[6]) ? 15'b000000000011111 : node15525;
															assign node15525 = (inp[0]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15529 = (inp[14]) ? node15539 : node15530;
													assign node15530 = (inp[0]) ? node15536 : node15531;
														assign node15531 = (inp[3]) ? node15533 : 15'b000000000111111;
															assign node15533 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
														assign node15536 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15539 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node15542 = (inp[3]) ? node15560 : node15543;
											assign node15543 = (inp[0]) ? node15553 : node15544;
												assign node15544 = (inp[6]) ? node15546 : 15'b000000000111111;
													assign node15546 = (inp[14]) ? node15548 : 15'b000000000111111;
														assign node15548 = (inp[8]) ? 15'b000000000011111 : node15549;
															assign node15549 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15553 = (inp[11]) ? node15557 : node15554;
													assign node15554 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15557 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15560 = (inp[0]) ? node15572 : node15561;
												assign node15561 = (inp[11]) ? node15569 : node15562;
													assign node15562 = (inp[8]) ? node15564 : 15'b000000000011111;
														assign node15564 = (inp[6]) ? node15566 : 15'b000000000011111;
															assign node15566 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15569 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node15572 = (inp[6]) ? node15574 : 15'b000000000001111;
													assign node15574 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node15577 = (inp[8]) ? node15623 : node15578;
									assign node15578 = (inp[14]) ? node15596 : node15579;
										assign node15579 = (inp[11]) ? node15585 : node15580;
											assign node15580 = (inp[2]) ? 15'b000000000111111 : node15581;
												assign node15581 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node15585 = (inp[3]) ? node15587 : 15'b000000000111111;
												assign node15587 = (inp[0]) ? node15593 : node15588;
													assign node15588 = (inp[6]) ? 15'b000000000011111 : node15589;
														assign node15589 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15593 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node15596 = (inp[13]) ? node15608 : node15597;
											assign node15597 = (inp[3]) ? node15603 : node15598;
												assign node15598 = (inp[0]) ? node15600 : 15'b000000001111111;
													assign node15600 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15603 = (inp[11]) ? node15605 : 15'b000000000011111;
													assign node15605 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15608 = (inp[6]) ? node15612 : node15609;
												assign node15609 = (inp[0]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15612 = (inp[3]) ? node15616 : node15613;
													assign node15613 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15616 = (inp[2]) ? 15'b000000000000111 : node15617;
														assign node15617 = (inp[0]) ? node15619 : 15'b000000000001111;
															assign node15619 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node15623 = (inp[6]) ? node15661 : node15624;
										assign node15624 = (inp[0]) ? node15642 : node15625;
											assign node15625 = (inp[3]) ? node15633 : node15626;
												assign node15626 = (inp[14]) ? 15'b000000000011111 : node15627;
													assign node15627 = (inp[13]) ? node15629 : 15'b000000001111111;
														assign node15629 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15633 = (inp[2]) ? node15637 : node15634;
													assign node15634 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15637 = (inp[11]) ? 15'b000000000001111 : node15638;
														assign node15638 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15642 = (inp[11]) ? node15652 : node15643;
												assign node15643 = (inp[3]) ? node15647 : node15644;
													assign node15644 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15647 = (inp[2]) ? node15649 : 15'b000000000011111;
														assign node15649 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node15652 = (inp[13]) ? node15656 : node15653;
													assign node15653 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node15656 = (inp[3]) ? node15658 : 15'b000000000001111;
														assign node15658 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node15661 = (inp[14]) ? node15677 : node15662;
											assign node15662 = (inp[2]) ? node15672 : node15663;
												assign node15663 = (inp[11]) ? node15665 : 15'b000000000111111;
													assign node15665 = (inp[0]) ? 15'b000000000001111 : node15666;
														assign node15666 = (inp[13]) ? node15668 : 15'b000000000011111;
															assign node15668 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node15672 = (inp[11]) ? 15'b000000000000111 : node15673;
													assign node15673 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node15677 = (inp[13]) ? node15685 : node15678;
												assign node15678 = (inp[11]) ? node15680 : 15'b000000000011111;
													assign node15680 = (inp[3]) ? 15'b000000000000111 : node15681;
														assign node15681 = (inp[0]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node15685 = (inp[2]) ? node15687 : 15'b000000000000111;
													assign node15687 = (inp[11]) ? 15'b000000000000001 : 15'b000000000000111;
					assign node15690 = (inp[0]) ? node16206 : node15691;
						assign node15691 = (inp[10]) ? node15937 : node15692;
							assign node15692 = (inp[5]) ? node15792 : node15693;
								assign node15693 = (inp[11]) ? node15747 : node15694;
									assign node15694 = (inp[9]) ? node15728 : node15695;
										assign node15695 = (inp[6]) ? node15713 : node15696;
											assign node15696 = (inp[14]) ? node15708 : node15697;
												assign node15697 = (inp[3]) ? node15705 : node15698;
													assign node15698 = (inp[13]) ? node15700 : 15'b000001111111111;
														assign node15700 = (inp[8]) ? 15'b000000111111111 : node15701;
															assign node15701 = (inp[2]) ? 15'b000000111111111 : 15'b000001111111111;
													assign node15705 = (inp[13]) ? 15'b000000001111111 : 15'b000000111111111;
												assign node15708 = (inp[8]) ? node15710 : 15'b000000011111111;
													assign node15710 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
											assign node15713 = (inp[8]) ? node15723 : node15714;
												assign node15714 = (inp[14]) ? 15'b000000011111111 : node15715;
													assign node15715 = (inp[2]) ? node15717 : 15'b000000111111111;
														assign node15717 = (inp[3]) ? 15'b000000011111111 : node15718;
															assign node15718 = (inp[13]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node15723 = (inp[2]) ? 15'b000000000111111 : node15724;
													assign node15724 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
										assign node15728 = (inp[14]) ? node15744 : node15729;
											assign node15729 = (inp[2]) ? node15737 : node15730;
												assign node15730 = (inp[3]) ? node15732 : 15'b000000111111111;
													assign node15732 = (inp[8]) ? 15'b000000011111111 : node15733;
														assign node15733 = (inp[6]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node15737 = (inp[6]) ? node15741 : node15738;
													assign node15738 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15741 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15744 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
									assign node15747 = (inp[13]) ? node15771 : node15748;
										assign node15748 = (inp[2]) ? node15758 : node15749;
											assign node15749 = (inp[3]) ? node15753 : node15750;
												assign node15750 = (inp[8]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node15753 = (inp[14]) ? node15755 : 15'b000000001111111;
													assign node15755 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15758 = (inp[6]) ? node15766 : node15759;
												assign node15759 = (inp[14]) ? 15'b000000001111111 : node15760;
													assign node15760 = (inp[9]) ? 15'b000000001111111 : node15761;
														assign node15761 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15766 = (inp[3]) ? node15768 : 15'b000000001111111;
													assign node15768 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node15771 = (inp[3]) ? node15783 : node15772;
											assign node15772 = (inp[8]) ? node15780 : node15773;
												assign node15773 = (inp[6]) ? node15777 : node15774;
													assign node15774 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15777 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15780 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node15783 = (inp[2]) ? node15789 : node15784;
												assign node15784 = (inp[8]) ? node15786 : 15'b000000000111111;
													assign node15786 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15789 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
								assign node15792 = (inp[2]) ? node15868 : node15793;
									assign node15793 = (inp[13]) ? node15829 : node15794;
										assign node15794 = (inp[8]) ? node15814 : node15795;
											assign node15795 = (inp[6]) ? node15807 : node15796;
												assign node15796 = (inp[9]) ? node15800 : node15797;
													assign node15797 = (inp[3]) ? 15'b000000011111111 : 15'b000000111111111;
													assign node15800 = (inp[14]) ? 15'b000000001111111 : node15801;
														assign node15801 = (inp[11]) ? node15803 : 15'b000000011111111;
															assign node15803 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node15807 = (inp[3]) ? 15'b000000001111111 : node15808;
													assign node15808 = (inp[9]) ? 15'b000000001111111 : node15809;
														assign node15809 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node15814 = (inp[9]) ? node15822 : node15815;
												assign node15815 = (inp[6]) ? node15819 : node15816;
													assign node15816 = (inp[14]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15819 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15822 = (inp[3]) ? 15'b000000000011111 : node15823;
													assign node15823 = (inp[6]) ? node15825 : 15'b000000001111111;
														assign node15825 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node15829 = (inp[14]) ? node15853 : node15830;
											assign node15830 = (inp[8]) ? node15846 : node15831;
												assign node15831 = (inp[11]) ? node15839 : node15832;
													assign node15832 = (inp[9]) ? node15834 : 15'b000000011111111;
														assign node15834 = (inp[6]) ? 15'b000000001111111 : node15835;
															assign node15835 = (inp[3]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15839 = (inp[6]) ? 15'b000000000011111 : node15840;
														assign node15840 = (inp[9]) ? node15842 : 15'b000000001111111;
															assign node15842 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15846 = (inp[9]) ? node15848 : 15'b000000000111111;
													assign node15848 = (inp[11]) ? 15'b000000000011111 : node15849;
														assign node15849 = (inp[6]) ? 15'b000000000011111 : 15'b000000001111111;
											assign node15853 = (inp[9]) ? node15859 : node15854;
												assign node15854 = (inp[3]) ? node15856 : 15'b000000000111111;
													assign node15856 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15859 = (inp[11]) ? node15865 : node15860;
													assign node15860 = (inp[6]) ? node15862 : 15'b000000000111111;
														assign node15862 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node15865 = (inp[3]) ? 15'b000000000000111 : 15'b000000000011111;
									assign node15868 = (inp[6]) ? node15912 : node15869;
										assign node15869 = (inp[8]) ? node15897 : node15870;
											assign node15870 = (inp[14]) ? node15890 : node15871;
												assign node15871 = (inp[3]) ? node15883 : node15872;
													assign node15872 = (inp[13]) ? node15878 : node15873;
														assign node15873 = (inp[9]) ? node15875 : 15'b000000011111111;
															assign node15875 = (inp[11]) ? 15'b000000001111111 : 15'b000000011111111;
														assign node15878 = (inp[9]) ? node15880 : 15'b000000001111111;
															assign node15880 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node15883 = (inp[11]) ? node15885 : 15'b000000001111111;
														assign node15885 = (inp[13]) ? node15887 : 15'b000000000111111;
															assign node15887 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15890 = (inp[3]) ? 15'b000000000011111 : node15891;
													assign node15891 = (inp[9]) ? node15893 : 15'b000000000111111;
														assign node15893 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node15897 = (inp[3]) ? node15905 : node15898;
												assign node15898 = (inp[9]) ? 15'b000000000011111 : node15899;
													assign node15899 = (inp[11]) ? node15901 : 15'b000000001111111;
														assign node15901 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15905 = (inp[14]) ? node15907 : 15'b000000000011111;
													assign node15907 = (inp[13]) ? 15'b000000000001111 : node15908;
														assign node15908 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node15912 = (inp[13]) ? node15920 : node15913;
											assign node15913 = (inp[8]) ? 15'b000000000011111 : node15914;
												assign node15914 = (inp[14]) ? node15916 : 15'b000000000111111;
													assign node15916 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node15920 = (inp[14]) ? node15928 : node15921;
												assign node15921 = (inp[8]) ? node15923 : 15'b000000000011111;
													assign node15923 = (inp[11]) ? 15'b000000000001111 : node15924;
														assign node15924 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node15928 = (inp[8]) ? 15'b000000000001111 : node15929;
													assign node15929 = (inp[3]) ? node15931 : 15'b000000000011111;
														assign node15931 = (inp[9]) ? 15'b000000000000111 : node15932;
															assign node15932 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
							assign node15937 = (inp[3]) ? node16059 : node15938;
								assign node15938 = (inp[8]) ? node15986 : node15939;
									assign node15939 = (inp[6]) ? node15961 : node15940;
										assign node15940 = (inp[9]) ? node15952 : node15941;
											assign node15941 = (inp[5]) ? node15945 : node15942;
												assign node15942 = (inp[11]) ? 15'b000000011111111 : 15'b000000111111111;
												assign node15945 = (inp[13]) ? node15949 : node15946;
													assign node15946 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15949 = (inp[11]) ? 15'b000000001111111 : 15'b000000000111111;
											assign node15952 = (inp[14]) ? 15'b000000000111111 : node15953;
												assign node15953 = (inp[13]) ? node15957 : node15954;
													assign node15954 = (inp[11]) ? 15'b000000001111111 : 15'b000000111111111;
													assign node15957 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
										assign node15961 = (inp[2]) ? node15973 : node15962;
											assign node15962 = (inp[11]) ? node15964 : 15'b000000001111111;
												assign node15964 = (inp[14]) ? 15'b000000000111111 : node15965;
													assign node15965 = (inp[13]) ? node15967 : 15'b000000001111111;
														assign node15967 = (inp[5]) ? 15'b000000000111111 : node15968;
															assign node15968 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
											assign node15973 = (inp[13]) ? node15981 : node15974;
												assign node15974 = (inp[9]) ? 15'b000000000011111 : node15975;
													assign node15975 = (inp[5]) ? node15977 : 15'b000000001111111;
														assign node15977 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node15981 = (inp[14]) ? 15'b000000000011111 : node15982;
													assign node15982 = (inp[9]) ? 15'b000000000001111 : 15'b000000000111111;
									assign node15986 = (inp[9]) ? node16028 : node15987;
										assign node15987 = (inp[6]) ? node16011 : node15988;
											assign node15988 = (inp[13]) ? node16002 : node15989;
												assign node15989 = (inp[2]) ? node15995 : node15990;
													assign node15990 = (inp[14]) ? node15992 : 15'b000000011111111;
														assign node15992 = (inp[5]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node15995 = (inp[5]) ? 15'b000000000111111 : node15996;
														assign node15996 = (inp[14]) ? node15998 : 15'b000000001111111;
															assign node15998 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node16002 = (inp[2]) ? node16008 : node16003;
													assign node16003 = (inp[5]) ? 15'b000000000111111 : node16004;
														assign node16004 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16008 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node16011 = (inp[5]) ? node16017 : node16012;
												assign node16012 = (inp[14]) ? 15'b000000000111111 : node16013;
													assign node16013 = (inp[13]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node16017 = (inp[14]) ? node16025 : node16018;
													assign node16018 = (inp[13]) ? node16020 : 15'b000000000111111;
														assign node16020 = (inp[11]) ? 15'b000000000011111 : node16021;
															assign node16021 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16025 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node16028 = (inp[2]) ? node16044 : node16029;
											assign node16029 = (inp[11]) ? node16037 : node16030;
												assign node16030 = (inp[14]) ? node16034 : node16031;
													assign node16031 = (inp[5]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16034 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16037 = (inp[13]) ? node16039 : 15'b000000000011111;
													assign node16039 = (inp[5]) ? node16041 : 15'b000000000011111;
														assign node16041 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node16044 = (inp[5]) ? node16054 : node16045;
												assign node16045 = (inp[6]) ? 15'b000000000001111 : node16046;
													assign node16046 = (inp[13]) ? node16048 : 15'b000000000011111;
														assign node16048 = (inp[11]) ? node16050 : 15'b000000000011111;
															assign node16050 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16054 = (inp[11]) ? node16056 : 15'b000000000001111;
													assign node16056 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node16059 = (inp[5]) ? node16135 : node16060;
									assign node16060 = (inp[8]) ? node16098 : node16061;
										assign node16061 = (inp[11]) ? node16075 : node16062;
											assign node16062 = (inp[14]) ? node16066 : node16063;
												assign node16063 = (inp[2]) ? 15'b000000001111111 : 15'b000000011111111;
												assign node16066 = (inp[2]) ? node16072 : node16067;
													assign node16067 = (inp[9]) ? 15'b000000000111111 : node16068;
														assign node16068 = (inp[13]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node16072 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node16075 = (inp[14]) ? node16091 : node16076;
												assign node16076 = (inp[2]) ? node16084 : node16077;
													assign node16077 = (inp[13]) ? 15'b000000000111111 : node16078;
														assign node16078 = (inp[9]) ? node16080 : 15'b000000001111111;
															assign node16080 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16084 = (inp[13]) ? 15'b000000000011111 : node16085;
														assign node16085 = (inp[6]) ? node16087 : 15'b000000000111111;
															assign node16087 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16091 = (inp[9]) ? node16095 : node16092;
													assign node16092 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16095 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node16098 = (inp[11]) ? node16118 : node16099;
											assign node16099 = (inp[13]) ? node16107 : node16100;
												assign node16100 = (inp[14]) ? node16104 : node16101;
													assign node16101 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16104 = (inp[2]) ? 15'b000000000111111 : 15'b000000000011111;
												assign node16107 = (inp[6]) ? node16115 : node16108;
													assign node16108 = (inp[14]) ? 15'b000000000011111 : node16109;
														assign node16109 = (inp[9]) ? node16111 : 15'b000000000111111;
															assign node16111 = (inp[2]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16115 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node16118 = (inp[6]) ? node16126 : node16119;
												assign node16119 = (inp[13]) ? node16123 : node16120;
													assign node16120 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16123 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16126 = (inp[13]) ? node16130 : node16127;
													assign node16127 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node16130 = (inp[2]) ? 15'b000000000000111 : node16131;
														assign node16131 = (inp[14]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node16135 = (inp[9]) ? node16177 : node16136;
										assign node16136 = (inp[6]) ? node16154 : node16137;
											assign node16137 = (inp[2]) ? node16147 : node16138;
												assign node16138 = (inp[11]) ? node16142 : node16139;
													assign node16139 = (inp[14]) ? 15'b000000000111111 : 15'b000000011111111;
													assign node16142 = (inp[8]) ? node16144 : 15'b000000000111111;
														assign node16144 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16147 = (inp[13]) ? node16151 : node16148;
													assign node16148 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16151 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node16154 = (inp[13]) ? node16168 : node16155;
												assign node16155 = (inp[2]) ? node16161 : node16156;
													assign node16156 = (inp[11]) ? 15'b000000000011111 : node16157;
														assign node16157 = (inp[8]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16161 = (inp[11]) ? node16163 : 15'b000000000011111;
														assign node16163 = (inp[14]) ? node16165 : 15'b000000000001111;
															assign node16165 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node16168 = (inp[14]) ? 15'b000000000000111 : node16169;
													assign node16169 = (inp[11]) ? node16171 : 15'b000000000001111;
														assign node16171 = (inp[2]) ? node16173 : 15'b000000000001111;
															assign node16173 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node16177 = (inp[13]) ? node16193 : node16178;
											assign node16178 = (inp[6]) ? node16184 : node16179;
												assign node16179 = (inp[11]) ? node16181 : 15'b000000000011111;
													assign node16181 = (inp[8]) ? 15'b000000000011111 : 15'b000000000001111;
												assign node16184 = (inp[11]) ? node16190 : node16185;
													assign node16185 = (inp[8]) ? 15'b000000000001111 : node16186;
														assign node16186 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node16190 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node16193 = (inp[6]) ? node16199 : node16194;
												assign node16194 = (inp[2]) ? node16196 : 15'b000000000001111;
													assign node16196 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node16199 = (inp[2]) ? node16203 : node16200;
													assign node16200 = (inp[8]) ? 15'b000000000000111 : 15'b000000000011111;
													assign node16203 = (inp[8]) ? 15'b000000000000001 : 15'b000000000000011;
						assign node16206 = (inp[5]) ? node16480 : node16207;
							assign node16207 = (inp[2]) ? node16333 : node16208;
								assign node16208 = (inp[13]) ? node16266 : node16209;
									assign node16209 = (inp[14]) ? node16241 : node16210;
										assign node16210 = (inp[11]) ? node16224 : node16211;
											assign node16211 = (inp[10]) ? node16213 : 15'b000000111111111;
												assign node16213 = (inp[3]) ? node16219 : node16214;
													assign node16214 = (inp[6]) ? node16216 : 15'b000000011111111;
														assign node16216 = (inp[9]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node16219 = (inp[8]) ? 15'b000000000111111 : node16220;
														assign node16220 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
											assign node16224 = (inp[6]) ? node16234 : node16225;
												assign node16225 = (inp[3]) ? node16229 : node16226;
													assign node16226 = (inp[8]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node16229 = (inp[8]) ? node16231 : 15'b000000001111111;
														assign node16231 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node16234 = (inp[3]) ? node16238 : node16235;
													assign node16235 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16238 = (inp[10]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node16241 = (inp[10]) ? node16255 : node16242;
											assign node16242 = (inp[8]) ? node16248 : node16243;
												assign node16243 = (inp[3]) ? node16245 : 15'b000000011111111;
													assign node16245 = (inp[9]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node16248 = (inp[9]) ? node16252 : node16249;
													assign node16249 = (inp[11]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16252 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node16255 = (inp[8]) ? node16261 : node16256;
												assign node16256 = (inp[6]) ? node16258 : 15'b000000000111111;
													assign node16258 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16261 = (inp[3]) ? 15'b000000000011111 : node16262;
													assign node16262 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
									assign node16266 = (inp[3]) ? node16306 : node16267;
										assign node16267 = (inp[8]) ? node16293 : node16268;
											assign node16268 = (inp[14]) ? node16282 : node16269;
												assign node16269 = (inp[11]) ? node16275 : node16270;
													assign node16270 = (inp[9]) ? 15'b000000001111111 : node16271;
														assign node16271 = (inp[10]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node16275 = (inp[6]) ? node16277 : 15'b000000001111111;
														assign node16277 = (inp[9]) ? 15'b000000000111111 : node16278;
															assign node16278 = (inp[10]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node16282 = (inp[9]) ? node16290 : node16283;
													assign node16283 = (inp[10]) ? node16285 : 15'b000000001111111;
														assign node16285 = (inp[6]) ? node16287 : 15'b000000000111111;
															assign node16287 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16290 = (inp[10]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node16293 = (inp[9]) ? node16301 : node16294;
												assign node16294 = (inp[6]) ? 15'b000000000011111 : node16295;
													assign node16295 = (inp[11]) ? node16297 : 15'b000000000111111;
														assign node16297 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16301 = (inp[14]) ? 15'b000000000011111 : node16302;
													assign node16302 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node16306 = (inp[10]) ? node16326 : node16307;
											assign node16307 = (inp[8]) ? node16317 : node16308;
												assign node16308 = (inp[6]) ? node16310 : 15'b000000000111111;
													assign node16310 = (inp[9]) ? 15'b000000000011111 : node16311;
														assign node16311 = (inp[14]) ? node16313 : 15'b000000000111111;
															assign node16313 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16317 = (inp[6]) ? node16321 : node16318;
													assign node16318 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16321 = (inp[11]) ? 15'b000000000001111 : node16322;
														assign node16322 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node16326 = (inp[14]) ? node16330 : node16327;
												assign node16327 = (inp[9]) ? 15'b000000000011111 : 15'b000000000001111;
												assign node16330 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
								assign node16333 = (inp[10]) ? node16411 : node16334;
									assign node16334 = (inp[13]) ? node16368 : node16335;
										assign node16335 = (inp[8]) ? node16355 : node16336;
											assign node16336 = (inp[3]) ? node16346 : node16337;
												assign node16337 = (inp[9]) ? node16341 : node16338;
													assign node16338 = (inp[6]) ? 15'b000000001111111 : 15'b000000011111111;
													assign node16341 = (inp[11]) ? node16343 : 15'b000000001111111;
														assign node16343 = (inp[6]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node16346 = (inp[9]) ? node16352 : node16347;
													assign node16347 = (inp[6]) ? node16349 : 15'b000000001111111;
														assign node16349 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16352 = (inp[6]) ? 15'b000000000011111 : 15'b000000000111111;
											assign node16355 = (inp[6]) ? node16361 : node16356;
												assign node16356 = (inp[9]) ? 15'b000000000111111 : node16357;
													assign node16357 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node16361 = (inp[3]) ? node16365 : node16362;
													assign node16362 = (inp[14]) ? 15'b000000000111111 : 15'b000000000011111;
													assign node16365 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node16368 = (inp[9]) ? node16390 : node16369;
											assign node16369 = (inp[14]) ? node16379 : node16370;
												assign node16370 = (inp[8]) ? node16372 : 15'b000000000111111;
													assign node16372 = (inp[6]) ? 15'b000000000011111 : node16373;
														assign node16373 = (inp[3]) ? node16375 : 15'b000000000111111;
															assign node16375 = (inp[11]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16379 = (inp[6]) ? node16385 : node16380;
													assign node16380 = (inp[8]) ? node16382 : 15'b000000000111111;
														assign node16382 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node16385 = (inp[3]) ? node16387 : 15'b000000000011111;
														assign node16387 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node16390 = (inp[14]) ? node16400 : node16391;
												assign node16391 = (inp[6]) ? node16395 : node16392;
													assign node16392 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16395 = (inp[3]) ? 15'b000000000001111 : node16396;
														assign node16396 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16400 = (inp[3]) ? node16404 : node16401;
													assign node16401 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node16404 = (inp[6]) ? node16406 : 15'b000000000001111;
														assign node16406 = (inp[8]) ? 15'b000000000000111 : node16407;
															assign node16407 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node16411 = (inp[11]) ? node16447 : node16412;
										assign node16412 = (inp[3]) ? node16428 : node16413;
											assign node16413 = (inp[13]) ? node16419 : node16414;
												assign node16414 = (inp[6]) ? node16416 : 15'b000000000111111;
													assign node16416 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16419 = (inp[9]) ? node16425 : node16420;
													assign node16420 = (inp[6]) ? 15'b000000000011111 : node16421;
														assign node16421 = (inp[14]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16425 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node16428 = (inp[13]) ? node16438 : node16429;
												assign node16429 = (inp[8]) ? 15'b000000000011111 : node16430;
													assign node16430 = (inp[14]) ? node16432 : 15'b000000000011111;
														assign node16432 = (inp[6]) ? node16434 : 15'b000000000011111;
															assign node16434 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16438 = (inp[9]) ? node16442 : node16439;
													assign node16439 = (inp[6]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node16442 = (inp[8]) ? 15'b000000000000011 : node16443;
														assign node16443 = (inp[6]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node16447 = (inp[3]) ? node16465 : node16448;
											assign node16448 = (inp[6]) ? node16454 : node16449;
												assign node16449 = (inp[9]) ? node16451 : 15'b000000000011111;
													assign node16451 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16454 = (inp[14]) ? node16458 : node16455;
													assign node16455 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node16458 = (inp[8]) ? node16460 : 15'b000000000011111;
														assign node16460 = (inp[9]) ? 15'b000000000000111 : node16461;
															assign node16461 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node16465 = (inp[13]) ? node16473 : node16466;
												assign node16466 = (inp[14]) ? 15'b000000000001111 : node16467;
													assign node16467 = (inp[8]) ? node16469 : 15'b000000000001111;
														assign node16469 = (inp[6]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node16473 = (inp[9]) ? 15'b000000000000011 : node16474;
													assign node16474 = (inp[14]) ? 15'b000000000000111 : node16475;
														assign node16475 = (inp[8]) ? 15'b000000000000111 : 15'b000000000001111;
							assign node16480 = (inp[6]) ? node16610 : node16481;
								assign node16481 = (inp[13]) ? node16545 : node16482;
									assign node16482 = (inp[11]) ? node16508 : node16483;
										assign node16483 = (inp[9]) ? node16491 : node16484;
											assign node16484 = (inp[14]) ? node16486 : 15'b000000001111111;
												assign node16486 = (inp[8]) ? node16488 : 15'b000000001111111;
													assign node16488 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node16491 = (inp[10]) ? node16503 : node16492;
												assign node16492 = (inp[8]) ? node16498 : node16493;
													assign node16493 = (inp[3]) ? 15'b000000000111111 : node16494;
														assign node16494 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16498 = (inp[14]) ? 15'b000000000011111 : node16499;
														assign node16499 = (inp[3]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node16503 = (inp[2]) ? 15'b000000000011111 : node16504;
													assign node16504 = (inp[8]) ? 15'b000000000011111 : 15'b000000000111111;
										assign node16508 = (inp[8]) ? node16526 : node16509;
											assign node16509 = (inp[10]) ? node16517 : node16510;
												assign node16510 = (inp[14]) ? node16514 : node16511;
													assign node16511 = (inp[2]) ? 15'b000000000111111 : 15'b000000001111111;
													assign node16514 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16517 = (inp[3]) ? node16521 : node16518;
													assign node16518 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16521 = (inp[2]) ? 15'b000000000000111 : node16522;
														assign node16522 = (inp[9]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node16526 = (inp[14]) ? node16536 : node16527;
												assign node16527 = (inp[10]) ? node16533 : node16528;
													assign node16528 = (inp[2]) ? 15'b000000000011111 : node16529;
														assign node16529 = (inp[3]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16533 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16536 = (inp[9]) ? node16542 : node16537;
													assign node16537 = (inp[10]) ? 15'b000000000001111 : node16538;
														assign node16538 = (inp[2]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node16542 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
									assign node16545 = (inp[9]) ? node16573 : node16546;
										assign node16546 = (inp[2]) ? node16558 : node16547;
											assign node16547 = (inp[11]) ? node16555 : node16548;
												assign node16548 = (inp[8]) ? 15'b000000000111111 : node16549;
													assign node16549 = (inp[3]) ? node16551 : 15'b000000001111111;
														assign node16551 = (inp[14]) ? 15'b000000000111111 : 15'b000000001111111;
												assign node16555 = (inp[3]) ? 15'b000000000001111 : 15'b000000001111111;
											assign node16558 = (inp[14]) ? node16568 : node16559;
												assign node16559 = (inp[8]) ? node16561 : 15'b000000000011111;
													assign node16561 = (inp[10]) ? node16563 : 15'b000000000011111;
														assign node16563 = (inp[11]) ? 15'b000000000001111 : node16564;
															assign node16564 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16568 = (inp[11]) ? 15'b000000000000111 : node16569;
													assign node16569 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
										assign node16573 = (inp[8]) ? node16589 : node16574;
											assign node16574 = (inp[10]) ? node16580 : node16575;
												assign node16575 = (inp[2]) ? node16577 : 15'b000000000011111;
													assign node16577 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16580 = (inp[11]) ? node16584 : node16581;
													assign node16581 = (inp[14]) ? 15'b000000000011111 : 15'b000000000001111;
													assign node16584 = (inp[2]) ? 15'b000000000000111 : node16585;
														assign node16585 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node16589 = (inp[2]) ? node16597 : node16590;
												assign node16590 = (inp[11]) ? 15'b000000000000111 : node16591;
													assign node16591 = (inp[10]) ? 15'b000000000001111 : node16592;
														assign node16592 = (inp[14]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16597 = (inp[3]) ? node16599 : 15'b000000000001111;
													assign node16599 = (inp[11]) ? node16605 : node16600;
														assign node16600 = (inp[14]) ? node16602 : 15'b000000000000111;
															assign node16602 = (inp[10]) ? 15'b000000000000011 : 15'b000000000000111;
														assign node16605 = (inp[14]) ? node16607 : 15'b000000000000011;
															assign node16607 = (inp[10]) ? 15'b000000000000001 : 15'b000000000000011;
								assign node16610 = (inp[14]) ? node16670 : node16611;
									assign node16611 = (inp[8]) ? node16639 : node16612;
										assign node16612 = (inp[11]) ? node16630 : node16613;
											assign node16613 = (inp[13]) ? node16623 : node16614;
												assign node16614 = (inp[2]) ? node16616 : 15'b000000001111111;
													assign node16616 = (inp[10]) ? node16618 : 15'b000000000111111;
														assign node16618 = (inp[3]) ? 15'b000000000011111 : node16619;
															assign node16619 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16623 = (inp[2]) ? node16627 : node16624;
													assign node16624 = (inp[9]) ? 15'b000000000011111 : 15'b000000000111111;
													assign node16627 = (inp[3]) ? 15'b000000000001111 : 15'b000000000011111;
											assign node16630 = (inp[2]) ? node16636 : node16631;
												assign node16631 = (inp[3]) ? 15'b000000000011111 : node16632;
													assign node16632 = (inp[13]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16636 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
										assign node16639 = (inp[3]) ? node16655 : node16640;
											assign node16640 = (inp[9]) ? node16644 : node16641;
												assign node16641 = (inp[13]) ? 15'b000000000011111 : 15'b000000000111111;
												assign node16644 = (inp[13]) ? node16650 : node16645;
													assign node16645 = (inp[2]) ? node16647 : 15'b000000000011111;
														assign node16647 = (inp[11]) ? 15'b000000000001111 : 15'b000000000011111;
													assign node16650 = (inp[2]) ? node16652 : 15'b000000000001111;
														assign node16652 = (inp[11]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node16655 = (inp[9]) ? node16661 : node16656;
												assign node16656 = (inp[11]) ? node16658 : 15'b000000000001111;
													assign node16658 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node16661 = (inp[2]) ? node16667 : node16662;
													assign node16662 = (inp[11]) ? 15'b000000000000111 : node16663;
														assign node16663 = (inp[13]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node16667 = (inp[11]) ? 15'b000000000000011 : 15'b000000000000111;
									assign node16670 = (inp[13]) ? node16702 : node16671;
										assign node16671 = (inp[2]) ? node16685 : node16672;
											assign node16672 = (inp[3]) ? node16678 : node16673;
												assign node16673 = (inp[9]) ? node16675 : 15'b000000000011111;
													assign node16675 = (inp[8]) ? 15'b000000000001111 : 15'b000000000011111;
												assign node16678 = (inp[10]) ? node16682 : node16679;
													assign node16679 = (inp[11]) ? 15'b000000000011111 : 15'b000000000001111;
													assign node16682 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
											assign node16685 = (inp[10]) ? node16691 : node16686;
												assign node16686 = (inp[11]) ? node16688 : 15'b000000000001111;
													assign node16688 = (inp[3]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node16691 = (inp[11]) ? node16695 : node16692;
													assign node16692 = (inp[9]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node16695 = (inp[9]) ? node16697 : 15'b000000000000111;
														assign node16697 = (inp[8]) ? node16699 : 15'b000000000000011;
															assign node16699 = (inp[3]) ? 15'b000000000000001 : 15'b000000000000011;
										assign node16702 = (inp[8]) ? node16722 : node16703;
											assign node16703 = (inp[9]) ? node16711 : node16704;
												assign node16704 = (inp[3]) ? node16708 : node16705;
													assign node16705 = (inp[11]) ? 15'b000000000001111 : 15'b000000000111111;
													assign node16708 = (inp[10]) ? 15'b000000000000111 : 15'b000000000001111;
												assign node16711 = (inp[3]) ? node16715 : node16712;
													assign node16712 = (inp[2]) ? 15'b000000000000111 : 15'b000000000001111;
													assign node16715 = (inp[10]) ? node16717 : 15'b000000000000111;
														assign node16717 = (inp[2]) ? node16719 : 15'b000000000000011;
															assign node16719 = (inp[11]) ? 15'b000000000000001 : 15'b000000000000011;
											assign node16722 = (inp[11]) ? node16728 : node16723;
												assign node16723 = (inp[10]) ? node16725 : 15'b000000000000111;
													assign node16725 = (inp[2]) ? 15'b000000000000011 : 15'b000000000000111;
												assign node16728 = (inp[3]) ? node16732 : node16729;
													assign node16729 = (inp[10]) ? 15'b000000000000011 : 15'b000000000000111;
													assign node16732 = (inp[2]) ? 15'b000000000000001 : node16733;
														assign node16733 = (inp[10]) ? 15'b000000000000001 : 15'b000000000000011;

endmodule