module dtc_split66_bm97 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node118;

	assign outp = (inp[3]) ? node28 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b000;
			assign node3 = (inp[9]) ? node5 : 3'b000;
				assign node5 = (inp[7]) ? node7 : 3'b001;
					assign node7 = (inp[10]) ? node9 : 3'b000;
						assign node9 = (inp[4]) ? node19 : node10;
							assign node10 = (inp[11]) ? node12 : 3'b000;
								assign node12 = (inp[5]) ? node16 : node13;
									assign node13 = (inp[8]) ? 3'b100 : 3'b000;
									assign node16 = (inp[8]) ? 3'b101 : 3'b001;
							assign node19 = (inp[11]) ? node21 : 3'b100;
								assign node21 = (inp[5]) ? node25 : node22;
									assign node22 = (inp[8]) ? 3'b100 : 3'b000;
									assign node25 = (inp[8]) ? 3'b110 : 3'b010;
		assign node28 = (inp[9]) ? node56 : node29;
			assign node29 = (inp[6]) ? 3'b000 : node30;
				assign node30 = (inp[7]) ? 3'b000 : node31;
					assign node31 = (inp[4]) ? node33 : 3'b100;
						assign node33 = (inp[11]) ? node41 : node34;
							assign node34 = (inp[8]) ? 3'b100 : node35;
								assign node35 = (inp[10]) ? node37 : 3'b100;
									assign node37 = (inp[1]) ? 3'b100 : 3'b000;
							assign node41 = (inp[5]) ? node49 : node42;
								assign node42 = (inp[10]) ? node46 : node43;
									assign node43 = (inp[1]) ? 3'b100 : 3'b100;
									assign node46 = (inp[8]) ? 3'b000 : 3'b100;
								assign node49 = (inp[0]) ? 3'b000 : node50;
									assign node50 = (inp[2]) ? 3'b000 : 3'b100;
			assign node56 = (inp[4]) ? node78 : node57;
				assign node57 = (inp[6]) ? node61 : node58;
					assign node58 = (inp[7]) ? 3'b110 : 3'b000;
					assign node61 = (inp[7]) ? node63 : 3'b110;
						assign node63 = (inp[10]) ? node65 : 3'b000;
							assign node65 = (inp[5]) ? node71 : node66;
								assign node66 = (inp[1]) ? node68 : 3'b010;
									assign node68 = (inp[0]) ? 3'b010 : 3'b010;
								assign node71 = (inp[11]) ? node75 : node72;
									assign node72 = (inp[2]) ? 3'b000 : 3'b000;
									assign node75 = (inp[2]) ? 3'b100 : 3'b100;
				assign node78 = (inp[6]) ? node112 : node79;
					assign node79 = (inp[7]) ? node101 : node80;
						assign node80 = (inp[10]) ? node90 : node81;
							assign node81 = (inp[11]) ? node83 : 3'b010;
								assign node83 = (inp[5]) ? node87 : node84;
									assign node84 = (inp[0]) ? 3'b010 : 3'b010;
									assign node87 = (inp[2]) ? 3'b110 : 3'b110;
							assign node90 = (inp[11]) ? node96 : node91;
								assign node91 = (inp[8]) ? 3'b001 : node92;
									assign node92 = (inp[1]) ? 3'b001 : 3'b101;
								assign node96 = (inp[8]) ? 3'b101 : node97;
									assign node97 = (inp[0]) ? 3'b101 : 3'b011;
						assign node101 = (inp[11]) ? node103 : 3'b001;
							assign node103 = (inp[10]) ? node105 : 3'b001;
								assign node105 = (inp[8]) ? node109 : node106;
									assign node106 = (inp[2]) ? 3'b001 : 3'b001;
									assign node109 = (inp[0]) ? 3'b110 : 3'b110;
					assign node112 = (inp[7]) ? 3'b000 : node113;
						assign node113 = (inp[11]) ? node115 : 3'b000;
							assign node115 = (inp[10]) ? node117 : 3'b000;
								assign node117 = (inp[8]) ? 3'b100 : node118;
									assign node118 = (inp[0]) ? 3'b010 : 3'b010;

endmodule