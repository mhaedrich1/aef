module dtc_split33_bm12 (
	input  wire [9-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node10;
	wire [1-1:0] node11;
	wire [1-1:0] node13;
	wire [1-1:0] node16;
	wire [1-1:0] node17;
	wire [1-1:0] node19;
	wire [1-1:0] node20;
	wire [1-1:0] node25;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node29;
	wire [1-1:0] node31;
	wire [1-1:0] node34;
	wire [1-1:0] node36;
	wire [1-1:0] node37;
	wire [1-1:0] node41;
	wire [1-1:0] node42;
	wire [1-1:0] node43;
	wire [1-1:0] node45;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node51;
	wire [1-1:0] node56;
	wire [1-1:0] node57;
	wire [1-1:0] node58;
	wire [1-1:0] node59;
	wire [1-1:0] node61;
	wire [1-1:0] node63;
	wire [1-1:0] node66;
	wire [1-1:0] node67;
	wire [1-1:0] node71;
	wire [1-1:0] node72;
	wire [1-1:0] node74;
	wire [1-1:0] node75;
	wire [1-1:0] node79;
	wire [1-1:0] node80;
	wire [1-1:0] node81;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node91;
	wire [1-1:0] node94;
	wire [1-1:0] node97;
	wire [1-1:0] node98;
	wire [1-1:0] node99;

	assign outp = (inp[5]) ? node56 : node1;
		assign node1 = (inp[6]) ? node25 : node2;
			assign node2 = (inp[1]) ? node10 : node3;
				assign node3 = (inp[7]) ? node5 : 1'b1;
					assign node5 = (inp[0]) ? node7 : 1'b1;
						assign node7 = (inp[2]) ? 1'b0 : 1'b1;
				assign node10 = (inp[8]) ? node16 : node11;
					assign node11 = (inp[3]) ? node13 : 1'b1;
						assign node13 = (inp[7]) ? 1'b0 : 1'b1;
					assign node16 = (inp[2]) ? 1'b0 : node17;
						assign node17 = (inp[3]) ? node19 : 1'b1;
							assign node19 = (inp[7]) ? 1'b0 : node20;
								assign node20 = (inp[4]) ? 1'b0 : 1'b1;
			assign node25 = (inp[8]) ? node41 : node26;
				assign node26 = (inp[1]) ? node34 : node27;
					assign node27 = (inp[0]) ? node29 : 1'b1;
						assign node29 = (inp[3]) ? node31 : 1'b1;
							assign node31 = (inp[7]) ? 1'b0 : 1'b1;
					assign node34 = (inp[4]) ? node36 : 1'b1;
						assign node36 = (inp[3]) ? 1'b0 : node37;
							assign node37 = (inp[7]) ? 1'b0 : 1'b1;
				assign node41 = (inp[4]) ? 1'b0 : node42;
					assign node42 = (inp[7]) ? node48 : node43;
						assign node43 = (inp[0]) ? node45 : 1'b1;
							assign node45 = (inp[2]) ? 1'b0 : 1'b1;
						assign node48 = (inp[2]) ? 1'b0 : node49;
							assign node49 = (inp[0]) ? node51 : 1'b1;
								assign node51 = (inp[3]) ? 1'b0 : 1'b1;
		assign node56 = (inp[8]) ? node86 : node57;
			assign node57 = (inp[7]) ? node71 : node58;
				assign node58 = (inp[6]) ? node66 : node59;
					assign node59 = (inp[2]) ? node61 : 1'b1;
						assign node61 = (inp[3]) ? node63 : 1'b1;
							assign node63 = (inp[0]) ? 1'b0 : 1'b1;
					assign node66 = (inp[1]) ? 1'b0 : node67;
						assign node67 = (inp[4]) ? 1'b0 : 1'b1;
				assign node71 = (inp[4]) ? node79 : node72;
					assign node72 = (inp[3]) ? node74 : 1'b1;
						assign node74 = (inp[0]) ? 1'b0 : node75;
							assign node75 = (inp[2]) ? 1'b0 : 1'b1;
					assign node79 = (inp[1]) ? 1'b0 : node80;
						assign node80 = (inp[2]) ? 1'b0 : node81;
							assign node81 = (inp[0]) ? 1'b0 : 1'b1;
			assign node86 = (inp[7]) ? 1'b0 : node87;
				assign node87 = (inp[2]) ? node97 : node88;
					assign node88 = (inp[4]) ? node94 : node89;
						assign node89 = (inp[6]) ? node91 : 1'b1;
							assign node91 = (inp[0]) ? 1'b0 : 1'b1;
						assign node94 = (inp[1]) ? 1'b0 : 1'b1;
					assign node97 = (inp[3]) ? 1'b0 : node98;
						assign node98 = (inp[0]) ? 1'b0 : node99;
							assign node99 = (inp[4]) ? 1'b0 : 1'b1;

endmodule