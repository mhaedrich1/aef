module dtc_split125_bm73 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node15;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node113;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node210;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node271;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node296;
	wire [3-1:0] node297;
	wire [3-1:0] node299;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node329;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node345;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node351;
	wire [3-1:0] node355;
	wire [3-1:0] node356;
	wire [3-1:0] node357;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node379;
	wire [3-1:0] node381;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node389;
	wire [3-1:0] node390;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node397;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node411;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node432;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node435;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node444;
	wire [3-1:0] node446;
	wire [3-1:0] node448;

	assign outp = (inp[9]) ? node158 : node1;
		assign node1 = (inp[3]) ? node117 : node2;
			assign node2 = (inp[6]) ? node76 : node3;
				assign node3 = (inp[7]) ? node41 : node4;
					assign node4 = (inp[4]) ? node30 : node5;
						assign node5 = (inp[10]) ? node23 : node6;
							assign node6 = (inp[0]) ? node18 : node7;
								assign node7 = (inp[2]) ? node9 : 3'b101;
									assign node9 = (inp[11]) ? node15 : node10;
										assign node10 = (inp[5]) ? 3'b001 : node11;
											assign node11 = (inp[8]) ? 3'b001 : 3'b101;
										assign node15 = (inp[8]) ? 3'b101 : 3'b011;
								assign node18 = (inp[11]) ? node20 : 3'b001;
									assign node20 = (inp[5]) ? 3'b001 : 3'b101;
							assign node23 = (inp[5]) ? node25 : 3'b111;
								assign node25 = (inp[8]) ? 3'b101 : node26;
									assign node26 = (inp[11]) ? 3'b111 : 3'b011;
						assign node30 = (inp[10]) ? node36 : node31;
							assign node31 = (inp[11]) ? node33 : 3'b010;
								assign node33 = (inp[8]) ? 3'b010 : 3'b110;
							assign node36 = (inp[2]) ? 3'b101 : node37;
								assign node37 = (inp[1]) ? 3'b001 : 3'b011;
					assign node41 = (inp[5]) ? node59 : node42;
						assign node42 = (inp[8]) ? node52 : node43;
							assign node43 = (inp[11]) ? node49 : node44;
								assign node44 = (inp[0]) ? 3'b110 : node45;
									assign node45 = (inp[4]) ? 3'b100 : 3'b110;
								assign node49 = (inp[4]) ? 3'b010 : 3'b011;
							assign node52 = (inp[2]) ? node54 : 3'b110;
								assign node54 = (inp[4]) ? node56 : 3'b101;
									assign node56 = (inp[10]) ? 3'b110 : 3'b100;
						assign node59 = (inp[10]) ? node67 : node60;
							assign node60 = (inp[4]) ? node64 : node61;
								assign node61 = (inp[0]) ? 3'b010 : 3'b100;
								assign node64 = (inp[11]) ? 3'b100 : 3'b000;
							assign node67 = (inp[1]) ? node69 : 3'b010;
								assign node69 = (inp[11]) ? 3'b110 : node70;
									assign node70 = (inp[8]) ? node72 : 3'b001;
										assign node72 = (inp[2]) ? 3'b100 : 3'b110;
				assign node76 = (inp[4]) ? node100 : node77;
					assign node77 = (inp[7]) ? 3'b000 : node78;
						assign node78 = (inp[5]) ? node88 : node79;
							assign node79 = (inp[8]) ? node83 : node80;
								assign node80 = (inp[10]) ? 3'b001 : 3'b010;
								assign node83 = (inp[11]) ? node85 : 3'b010;
									assign node85 = (inp[10]) ? 3'b110 : 3'b100;
							assign node88 = (inp[8]) ? node92 : node89;
								assign node89 = (inp[2]) ? 3'b110 : 3'b100;
								assign node92 = (inp[11]) ? node96 : node93;
									assign node93 = (inp[10]) ? 3'b100 : 3'b000;
									assign node96 = (inp[10]) ? 3'b010 : 3'b000;
					assign node100 = (inp[7]) ? 3'b000 : node101;
						assign node101 = (inp[2]) ? node107 : node102;
							assign node102 = (inp[0]) ? node104 : 3'b000;
								assign node104 = (inp[11]) ? 3'b010 : 3'b000;
							assign node107 = (inp[11]) ? node109 : 3'b000;
								assign node109 = (inp[10]) ? node111 : 3'b000;
									assign node111 = (inp[0]) ? node113 : 3'b100;
										assign node113 = (inp[8]) ? 3'b000 : 3'b100;
			assign node117 = (inp[6]) ? 3'b000 : node118;
				assign node118 = (inp[11]) ? node132 : node119;
					assign node119 = (inp[10]) ? node121 : 3'b000;
						assign node121 = (inp[7]) ? node125 : node122;
							assign node122 = (inp[0]) ? 3'b000 : 3'b100;
							assign node125 = (inp[2]) ? 3'b000 : node126;
								assign node126 = (inp[1]) ? node128 : 3'b000;
									assign node128 = (inp[0]) ? 3'b000 : 3'b100;
					assign node132 = (inp[4]) ? node148 : node133;
						assign node133 = (inp[7]) ? node141 : node134;
							assign node134 = (inp[5]) ? 3'b010 : node135;
								assign node135 = (inp[10]) ? 3'b001 : node136;
									assign node136 = (inp[8]) ? 3'b100 : 3'b010;
							assign node141 = (inp[8]) ? node145 : node142;
								assign node142 = (inp[10]) ? 3'b010 : 3'b000;
								assign node145 = (inp[5]) ? 3'b000 : 3'b100;
						assign node148 = (inp[7]) ? 3'b000 : node149;
							assign node149 = (inp[0]) ? node151 : 3'b010;
								assign node151 = (inp[5]) ? 3'b000 : node152;
									assign node152 = (inp[1]) ? 3'b100 : 3'b000;
		assign node158 = (inp[6]) ? node314 : node159;
			assign node159 = (inp[3]) ? node201 : node160;
				assign node160 = (inp[10]) ? node192 : node161;
					assign node161 = (inp[7]) ? node173 : node162;
						assign node162 = (inp[4]) ? node164 : 3'b111;
							assign node164 = (inp[5]) ? node168 : node165;
								assign node165 = (inp[11]) ? 3'b111 : 3'b011;
								assign node168 = (inp[2]) ? 3'b011 : node169;
									assign node169 = (inp[8]) ? 3'b101 : 3'b011;
						assign node173 = (inp[8]) ? node183 : node174;
							assign node174 = (inp[4]) ? node180 : node175;
								assign node175 = (inp[11]) ? 3'b111 : node176;
									assign node176 = (inp[5]) ? 3'b011 : 3'b111;
								assign node180 = (inp[0]) ? 3'b101 : 3'b111;
							assign node183 = (inp[11]) ? node189 : node184;
								assign node184 = (inp[5]) ? 3'b101 : node185;
									assign node185 = (inp[4]) ? 3'b001 : 3'b011;
								assign node189 = (inp[1]) ? 3'b001 : 3'b011;
					assign node192 = (inp[1]) ? 3'b111 : node193;
						assign node193 = (inp[7]) ? node195 : 3'b111;
							assign node195 = (inp[8]) ? node197 : 3'b111;
								assign node197 = (inp[2]) ? 3'b111 : 3'b011;
				assign node201 = (inp[10]) ? node255 : node202;
					assign node202 = (inp[4]) ? node238 : node203;
						assign node203 = (inp[1]) ? node217 : node204;
							assign node204 = (inp[11]) ? node206 : 3'b101;
								assign node206 = (inp[7]) ? node210 : node207;
									assign node207 = (inp[2]) ? 3'b001 : 3'b011;
									assign node210 = (inp[5]) ? 3'b110 : node211;
										assign node211 = (inp[8]) ? 3'b001 : node212;
											assign node212 = (inp[0]) ? 3'b001 : 3'b101;
							assign node217 = (inp[7]) ? node227 : node218;
								assign node218 = (inp[0]) ? node224 : node219;
									assign node219 = (inp[11]) ? node221 : 3'b101;
										assign node221 = (inp[5]) ? 3'b001 : 3'b011;
									assign node224 = (inp[8]) ? 3'b110 : 3'b101;
								assign node227 = (inp[0]) ? node231 : node228;
									assign node228 = (inp[11]) ? 3'b110 : 3'b100;
									assign node231 = (inp[11]) ? node233 : 3'b010;
										assign node233 = (inp[5]) ? 3'b110 : node234;
											assign node234 = (inp[8]) ? 3'b110 : 3'b001;
						assign node238 = (inp[7]) ? node248 : node239;
							assign node239 = (inp[8]) ? 3'b010 : node240;
								assign node240 = (inp[5]) ? node244 : node241;
									assign node241 = (inp[11]) ? 3'b001 : 3'b110;
									assign node244 = (inp[11]) ? 3'b110 : 3'b010;
							assign node248 = (inp[5]) ? node252 : node249;
								assign node249 = (inp[11]) ? 3'b010 : 3'b100;
								assign node252 = (inp[8]) ? 3'b000 : 3'b100;
					assign node255 = (inp[4]) ? node287 : node256;
						assign node256 = (inp[7]) ? node266 : node257;
							assign node257 = (inp[11]) ? 3'b111 : node258;
								assign node258 = (inp[1]) ? 3'b011 : node259;
									assign node259 = (inp[8]) ? node261 : 3'b111;
										assign node261 = (inp[0]) ? 3'b101 : 3'b011;
							assign node266 = (inp[2]) ? node276 : node267;
								assign node267 = (inp[0]) ? 3'b110 : node268;
									assign node268 = (inp[8]) ? 3'b011 : node269;
										assign node269 = (inp[11]) ? node271 : 3'b011;
											assign node271 = (inp[5]) ? 3'b011 : 3'b111;
								assign node276 = (inp[8]) ? node280 : node277;
									assign node277 = (inp[11]) ? 3'b011 : 3'b001;
									assign node280 = (inp[11]) ? node284 : node281;
										assign node281 = (inp[5]) ? 3'b110 : 3'b001;
										assign node284 = (inp[0]) ? 3'b001 : 3'b101;
						assign node287 = (inp[8]) ? node305 : node288;
							assign node288 = (inp[1]) ? node296 : node289;
								assign node289 = (inp[5]) ? 3'b001 : node290;
									assign node290 = (inp[7]) ? 3'b110 : node291;
										assign node291 = (inp[2]) ? 3'b101 : 3'b111;
								assign node296 = (inp[2]) ? node302 : node297;
									assign node297 = (inp[7]) ? node299 : 3'b101;
										assign node299 = (inp[11]) ? 3'b101 : 3'b001;
									assign node302 = (inp[0]) ? 3'b001 : 3'b011;
							assign node305 = (inp[11]) ? node309 : node306;
								assign node306 = (inp[5]) ? 3'b100 : 3'b010;
								assign node309 = (inp[0]) ? 3'b001 : node310;
									assign node310 = (inp[5]) ? 3'b110 : 3'b001;
			assign node314 = (inp[3]) ? node402 : node315;
				assign node315 = (inp[10]) ? node355 : node316;
					assign node316 = (inp[7]) ? node338 : node317;
						assign node317 = (inp[11]) ? node325 : node318;
							assign node318 = (inp[1]) ? node322 : node319;
								assign node319 = (inp[4]) ? 3'b010 : 3'b110;
								assign node322 = (inp[4]) ? 3'b110 : 3'b001;
							assign node325 = (inp[2]) ? node335 : node326;
								assign node326 = (inp[4]) ? 3'b001 : node327;
									assign node327 = (inp[0]) ? node329 : 3'b101;
										assign node329 = (inp[5]) ? node331 : 3'b101;
											assign node331 = (inp[8]) ? 3'b001 : 3'b101;
								assign node335 = (inp[5]) ? 3'b110 : 3'b101;
						assign node338 = (inp[4]) ? node348 : node339;
							assign node339 = (inp[5]) ? node345 : node340;
								assign node340 = (inp[11]) ? node342 : 3'b110;
									assign node342 = (inp[2]) ? 3'b001 : 3'b101;
								assign node345 = (inp[8]) ? 3'b010 : 3'b110;
							assign node348 = (inp[5]) ? 3'b000 : node349;
								assign node349 = (inp[0]) ? node351 : 3'b010;
									assign node351 = (inp[1]) ? 3'b010 : 3'b100;
					assign node355 = (inp[5]) ? node375 : node356;
						assign node356 = (inp[0]) ? node362 : node357;
							assign node357 = (inp[2]) ? node359 : 3'b011;
								assign node359 = (inp[11]) ? 3'b111 : 3'b011;
							assign node362 = (inp[4]) ? node366 : node363;
								assign node363 = (inp[2]) ? 3'b101 : 3'b111;
								assign node366 = (inp[8]) ? node370 : node367;
									assign node367 = (inp[11]) ? 3'b011 : 3'b101;
									assign node370 = (inp[2]) ? 3'b001 : node371;
										assign node371 = (inp[1]) ? 3'b101 : 3'b001;
						assign node375 = (inp[0]) ? node389 : node376;
							assign node376 = (inp[1]) ? node384 : node377;
								assign node377 = (inp[7]) ? node379 : 3'b011;
									assign node379 = (inp[4]) ? node381 : 3'b001;
										assign node381 = (inp[11]) ? 3'b001 : 3'b010;
								assign node384 = (inp[8]) ? 3'b001 : node385;
									assign node385 = (inp[11]) ? 3'b001 : 3'b110;
							assign node389 = (inp[4]) ? node395 : node390;
								assign node390 = (inp[11]) ? node392 : 3'b110;
									assign node392 = (inp[7]) ? 3'b001 : 3'b011;
								assign node395 = (inp[2]) ? node397 : 3'b110;
									assign node397 = (inp[8]) ? node399 : 3'b001;
										assign node399 = (inp[11]) ? 3'b010 : 3'b110;
				assign node402 = (inp[10]) ? node422 : node403;
					assign node403 = (inp[11]) ? node405 : 3'b000;
						assign node405 = (inp[4]) ? 3'b000 : node406;
							assign node406 = (inp[0]) ? node416 : node407;
								assign node407 = (inp[7]) ? 3'b100 : node408;
									assign node408 = (inp[5]) ? 3'b100 : node409;
										assign node409 = (inp[8]) ? node411 : 3'b010;
											assign node411 = (inp[1]) ? 3'b100 : 3'b010;
								assign node416 = (inp[7]) ? 3'b000 : node417;
									assign node417 = (inp[2]) ? 3'b000 : 3'b100;
					assign node422 = (inp[5]) ? node432 : node423;
						assign node423 = (inp[4]) ? node425 : 3'b001;
							assign node425 = (inp[11]) ? node427 : 3'b100;
								assign node427 = (inp[1]) ? 3'b010 : node428;
									assign node428 = (inp[8]) ? 3'b000 : 3'b100;
						assign node432 = (inp[7]) ? node444 : node433;
							assign node433 = (inp[4]) ? 3'b100 : node434;
								assign node434 = (inp[11]) ? 3'b110 : node435;
									assign node435 = (inp[8]) ? node439 : node436;
										assign node436 = (inp[0]) ? 3'b010 : 3'b110;
										assign node439 = (inp[0]) ? 3'b100 : 3'b010;
							assign node444 = (inp[8]) ? node446 : 3'b010;
								assign node446 = (inp[2]) ? node448 : 3'b000;
									assign node448 = (inp[0]) ? 3'b000 : 3'b100;

endmodule