module dtc_split5_bm47 (
	input  wire [16-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node3;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node6;
	wire [1-1:0] node8;
	wire [1-1:0] node9;
	wire [1-1:0] node10;
	wire [1-1:0] node12;
	wire [1-1:0] node15;
	wire [1-1:0] node16;
	wire [1-1:0] node20;
	wire [1-1:0] node22;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node28;
	wire [1-1:0] node29;
	wire [1-1:0] node30;
	wire [1-1:0] node32;
	wire [1-1:0] node35;
	wire [1-1:0] node36;
	wire [1-1:0] node37;
	wire [1-1:0] node41;
	wire [1-1:0] node43;
	wire [1-1:0] node47;
	wire [1-1:0] node48;
	wire [1-1:0] node49;
	wire [1-1:0] node51;
	wire [1-1:0] node54;
	wire [1-1:0] node56;
	wire [1-1:0] node59;
	wire [1-1:0] node61;
	wire [1-1:0] node64;
	wire [1-1:0] node65;
	wire [1-1:0] node67;
	wire [1-1:0] node68;
	wire [1-1:0] node69;
	wire [1-1:0] node71;
	wire [1-1:0] node74;
	wire [1-1:0] node76;
	wire [1-1:0] node79;
	wire [1-1:0] node80;
	wire [1-1:0] node85;
	wire [1-1:0] node86;
	wire [1-1:0] node87;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node91;
	wire [1-1:0] node92;
	wire [1-1:0] node93;
	wire [1-1:0] node94;
	wire [1-1:0] node95;
	wire [1-1:0] node99;
	wire [1-1:0] node101;
	wire [1-1:0] node104;
	wire [1-1:0] node106;
	wire [1-1:0] node110;
	wire [1-1:0] node111;
	wire [1-1:0] node112;
	wire [1-1:0] node113;
	wire [1-1:0] node114;
	wire [1-1:0] node118;
	wire [1-1:0] node120;
	wire [1-1:0] node124;
	wire [1-1:0] node125;
	wire [1-1:0] node126;
	wire [1-1:0] node127;
	wire [1-1:0] node131;
	wire [1-1:0] node133;
	wire [1-1:0] node136;
	wire [1-1:0] node138;
	wire [1-1:0] node141;
	wire [1-1:0] node142;
	wire [1-1:0] node144;
	wire [1-1:0] node145;
	wire [1-1:0] node146;
	wire [1-1:0] node148;
	wire [1-1:0] node151;
	wire [1-1:0] node152;
	wire [1-1:0] node156;
	wire [1-1:0] node158;
	wire [1-1:0] node162;
	wire [1-1:0] node163;
	wire [1-1:0] node164;
	wire [1-1:0] node165;
	wire [1-1:0] node167;
	wire [1-1:0] node168;
	wire [1-1:0] node169;
	wire [1-1:0] node171;
	wire [1-1:0] node174;
	wire [1-1:0] node175;
	wire [1-1:0] node176;
	wire [1-1:0] node180;
	wire [1-1:0] node184;
	wire [1-1:0] node185;
	wire [1-1:0] node186;
	wire [1-1:0] node187;
	wire [1-1:0] node188;
	wire [1-1:0] node190;
	wire [1-1:0] node191;
	wire [1-1:0] node195;
	wire [1-1:0] node198;
	wire [1-1:0] node199;
	wire [1-1:0] node200;
	wire [1-1:0] node201;
	wire [1-1:0] node204;
	wire [1-1:0] node209;
	wire [1-1:0] node210;
	wire [1-1:0] node214;
	wire [1-1:0] node216;
	wire [1-1:0] node217;
	wire [1-1:0] node218;
	wire [1-1:0] node222;
	wire [1-1:0] node224;
	wire [1-1:0] node225;
	wire [1-1:0] node228;
	wire [1-1:0] node231;
	wire [1-1:0] node232;
	wire [1-1:0] node234;
	wire [1-1:0] node235;
	wire [1-1:0] node237;
	wire [1-1:0] node240;
	wire [1-1:0] node241;
	wire [1-1:0] node243;
	wire [1-1:0] node246;
	wire [1-1:0] node248;
	wire [1-1:0] node252;
	wire [1-1:0] node253;
	wire [1-1:0] node254;
	wire [1-1:0] node256;
	wire [1-1:0] node257;
	wire [1-1:0] node258;
	wire [1-1:0] node259;
	wire [1-1:0] node263;
	wire [1-1:0] node264;
	wire [1-1:0] node265;
	wire [1-1:0] node268;
	wire [1-1:0] node273;
	wire [1-1:0] node274;
	wire [1-1:0] node275;
	wire [1-1:0] node276;
	wire [1-1:0] node279;
	wire [1-1:0] node280;
	wire [1-1:0] node284;
	wire [1-1:0] node285;
	wire [1-1:0] node287;
	wire [1-1:0] node291;
	wire [1-1:0] node292;
	wire [1-1:0] node293;
	wire [1-1:0] node294;
	wire [1-1:0] node299;
	wire [1-1:0] node300;
	wire [1-1:0] node304;
	wire [1-1:0] node306;
	wire [1-1:0] node307;
	wire [1-1:0] node308;
	wire [1-1:0] node309;
	wire [1-1:0] node313;
	wire [1-1:0] node314;
	wire [1-1:0] node316;
	wire [1-1:0] node319;
	wire [1-1:0] node321;
	wire [1-1:0] node325;
	wire [1-1:0] node326;
	wire [1-1:0] node327;
	wire [1-1:0] node328;
	wire [1-1:0] node329;
	wire [1-1:0] node330;
	wire [1-1:0] node332;
	wire [1-1:0] node333;
	wire [1-1:0] node334;
	wire [1-1:0] node338;
	wire [1-1:0] node340;
	wire [1-1:0] node344;
	wire [1-1:0] node345;
	wire [1-1:0] node346;
	wire [1-1:0] node347;
	wire [1-1:0] node350;
	wire [1-1:0] node351;
	wire [1-1:0] node355;
	wire [1-1:0] node357;
	wire [1-1:0] node360;
	wire [1-1:0] node361;
	wire [1-1:0] node363;
	wire [1-1:0] node366;
	wire [1-1:0] node368;
	wire [1-1:0] node370;
	wire [1-1:0] node373;
	wire [1-1:0] node375;
	wire [1-1:0] node376;
	wire [1-1:0] node377;
	wire [1-1:0] node378;
	wire [1-1:0] node380;
	wire [1-1:0] node383;
	wire [1-1:0] node385;
	wire [1-1:0] node388;
	wire [1-1:0] node390;
	wire [1-1:0] node394;
	wire [1-1:0] node395;
	wire [1-1:0] node396;
	wire [1-1:0] node398;
	wire [1-1:0] node399;
	wire [1-1:0] node400;
	wire [1-1:0] node402;
	wire [1-1:0] node405;
	wire [1-1:0] node406;
	wire [1-1:0] node407;
	wire [1-1:0] node411;
	wire [1-1:0] node415;
	wire [1-1:0] node416;
	wire [1-1:0] node417;
	wire [1-1:0] node418;
	wire [1-1:0] node419;
	wire [1-1:0] node420;
	wire [1-1:0] node421;
	wire [1-1:0] node428;
	wire [1-1:0] node429;
	wire [1-1:0] node431;
	wire [1-1:0] node434;
	wire [1-1:0] node435;
	wire [1-1:0] node436;
	wire [1-1:0] node440;
	wire [1-1:0] node441;
	wire [1-1:0] node445;
	wire [1-1:0] node446;
	wire [1-1:0] node448;
	wire [1-1:0] node449;
	wire [1-1:0] node451;
	wire [1-1:0] node454;
	wire [1-1:0] node455;
	wire [1-1:0] node457;
	wire [1-1:0] node460;
	wire [1-1:0] node464;
	wire [1-1:0] node465;
	wire [1-1:0] node466;
	wire [1-1:0] node468;
	wire [1-1:0] node469;
	wire [1-1:0] node470;
	wire [1-1:0] node471;
	wire [1-1:0] node472;
	wire [1-1:0] node477;
	wire [1-1:0] node478;
	wire [1-1:0] node483;
	wire [1-1:0] node484;
	wire [1-1:0] node485;
	wire [1-1:0] node486;
	wire [1-1:0] node489;
	wire [1-1:0] node493;
	wire [1-1:0] node494;
	wire [1-1:0] node496;
	wire [1-1:0] node497;
	wire [1-1:0] node501;
	wire [1-1:0] node502;
	wire [1-1:0] node506;
	wire [1-1:0] node507;
	wire [1-1:0] node509;
	wire [1-1:0] node510;
	wire [1-1:0] node511;
	wire [1-1:0] node512;
	wire [1-1:0] node517;
	wire [1-1:0] node518;
	wire [1-1:0] node523;
	wire [1-1:0] node524;
	wire [1-1:0] node525;
	wire [1-1:0] node526;
	wire [1-1:0] node527;
	wire [1-1:0] node529;
	wire [1-1:0] node530;
	wire [1-1:0] node532;
	wire [1-1:0] node533;
	wire [1-1:0] node536;
	wire [1-1:0] node537;
	wire [1-1:0] node542;
	wire [1-1:0] node543;
	wire [1-1:0] node544;
	wire [1-1:0] node545;
	wire [1-1:0] node546;
	wire [1-1:0] node552;
	wire [1-1:0] node553;
	wire [1-1:0] node555;
	wire [1-1:0] node556;
	wire [1-1:0] node560;
	wire [1-1:0] node561;
	wire [1-1:0] node562;
	wire [1-1:0] node563;
	wire [1-1:0] node568;
	wire [1-1:0] node569;
	wire [1-1:0] node573;
	wire [1-1:0] node575;
	wire [1-1:0] node576;
	wire [1-1:0] node578;
	wire [1-1:0] node579;
	wire [1-1:0] node580;
	wire [1-1:0] node584;
	wire [1-1:0] node586;
	wire [1-1:0] node590;
	wire [1-1:0] node591;
	wire [1-1:0] node592;
	wire [1-1:0] node594;
	wire [1-1:0] node595;
	wire [1-1:0] node597;
	wire [1-1:0] node598;
	wire [1-1:0] node599;
	wire [1-1:0] node602;
	wire [1-1:0] node607;
	wire [1-1:0] node608;
	wire [1-1:0] node609;
	wire [1-1:0] node611;
	wire [1-1:0] node613;
	wire [1-1:0] node616;
	wire [1-1:0] node617;
	wire [1-1:0] node618;
	wire [1-1:0] node622;
	wire [1-1:0] node625;
	wire [1-1:0] node627;
	wire [1-1:0] node628;
	wire [1-1:0] node630;
	wire [1-1:0] node633;
	wire [1-1:0] node635;
	wire [1-1:0] node636;
	wire [1-1:0] node639;
	wire [1-1:0] node642;
	wire [1-1:0] node643;
	wire [1-1:0] node645;
	wire [1-1:0] node646;
	wire [1-1:0] node647;
	wire [1-1:0] node651;
	wire [1-1:0] node655;
	wire [1-1:0] node656;
	wire [1-1:0] node657;
	wire [1-1:0] node659;
	wire [1-1:0] node660;
	wire [1-1:0] node662;
	wire [1-1:0] node666;
	wire [1-1:0] node667;
	wire [1-1:0] node668;
	wire [1-1:0] node669;
	wire [1-1:0] node673;
	wire [1-1:0] node674;
	wire [1-1:0] node675;
	wire [1-1:0] node680;
	wire [1-1:0] node682;
	wire [1-1:0] node683;
	wire [1-1:0] node684;
	wire [1-1:0] node686;
	wire [1-1:0] node689;
	wire [1-1:0] node691;
	wire [1-1:0] node694;
	wire [1-1:0] node695;
	wire [1-1:0] node699;
	wire [1-1:0] node701;
	wire [1-1:0] node702;
	wire [1-1:0] node703;
	wire [1-1:0] node705;
	wire [1-1:0] node708;
	wire [1-1:0] node710;
	wire [1-1:0] node714;
	wire [1-1:0] node715;
	wire [1-1:0] node716;
	wire [1-1:0] node718;
	wire [1-1:0] node719;
	wire [1-1:0] node720;
	wire [1-1:0] node722;
	wire [1-1:0] node725;
	wire [1-1:0] node726;
	wire [1-1:0] node730;
	wire [1-1:0] node731;
	wire [1-1:0] node736;
	wire [1-1:0] node737;
	wire [1-1:0] node738;
	wire [1-1:0] node739;
	wire [1-1:0] node741;
	wire [1-1:0] node744;
	wire [1-1:0] node745;
	wire [1-1:0] node747;
	wire [1-1:0] node750;
	wire [1-1:0] node752;
	wire [1-1:0] node755;
	wire [1-1:0] node757;
	wire [1-1:0] node758;
	wire [1-1:0] node759;
	wire [1-1:0] node760;
	wire [1-1:0] node764;
	wire [1-1:0] node765;
	wire [1-1:0] node769;
	wire [1-1:0] node770;
	wire [1-1:0] node774;
	wire [1-1:0] node776;
	wire [1-1:0] node777;
	wire [1-1:0] node778;
	wire [1-1:0] node779;
	wire [1-1:0] node780;
	wire [1-1:0] node784;
	wire [1-1:0] node786;
	wire [1-1:0] node789;
	wire [1-1:0] node791;
	wire [1-1:0] node795;
	wire [1-1:0] node796;
	wire [1-1:0] node797;
	wire [1-1:0] node798;
	wire [1-1:0] node799;
	wire [1-1:0] node800;
	wire [1-1:0] node801;
	wire [1-1:0] node802;
	wire [1-1:0] node804;
	wire [1-1:0] node805;
	wire [1-1:0] node806;
	wire [1-1:0] node810;
	wire [1-1:0] node811;
	wire [1-1:0] node813;
	wire [1-1:0] node816;
	wire [1-1:0] node817;
	wire [1-1:0] node822;
	wire [1-1:0] node823;
	wire [1-1:0] node824;
	wire [1-1:0] node825;
	wire [1-1:0] node826;
	wire [1-1:0] node828;
	wire [1-1:0] node831;
	wire [1-1:0] node835;
	wire [1-1:0] node836;
	wire [1-1:0] node837;
	wire [1-1:0] node841;
	wire [1-1:0] node842;
	wire [1-1:0] node844;
	wire [1-1:0] node847;
	wire [1-1:0] node849;
	wire [1-1:0] node852;
	wire [1-1:0] node853;
	wire [1-1:0] node855;
	wire [1-1:0] node856;
	wire [1-1:0] node857;
	wire [1-1:0] node858;
	wire [1-1:0] node860;
	wire [1-1:0] node863;
	wire [1-1:0] node865;
	wire [1-1:0] node869;
	wire [1-1:0] node871;
	wire [1-1:0] node875;
	wire [1-1:0] node876;
	wire [1-1:0] node877;
	wire [1-1:0] node879;
	wire [1-1:0] node880;
	wire [1-1:0] node881;
	wire [1-1:0] node882;
	wire [1-1:0] node886;
	wire [1-1:0] node888;
	wire [1-1:0] node891;
	wire [1-1:0] node892;
	wire [1-1:0] node897;
	wire [1-1:0] node898;
	wire [1-1:0] node899;
	wire [1-1:0] node900;
	wire [1-1:0] node901;
	wire [1-1:0] node902;
	wire [1-1:0] node906;
	wire [1-1:0] node907;
	wire [1-1:0] node909;
	wire [1-1:0] node914;
	wire [1-1:0] node915;
	wire [1-1:0] node916;
	wire [1-1:0] node918;
	wire [1-1:0] node921;
	wire [1-1:0] node922;
	wire [1-1:0] node926;
	wire [1-1:0] node928;
	wire [1-1:0] node931;
	wire [1-1:0] node933;
	wire [1-1:0] node934;
	wire [1-1:0] node935;
	wire [1-1:0] node936;
	wire [1-1:0] node937;
	wire [1-1:0] node941;
	wire [1-1:0] node946;
	wire [1-1:0] node947;
	wire [1-1:0] node949;
	wire [1-1:0] node950;
	wire [1-1:0] node951;
	wire [1-1:0] node952;
	wire [1-1:0] node956;
	wire [1-1:0] node957;
	wire [1-1:0] node959;
	wire [1-1:0] node962;
	wire [1-1:0] node964;
	wire [1-1:0] node968;
	wire [1-1:0] node969;
	wire [1-1:0] node970;
	wire [1-1:0] node971;
	wire [1-1:0] node972;
	wire [1-1:0] node973;
	wire [1-1:0] node977;
	wire [1-1:0] node978;
	wire [1-1:0] node979;
	wire [1-1:0] node980;
	wire [1-1:0] node984;
	wire [1-1:0] node985;
	wire [1-1:0] node989;
	wire [1-1:0] node990;
	wire [1-1:0] node992;
	wire [1-1:0] node997;
	wire [1-1:0] node998;
	wire [1-1:0] node999;
	wire [1-1:0] node1001;
	wire [1-1:0] node1004;
	wire [1-1:0] node1006;
	wire [1-1:0] node1009;
	wire [1-1:0] node1010;
	wire [1-1:0] node1014;
	wire [1-1:0] node1015;
	wire [1-1:0] node1017;
	wire [1-1:0] node1018;
	wire [1-1:0] node1019;
	wire [1-1:0] node1023;
	wire [1-1:0] node1024;
	wire [1-1:0] node1025;
	wire [1-1:0] node1029;
	wire [1-1:0] node1031;
	wire [1-1:0] node1035;
	wire [1-1:0] node1036;
	wire [1-1:0] node1037;
	wire [1-1:0] node1038;
	wire [1-1:0] node1039;
	wire [1-1:0] node1040;
	wire [1-1:0] node1042;
	wire [1-1:0] node1043;
	wire [1-1:0] node1044;
	wire [1-1:0] node1045;
	wire [1-1:0] node1049;
	wire [1-1:0] node1051;
	wire [1-1:0] node1054;
	wire [1-1:0] node1056;
	wire [1-1:0] node1060;
	wire [1-1:0] node1061;
	wire [1-1:0] node1062;
	wire [1-1:0] node1063;
	wire [1-1:0] node1065;
	wire [1-1:0] node1067;
	wire [1-1:0] node1068;
	wire [1-1:0] node1071;
	wire [1-1:0] node1074;
	wire [1-1:0] node1078;
	wire [1-1:0] node1079;
	wire [1-1:0] node1080;
	wire [1-1:0] node1082;
	wire [1-1:0] node1085;
	wire [1-1:0] node1088;
	wire [1-1:0] node1090;
	wire [1-1:0] node1093;
	wire [1-1:0] node1095;
	wire [1-1:0] node1096;
	wire [1-1:0] node1097;
	wire [1-1:0] node1098;
	wire [1-1:0] node1100;
	wire [1-1:0] node1103;
	wire [1-1:0] node1104;
	wire [1-1:0] node1108;
	wire [1-1:0] node1110;
	wire [1-1:0] node1114;
	wire [1-1:0] node1115;
	wire [1-1:0] node1117;
	wire [1-1:0] node1118;
	wire [1-1:0] node1119;
	wire [1-1:0] node1121;
	wire [1-1:0] node1124;
	wire [1-1:0] node1125;
	wire [1-1:0] node1126;
	wire [1-1:0] node1130;
	wire [1-1:0] node1131;
	wire [1-1:0] node1136;
	wire [1-1:0] node1137;
	wire [1-1:0] node1138;
	wire [1-1:0] node1139;
	wire [1-1:0] node1140;
	wire [1-1:0] node1141;
	wire [1-1:0] node1142;
	wire [1-1:0] node1146;
	wire [1-1:0] node1149;
	wire [1-1:0] node1150;
	wire [1-1:0] node1155;
	wire [1-1:0] node1156;
	wire [1-1:0] node1157;
	wire [1-1:0] node1161;
	wire [1-1:0] node1162;
	wire [1-1:0] node1163;
	wire [1-1:0] node1167;
	wire [1-1:0] node1168;
	wire [1-1:0] node1172;
	wire [1-1:0] node1174;
	wire [1-1:0] node1175;
	wire [1-1:0] node1176;
	wire [1-1:0] node1178;
	wire [1-1:0] node1180;
	wire [1-1:0] node1183;
	wire [1-1:0] node1185;
	wire [1-1:0] node1186;
	wire [1-1:0] node1191;
	wire [1-1:0] node1192;
	wire [1-1:0] node1193;
	wire [1-1:0] node1195;
	wire [1-1:0] node1196;
	wire [1-1:0] node1198;
	wire [1-1:0] node1201;
	wire [1-1:0] node1202;
	wire [1-1:0] node1204;
	wire [1-1:0] node1207;
	wire [1-1:0] node1208;
	wire [1-1:0] node1213;
	wire [1-1:0] node1214;
	wire [1-1:0] node1215;
	wire [1-1:0] node1216;
	wire [1-1:0] node1217;
	wire [1-1:0] node1219;
	wire [1-1:0] node1223;
	wire [1-1:0] node1224;
	wire [1-1:0] node1228;
	wire [1-1:0] node1229;
	wire [1-1:0] node1231;
	wire [1-1:0] node1232;
	wire [1-1:0] node1233;
	wire [1-1:0] node1238;
	wire [1-1:0] node1239;
	wire [1-1:0] node1241;
	wire [1-1:0] node1244;
	wire [1-1:0] node1246;
	wire [1-1:0] node1247;
	wire [1-1:0] node1251;
	wire [1-1:0] node1253;
	wire [1-1:0] node1254;
	wire [1-1:0] node1255;
	wire [1-1:0] node1256;
	wire [1-1:0] node1260;
	wire [1-1:0] node1261;
	wire [1-1:0] node1263;
	wire [1-1:0] node1266;
	wire [1-1:0] node1268;
	wire [1-1:0] node1272;
	wire [1-1:0] node1273;
	wire [1-1:0] node1274;
	wire [1-1:0] node1276;
	wire [1-1:0] node1277;
	wire [1-1:0] node1278;
	wire [1-1:0] node1280;
	wire [1-1:0] node1283;
	wire [1-1:0] node1284;
	wire [1-1:0] node1286;
	wire [1-1:0] node1289;
	wire [1-1:0] node1291;
	wire [1-1:0] node1295;
	wire [1-1:0] node1296;
	wire [1-1:0] node1297;
	wire [1-1:0] node1298;
	wire [1-1:0] node1299;
	wire [1-1:0] node1303;
	wire [1-1:0] node1304;
	wire [1-1:0] node1305;
	wire [1-1:0] node1309;
	wire [1-1:0] node1310;
	wire [1-1:0] node1314;
	wire [1-1:0] node1316;
	wire [1-1:0] node1317;
	wire [1-1:0] node1318;
	wire [1-1:0] node1320;
	wire [1-1:0] node1323;
	wire [1-1:0] node1325;
	wire [1-1:0] node1328;
	wire [1-1:0] node1329;
	wire [1-1:0] node1333;
	wire [1-1:0] node1334;
	wire [1-1:0] node1336;
	wire [1-1:0] node1337;
	wire [1-1:0] node1339;
	wire [1-1:0] node1342;
	wire [1-1:0] node1343;
	wire [1-1:0] node1345;
	wire [1-1:0] node1348;
	wire [1-1:0] node1350;
	wire [1-1:0] node1354;
	wire [1-1:0] node1355;
	wire [1-1:0] node1356;
	wire [1-1:0] node1357;
	wire [1-1:0] node1359;
	wire [1-1:0] node1360;
	wire [1-1:0] node1361;
	wire [1-1:0] node1362;
	wire [1-1:0] node1363;
	wire [1-1:0] node1367;
	wire [1-1:0] node1369;
	wire [1-1:0] node1372;
	wire [1-1:0] node1374;
	wire [1-1:0] node1378;
	wire [1-1:0] node1379;
	wire [1-1:0] node1380;
	wire [1-1:0] node1381;
	wire [1-1:0] node1383;
	wire [1-1:0] node1386;
	wire [1-1:0] node1387;
	wire [1-1:0] node1390;
	wire [1-1:0] node1394;
	wire [1-1:0] node1395;
	wire [1-1:0] node1396;
	wire [1-1:0] node1398;
	wire [1-1:0] node1401;
	wire [1-1:0] node1402;
	wire [1-1:0] node1406;
	wire [1-1:0] node1408;
	wire [1-1:0] node1411;
	wire [1-1:0] node1413;
	wire [1-1:0] node1414;
	wire [1-1:0] node1415;
	wire [1-1:0] node1416;
	wire [1-1:0] node1420;
	wire [1-1:0] node1421;
	wire [1-1:0] node1422;
	wire [1-1:0] node1426;
	wire [1-1:0] node1427;
	wire [1-1:0] node1432;
	wire [1-1:0] node1433;
	wire [1-1:0] node1434;
	wire [1-1:0] node1436;
	wire [1-1:0] node1437;
	wire [1-1:0] node1438;
	wire [1-1:0] node1440;
	wire [1-1:0] node1443;
	wire [1-1:0] node1444;
	wire [1-1:0] node1445;
	wire [1-1:0] node1449;
	wire [1-1:0] node1451;
	wire [1-1:0] node1455;
	wire [1-1:0] node1456;
	wire [1-1:0] node1457;
	wire [1-1:0] node1458;
	wire [1-1:0] node1459;
	wire [1-1:0] node1460;
	wire [1-1:0] node1463;
	wire [1-1:0] node1466;
	wire [1-1:0] node1469;
	wire [1-1:0] node1471;
	wire [1-1:0] node1475;
	wire [1-1:0] node1476;
	wire [1-1:0] node1477;
	wire [1-1:0] node1478;
	wire [1-1:0] node1482;
	wire [1-1:0] node1483;
	wire [1-1:0] node1487;
	wire [1-1:0] node1489;
	wire [1-1:0] node1492;
	wire [1-1:0] node1494;
	wire [1-1:0] node1495;
	wire [1-1:0] node1496;
	wire [1-1:0] node1497;
	wire [1-1:0] node1498;
	wire [1-1:0] node1502;
	wire [1-1:0] node1504;
	wire [1-1:0] node1507;
	wire [1-1:0] node1509;
	wire [1-1:0] node1513;
	wire [1-1:0] node1514;
	wire [1-1:0] node1515;
	wire [1-1:0] node1517;
	wire [1-1:0] node1518;
	wire [1-1:0] node1519;
	wire [1-1:0] node1520;
	wire [1-1:0] node1522;
	wire [1-1:0] node1525;
	wire [1-1:0] node1527;
	wire [1-1:0] node1530;
	wire [1-1:0] node1531;
	wire [1-1:0] node1536;
	wire [1-1:0] node1537;
	wire [1-1:0] node1538;
	wire [1-1:0] node1539;
	wire [1-1:0] node1540;
	wire [1-1:0] node1544;
	wire [1-1:0] node1545;
	wire [1-1:0] node1547;
	wire [1-1:0] node1550;
	wire [1-1:0] node1551;
	wire [1-1:0] node1555;
	wire [1-1:0] node1557;
	wire [1-1:0] node1558;
	wire [1-1:0] node1559;
	wire [1-1:0] node1560;
	wire [1-1:0] node1564;
	wire [1-1:0] node1566;
	wire [1-1:0] node1569;
	wire [1-1:0] node1571;
	wire [1-1:0] node1574;
	wire [1-1:0] node1576;
	wire [1-1:0] node1577;
	wire [1-1:0] node1578;
	wire [1-1:0] node1579;
	wire [1-1:0] node1583;
	wire [1-1:0] node1584;
	wire [1-1:0] node1586;
	wire [1-1:0] node1589;
	wire [1-1:0] node1591;
	wire [1-1:0] node1595;
	wire [1-1:0] node1596;
	wire [1-1:0] node1597;
	wire [1-1:0] node1598;
	wire [1-1:0] node1599;
	wire [1-1:0] node1601;
	wire [1-1:0] node1602;
	wire [1-1:0] node1603;
	wire [1-1:0] node1604;
	wire [1-1:0] node1607;
	wire [1-1:0] node1609;
	wire [1-1:0] node1612;
	wire [1-1:0] node1614;
	wire [1-1:0] node1618;
	wire [1-1:0] node1619;
	wire [1-1:0] node1620;
	wire [1-1:0] node1621;
	wire [1-1:0] node1622;
	wire [1-1:0] node1626;
	wire [1-1:0] node1627;
	wire [1-1:0] node1628;
	wire [1-1:0] node1632;
	wire [1-1:0] node1633;
	wire [1-1:0] node1638;
	wire [1-1:0] node1639;
	wire [1-1:0] node1640;
	wire [1-1:0] node1644;
	wire [1-1:0] node1645;
	wire [1-1:0] node1647;
	wire [1-1:0] node1650;
	wire [1-1:0] node1652;
	wire [1-1:0] node1655;
	wire [1-1:0] node1657;
	wire [1-1:0] node1658;
	wire [1-1:0] node1659;
	wire [1-1:0] node1661;
	wire [1-1:0] node1664;
	wire [1-1:0] node1665;
	wire [1-1:0] node1667;
	wire [1-1:0] node1670;
	wire [1-1:0] node1672;
	wire [1-1:0] node1676;
	wire [1-1:0] node1677;
	wire [1-1:0] node1678;
	wire [1-1:0] node1680;
	wire [1-1:0] node1681;
	wire [1-1:0] node1682;
	wire [1-1:0] node1683;
	wire [1-1:0] node1687;
	wire [1-1:0] node1689;
	wire [1-1:0] node1691;
	wire [1-1:0] node1695;
	wire [1-1:0] node1696;
	wire [1-1:0] node1697;
	wire [1-1:0] node1698;
	wire [1-1:0] node1700;
	wire [1-1:0] node1703;
	wire [1-1:0] node1704;
	wire [1-1:0] node1705;
	wire [1-1:0] node1709;
	wire [1-1:0] node1710;
	wire [1-1:0] node1714;
	wire [1-1:0] node1716;
	wire [1-1:0] node1717;
	wire [1-1:0] node1719;
	wire [1-1:0] node1722;
	wire [1-1:0] node1723;
	wire [1-1:0] node1724;
	wire [1-1:0] node1728;
	wire [1-1:0] node1730;
	wire [1-1:0] node1733;
	wire [1-1:0] node1735;
	wire [1-1:0] node1736;
	wire [1-1:0] node1737;
	wire [1-1:0] node1738;
	wire [1-1:0] node1739;
	wire [1-1:0] node1743;
	wire [1-1:0] node1745;
	wire [1-1:0] node1750;
	wire [1-1:0] node1751;
	wire [1-1:0] node1752;
	wire [1-1:0] node1754;
	wire [1-1:0] node1755;
	wire [1-1:0] node1757;
	wire [1-1:0] node1760;
	wire [1-1:0] node1761;
	wire [1-1:0] node1763;
	wire [1-1:0] node1766;
	wire [1-1:0] node1767;
	wire [1-1:0] node1772;
	wire [1-1:0] node1773;
	wire [1-1:0] node1774;
	wire [1-1:0] node1775;
	wire [1-1:0] node1776;
	wire [1-1:0] node1777;
	wire [1-1:0] node1781;
	wire [1-1:0] node1783;
	wire [1-1:0] node1786;
	wire [1-1:0] node1788;
	wire [1-1:0] node1789;
	wire [1-1:0] node1791;
	wire [1-1:0] node1795;
	wire [1-1:0] node1796;
	wire [1-1:0] node1799;
	wire [1-1:0] node1800;
	wire [1-1:0] node1804;
	wire [1-1:0] node1806;
	wire [1-1:0] node1807;
	wire [1-1:0] node1808;
	wire [1-1:0] node1809;
	wire [1-1:0] node1810;
	wire [1-1:0] node1815;
	wire [1-1:0] node1817;
	wire [1-1:0] node1821;
	wire [1-1:0] node1822;
	wire [1-1:0] node1823;
	wire [1-1:0] node1824;
	wire [1-1:0] node1825;
	wire [1-1:0] node1826;
	wire [1-1:0] node1828;
	wire [1-1:0] node1829;
	wire [1-1:0] node1830;
	wire [1-1:0] node1834;
	wire [1-1:0] node1835;
	wire [1-1:0] node1840;
	wire [1-1:0] node1841;
	wire [1-1:0] node1842;
	wire [1-1:0] node1843;
	wire [1-1:0] node1844;
	wire [1-1:0] node1846;
	wire [1-1:0] node1849;
	wire [1-1:0] node1851;
	wire [1-1:0] node1854;
	wire [1-1:0] node1855;
	wire [1-1:0] node1860;
	wire [1-1:0] node1861;
	wire [1-1:0] node1862;
	wire [1-1:0] node1866;
	wire [1-1:0] node1867;
	wire [1-1:0] node1869;
	wire [1-1:0] node1872;
	wire [1-1:0] node1874;
	wire [1-1:0] node1877;
	wire [1-1:0] node1878;
	wire [1-1:0] node1880;
	wire [1-1:0] node1881;
	wire [1-1:0] node1883;
	wire [1-1:0] node1886;
	wire [1-1:0] node1888;
	wire [1-1:0] node1890;
	wire [1-1:0] node1891;
	wire [1-1:0] node1894;
	wire [1-1:0] node1898;
	wire [1-1:0] node1899;
	wire [1-1:0] node1900;
	wire [1-1:0] node1901;
	wire [1-1:0] node1902;
	wire [1-1:0] node1904;
	wire [1-1:0] node1905;
	wire [1-1:0] node1908;
	wire [1-1:0] node1909;
	wire [1-1:0] node1914;
	wire [1-1:0] node1915;
	wire [1-1:0] node1916;
	wire [1-1:0] node1918;
	wire [1-1:0] node1919;
	wire [1-1:0] node1922;
	wire [1-1:0] node1923;
	wire [1-1:0] node1927;
	wire [1-1:0] node1928;
	wire [1-1:0] node1930;
	wire [1-1:0] node1932;
	wire [1-1:0] node1935;
	wire [1-1:0] node1938;
	wire [1-1:0] node1940;
	wire [1-1:0] node1941;
	wire [1-1:0] node1942;
	wire [1-1:0] node1947;
	wire [1-1:0] node1948;
	wire [1-1:0] node1950;
	wire [1-1:0] node1952;
	wire [1-1:0] node1953;
	wire [1-1:0] node1958;
	wire [1-1:0] node1959;
	wire [1-1:0] node1960;
	wire [1-1:0] node1961;
	wire [1-1:0] node1963;
	wire [1-1:0] node1964;
	wire [1-1:0] node1965;
	wire [1-1:0] node1969;
	wire [1-1:0] node1970;
	wire [1-1:0] node1975;
	wire [1-1:0] node1976;
	wire [1-1:0] node1977;
	wire [1-1:0] node1979;
	wire [1-1:0] node1981;
	wire [1-1:0] node1985;
	wire [1-1:0] node1986;
	wire [1-1:0] node1988;
	wire [1-1:0] node1989;
	wire [1-1:0] node1994;
	wire [1-1:0] node1996;
	wire [1-1:0] node1997;
	wire [1-1:0] node1999;
	wire [1-1:0] node2003;
	wire [1-1:0] node2004;
	wire [1-1:0] node2005;
	wire [1-1:0] node2006;
	wire [1-1:0] node2007;
	wire [1-1:0] node2008;
	wire [1-1:0] node2010;
	wire [1-1:0] node2011;
	wire [1-1:0] node2012;
	wire [1-1:0] node2017;
	wire [1-1:0] node2018;
	wire [1-1:0] node2019;
	wire [1-1:0] node2021;
	wire [1-1:0] node2024;
	wire [1-1:0] node2027;
	wire [1-1:0] node2028;
	wire [1-1:0] node2032;
	wire [1-1:0] node2033;
	wire [1-1:0] node2034;
	wire [1-1:0] node2035;
	wire [1-1:0] node2037;
	wire [1-1:0] node2040;
	wire [1-1:0] node2042;
	wire [1-1:0] node2043;
	wire [1-1:0] node2046;
	wire [1-1:0] node2050;
	wire [1-1:0] node2051;
	wire [1-1:0] node2053;
	wire [1-1:0] node2057;
	wire [1-1:0] node2059;
	wire [1-1:0] node2060;
	wire [1-1:0] node2061;
	wire [1-1:0] node2063;
	wire [1-1:0] node2066;
	wire [1-1:0] node2067;
	wire [1-1:0] node2070;
	wire [1-1:0] node2074;
	wire [1-1:0] node2075;
	wire [1-1:0] node2076;
	wire [1-1:0] node2077;
	wire [1-1:0] node2079;
	wire [1-1:0] node2080;
	wire [1-1:0] node2082;
	wire [1-1:0] node2086;
	wire [1-1:0] node2087;
	wire [1-1:0] node2088;
	wire [1-1:0] node2090;
	wire [1-1:0] node2094;
	wire [1-1:0] node2095;
	wire [1-1:0] node2099;
	wire [1-1:0] node2101;
	wire [1-1:0] node2102;
	wire [1-1:0] node2104;
	wire [1-1:0] node2105;
	wire [1-1:0] node2109;
	wire [1-1:0] node2111;
	wire [1-1:0] node2113;
	wire [1-1:0] node2116;
	wire [1-1:0] node2118;
	wire [1-1:0] node2119;
	wire [1-1:0] node2120;
	wire [1-1:0] node2121;
	wire [1-1:0] node2125;
	wire [1-1:0] node2126;
	wire [1-1:0] node2127;
	wire [1-1:0] node2130;
	wire [1-1:0] node2135;
	wire [1-1:0] node2136;
	wire [1-1:0] node2137;
	wire [1-1:0] node2139;
	wire [1-1:0] node2140;
	wire [1-1:0] node2141;
	wire [1-1:0] node2144;
	wire [1-1:0] node2145;
	wire [1-1:0] node2148;
	wire [1-1:0] node2151;
	wire [1-1:0] node2152;
	wire [1-1:0] node2157;
	wire [1-1:0] node2158;
	wire [1-1:0] node2159;
	wire [1-1:0] node2160;
	wire [1-1:0] node2161;
	wire [1-1:0] node2162;
	wire [1-1:0] node2163;
	wire [1-1:0] node2167;
	wire [1-1:0] node2168;
	wire [1-1:0] node2172;
	wire [1-1:0] node2174;
	wire [1-1:0] node2178;
	wire [1-1:0] node2179;
	wire [1-1:0] node2181;
	wire [1-1:0] node2184;
	wire [1-1:0] node2185;
	wire [1-1:0] node2188;
	wire [1-1:0] node2189;
	wire [1-1:0] node2193;
	wire [1-1:0] node2195;
	wire [1-1:0] node2196;
	wire [1-1:0] node2197;
	wire [1-1:0] node2198;
	wire [1-1:0] node2200;
	wire [1-1:0] node2201;
	wire [1-1:0] node2204;
	wire [1-1:0] node2208;
	wire [1-1:0] node2210;
	wire [1-1:0] node2214;
	wire [1-1:0] node2215;
	wire [1-1:0] node2216;
	wire [1-1:0] node2217;
	wire [1-1:0] node2219;
	wire [1-1:0] node2220;
	wire [1-1:0] node2221;
	wire [1-1:0] node2225;
	wire [1-1:0] node2226;
	wire [1-1:0] node2228;
	wire [1-1:0] node2231;
	wire [1-1:0] node2233;
	wire [1-1:0] node2237;
	wire [1-1:0] node2238;
	wire [1-1:0] node2239;
	wire [1-1:0] node2240;
	wire [1-1:0] node2241;
	wire [1-1:0] node2243;
	wire [1-1:0] node2246;
	wire [1-1:0] node2248;
	wire [1-1:0] node2251;
	wire [1-1:0] node2252;
	wire [1-1:0] node2256;
	wire [1-1:0] node2258;
	wire [1-1:0] node2259;
	wire [1-1:0] node2260;
	wire [1-1:0] node2261;
	wire [1-1:0] node2265;
	wire [1-1:0] node2266;
	wire [1-1:0] node2270;
	wire [1-1:0] node2272;
	wire [1-1:0] node2275;
	wire [1-1:0] node2276;
	wire [1-1:0] node2278;
	wire [1-1:0] node2279;
	wire [1-1:0] node2280;
	wire [1-1:0] node2282;
	wire [1-1:0] node2285;
	wire [1-1:0] node2287;
	wire [1-1:0] node2290;
	wire [1-1:0] node2291;
	wire [1-1:0] node2296;
	wire [1-1:0] node2297;
	wire [1-1:0] node2298;
	wire [1-1:0] node2299;
	wire [1-1:0] node2300;
	wire [1-1:0] node2301;
	wire [1-1:0] node2302;
	wire [1-1:0] node2303;
	wire [1-1:0] node2304;
	wire [1-1:0] node2306;
	wire [1-1:0] node2307;
	wire [1-1:0] node2309;
	wire [1-1:0] node2312;
	wire [1-1:0] node2314;
	wire [1-1:0] node2316;
	wire [1-1:0] node2320;
	wire [1-1:0] node2321;
	wire [1-1:0] node2322;
	wire [1-1:0] node2323;
	wire [1-1:0] node2326;
	wire [1-1:0] node2327;
	wire [1-1:0] node2331;
	wire [1-1:0] node2332;
	wire [1-1:0] node2336;
	wire [1-1:0] node2338;
	wire [1-1:0] node2340;
	wire [1-1:0] node2341;
	wire [1-1:0] node2342;
	wire [1-1:0] node2346;
	wire [1-1:0] node2347;
	wire [1-1:0] node2351;
	wire [1-1:0] node2353;
	wire [1-1:0] node2354;
	wire [1-1:0] node2355;
	wire [1-1:0] node2356;
	wire [1-1:0] node2360;
	wire [1-1:0] node2361;
	wire [1-1:0] node2362;
	wire [1-1:0] node2366;
	wire [1-1:0] node2368;
	wire [1-1:0] node2372;
	wire [1-1:0] node2373;
	wire [1-1:0] node2374;
	wire [1-1:0] node2376;
	wire [1-1:0] node2377;
	wire [1-1:0] node2378;
	wire [1-1:0] node2380;
	wire [1-1:0] node2384;
	wire [1-1:0] node2386;
	wire [1-1:0] node2390;
	wire [1-1:0] node2391;
	wire [1-1:0] node2392;
	wire [1-1:0] node2393;
	wire [1-1:0] node2396;
	wire [1-1:0] node2397;
	wire [1-1:0] node2399;
	wire [1-1:0] node2403;
	wire [1-1:0] node2404;
	wire [1-1:0] node2405;
	wire [1-1:0] node2409;
	wire [1-1:0] node2411;
	wire [1-1:0] node2412;
	wire [1-1:0] node2416;
	wire [1-1:0] node2417;
	wire [1-1:0] node2419;
	wire [1-1:0] node2420;
	wire [1-1:0] node2421;
	wire [1-1:0] node2422;
	wire [1-1:0] node2426;
	wire [1-1:0] node2429;
	wire [1-1:0] node2430;
	wire [1-1:0] node2435;
	wire [1-1:0] node2436;
	wire [1-1:0] node2437;
	wire [1-1:0] node2439;
	wire [1-1:0] node2440;
	wire [1-1:0] node2441;
	wire [1-1:0] node2442;
	wire [1-1:0] node2444;
	wire [1-1:0] node2447;
	wire [1-1:0] node2449;
	wire [1-1:0] node2452;
	wire [1-1:0] node2453;
	wire [1-1:0] node2458;
	wire [1-1:0] node2459;
	wire [1-1:0] node2460;
	wire [1-1:0] node2461;
	wire [1-1:0] node2463;
	wire [1-1:0] node2466;
	wire [1-1:0] node2467;
	wire [1-1:0] node2469;
	wire [1-1:0] node2472;
	wire [1-1:0] node2474;
	wire [1-1:0] node2478;
	wire [1-1:0] node2479;
	wire [1-1:0] node2480;
	wire [1-1:0] node2484;
	wire [1-1:0] node2485;
	wire [1-1:0] node2486;
	wire [1-1:0] node2490;
	wire [1-1:0] node2491;
	wire [1-1:0] node2495;
	wire [1-1:0] node2496;
	wire [1-1:0] node2498;
	wire [1-1:0] node2499;
	wire [1-1:0] node2500;
	wire [1-1:0] node2504;
	wire [1-1:0] node2505;
	wire [1-1:0] node2506;
	wire [1-1:0] node2510;
	wire [1-1:0] node2511;
	wire [1-1:0] node2516;
	wire [1-1:0] node2517;
	wire [1-1:0] node2518;
	wire [1-1:0] node2519;
	wire [1-1:0] node2521;
	wire [1-1:0] node2522;
	wire [1-1:0] node2523;
	wire [1-1:0] node2524;
	wire [1-1:0] node2525;
	wire [1-1:0] node2530;
	wire [1-1:0] node2531;
	wire [1-1:0] node2536;
	wire [1-1:0] node2537;
	wire [1-1:0] node2538;
	wire [1-1:0] node2539;
	wire [1-1:0] node2540;
	wire [1-1:0] node2544;
	wire [1-1:0] node2545;
	wire [1-1:0] node2547;
	wire [1-1:0] node2550;
	wire [1-1:0] node2551;
	wire [1-1:0] node2555;
	wire [1-1:0] node2557;
	wire [1-1:0] node2558;
	wire [1-1:0] node2560;
	wire [1-1:0] node2563;
	wire [1-1:0] node2564;
	wire [1-1:0] node2567;
	wire [1-1:0] node2569;
	wire [1-1:0] node2572;
	wire [1-1:0] node2574;
	wire [1-1:0] node2575;
	wire [1-1:0] node2576;
	wire [1-1:0] node2579;
	wire [1-1:0] node2581;
	wire [1-1:0] node2582;
	wire [1-1:0] node2587;
	wire [1-1:0] node2588;
	wire [1-1:0] node2589;
	wire [1-1:0] node2591;
	wire [1-1:0] node2592;
	wire [1-1:0] node2594;
	wire [1-1:0] node2597;
	wire [1-1:0] node2598;
	wire [1-1:0] node2600;
	wire [1-1:0] node2603;
	wire [1-1:0] node2604;
	wire [1-1:0] node2609;
	wire [1-1:0] node2610;
	wire [1-1:0] node2611;
	wire [1-1:0] node2612;
	wire [1-1:0] node2613;
	wire [1-1:0] node2614;
	wire [1-1:0] node2618;
	wire [1-1:0] node2620;
	wire [1-1:0] node2624;
	wire [1-1:0] node2625;
	wire [1-1:0] node2626;
	wire [1-1:0] node2629;
	wire [1-1:0] node2631;
	wire [1-1:0] node2634;
	wire [1-1:0] node2635;
	wire [1-1:0] node2639;
	wire [1-1:0] node2641;
	wire [1-1:0] node2642;
	wire [1-1:0] node2643;
	wire [1-1:0] node2644;
	wire [1-1:0] node2648;
	wire [1-1:0] node2649;
	wire [1-1:0] node2650;
	wire [1-1:0] node2653;
	wire [1-1:0] node2656;
	wire [1-1:0] node2660;
	wire [1-1:0] node2661;
	wire [1-1:0] node2662;
	wire [1-1:0] node2664;
	wire [1-1:0] node2665;
	wire [1-1:0] node2666;
	wire [1-1:0] node2667;
	wire [1-1:0] node2671;
	wire [1-1:0] node2672;
	wire [1-1:0] node2674;
	wire [1-1:0] node2677;
	wire [1-1:0] node2679;
	wire [1-1:0] node2683;
	wire [1-1:0] node2684;
	wire [1-1:0] node2685;
	wire [1-1:0] node2686;
	wire [1-1:0] node2688;
	wire [1-1:0] node2691;
	wire [1-1:0] node2692;
	wire [1-1:0] node2694;
	wire [1-1:0] node2699;
	wire [1-1:0] node2700;
	wire [1-1:0] node2701;
	wire [1-1:0] node2703;
	wire [1-1:0] node2706;
	wire [1-1:0] node2708;
	wire [1-1:0] node2711;
	wire [1-1:0] node2713;
	wire [1-1:0] node2716;
	wire [1-1:0] node2717;
	wire [1-1:0] node2719;
	wire [1-1:0] node2720;
	wire [1-1:0] node2721;
	wire [1-1:0] node2722;
	wire [1-1:0] node2726;
	wire [1-1:0] node2728;
	wire [1-1:0] node2731;
	wire [1-1:0] node2732;
	wire [1-1:0] node2737;
	wire [1-1:0] node2738;
	wire [1-1:0] node2739;
	wire [1-1:0] node2740;
	wire [1-1:0] node2741;
	wire [1-1:0] node2743;
	wire [1-1:0] node2744;
	wire [1-1:0] node2745;
	wire [1-1:0] node2749;
	wire [1-1:0] node2750;
	wire [1-1:0] node2751;
	wire [1-1:0] node2755;
	wire [1-1:0] node2757;
	wire [1-1:0] node2761;
	wire [1-1:0] node2762;
	wire [1-1:0] node2763;
	wire [1-1:0] node2764;
	wire [1-1:0] node2765;
	wire [1-1:0] node2766;
	wire [1-1:0] node2770;
	wire [1-1:0] node2772;
	wire [1-1:0] node2774;
	wire [1-1:0] node2777;
	wire [1-1:0] node2778;
	wire [1-1:0] node2780;
	wire [1-1:0] node2784;
	wire [1-1:0] node2785;
	wire [1-1:0] node2786;
	wire [1-1:0] node2790;
	wire [1-1:0] node2792;
	wire [1-1:0] node2794;
	wire [1-1:0] node2797;
	wire [1-1:0] node2799;
	wire [1-1:0] node2800;
	wire [1-1:0] node2801;
	wire [1-1:0] node2803;
	wire [1-1:0] node2806;
	wire [1-1:0] node2807;
	wire [1-1:0] node2808;
	wire [1-1:0] node2812;
	wire [1-1:0] node2814;
	wire [1-1:0] node2815;
	wire [1-1:0] node2820;
	wire [1-1:0] node2821;
	wire [1-1:0] node2822;
	wire [1-1:0] node2823;
	wire [1-1:0] node2825;
	wire [1-1:0] node2826;
	wire [1-1:0] node2828;
	wire [1-1:0] node2831;
	wire [1-1:0] node2832;
	wire [1-1:0] node2834;
	wire [1-1:0] node2837;
	wire [1-1:0] node2838;
	wire [1-1:0] node2843;
	wire [1-1:0] node2844;
	wire [1-1:0] node2845;
	wire [1-1:0] node2846;
	wire [1-1:0] node2847;
	wire [1-1:0] node2848;
	wire [1-1:0] node2852;
	wire [1-1:0] node2854;
	wire [1-1:0] node2857;
	wire [1-1:0] node2859;
	wire [1-1:0] node2863;
	wire [1-1:0] node2864;
	wire [1-1:0] node2865;
	wire [1-1:0] node2869;
	wire [1-1:0] node2870;
	wire [1-1:0] node2872;
	wire [1-1:0] node2875;
	wire [1-1:0] node2876;
	wire [1-1:0] node2880;
	wire [1-1:0] node2882;
	wire [1-1:0] node2883;
	wire [1-1:0] node2884;
	wire [1-1:0] node2885;
	wire [1-1:0] node2887;
	wire [1-1:0] node2890;
	wire [1-1:0] node2891;
	wire [1-1:0] node2895;
	wire [1-1:0] node2897;
	wire [1-1:0] node2901;
	wire [1-1:0] node2902;
	wire [1-1:0] node2903;
	wire [1-1:0] node2904;
	wire [1-1:0] node2906;
	wire [1-1:0] node2907;
	wire [1-1:0] node2908;
	wire [1-1:0] node2910;
	wire [1-1:0] node2913;
	wire [1-1:0] node2914;
	wire [1-1:0] node2918;
	wire [1-1:0] node2920;
	wire [1-1:0] node2924;
	wire [1-1:0] node2925;
	wire [1-1:0] node2926;
	wire [1-1:0] node2927;
	wire [1-1:0] node2928;
	wire [1-1:0] node2929;
	wire [1-1:0] node2933;
	wire [1-1:0] node2934;
	wire [1-1:0] node2938;
	wire [1-1:0] node2940;
	wire [1-1:0] node2944;
	wire [1-1:0] node2945;
	wire [1-1:0] node2946;
	wire [1-1:0] node2948;
	wire [1-1:0] node2951;
	wire [1-1:0] node2952;
	wire [1-1:0] node2956;
	wire [1-1:0] node2957;
	wire [1-1:0] node2961;
	wire [1-1:0] node2963;
	wire [1-1:0] node2964;
	wire [1-1:0] node2965;
	wire [1-1:0] node2966;
	wire [1-1:0] node2967;
	wire [1-1:0] node2971;
	wire [1-1:0] node2972;
	wire [1-1:0] node2976;
	wire [1-1:0] node2977;
	wire [1-1:0] node2982;
	wire [1-1:0] node2983;
	wire [1-1:0] node2985;
	wire [1-1:0] node2986;
	wire [1-1:0] node2987;
	wire [1-1:0] node2989;
	wire [1-1:0] node2992;
	wire [1-1:0] node2993;
	wire [1-1:0] node2995;
	wire [1-1:0] node2998;
	wire [1-1:0] node3000;
	wire [1-1:0] node3004;
	wire [1-1:0] node3005;
	wire [1-1:0] node3006;
	wire [1-1:0] node3007;
	wire [1-1:0] node3008;
	wire [1-1:0] node3010;
	wire [1-1:0] node3013;
	wire [1-1:0] node3015;
	wire [1-1:0] node3018;
	wire [1-1:0] node3020;
	wire [1-1:0] node3023;
	wire [1-1:0] node3025;
	wire [1-1:0] node3026;
	wire [1-1:0] node3027;
	wire [1-1:0] node3028;
	wire [1-1:0] node3032;
	wire [1-1:0] node3033;
	wire [1-1:0] node3037;
	wire [1-1:0] node3039;
	wire [1-1:0] node3042;
	wire [1-1:0] node3044;
	wire [1-1:0] node3045;
	wire [1-1:0] node3046;
	wire [1-1:0] node3048;
	wire [1-1:0] node3051;
	wire [1-1:0] node3052;
	wire [1-1:0] node3054;
	wire [1-1:0] node3057;
	wire [1-1:0] node3059;

	assign outp = (inp[4]) ? node2214 : node1;
		assign node1 = (inp[0]) ? node795 : node2;
			assign node2 = (inp[8]) ? node714 : node3;
				assign node3 = (inp[1]) ? node85 : node4;
					assign node4 = (inp[6]) ? node26 : node5;
						assign node5 = (inp[15]) ? 1'b1 : node6;
							assign node6 = (inp[12]) ? node8 : 1'b1;
								assign node8 = (inp[7]) ? node20 : node9;
									assign node9 = (inp[3]) ? node15 : node10;
										assign node10 = (inp[9]) ? node12 : 1'b0;
											assign node12 = (inp[10]) ? 1'b0 : 1'b1;
										assign node15 = (inp[10]) ? 1'b1 : node16;
											assign node16 = (inp[9]) ? 1'b0 : 1'b1;
									assign node20 = (inp[9]) ? node22 : 1'b0;
										assign node22 = (inp[10]) ? 1'b0 : 1'b1;
						assign node26 = (inp[5]) ? node64 : node27;
							assign node27 = (inp[15]) ? node47 : node28;
								assign node28 = (inp[12]) ? 1'b1 : node29;
									assign node29 = (inp[3]) ? node35 : node30;
										assign node30 = (inp[9]) ? node32 : 1'b0;
											assign node32 = (inp[10]) ? 1'b0 : 1'b1;
										assign node35 = (inp[7]) ? node41 : node36;
											assign node36 = (inp[10]) ? 1'b1 : node37;
												assign node37 = (inp[9]) ? 1'b0 : 1'b1;
											assign node41 = (inp[9]) ? node43 : 1'b0;
												assign node43 = (inp[10]) ? 1'b0 : 1'b1;
								assign node47 = (inp[10]) ? node59 : node48;
									assign node48 = (inp[9]) ? node54 : node49;
										assign node49 = (inp[3]) ? node51 : 1'b0;
											assign node51 = (inp[7]) ? 1'b0 : 1'b1;
										assign node54 = (inp[3]) ? node56 : 1'b1;
											assign node56 = (inp[7]) ? 1'b1 : 1'b0;
									assign node59 = (inp[3]) ? node61 : 1'b0;
										assign node61 = (inp[7]) ? 1'b0 : 1'b1;
							assign node64 = (inp[15]) ? 1'b1 : node65;
								assign node65 = (inp[12]) ? node67 : 1'b1;
									assign node67 = (inp[7]) ? node79 : node68;
										assign node68 = (inp[3]) ? node74 : node69;
											assign node69 = (inp[9]) ? node71 : 1'b0;
												assign node71 = (inp[10]) ? 1'b0 : 1'b1;
											assign node74 = (inp[9]) ? node76 : 1'b1;
												assign node76 = (inp[10]) ? 1'b1 : 1'b0;
										assign node79 = (inp[10]) ? 1'b0 : node80;
											assign node80 = (inp[9]) ? 1'b1 : 1'b0;
					assign node85 = (inp[14]) ? node325 : node86;
						assign node86 = (inp[13]) ? node162 : node87;
							assign node87 = (inp[15]) ? node141 : node88;
								assign node88 = (inp[12]) ? node110 : node89;
									assign node89 = (inp[6]) ? node91 : 1'b0;
										assign node91 = (inp[5]) ? 1'b0 : node92;
											assign node92 = (inp[10]) ? node104 : node93;
												assign node93 = (inp[9]) ? node99 : node94;
													assign node94 = (inp[2]) ? 1'b1 : node95;
														assign node95 = (inp[7]) ? 1'b1 : 1'b0;
													assign node99 = (inp[3]) ? node101 : 1'b0;
														assign node101 = (inp[7]) ? 1'b0 : 1'b1;
												assign node104 = (inp[3]) ? node106 : 1'b1;
													assign node106 = (inp[7]) ? 1'b1 : 1'b0;
									assign node110 = (inp[5]) ? node124 : node111;
										assign node111 = (inp[6]) ? 1'b0 : node112;
											assign node112 = (inp[10]) ? node118 : node113;
												assign node113 = (inp[9]) ? 1'b0 : node114;
													assign node114 = (inp[3]) ? 1'b0 : 1'b1;
												assign node118 = (inp[3]) ? node120 : 1'b1;
													assign node120 = (inp[7]) ? 1'b1 : 1'b0;
										assign node124 = (inp[7]) ? node136 : node125;
											assign node125 = (inp[3]) ? node131 : node126;
												assign node126 = (inp[10]) ? 1'b1 : node127;
													assign node127 = (inp[9]) ? 1'b0 : 1'b1;
												assign node131 = (inp[9]) ? node133 : 1'b0;
													assign node133 = (inp[10]) ? 1'b0 : 1'b1;
											assign node136 = (inp[9]) ? node138 : 1'b1;
												assign node138 = (inp[10]) ? 1'b1 : 1'b0;
								assign node141 = (inp[5]) ? 1'b0 : node142;
									assign node142 = (inp[6]) ? node144 : 1'b0;
										assign node144 = (inp[7]) ? node156 : node145;
											assign node145 = (inp[3]) ? node151 : node146;
												assign node146 = (inp[9]) ? node148 : 1'b1;
													assign node148 = (inp[10]) ? 1'b1 : 1'b0;
												assign node151 = (inp[10]) ? 1'b0 : node152;
													assign node152 = (inp[9]) ? 1'b1 : 1'b0;
											assign node156 = (inp[9]) ? node158 : 1'b1;
												assign node158 = (inp[10]) ? 1'b1 : 1'b0;
							assign node162 = (inp[11]) ? node252 : node163;
								assign node163 = (inp[5]) ? node231 : node164;
									assign node164 = (inp[6]) ? node184 : node165;
										assign node165 = (inp[12]) ? node167 : 1'b1;
											assign node167 = (inp[15]) ? 1'b1 : node168;
												assign node168 = (inp[9]) ? node174 : node169;
													assign node169 = (inp[3]) ? node171 : 1'b0;
														assign node171 = (inp[7]) ? 1'b0 : 1'b1;
													assign node174 = (inp[10]) ? node180 : node175;
														assign node175 = (inp[7]) ? 1'b1 : node176;
															assign node176 = (inp[3]) ? 1'b0 : 1'b1;
														assign node180 = (inp[7]) ? 1'b0 : 1'b1;
										assign node184 = (inp[12]) ? node214 : node185;
											assign node185 = (inp[10]) ? node209 : node186;
												assign node186 = (inp[2]) ? node198 : node187;
													assign node187 = (inp[9]) ? node195 : node188;
														assign node188 = (inp[15]) ? node190 : 1'b1;
															assign node190 = (inp[7]) ? 1'b0 : node191;
																assign node191 = (inp[3]) ? 1'b1 : 1'b0;
														assign node195 = (inp[7]) ? 1'b1 : 1'b0;
													assign node198 = (inp[15]) ? 1'b1 : node199;
														assign node199 = (inp[7]) ? 1'b1 : node200;
															assign node200 = (inp[9]) ? node204 : node201;
																assign node201 = (inp[3]) ? 1'b1 : 1'b0;
																assign node204 = (inp[3]) ? 1'b0 : 1'b1;
												assign node209 = (inp[7]) ? 1'b0 : node210;
													assign node210 = (inp[3]) ? 1'b1 : 1'b0;
											assign node214 = (inp[15]) ? node216 : 1'b1;
												assign node216 = (inp[3]) ? node222 : node217;
													assign node217 = (inp[10]) ? 1'b0 : node218;
														assign node218 = (inp[9]) ? 1'b1 : 1'b0;
													assign node222 = (inp[9]) ? node224 : 1'b1;
														assign node224 = (inp[7]) ? node228 : node225;
															assign node225 = (inp[10]) ? 1'b1 : 1'b0;
															assign node228 = (inp[10]) ? 1'b0 : 1'b1;
									assign node231 = (inp[15]) ? 1'b1 : node232;
										assign node232 = (inp[12]) ? node234 : 1'b1;
											assign node234 = (inp[9]) ? node240 : node235;
												assign node235 = (inp[3]) ? node237 : 1'b0;
													assign node237 = (inp[7]) ? 1'b0 : 1'b1;
												assign node240 = (inp[10]) ? node246 : node241;
													assign node241 = (inp[3]) ? node243 : 1'b1;
														assign node243 = (inp[7]) ? 1'b1 : 1'b0;
													assign node246 = (inp[3]) ? node248 : 1'b0;
														assign node248 = (inp[7]) ? 1'b0 : 1'b1;
								assign node252 = (inp[15]) ? node304 : node253;
									assign node253 = (inp[12]) ? node273 : node254;
										assign node254 = (inp[6]) ? node256 : 1'b0;
											assign node256 = (inp[5]) ? 1'b0 : node257;
												assign node257 = (inp[3]) ? node263 : node258;
													assign node258 = (inp[10]) ? 1'b1 : node259;
														assign node259 = (inp[9]) ? 1'b0 : 1'b1;
													assign node263 = (inp[10]) ? 1'b0 : node264;
														assign node264 = (inp[9]) ? node268 : node265;
															assign node265 = (inp[7]) ? 1'b1 : 1'b0;
															assign node268 = (inp[7]) ? 1'b0 : 1'b1;
										assign node273 = (inp[7]) ? node291 : node274;
											assign node274 = (inp[3]) ? node284 : node275;
												assign node275 = (inp[10]) ? node279 : node276;
													assign node276 = (inp[9]) ? 1'b0 : 1'b1;
													assign node279 = (inp[5]) ? 1'b1 : node280;
														assign node280 = (inp[6]) ? 1'b0 : 1'b1;
												assign node284 = (inp[10]) ? 1'b0 : node285;
													assign node285 = (inp[9]) ? node287 : 1'b0;
														assign node287 = (inp[6]) ? 1'b0 : 1'b1;
											assign node291 = (inp[5]) ? node299 : node292;
												assign node292 = (inp[6]) ? 1'b0 : node293;
													assign node293 = (inp[10]) ? 1'b1 : node294;
														assign node294 = (inp[9]) ? 1'b0 : 1'b1;
												assign node299 = (inp[10]) ? 1'b1 : node300;
													assign node300 = (inp[9]) ? 1'b0 : 1'b1;
									assign node304 = (inp[6]) ? node306 : 1'b0;
										assign node306 = (inp[5]) ? 1'b0 : node307;
											assign node307 = (inp[9]) ? node313 : node308;
												assign node308 = (inp[7]) ? 1'b1 : node309;
													assign node309 = (inp[3]) ? 1'b0 : 1'b1;
												assign node313 = (inp[10]) ? node319 : node314;
													assign node314 = (inp[3]) ? node316 : 1'b0;
														assign node316 = (inp[7]) ? 1'b0 : 1'b1;
													assign node319 = (inp[3]) ? node321 : 1'b1;
														assign node321 = (inp[7]) ? 1'b1 : 1'b0;
						assign node325 = (inp[2]) ? node523 : node326;
							assign node326 = (inp[13]) ? node394 : node327;
								assign node327 = (inp[5]) ? node373 : node328;
									assign node328 = (inp[6]) ? node344 : node329;
										assign node329 = (inp[15]) ? 1'b1 : node330;
											assign node330 = (inp[12]) ? node332 : 1'b1;
												assign node332 = (inp[7]) ? node338 : node333;
													assign node333 = (inp[3]) ? 1'b1 : node334;
														assign node334 = (inp[9]) ? 1'b1 : 1'b0;
													assign node338 = (inp[9]) ? node340 : 1'b0;
														assign node340 = (inp[10]) ? 1'b0 : 1'b1;
										assign node344 = (inp[10]) ? node360 : node345;
											assign node345 = (inp[9]) ? node355 : node346;
												assign node346 = (inp[15]) ? node350 : node347;
													assign node347 = (inp[12]) ? 1'b1 : 1'b0;
													assign node350 = (inp[7]) ? 1'b0 : node351;
														assign node351 = (inp[3]) ? 1'b1 : 1'b0;
												assign node355 = (inp[3]) ? node357 : 1'b1;
													assign node357 = (inp[7]) ? 1'b1 : 1'b0;
											assign node360 = (inp[3]) ? node366 : node361;
												assign node361 = (inp[12]) ? node363 : 1'b0;
													assign node363 = (inp[15]) ? 1'b0 : 1'b1;
												assign node366 = (inp[7]) ? node368 : 1'b1;
													assign node368 = (inp[12]) ? node370 : 1'b0;
														assign node370 = (inp[15]) ? 1'b0 : 1'b1;
									assign node373 = (inp[12]) ? node375 : 1'b1;
										assign node375 = (inp[15]) ? 1'b1 : node376;
											assign node376 = (inp[7]) ? node388 : node377;
												assign node377 = (inp[3]) ? node383 : node378;
													assign node378 = (inp[6]) ? node380 : 1'b0;
														assign node380 = (inp[9]) ? 1'b1 : 1'b0;
													assign node383 = (inp[9]) ? node385 : 1'b1;
														assign node385 = (inp[10]) ? 1'b1 : 1'b0;
												assign node388 = (inp[9]) ? node390 : 1'b0;
													assign node390 = (inp[10]) ? 1'b0 : 1'b1;
								assign node394 = (inp[11]) ? node464 : node395;
									assign node395 = (inp[6]) ? node415 : node396;
										assign node396 = (inp[12]) ? node398 : 1'b0;
											assign node398 = (inp[15]) ? 1'b0 : node399;
												assign node399 = (inp[9]) ? node405 : node400;
													assign node400 = (inp[3]) ? node402 : 1'b1;
														assign node402 = (inp[7]) ? 1'b1 : 1'b0;
													assign node405 = (inp[10]) ? node411 : node406;
														assign node406 = (inp[7]) ? 1'b0 : node407;
															assign node407 = (inp[3]) ? 1'b1 : 1'b0;
														assign node411 = (inp[3]) ? 1'b0 : 1'b1;
										assign node415 = (inp[5]) ? node445 : node416;
											assign node416 = (inp[15]) ? node428 : node417;
												assign node417 = (inp[12]) ? 1'b0 : node418;
													assign node418 = (inp[10]) ? 1'b1 : node419;
														assign node419 = (inp[9]) ? 1'b0 : node420;
															assign node420 = (inp[7]) ? 1'b1 : node421;
																assign node421 = (inp[3]) ? 1'b0 : 1'b1;
												assign node428 = (inp[9]) ? node434 : node429;
													assign node429 = (inp[3]) ? node431 : 1'b1;
														assign node431 = (inp[7]) ? 1'b1 : 1'b0;
													assign node434 = (inp[10]) ? node440 : node435;
														assign node435 = (inp[7]) ? 1'b0 : node436;
															assign node436 = (inp[3]) ? 1'b1 : 1'b0;
														assign node440 = (inp[7]) ? 1'b1 : node441;
															assign node441 = (inp[3]) ? 1'b0 : 1'b1;
											assign node445 = (inp[15]) ? 1'b0 : node446;
												assign node446 = (inp[12]) ? node448 : 1'b0;
													assign node448 = (inp[3]) ? node454 : node449;
														assign node449 = (inp[9]) ? node451 : 1'b1;
															assign node451 = (inp[10]) ? 1'b1 : 1'b0;
														assign node454 = (inp[7]) ? node460 : node455;
															assign node455 = (inp[9]) ? node457 : 1'b0;
																assign node457 = (inp[10]) ? 1'b0 : 1'b1;
															assign node460 = (inp[9]) ? 1'b0 : 1'b1;
									assign node464 = (inp[5]) ? node506 : node465;
										assign node465 = (inp[6]) ? node483 : node466;
											assign node466 = (inp[12]) ? node468 : 1'b1;
												assign node468 = (inp[15]) ? 1'b1 : node469;
													assign node469 = (inp[7]) ? node477 : node470;
														assign node470 = (inp[10]) ? 1'b1 : node471;
															assign node471 = (inp[3]) ? 1'b0 : node472;
																assign node472 = (inp[9]) ? 1'b1 : 1'b0;
														assign node477 = (inp[10]) ? 1'b0 : node478;
															assign node478 = (inp[9]) ? 1'b1 : 1'b0;
											assign node483 = (inp[15]) ? node493 : node484;
												assign node484 = (inp[12]) ? 1'b1 : node485;
													assign node485 = (inp[10]) ? node489 : node486;
														assign node486 = (inp[9]) ? 1'b1 : 1'b0;
														assign node489 = (inp[9]) ? 1'b0 : 1'b1;
												assign node493 = (inp[10]) ? node501 : node494;
													assign node494 = (inp[9]) ? node496 : 1'b0;
														assign node496 = (inp[7]) ? 1'b1 : node497;
															assign node497 = (inp[3]) ? 1'b0 : 1'b1;
													assign node501 = (inp[7]) ? 1'b0 : node502;
														assign node502 = (inp[3]) ? 1'b1 : 1'b0;
										assign node506 = (inp[15]) ? 1'b1 : node507;
											assign node507 = (inp[12]) ? node509 : 1'b1;
												assign node509 = (inp[7]) ? node517 : node510;
													assign node510 = (inp[6]) ? 1'b1 : node511;
														assign node511 = (inp[9]) ? 1'b0 : node512;
															assign node512 = (inp[3]) ? 1'b1 : 1'b0;
													assign node517 = (inp[6]) ? 1'b0 : node518;
														assign node518 = (inp[10]) ? 1'b0 : 1'b1;
							assign node523 = (inp[11]) ? node655 : node524;
								assign node524 = (inp[13]) ? node590 : node525;
									assign node525 = (inp[5]) ? node573 : node526;
										assign node526 = (inp[6]) ? node542 : node527;
											assign node527 = (inp[12]) ? node529 : 1'b0;
												assign node529 = (inp[15]) ? 1'b0 : node530;
													assign node530 = (inp[9]) ? node532 : 1'b1;
														assign node532 = (inp[3]) ? node536 : node533;
															assign node533 = (inp[10]) ? 1'b1 : 1'b0;
															assign node536 = (inp[10]) ? 1'b0 : node537;
																assign node537 = (inp[7]) ? 1'b0 : 1'b1;
											assign node542 = (inp[9]) ? node552 : node543;
												assign node543 = (inp[15]) ? 1'b1 : node544;
													assign node544 = (inp[12]) ? 1'b0 : node545;
														assign node545 = (inp[7]) ? 1'b1 : node546;
															assign node546 = (inp[3]) ? 1'b0 : 1'b1;
												assign node552 = (inp[10]) ? node560 : node553;
													assign node553 = (inp[3]) ? node555 : 1'b0;
														assign node555 = (inp[7]) ? 1'b0 : node556;
															assign node556 = (inp[12]) ? 1'b0 : 1'b1;
													assign node560 = (inp[7]) ? node568 : node561;
														assign node561 = (inp[3]) ? 1'b0 : node562;
															assign node562 = (inp[15]) ? 1'b1 : node563;
																assign node563 = (inp[12]) ? 1'b0 : 1'b1;
														assign node568 = (inp[15]) ? 1'b1 : node569;
															assign node569 = (inp[3]) ? 1'b1 : 1'b0;
										assign node573 = (inp[12]) ? node575 : 1'b0;
											assign node575 = (inp[15]) ? 1'b0 : node576;
												assign node576 = (inp[9]) ? node578 : 1'b1;
													assign node578 = (inp[10]) ? node584 : node579;
														assign node579 = (inp[7]) ? 1'b0 : node580;
															assign node580 = (inp[3]) ? 1'b1 : 1'b0;
														assign node584 = (inp[3]) ? node586 : 1'b1;
															assign node586 = (inp[7]) ? 1'b1 : 1'b0;
									assign node590 = (inp[15]) ? node642 : node591;
										assign node591 = (inp[12]) ? node607 : node592;
											assign node592 = (inp[6]) ? node594 : 1'b1;
												assign node594 = (inp[5]) ? 1'b1 : node595;
													assign node595 = (inp[9]) ? node597 : 1'b0;
														assign node597 = (inp[7]) ? 1'b0 : node598;
															assign node598 = (inp[10]) ? node602 : node599;
																assign node599 = (inp[3]) ? 1'b0 : 1'b1;
																assign node602 = (inp[3]) ? 1'b1 : 1'b0;
											assign node607 = (inp[6]) ? node625 : node608;
												assign node608 = (inp[3]) ? node616 : node609;
													assign node609 = (inp[5]) ? node611 : 1'b0;
														assign node611 = (inp[9]) ? node613 : 1'b0;
															assign node613 = (inp[10]) ? 1'b0 : 1'b1;
													assign node616 = (inp[7]) ? node622 : node617;
														assign node617 = (inp[10]) ? 1'b1 : node618;
															assign node618 = (inp[9]) ? 1'b0 : 1'b1;
														assign node622 = (inp[10]) ? 1'b0 : 1'b1;
												assign node625 = (inp[5]) ? node627 : 1'b1;
													assign node627 = (inp[9]) ? node633 : node628;
														assign node628 = (inp[3]) ? node630 : 1'b0;
															assign node630 = (inp[7]) ? 1'b0 : 1'b1;
														assign node633 = (inp[3]) ? node635 : 1'b1;
															assign node635 = (inp[10]) ? node639 : node636;
																assign node636 = (inp[7]) ? 1'b1 : 1'b0;
																assign node639 = (inp[7]) ? 1'b0 : 1'b1;
										assign node642 = (inp[5]) ? 1'b1 : node643;
											assign node643 = (inp[6]) ? node645 : 1'b1;
												assign node645 = (inp[7]) ? node651 : node646;
													assign node646 = (inp[10]) ? 1'b1 : node647;
														assign node647 = (inp[12]) ? 1'b1 : 1'b0;
													assign node651 = (inp[10]) ? 1'b0 : 1'b1;
								assign node655 = (inp[15]) ? node699 : node656;
									assign node656 = (inp[12]) ? node666 : node657;
										assign node657 = (inp[6]) ? node659 : 1'b0;
											assign node659 = (inp[5]) ? 1'b0 : node660;
												assign node660 = (inp[9]) ? node662 : 1'b1;
													assign node662 = (inp[7]) ? 1'b1 : 1'b0;
										assign node666 = (inp[6]) ? node680 : node667;
											assign node667 = (inp[9]) ? node673 : node668;
												assign node668 = (inp[7]) ? 1'b1 : node669;
													assign node669 = (inp[3]) ? 1'b0 : 1'b1;
												assign node673 = (inp[10]) ? 1'b1 : node674;
													assign node674 = (inp[7]) ? 1'b0 : node675;
														assign node675 = (inp[3]) ? 1'b1 : 1'b0;
											assign node680 = (inp[5]) ? node682 : 1'b0;
												assign node682 = (inp[7]) ? node694 : node683;
													assign node683 = (inp[3]) ? node689 : node684;
														assign node684 = (inp[9]) ? node686 : 1'b1;
															assign node686 = (inp[10]) ? 1'b1 : 1'b0;
														assign node689 = (inp[9]) ? node691 : 1'b0;
															assign node691 = (inp[10]) ? 1'b0 : 1'b1;
													assign node694 = (inp[10]) ? 1'b1 : node695;
														assign node695 = (inp[13]) ? 1'b1 : 1'b0;
									assign node699 = (inp[6]) ? node701 : 1'b0;
										assign node701 = (inp[5]) ? 1'b0 : node702;
											assign node702 = (inp[10]) ? node708 : node703;
												assign node703 = (inp[7]) ? node705 : 1'b0;
													assign node705 = (inp[9]) ? 1'b0 : 1'b1;
												assign node708 = (inp[3]) ? node710 : 1'b1;
													assign node710 = (inp[7]) ? 1'b1 : 1'b0;
				assign node714 = (inp[12]) ? node736 : node715;
					assign node715 = (inp[5]) ? 1'b1 : node716;
						assign node716 = (inp[6]) ? node718 : 1'b1;
							assign node718 = (inp[7]) ? node730 : node719;
								assign node719 = (inp[3]) ? node725 : node720;
									assign node720 = (inp[9]) ? node722 : 1'b0;
										assign node722 = (inp[10]) ? 1'b0 : 1'b1;
									assign node725 = (inp[10]) ? 1'b1 : node726;
										assign node726 = (inp[9]) ? 1'b0 : 1'b1;
								assign node730 = (inp[10]) ? 1'b0 : node731;
									assign node731 = (inp[9]) ? 1'b1 : 1'b0;
					assign node736 = (inp[15]) ? node774 : node737;
						assign node737 = (inp[6]) ? node755 : node738;
							assign node738 = (inp[3]) ? node744 : node739;
								assign node739 = (inp[9]) ? node741 : 1'b0;
									assign node741 = (inp[10]) ? 1'b0 : 1'b1;
								assign node744 = (inp[7]) ? node750 : node745;
									assign node745 = (inp[9]) ? node747 : 1'b1;
										assign node747 = (inp[10]) ? 1'b1 : 1'b0;
									assign node750 = (inp[9]) ? node752 : 1'b0;
										assign node752 = (inp[10]) ? 1'b0 : 1'b1;
							assign node755 = (inp[5]) ? node757 : 1'b1;
								assign node757 = (inp[10]) ? node769 : node758;
									assign node758 = (inp[9]) ? node764 : node759;
										assign node759 = (inp[7]) ? 1'b0 : node760;
											assign node760 = (inp[3]) ? 1'b1 : 1'b0;
										assign node764 = (inp[7]) ? 1'b1 : node765;
											assign node765 = (inp[3]) ? 1'b0 : 1'b1;
									assign node769 = (inp[7]) ? 1'b0 : node770;
										assign node770 = (inp[3]) ? 1'b1 : 1'b0;
						assign node774 = (inp[6]) ? node776 : 1'b1;
							assign node776 = (inp[5]) ? 1'b1 : node777;
								assign node777 = (inp[10]) ? node789 : node778;
									assign node778 = (inp[9]) ? node784 : node779;
										assign node779 = (inp[7]) ? 1'b0 : node780;
											assign node780 = (inp[3]) ? 1'b1 : 1'b0;
										assign node784 = (inp[3]) ? node786 : 1'b1;
											assign node786 = (inp[7]) ? 1'b1 : 1'b0;
									assign node789 = (inp[3]) ? node791 : 1'b0;
										assign node791 = (inp[7]) ? 1'b0 : 1'b1;
			assign node795 = (inp[1]) ? node1513 : node796;
				assign node796 = (inp[2]) ? node1272 : node797;
					assign node797 = (inp[14]) ? node1035 : node798;
						assign node798 = (inp[11]) ? node946 : node799;
							assign node799 = (inp[13]) ? node875 : node800;
								assign node800 = (inp[6]) ? node822 : node801;
									assign node801 = (inp[15]) ? 1'b0 : node802;
										assign node802 = (inp[12]) ? node804 : 1'b0;
											assign node804 = (inp[9]) ? node810 : node805;
												assign node805 = (inp[7]) ? 1'b1 : node806;
													assign node806 = (inp[3]) ? 1'b0 : 1'b1;
												assign node810 = (inp[10]) ? node816 : node811;
													assign node811 = (inp[3]) ? node813 : 1'b0;
														assign node813 = (inp[7]) ? 1'b0 : 1'b1;
													assign node816 = (inp[7]) ? 1'b1 : node817;
														assign node817 = (inp[3]) ? 1'b0 : 1'b1;
									assign node822 = (inp[5]) ? node852 : node823;
										assign node823 = (inp[15]) ? node835 : node824;
											assign node824 = (inp[12]) ? 1'b0 : node825;
												assign node825 = (inp[3]) ? node831 : node826;
													assign node826 = (inp[9]) ? node828 : 1'b1;
														assign node828 = (inp[10]) ? 1'b1 : 1'b0;
													assign node831 = (inp[7]) ? 1'b1 : 1'b0;
											assign node835 = (inp[3]) ? node841 : node836;
												assign node836 = (inp[10]) ? 1'b1 : node837;
													assign node837 = (inp[9]) ? 1'b0 : 1'b1;
												assign node841 = (inp[7]) ? node847 : node842;
													assign node842 = (inp[9]) ? node844 : 1'b0;
														assign node844 = (inp[10]) ? 1'b0 : 1'b1;
													assign node847 = (inp[9]) ? node849 : 1'b1;
														assign node849 = (inp[8]) ? 1'b1 : 1'b0;
										assign node852 = (inp[15]) ? 1'b0 : node853;
											assign node853 = (inp[12]) ? node855 : 1'b0;
												assign node855 = (inp[7]) ? node869 : node856;
													assign node856 = (inp[10]) ? 1'b0 : node857;
														assign node857 = (inp[8]) ? node863 : node858;
															assign node858 = (inp[9]) ? node860 : 1'b1;
																assign node860 = (inp[3]) ? 1'b1 : 1'b0;
															assign node863 = (inp[3]) ? node865 : 1'b0;
																assign node865 = (inp[9]) ? 1'b1 : 1'b0;
													assign node869 = (inp[9]) ? node871 : 1'b1;
														assign node871 = (inp[10]) ? 1'b1 : 1'b0;
								assign node875 = (inp[6]) ? node897 : node876;
									assign node876 = (inp[15]) ? 1'b1 : node877;
										assign node877 = (inp[12]) ? node879 : 1'b1;
											assign node879 = (inp[7]) ? node891 : node880;
												assign node880 = (inp[3]) ? node886 : node881;
													assign node881 = (inp[10]) ? 1'b0 : node882;
														assign node882 = (inp[9]) ? 1'b1 : 1'b0;
													assign node886 = (inp[9]) ? node888 : 1'b1;
														assign node888 = (inp[10]) ? 1'b1 : 1'b0;
												assign node891 = (inp[10]) ? 1'b0 : node892;
													assign node892 = (inp[9]) ? 1'b1 : 1'b0;
									assign node897 = (inp[5]) ? node931 : node898;
										assign node898 = (inp[15]) ? node914 : node899;
											assign node899 = (inp[12]) ? 1'b1 : node900;
												assign node900 = (inp[9]) ? node906 : node901;
													assign node901 = (inp[7]) ? 1'b0 : node902;
														assign node902 = (inp[3]) ? 1'b1 : 1'b0;
													assign node906 = (inp[10]) ? 1'b0 : node907;
														assign node907 = (inp[3]) ? node909 : 1'b1;
															assign node909 = (inp[7]) ? 1'b1 : 1'b0;
											assign node914 = (inp[7]) ? node926 : node915;
												assign node915 = (inp[3]) ? node921 : node916;
													assign node916 = (inp[9]) ? node918 : 1'b0;
														assign node918 = (inp[10]) ? 1'b0 : 1'b1;
													assign node921 = (inp[10]) ? 1'b1 : node922;
														assign node922 = (inp[9]) ? 1'b0 : 1'b1;
												assign node926 = (inp[9]) ? node928 : 1'b0;
													assign node928 = (inp[10]) ? 1'b0 : 1'b1;
										assign node931 = (inp[12]) ? node933 : 1'b1;
											assign node933 = (inp[15]) ? 1'b1 : node934;
												assign node934 = (inp[7]) ? 1'b0 : node935;
													assign node935 = (inp[3]) ? node941 : node936;
														assign node936 = (inp[10]) ? 1'b0 : node937;
															assign node937 = (inp[9]) ? 1'b1 : 1'b0;
														assign node941 = (inp[9]) ? 1'b0 : 1'b1;
							assign node946 = (inp[6]) ? node968 : node947;
								assign node947 = (inp[12]) ? node949 : 1'b0;
									assign node949 = (inp[15]) ? 1'b0 : node950;
										assign node950 = (inp[3]) ? node956 : node951;
											assign node951 = (inp[10]) ? 1'b1 : node952;
												assign node952 = (inp[9]) ? 1'b0 : 1'b1;
											assign node956 = (inp[7]) ? node962 : node957;
												assign node957 = (inp[9]) ? node959 : 1'b0;
													assign node959 = (inp[10]) ? 1'b0 : 1'b1;
												assign node962 = (inp[9]) ? node964 : 1'b1;
													assign node964 = (inp[10]) ? 1'b1 : 1'b0;
								assign node968 = (inp[5]) ? node1014 : node969;
									assign node969 = (inp[15]) ? node997 : node970;
										assign node970 = (inp[12]) ? 1'b0 : node971;
											assign node971 = (inp[3]) ? node977 : node972;
												assign node972 = (inp[10]) ? 1'b1 : node973;
													assign node973 = (inp[9]) ? 1'b0 : 1'b1;
												assign node977 = (inp[8]) ? node989 : node978;
													assign node978 = (inp[7]) ? node984 : node979;
														assign node979 = (inp[10]) ? 1'b0 : node980;
															assign node980 = (inp[9]) ? 1'b1 : 1'b0;
														assign node984 = (inp[10]) ? 1'b1 : node985;
															assign node985 = (inp[9]) ? 1'b0 : 1'b1;
													assign node989 = (inp[10]) ? 1'b0 : node990;
														assign node990 = (inp[9]) ? node992 : 1'b0;
															assign node992 = (inp[13]) ? 1'b1 : 1'b0;
										assign node997 = (inp[10]) ? node1009 : node998;
											assign node998 = (inp[9]) ? node1004 : node999;
												assign node999 = (inp[3]) ? node1001 : 1'b1;
													assign node1001 = (inp[7]) ? 1'b1 : 1'b0;
												assign node1004 = (inp[3]) ? node1006 : 1'b0;
													assign node1006 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1009 = (inp[7]) ? 1'b1 : node1010;
												assign node1010 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1014 = (inp[15]) ? 1'b0 : node1015;
										assign node1015 = (inp[12]) ? node1017 : 1'b0;
											assign node1017 = (inp[3]) ? node1023 : node1018;
												assign node1018 = (inp[10]) ? 1'b1 : node1019;
													assign node1019 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1023 = (inp[7]) ? node1029 : node1024;
													assign node1024 = (inp[10]) ? 1'b0 : node1025;
														assign node1025 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1029 = (inp[9]) ? node1031 : 1'b1;
														assign node1031 = (inp[10]) ? 1'b1 : 1'b0;
						assign node1035 = (inp[11]) ? node1191 : node1036;
							assign node1036 = (inp[13]) ? node1114 : node1037;
								assign node1037 = (inp[5]) ? node1093 : node1038;
									assign node1038 = (inp[6]) ? node1060 : node1039;
										assign node1039 = (inp[15]) ? 1'b1 : node1040;
											assign node1040 = (inp[12]) ? node1042 : 1'b1;
												assign node1042 = (inp[10]) ? node1054 : node1043;
													assign node1043 = (inp[9]) ? node1049 : node1044;
														assign node1044 = (inp[7]) ? 1'b0 : node1045;
															assign node1045 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1049 = (inp[3]) ? node1051 : 1'b1;
															assign node1051 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1054 = (inp[3]) ? node1056 : 1'b0;
														assign node1056 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1060 = (inp[15]) ? node1078 : node1061;
											assign node1061 = (inp[12]) ? 1'b1 : node1062;
												assign node1062 = (inp[10]) ? node1074 : node1063;
													assign node1063 = (inp[3]) ? node1065 : 1'b1;
														assign node1065 = (inp[8]) ? node1067 : 1'b0;
															assign node1067 = (inp[7]) ? node1071 : node1068;
																assign node1068 = (inp[9]) ? 1'b0 : 1'b1;
																assign node1071 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1074 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1078 = (inp[7]) ? node1088 : node1079;
												assign node1079 = (inp[3]) ? node1085 : node1080;
													assign node1080 = (inp[9]) ? node1082 : 1'b0;
														assign node1082 = (inp[8]) ? 1'b0 : 1'b1;
													assign node1085 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1088 = (inp[9]) ? node1090 : 1'b0;
													assign node1090 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1093 = (inp[12]) ? node1095 : 1'b1;
										assign node1095 = (inp[15]) ? 1'b1 : node1096;
											assign node1096 = (inp[7]) ? node1108 : node1097;
												assign node1097 = (inp[3]) ? node1103 : node1098;
													assign node1098 = (inp[6]) ? node1100 : 1'b0;
														assign node1100 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1103 = (inp[10]) ? 1'b1 : node1104;
														assign node1104 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1108 = (inp[9]) ? node1110 : 1'b0;
													assign node1110 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1114 = (inp[6]) ? node1136 : node1115;
									assign node1115 = (inp[12]) ? node1117 : 1'b0;
										assign node1117 = (inp[15]) ? 1'b0 : node1118;
											assign node1118 = (inp[9]) ? node1124 : node1119;
												assign node1119 = (inp[3]) ? node1121 : 1'b1;
													assign node1121 = (inp[7]) ? 1'b1 : 1'b0;
												assign node1124 = (inp[10]) ? node1130 : node1125;
													assign node1125 = (inp[7]) ? 1'b0 : node1126;
														assign node1126 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1130 = (inp[7]) ? 1'b1 : node1131;
														assign node1131 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1136 = (inp[5]) ? node1172 : node1137;
										assign node1137 = (inp[15]) ? node1155 : node1138;
											assign node1138 = (inp[12]) ? 1'b0 : node1139;
												assign node1139 = (inp[7]) ? node1149 : node1140;
													assign node1140 = (inp[3]) ? node1146 : node1141;
														assign node1141 = (inp[10]) ? 1'b1 : node1142;
															assign node1142 = (inp[9]) ? 1'b0 : 1'b1;
														assign node1146 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1149 = (inp[10]) ? 1'b1 : node1150;
														assign node1150 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1155 = (inp[3]) ? node1161 : node1156;
												assign node1156 = (inp[10]) ? 1'b1 : node1157;
													assign node1157 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1161 = (inp[7]) ? node1167 : node1162;
													assign node1162 = (inp[10]) ? 1'b0 : node1163;
														assign node1163 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1167 = (inp[10]) ? 1'b1 : node1168;
														assign node1168 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1172 = (inp[12]) ? node1174 : 1'b0;
											assign node1174 = (inp[15]) ? 1'b0 : node1175;
												assign node1175 = (inp[3]) ? node1183 : node1176;
													assign node1176 = (inp[8]) ? node1178 : 1'b1;
														assign node1178 = (inp[7]) ? node1180 : 1'b1;
															assign node1180 = (inp[9]) ? 1'b0 : 1'b1;
													assign node1183 = (inp[7]) ? node1185 : 1'b0;
														assign node1185 = (inp[10]) ? 1'b1 : node1186;
															assign node1186 = (inp[9]) ? 1'b0 : 1'b1;
							assign node1191 = (inp[12]) ? node1213 : node1192;
								assign node1192 = (inp[5]) ? 1'b1 : node1193;
									assign node1193 = (inp[6]) ? node1195 : 1'b1;
										assign node1195 = (inp[3]) ? node1201 : node1196;
											assign node1196 = (inp[9]) ? node1198 : 1'b0;
												assign node1198 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1201 = (inp[7]) ? node1207 : node1202;
												assign node1202 = (inp[9]) ? node1204 : 1'b1;
													assign node1204 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1207 = (inp[10]) ? 1'b0 : node1208;
													assign node1208 = (inp[9]) ? 1'b1 : 1'b0;
								assign node1213 = (inp[15]) ? node1251 : node1214;
									assign node1214 = (inp[9]) ? node1228 : node1215;
										assign node1215 = (inp[5]) ? node1223 : node1216;
											assign node1216 = (inp[6]) ? 1'b1 : node1217;
												assign node1217 = (inp[3]) ? node1219 : 1'b0;
													assign node1219 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1223 = (inp[7]) ? 1'b0 : node1224;
												assign node1224 = (inp[3]) ? 1'b1 : 1'b0;
										assign node1228 = (inp[10]) ? node1238 : node1229;
											assign node1229 = (inp[3]) ? node1231 : 1'b1;
												assign node1231 = (inp[7]) ? 1'b1 : node1232;
													assign node1232 = (inp[5]) ? 1'b0 : node1233;
														assign node1233 = (inp[6]) ? 1'b1 : 1'b0;
											assign node1238 = (inp[3]) ? node1244 : node1239;
												assign node1239 = (inp[6]) ? node1241 : 1'b0;
													assign node1241 = (inp[5]) ? 1'b0 : 1'b1;
												assign node1244 = (inp[7]) ? node1246 : 1'b1;
													assign node1246 = (inp[5]) ? 1'b0 : node1247;
														assign node1247 = (inp[6]) ? 1'b1 : 1'b0;
									assign node1251 = (inp[6]) ? node1253 : 1'b1;
										assign node1253 = (inp[5]) ? 1'b1 : node1254;
											assign node1254 = (inp[3]) ? node1260 : node1255;
												assign node1255 = (inp[10]) ? 1'b0 : node1256;
													assign node1256 = (inp[9]) ? 1'b1 : 1'b0;
												assign node1260 = (inp[7]) ? node1266 : node1261;
													assign node1261 = (inp[9]) ? node1263 : 1'b1;
														assign node1263 = (inp[10]) ? 1'b1 : 1'b0;
													assign node1266 = (inp[9]) ? node1268 : 1'b0;
														assign node1268 = (inp[13]) ? 1'b0 : 1'b1;
					assign node1272 = (inp[13]) ? node1354 : node1273;
						assign node1273 = (inp[12]) ? node1295 : node1274;
							assign node1274 = (inp[6]) ? node1276 : 1'b0;
								assign node1276 = (inp[5]) ? 1'b0 : node1277;
									assign node1277 = (inp[3]) ? node1283 : node1278;
										assign node1278 = (inp[9]) ? node1280 : 1'b1;
											assign node1280 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1283 = (inp[7]) ? node1289 : node1284;
											assign node1284 = (inp[9]) ? node1286 : 1'b0;
												assign node1286 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1289 = (inp[9]) ? node1291 : 1'b1;
												assign node1291 = (inp[10]) ? 1'b1 : 1'b0;
							assign node1295 = (inp[15]) ? node1333 : node1296;
								assign node1296 = (inp[6]) ? node1314 : node1297;
									assign node1297 = (inp[9]) ? node1303 : node1298;
										assign node1298 = (inp[7]) ? 1'b1 : node1299;
											assign node1299 = (inp[3]) ? 1'b0 : 1'b1;
										assign node1303 = (inp[10]) ? node1309 : node1304;
											assign node1304 = (inp[7]) ? 1'b0 : node1305;
												assign node1305 = (inp[3]) ? 1'b1 : 1'b0;
											assign node1309 = (inp[7]) ? 1'b1 : node1310;
												assign node1310 = (inp[3]) ? 1'b0 : 1'b1;
									assign node1314 = (inp[5]) ? node1316 : 1'b0;
										assign node1316 = (inp[7]) ? node1328 : node1317;
											assign node1317 = (inp[3]) ? node1323 : node1318;
												assign node1318 = (inp[9]) ? node1320 : 1'b1;
													assign node1320 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1323 = (inp[9]) ? node1325 : 1'b0;
													assign node1325 = (inp[10]) ? 1'b0 : 1'b1;
											assign node1328 = (inp[10]) ? 1'b1 : node1329;
												assign node1329 = (inp[9]) ? 1'b0 : 1'b1;
								assign node1333 = (inp[5]) ? 1'b0 : node1334;
									assign node1334 = (inp[6]) ? node1336 : 1'b0;
										assign node1336 = (inp[3]) ? node1342 : node1337;
											assign node1337 = (inp[9]) ? node1339 : 1'b1;
												assign node1339 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1342 = (inp[7]) ? node1348 : node1343;
												assign node1343 = (inp[9]) ? node1345 : 1'b0;
													assign node1345 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1348 = (inp[9]) ? node1350 : 1'b1;
													assign node1350 = (inp[10]) ? 1'b1 : 1'b0;
						assign node1354 = (inp[11]) ? node1432 : node1355;
							assign node1355 = (inp[15]) ? node1411 : node1356;
								assign node1356 = (inp[12]) ? node1378 : node1357;
									assign node1357 = (inp[6]) ? node1359 : 1'b1;
										assign node1359 = (inp[5]) ? 1'b1 : node1360;
											assign node1360 = (inp[7]) ? node1372 : node1361;
												assign node1361 = (inp[3]) ? node1367 : node1362;
													assign node1362 = (inp[10]) ? 1'b0 : node1363;
														assign node1363 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1367 = (inp[9]) ? node1369 : 1'b1;
														assign node1369 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1372 = (inp[9]) ? node1374 : 1'b0;
													assign node1374 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1378 = (inp[5]) ? node1394 : node1379;
										assign node1379 = (inp[6]) ? 1'b1 : node1380;
											assign node1380 = (inp[3]) ? node1386 : node1381;
												assign node1381 = (inp[9]) ? node1383 : 1'b0;
													assign node1383 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1386 = (inp[7]) ? node1390 : node1387;
													assign node1387 = (inp[10]) ? 1'b1 : 1'b0;
													assign node1390 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1394 = (inp[10]) ? node1406 : node1395;
											assign node1395 = (inp[9]) ? node1401 : node1396;
												assign node1396 = (inp[3]) ? node1398 : 1'b0;
													assign node1398 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1401 = (inp[7]) ? 1'b1 : node1402;
													assign node1402 = (inp[3]) ? 1'b0 : 1'b1;
											assign node1406 = (inp[3]) ? node1408 : 1'b0;
												assign node1408 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1411 = (inp[6]) ? node1413 : 1'b1;
									assign node1413 = (inp[5]) ? 1'b1 : node1414;
										assign node1414 = (inp[3]) ? node1420 : node1415;
											assign node1415 = (inp[10]) ? 1'b0 : node1416;
												assign node1416 = (inp[9]) ? 1'b1 : 1'b0;
											assign node1420 = (inp[7]) ? node1426 : node1421;
												assign node1421 = (inp[10]) ? 1'b1 : node1422;
													assign node1422 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1426 = (inp[10]) ? 1'b0 : node1427;
													assign node1427 = (inp[9]) ? 1'b1 : 1'b0;
							assign node1432 = (inp[5]) ? node1492 : node1433;
								assign node1433 = (inp[6]) ? node1455 : node1434;
									assign node1434 = (inp[12]) ? node1436 : 1'b0;
										assign node1436 = (inp[15]) ? 1'b0 : node1437;
											assign node1437 = (inp[9]) ? node1443 : node1438;
												assign node1438 = (inp[3]) ? node1440 : 1'b1;
													assign node1440 = (inp[7]) ? 1'b1 : 1'b0;
												assign node1443 = (inp[10]) ? node1449 : node1444;
													assign node1444 = (inp[7]) ? 1'b0 : node1445;
														assign node1445 = (inp[3]) ? 1'b1 : 1'b0;
													assign node1449 = (inp[3]) ? node1451 : 1'b1;
														assign node1451 = (inp[7]) ? 1'b1 : 1'b0;
									assign node1455 = (inp[15]) ? node1475 : node1456;
										assign node1456 = (inp[12]) ? 1'b0 : node1457;
											assign node1457 = (inp[7]) ? node1469 : node1458;
												assign node1458 = (inp[10]) ? node1466 : node1459;
													assign node1459 = (inp[3]) ? node1463 : node1460;
														assign node1460 = (inp[14]) ? 1'b0 : 1'b1;
														assign node1463 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1466 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1469 = (inp[9]) ? node1471 : 1'b1;
													assign node1471 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1475 = (inp[10]) ? node1487 : node1476;
											assign node1476 = (inp[9]) ? node1482 : node1477;
												assign node1477 = (inp[7]) ? 1'b1 : node1478;
													assign node1478 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1482 = (inp[7]) ? 1'b0 : node1483;
													assign node1483 = (inp[3]) ? 1'b1 : 1'b0;
											assign node1487 = (inp[3]) ? node1489 : 1'b1;
												assign node1489 = (inp[7]) ? 1'b1 : 1'b0;
								assign node1492 = (inp[12]) ? node1494 : 1'b0;
									assign node1494 = (inp[15]) ? 1'b0 : node1495;
										assign node1495 = (inp[10]) ? node1507 : node1496;
											assign node1496 = (inp[9]) ? node1502 : node1497;
												assign node1497 = (inp[7]) ? 1'b1 : node1498;
													assign node1498 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1502 = (inp[3]) ? node1504 : 1'b0;
													assign node1504 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1507 = (inp[3]) ? node1509 : 1'b1;
												assign node1509 = (inp[7]) ? 1'b1 : 1'b0;
				assign node1513 = (inp[8]) ? node1595 : node1514;
					assign node1514 = (inp[6]) ? node1536 : node1515;
						assign node1515 = (inp[12]) ? node1517 : 1'b1;
							assign node1517 = (inp[15]) ? 1'b1 : node1518;
								assign node1518 = (inp[10]) ? node1530 : node1519;
									assign node1519 = (inp[9]) ? node1525 : node1520;
										assign node1520 = (inp[3]) ? node1522 : 1'b0;
											assign node1522 = (inp[7]) ? 1'b0 : 1'b1;
										assign node1525 = (inp[3]) ? node1527 : 1'b1;
											assign node1527 = (inp[7]) ? 1'b1 : 1'b0;
									assign node1530 = (inp[7]) ? 1'b0 : node1531;
										assign node1531 = (inp[3]) ? 1'b1 : 1'b0;
						assign node1536 = (inp[5]) ? node1574 : node1537;
							assign node1537 = (inp[12]) ? node1555 : node1538;
								assign node1538 = (inp[3]) ? node1544 : node1539;
									assign node1539 = (inp[10]) ? 1'b0 : node1540;
										assign node1540 = (inp[9]) ? 1'b1 : 1'b0;
									assign node1544 = (inp[7]) ? node1550 : node1545;
										assign node1545 = (inp[9]) ? node1547 : 1'b1;
											assign node1547 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1550 = (inp[10]) ? 1'b0 : node1551;
											assign node1551 = (inp[9]) ? 1'b1 : 1'b0;
								assign node1555 = (inp[15]) ? node1557 : 1'b1;
									assign node1557 = (inp[7]) ? node1569 : node1558;
										assign node1558 = (inp[3]) ? node1564 : node1559;
											assign node1559 = (inp[10]) ? 1'b0 : node1560;
												assign node1560 = (inp[9]) ? 1'b1 : 1'b0;
											assign node1564 = (inp[9]) ? node1566 : 1'b1;
												assign node1566 = (inp[10]) ? 1'b1 : 1'b0;
										assign node1569 = (inp[9]) ? node1571 : 1'b0;
											assign node1571 = (inp[10]) ? 1'b0 : 1'b1;
							assign node1574 = (inp[12]) ? node1576 : 1'b1;
								assign node1576 = (inp[15]) ? 1'b1 : node1577;
									assign node1577 = (inp[3]) ? node1583 : node1578;
										assign node1578 = (inp[10]) ? 1'b0 : node1579;
											assign node1579 = (inp[9]) ? 1'b1 : 1'b0;
										assign node1583 = (inp[7]) ? node1589 : node1584;
											assign node1584 = (inp[9]) ? node1586 : 1'b1;
												assign node1586 = (inp[10]) ? 1'b1 : 1'b0;
											assign node1589 = (inp[9]) ? node1591 : 1'b0;
												assign node1591 = (inp[10]) ? 1'b0 : 1'b1;
					assign node1595 = (inp[13]) ? node1821 : node1596;
						assign node1596 = (inp[14]) ? node1676 : node1597;
							assign node1597 = (inp[15]) ? node1655 : node1598;
								assign node1598 = (inp[12]) ? node1618 : node1599;
									assign node1599 = (inp[6]) ? node1601 : 1'b0;
										assign node1601 = (inp[5]) ? 1'b0 : node1602;
											assign node1602 = (inp[10]) ? node1612 : node1603;
												assign node1603 = (inp[9]) ? node1607 : node1604;
													assign node1604 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1607 = (inp[3]) ? node1609 : 1'b0;
														assign node1609 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1612 = (inp[3]) ? node1614 : 1'b1;
													assign node1614 = (inp[7]) ? 1'b1 : 1'b0;
									assign node1618 = (inp[5]) ? node1638 : node1619;
										assign node1619 = (inp[6]) ? 1'b0 : node1620;
											assign node1620 = (inp[3]) ? node1626 : node1621;
												assign node1621 = (inp[10]) ? 1'b1 : node1622;
													assign node1622 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1626 = (inp[7]) ? node1632 : node1627;
													assign node1627 = (inp[10]) ? 1'b0 : node1628;
														assign node1628 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1632 = (inp[2]) ? 1'b1 : node1633;
														assign node1633 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1638 = (inp[3]) ? node1644 : node1639;
											assign node1639 = (inp[10]) ? 1'b1 : node1640;
												assign node1640 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1644 = (inp[7]) ? node1650 : node1645;
												assign node1645 = (inp[9]) ? node1647 : 1'b0;
													assign node1647 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1650 = (inp[9]) ? node1652 : 1'b1;
													assign node1652 = (inp[10]) ? 1'b1 : 1'b0;
								assign node1655 = (inp[6]) ? node1657 : 1'b0;
									assign node1657 = (inp[5]) ? 1'b0 : node1658;
										assign node1658 = (inp[9]) ? node1664 : node1659;
											assign node1659 = (inp[3]) ? node1661 : 1'b1;
												assign node1661 = (inp[7]) ? 1'b1 : 1'b0;
											assign node1664 = (inp[10]) ? node1670 : node1665;
												assign node1665 = (inp[3]) ? node1667 : 1'b0;
													assign node1667 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1670 = (inp[3]) ? node1672 : 1'b1;
													assign node1672 = (inp[7]) ? 1'b1 : 1'b0;
							assign node1676 = (inp[2]) ? node1750 : node1677;
								assign node1677 = (inp[6]) ? node1695 : node1678;
									assign node1678 = (inp[12]) ? node1680 : 1'b1;
										assign node1680 = (inp[15]) ? 1'b1 : node1681;
											assign node1681 = (inp[3]) ? node1687 : node1682;
												assign node1682 = (inp[10]) ? 1'b0 : node1683;
													assign node1683 = (inp[9]) ? 1'b1 : 1'b0;
												assign node1687 = (inp[7]) ? node1689 : 1'b1;
													assign node1689 = (inp[9]) ? node1691 : 1'b0;
														assign node1691 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1695 = (inp[5]) ? node1733 : node1696;
										assign node1696 = (inp[12]) ? node1714 : node1697;
											assign node1697 = (inp[9]) ? node1703 : node1698;
												assign node1698 = (inp[3]) ? node1700 : 1'b0;
													assign node1700 = (inp[7]) ? 1'b0 : 1'b1;
												assign node1703 = (inp[10]) ? node1709 : node1704;
													assign node1704 = (inp[7]) ? 1'b1 : node1705;
														assign node1705 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1709 = (inp[7]) ? 1'b0 : node1710;
														assign node1710 = (inp[3]) ? 1'b1 : 1'b0;
											assign node1714 = (inp[15]) ? node1716 : 1'b1;
												assign node1716 = (inp[3]) ? node1722 : node1717;
													assign node1717 = (inp[9]) ? node1719 : 1'b0;
														assign node1719 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1722 = (inp[7]) ? node1728 : node1723;
														assign node1723 = (inp[10]) ? 1'b1 : node1724;
															assign node1724 = (inp[9]) ? 1'b0 : 1'b1;
														assign node1728 = (inp[9]) ? node1730 : 1'b0;
															assign node1730 = (inp[10]) ? 1'b0 : 1'b1;
										assign node1733 = (inp[12]) ? node1735 : 1'b1;
											assign node1735 = (inp[15]) ? 1'b1 : node1736;
												assign node1736 = (inp[11]) ? 1'b0 : node1737;
													assign node1737 = (inp[10]) ? node1743 : node1738;
														assign node1738 = (inp[9]) ? 1'b1 : node1739;
															assign node1739 = (inp[3]) ? 1'b1 : 1'b0;
														assign node1743 = (inp[3]) ? node1745 : 1'b0;
															assign node1745 = (inp[7]) ? 1'b0 : 1'b1;
								assign node1750 = (inp[6]) ? node1772 : node1751;
									assign node1751 = (inp[15]) ? 1'b0 : node1752;
										assign node1752 = (inp[12]) ? node1754 : 1'b0;
											assign node1754 = (inp[3]) ? node1760 : node1755;
												assign node1755 = (inp[9]) ? node1757 : 1'b1;
													assign node1757 = (inp[10]) ? 1'b1 : 1'b0;
												assign node1760 = (inp[7]) ? node1766 : node1761;
													assign node1761 = (inp[9]) ? node1763 : 1'b0;
														assign node1763 = (inp[10]) ? 1'b0 : 1'b1;
													assign node1766 = (inp[10]) ? 1'b1 : node1767;
														assign node1767 = (inp[9]) ? 1'b0 : 1'b1;
									assign node1772 = (inp[5]) ? node1804 : node1773;
										assign node1773 = (inp[10]) ? node1795 : node1774;
											assign node1774 = (inp[9]) ? node1786 : node1775;
												assign node1775 = (inp[15]) ? node1781 : node1776;
													assign node1776 = (inp[12]) ? 1'b0 : node1777;
														assign node1777 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1781 = (inp[3]) ? node1783 : 1'b1;
														assign node1783 = (inp[11]) ? 1'b1 : 1'b0;
												assign node1786 = (inp[3]) ? node1788 : 1'b0;
													assign node1788 = (inp[7]) ? 1'b0 : node1789;
														assign node1789 = (inp[11]) ? node1791 : 1'b1;
															assign node1791 = (inp[12]) ? 1'b0 : 1'b1;
											assign node1795 = (inp[7]) ? node1799 : node1796;
												assign node1796 = (inp[3]) ? 1'b0 : 1'b1;
												assign node1799 = (inp[15]) ? 1'b1 : node1800;
													assign node1800 = (inp[12]) ? 1'b0 : 1'b1;
										assign node1804 = (inp[12]) ? node1806 : 1'b0;
											assign node1806 = (inp[15]) ? 1'b0 : node1807;
												assign node1807 = (inp[10]) ? node1815 : node1808;
													assign node1808 = (inp[9]) ? 1'b0 : node1809;
														assign node1809 = (inp[7]) ? 1'b1 : node1810;
															assign node1810 = (inp[11]) ? 1'b0 : 1'b1;
													assign node1815 = (inp[3]) ? node1817 : 1'b1;
														assign node1817 = (inp[7]) ? 1'b1 : 1'b0;
						assign node1821 = (inp[11]) ? node2003 : node1822;
							assign node1822 = (inp[14]) ? node1898 : node1823;
								assign node1823 = (inp[15]) ? node1877 : node1824;
									assign node1824 = (inp[12]) ? node1840 : node1825;
										assign node1825 = (inp[5]) ? 1'b1 : node1826;
											assign node1826 = (inp[6]) ? node1828 : 1'b1;
												assign node1828 = (inp[3]) ? node1834 : node1829;
													assign node1829 = (inp[10]) ? 1'b0 : node1830;
														assign node1830 = (inp[9]) ? 1'b1 : 1'b0;
													assign node1834 = (inp[10]) ? 1'b1 : node1835;
														assign node1835 = (inp[9]) ? 1'b1 : 1'b0;
										assign node1840 = (inp[5]) ? node1860 : node1841;
											assign node1841 = (inp[6]) ? 1'b1 : node1842;
												assign node1842 = (inp[10]) ? node1854 : node1843;
													assign node1843 = (inp[9]) ? node1849 : node1844;
														assign node1844 = (inp[3]) ? node1846 : 1'b0;
															assign node1846 = (inp[7]) ? 1'b0 : 1'b1;
														assign node1849 = (inp[3]) ? node1851 : 1'b1;
															assign node1851 = (inp[7]) ? 1'b1 : 1'b0;
													assign node1854 = (inp[2]) ? 1'b0 : node1855;
														assign node1855 = (inp[7]) ? 1'b0 : 1'b1;
											assign node1860 = (inp[3]) ? node1866 : node1861;
												assign node1861 = (inp[10]) ? 1'b0 : node1862;
													assign node1862 = (inp[9]) ? 1'b1 : 1'b0;
												assign node1866 = (inp[7]) ? node1872 : node1867;
													assign node1867 = (inp[9]) ? node1869 : 1'b1;
														assign node1869 = (inp[10]) ? 1'b1 : 1'b0;
													assign node1872 = (inp[9]) ? node1874 : 1'b0;
														assign node1874 = (inp[10]) ? 1'b0 : 1'b1;
									assign node1877 = (inp[5]) ? 1'b1 : node1878;
										assign node1878 = (inp[6]) ? node1880 : 1'b1;
											assign node1880 = (inp[3]) ? node1886 : node1881;
												assign node1881 = (inp[9]) ? node1883 : 1'b0;
													assign node1883 = (inp[10]) ? 1'b0 : 1'b1;
												assign node1886 = (inp[2]) ? node1888 : 1'b1;
													assign node1888 = (inp[9]) ? node1890 : 1'b1;
														assign node1890 = (inp[7]) ? node1894 : node1891;
															assign node1891 = (inp[10]) ? 1'b1 : 1'b0;
															assign node1894 = (inp[10]) ? 1'b0 : 1'b1;
								assign node1898 = (inp[2]) ? node1958 : node1899;
									assign node1899 = (inp[5]) ? node1947 : node1900;
										assign node1900 = (inp[6]) ? node1914 : node1901;
											assign node1901 = (inp[15]) ? 1'b0 : node1902;
												assign node1902 = (inp[12]) ? node1904 : 1'b0;
													assign node1904 = (inp[7]) ? node1908 : node1905;
														assign node1905 = (inp[3]) ? 1'b0 : 1'b1;
														assign node1908 = (inp[3]) ? 1'b1 : node1909;
															assign node1909 = (inp[9]) ? 1'b0 : 1'b1;
											assign node1914 = (inp[12]) ? node1938 : node1915;
												assign node1915 = (inp[15]) ? node1927 : node1916;
													assign node1916 = (inp[9]) ? node1918 : 1'b1;
														assign node1918 = (inp[10]) ? node1922 : node1919;
															assign node1919 = (inp[7]) ? 1'b0 : 1'b1;
															assign node1922 = (inp[7]) ? 1'b1 : node1923;
																assign node1923 = (inp[3]) ? 1'b0 : 1'b1;
													assign node1927 = (inp[7]) ? node1935 : node1928;
														assign node1928 = (inp[9]) ? node1930 : 1'b0;
															assign node1930 = (inp[10]) ? node1932 : 1'b1;
																assign node1932 = (inp[3]) ? 1'b0 : 1'b1;
														assign node1935 = (inp[9]) ? 1'b0 : 1'b1;
												assign node1938 = (inp[15]) ? node1940 : 1'b0;
													assign node1940 = (inp[10]) ? 1'b1 : node1941;
														assign node1941 = (inp[3]) ? 1'b0 : node1942;
															assign node1942 = (inp[9]) ? 1'b0 : 1'b1;
										assign node1947 = (inp[15]) ? 1'b0 : node1948;
											assign node1948 = (inp[12]) ? node1950 : 1'b0;
												assign node1950 = (inp[9]) ? node1952 : 1'b1;
													assign node1952 = (inp[6]) ? 1'b0 : node1953;
														assign node1953 = (inp[7]) ? 1'b0 : 1'b1;
									assign node1958 = (inp[5]) ? node1994 : node1959;
										assign node1959 = (inp[6]) ? node1975 : node1960;
											assign node1960 = (inp[15]) ? 1'b1 : node1961;
												assign node1961 = (inp[12]) ? node1963 : 1'b1;
													assign node1963 = (inp[7]) ? node1969 : node1964;
														assign node1964 = (inp[10]) ? 1'b1 : node1965;
															assign node1965 = (inp[9]) ? 1'b1 : 1'b0;
														assign node1969 = (inp[10]) ? 1'b0 : node1970;
															assign node1970 = (inp[9]) ? 1'b1 : 1'b0;
											assign node1975 = (inp[9]) ? node1985 : node1976;
												assign node1976 = (inp[7]) ? 1'b0 : node1977;
													assign node1977 = (inp[12]) ? node1979 : 1'b0;
														assign node1979 = (inp[15]) ? node1981 : 1'b1;
															assign node1981 = (inp[3]) ? 1'b1 : 1'b0;
												assign node1985 = (inp[12]) ? 1'b1 : node1986;
													assign node1986 = (inp[10]) ? node1988 : 1'b1;
														assign node1988 = (inp[7]) ? 1'b0 : node1989;
															assign node1989 = (inp[3]) ? 1'b1 : 1'b0;
										assign node1994 = (inp[12]) ? node1996 : 1'b1;
											assign node1996 = (inp[15]) ? 1'b1 : node1997;
												assign node1997 = (inp[9]) ? node1999 : 1'b0;
													assign node1999 = (inp[10]) ? 1'b0 : 1'b1;
							assign node2003 = (inp[2]) ? node2135 : node2004;
								assign node2004 = (inp[14]) ? node2074 : node2005;
									assign node2005 = (inp[15]) ? node2057 : node2006;
										assign node2006 = (inp[7]) ? node2032 : node2007;
											assign node2007 = (inp[12]) ? node2017 : node2008;
												assign node2008 = (inp[6]) ? node2010 : 1'b0;
													assign node2010 = (inp[3]) ? 1'b0 : node2011;
														assign node2011 = (inp[5]) ? 1'b0 : node2012;
															assign node2012 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2017 = (inp[3]) ? node2027 : node2018;
													assign node2018 = (inp[10]) ? node2024 : node2019;
														assign node2019 = (inp[5]) ? node2021 : 1'b0;
															assign node2021 = (inp[9]) ? 1'b0 : 1'b1;
														assign node2024 = (inp[6]) ? 1'b0 : 1'b1;
													assign node2027 = (inp[10]) ? 1'b0 : node2028;
														assign node2028 = (inp[9]) ? 1'b1 : 1'b0;
											assign node2032 = (inp[10]) ? node2050 : node2033;
												assign node2033 = (inp[9]) ? 1'b0 : node2034;
													assign node2034 = (inp[3]) ? node2040 : node2035;
														assign node2035 = (inp[6]) ? node2037 : 1'b0;
															assign node2037 = (inp[12]) ? 1'b0 : 1'b1;
														assign node2040 = (inp[6]) ? node2042 : 1'b1;
															assign node2042 = (inp[12]) ? node2046 : node2043;
																assign node2043 = (inp[5]) ? 1'b0 : 1'b1;
																assign node2046 = (inp[5]) ? 1'b1 : 1'b0;
												assign node2050 = (inp[12]) ? 1'b1 : node2051;
													assign node2051 = (inp[6]) ? node2053 : 1'b0;
														assign node2053 = (inp[5]) ? 1'b0 : 1'b1;
										assign node2057 = (inp[6]) ? node2059 : 1'b0;
											assign node2059 = (inp[5]) ? 1'b0 : node2060;
												assign node2060 = (inp[3]) ? node2066 : node2061;
													assign node2061 = (inp[7]) ? node2063 : 1'b1;
														assign node2063 = (inp[9]) ? 1'b0 : 1'b1;
													assign node2066 = (inp[7]) ? node2070 : node2067;
														assign node2067 = (inp[9]) ? 1'b1 : 1'b0;
														assign node2070 = (inp[9]) ? 1'b0 : 1'b1;
									assign node2074 = (inp[15]) ? node2116 : node2075;
										assign node2075 = (inp[3]) ? node2099 : node2076;
											assign node2076 = (inp[12]) ? node2086 : node2077;
												assign node2077 = (inp[6]) ? node2079 : 1'b1;
													assign node2079 = (inp[5]) ? 1'b1 : node2080;
														assign node2080 = (inp[9]) ? node2082 : 1'b0;
															assign node2082 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2086 = (inp[10]) ? node2094 : node2087;
													assign node2087 = (inp[9]) ? 1'b1 : node2088;
														assign node2088 = (inp[6]) ? node2090 : 1'b0;
															assign node2090 = (inp[5]) ? 1'b0 : 1'b1;
													assign node2094 = (inp[5]) ? 1'b0 : node2095;
														assign node2095 = (inp[6]) ? 1'b1 : 1'b0;
											assign node2099 = (inp[7]) ? node2101 : 1'b1;
												assign node2101 = (inp[9]) ? node2109 : node2102;
													assign node2102 = (inp[6]) ? node2104 : 1'b0;
														assign node2104 = (inp[5]) ? 1'b1 : node2105;
															assign node2105 = (inp[12]) ? 1'b1 : 1'b0;
													assign node2109 = (inp[10]) ? node2111 : 1'b1;
														assign node2111 = (inp[12]) ? node2113 : 1'b1;
															assign node2113 = (inp[6]) ? 1'b1 : 1'b0;
										assign node2116 = (inp[6]) ? node2118 : 1'b1;
											assign node2118 = (inp[5]) ? 1'b1 : node2119;
												assign node2119 = (inp[9]) ? node2125 : node2120;
													assign node2120 = (inp[7]) ? 1'b0 : node2121;
														assign node2121 = (inp[3]) ? 1'b1 : 1'b0;
													assign node2125 = (inp[12]) ? 1'b1 : node2126;
														assign node2126 = (inp[3]) ? node2130 : node2127;
															assign node2127 = (inp[10]) ? 1'b0 : 1'b1;
															assign node2130 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2135 = (inp[6]) ? node2157 : node2136;
									assign node2136 = (inp[15]) ? 1'b0 : node2137;
										assign node2137 = (inp[12]) ? node2139 : 1'b0;
											assign node2139 = (inp[10]) ? node2151 : node2140;
												assign node2140 = (inp[3]) ? node2144 : node2141;
													assign node2141 = (inp[9]) ? 1'b0 : 1'b1;
													assign node2144 = (inp[9]) ? node2148 : node2145;
														assign node2145 = (inp[7]) ? 1'b1 : 1'b0;
														assign node2148 = (inp[5]) ? 1'b0 : 1'b1;
												assign node2151 = (inp[7]) ? 1'b1 : node2152;
													assign node2152 = (inp[3]) ? 1'b0 : 1'b1;
									assign node2157 = (inp[5]) ? node2193 : node2158;
										assign node2158 = (inp[15]) ? node2178 : node2159;
											assign node2159 = (inp[12]) ? 1'b0 : node2160;
												assign node2160 = (inp[7]) ? node2172 : node2161;
													assign node2161 = (inp[14]) ? node2167 : node2162;
														assign node2162 = (inp[3]) ? 1'b0 : node2163;
															assign node2163 = (inp[10]) ? 1'b1 : 1'b0;
														assign node2167 = (inp[3]) ? 1'b1 : node2168;
															assign node2168 = (inp[10]) ? 1'b1 : 1'b0;
													assign node2172 = (inp[9]) ? node2174 : 1'b1;
														assign node2174 = (inp[10]) ? 1'b1 : 1'b0;
											assign node2178 = (inp[9]) ? node2184 : node2179;
												assign node2179 = (inp[3]) ? node2181 : 1'b1;
													assign node2181 = (inp[12]) ? 1'b1 : 1'b0;
												assign node2184 = (inp[10]) ? node2188 : node2185;
													assign node2185 = (inp[3]) ? 1'b1 : 1'b0;
													assign node2188 = (inp[7]) ? 1'b1 : node2189;
														assign node2189 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2193 = (inp[12]) ? node2195 : 1'b0;
											assign node2195 = (inp[15]) ? 1'b0 : node2196;
												assign node2196 = (inp[10]) ? node2208 : node2197;
													assign node2197 = (inp[7]) ? 1'b0 : node2198;
														assign node2198 = (inp[14]) ? node2200 : 1'b1;
															assign node2200 = (inp[9]) ? node2204 : node2201;
																assign node2201 = (inp[3]) ? 1'b0 : 1'b1;
																assign node2204 = (inp[3]) ? 1'b1 : 1'b0;
													assign node2208 = (inp[3]) ? node2210 : 1'b1;
														assign node2210 = (inp[7]) ? 1'b1 : 1'b0;
		assign node2214 = (inp[1]) ? node2296 : node2215;
			assign node2215 = (inp[6]) ? node2237 : node2216;
				assign node2216 = (inp[15]) ? 1'b1 : node2217;
					assign node2217 = (inp[12]) ? node2219 : 1'b1;
						assign node2219 = (inp[3]) ? node2225 : node2220;
							assign node2220 = (inp[10]) ? 1'b0 : node2221;
								assign node2221 = (inp[9]) ? 1'b1 : 1'b0;
							assign node2225 = (inp[7]) ? node2231 : node2226;
								assign node2226 = (inp[9]) ? node2228 : 1'b1;
									assign node2228 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2231 = (inp[9]) ? node2233 : 1'b0;
									assign node2233 = (inp[10]) ? 1'b0 : 1'b1;
				assign node2237 = (inp[5]) ? node2275 : node2238;
					assign node2238 = (inp[12]) ? node2256 : node2239;
						assign node2239 = (inp[10]) ? node2251 : node2240;
							assign node2240 = (inp[9]) ? node2246 : node2241;
								assign node2241 = (inp[3]) ? node2243 : 1'b0;
									assign node2243 = (inp[7]) ? 1'b0 : 1'b1;
								assign node2246 = (inp[3]) ? node2248 : 1'b1;
									assign node2248 = (inp[7]) ? 1'b1 : 1'b0;
							assign node2251 = (inp[7]) ? 1'b0 : node2252;
								assign node2252 = (inp[3]) ? 1'b1 : 1'b0;
						assign node2256 = (inp[15]) ? node2258 : 1'b1;
							assign node2258 = (inp[10]) ? node2270 : node2259;
								assign node2259 = (inp[9]) ? node2265 : node2260;
									assign node2260 = (inp[7]) ? 1'b0 : node2261;
										assign node2261 = (inp[3]) ? 1'b1 : 1'b0;
									assign node2265 = (inp[7]) ? 1'b1 : node2266;
										assign node2266 = (inp[3]) ? 1'b0 : 1'b1;
								assign node2270 = (inp[3]) ? node2272 : 1'b0;
									assign node2272 = (inp[7]) ? 1'b0 : 1'b1;
					assign node2275 = (inp[15]) ? 1'b1 : node2276;
						assign node2276 = (inp[12]) ? node2278 : 1'b1;
							assign node2278 = (inp[7]) ? node2290 : node2279;
								assign node2279 = (inp[3]) ? node2285 : node2280;
									assign node2280 = (inp[9]) ? node2282 : 1'b0;
										assign node2282 = (inp[10]) ? 1'b0 : 1'b1;
									assign node2285 = (inp[9]) ? node2287 : 1'b1;
										assign node2287 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2290 = (inp[10]) ? 1'b0 : node2291;
									assign node2291 = (inp[9]) ? 1'b1 : 1'b0;
			assign node2296 = (inp[8]) ? node2982 : node2297;
				assign node2297 = (inp[11]) ? node2737 : node2298;
					assign node2298 = (inp[13]) ? node2516 : node2299;
						assign node2299 = (inp[2]) ? node2435 : node2300;
							assign node2300 = (inp[14]) ? node2372 : node2301;
								assign node2301 = (inp[15]) ? node2351 : node2302;
									assign node2302 = (inp[12]) ? node2320 : node2303;
										assign node2303 = (inp[5]) ? 1'b0 : node2304;
											assign node2304 = (inp[6]) ? node2306 : 1'b0;
												assign node2306 = (inp[3]) ? node2312 : node2307;
													assign node2307 = (inp[9]) ? node2309 : 1'b1;
														assign node2309 = (inp[10]) ? 1'b1 : 1'b0;
													assign node2312 = (inp[7]) ? node2314 : 1'b0;
														assign node2314 = (inp[9]) ? node2316 : 1'b1;
															assign node2316 = (inp[10]) ? 1'b1 : 1'b0;
										assign node2320 = (inp[6]) ? node2336 : node2321;
											assign node2321 = (inp[10]) ? node2331 : node2322;
												assign node2322 = (inp[3]) ? node2326 : node2323;
													assign node2323 = (inp[9]) ? 1'b0 : 1'b1;
													assign node2326 = (inp[5]) ? 1'b0 : node2327;
														assign node2327 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2331 = (inp[7]) ? 1'b1 : node2332;
													assign node2332 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2336 = (inp[5]) ? node2338 : 1'b0;
												assign node2338 = (inp[3]) ? node2340 : 1'b1;
													assign node2340 = (inp[7]) ? node2346 : node2341;
														assign node2341 = (inp[10]) ? 1'b0 : node2342;
															assign node2342 = (inp[9]) ? 1'b1 : 1'b0;
														assign node2346 = (inp[10]) ? 1'b1 : node2347;
															assign node2347 = (inp[0]) ? 1'b1 : 1'b0;
									assign node2351 = (inp[6]) ? node2353 : 1'b0;
										assign node2353 = (inp[5]) ? 1'b0 : node2354;
											assign node2354 = (inp[3]) ? node2360 : node2355;
												assign node2355 = (inp[10]) ? 1'b1 : node2356;
													assign node2356 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2360 = (inp[7]) ? node2366 : node2361;
													assign node2361 = (inp[10]) ? 1'b0 : node2362;
														assign node2362 = (inp[9]) ? 1'b1 : 1'b0;
													assign node2366 = (inp[9]) ? node2368 : 1'b1;
														assign node2368 = (inp[10]) ? 1'b1 : 1'b0;
								assign node2372 = (inp[12]) ? node2390 : node2373;
									assign node2373 = (inp[5]) ? 1'b1 : node2374;
										assign node2374 = (inp[6]) ? node2376 : 1'b1;
											assign node2376 = (inp[10]) ? node2384 : node2377;
												assign node2377 = (inp[9]) ? 1'b1 : node2378;
													assign node2378 = (inp[15]) ? node2380 : 1'b0;
														assign node2380 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2384 = (inp[3]) ? node2386 : 1'b0;
													assign node2386 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2390 = (inp[15]) ? node2416 : node2391;
										assign node2391 = (inp[7]) ? node2403 : node2392;
											assign node2392 = (inp[3]) ? node2396 : node2393;
												assign node2393 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2396 = (inp[10]) ? 1'b1 : node2397;
													assign node2397 = (inp[9]) ? node2399 : 1'b1;
														assign node2399 = (inp[0]) ? 1'b1 : 1'b0;
											assign node2403 = (inp[9]) ? node2409 : node2404;
												assign node2404 = (inp[5]) ? 1'b0 : node2405;
													assign node2405 = (inp[6]) ? 1'b1 : 1'b0;
												assign node2409 = (inp[10]) ? node2411 : 1'b1;
													assign node2411 = (inp[5]) ? 1'b0 : node2412;
														assign node2412 = (inp[6]) ? 1'b1 : 1'b0;
										assign node2416 = (inp[5]) ? 1'b1 : node2417;
											assign node2417 = (inp[6]) ? node2419 : 1'b1;
												assign node2419 = (inp[10]) ? node2429 : node2420;
													assign node2420 = (inp[9]) ? node2426 : node2421;
														assign node2421 = (inp[7]) ? 1'b0 : node2422;
															assign node2422 = (inp[3]) ? 1'b1 : 1'b0;
														assign node2426 = (inp[7]) ? 1'b1 : 1'b0;
													assign node2429 = (inp[7]) ? 1'b0 : node2430;
														assign node2430 = (inp[9]) ? 1'b0 : 1'b1;
							assign node2435 = (inp[15]) ? node2495 : node2436;
								assign node2436 = (inp[12]) ? node2458 : node2437;
									assign node2437 = (inp[6]) ? node2439 : 1'b0;
										assign node2439 = (inp[5]) ? 1'b0 : node2440;
											assign node2440 = (inp[7]) ? node2452 : node2441;
												assign node2441 = (inp[3]) ? node2447 : node2442;
													assign node2442 = (inp[9]) ? node2444 : 1'b1;
														assign node2444 = (inp[10]) ? 1'b1 : 1'b0;
													assign node2447 = (inp[9]) ? node2449 : 1'b0;
														assign node2449 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2452 = (inp[10]) ? 1'b1 : node2453;
													assign node2453 = (inp[9]) ? 1'b0 : 1'b1;
									assign node2458 = (inp[5]) ? node2478 : node2459;
										assign node2459 = (inp[6]) ? 1'b0 : node2460;
											assign node2460 = (inp[3]) ? node2466 : node2461;
												assign node2461 = (inp[9]) ? node2463 : 1'b1;
													assign node2463 = (inp[10]) ? 1'b1 : 1'b0;
												assign node2466 = (inp[7]) ? node2472 : node2467;
													assign node2467 = (inp[9]) ? node2469 : 1'b0;
														assign node2469 = (inp[10]) ? 1'b0 : 1'b1;
													assign node2472 = (inp[9]) ? node2474 : 1'b1;
														assign node2474 = (inp[10]) ? 1'b1 : 1'b0;
										assign node2478 = (inp[9]) ? node2484 : node2479;
											assign node2479 = (inp[7]) ? 1'b1 : node2480;
												assign node2480 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2484 = (inp[10]) ? node2490 : node2485;
												assign node2485 = (inp[7]) ? 1'b0 : node2486;
													assign node2486 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2490 = (inp[7]) ? 1'b1 : node2491;
													assign node2491 = (inp[3]) ? 1'b0 : 1'b1;
								assign node2495 = (inp[5]) ? 1'b0 : node2496;
									assign node2496 = (inp[6]) ? node2498 : 1'b0;
										assign node2498 = (inp[3]) ? node2504 : node2499;
											assign node2499 = (inp[10]) ? 1'b1 : node2500;
												assign node2500 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2504 = (inp[7]) ? node2510 : node2505;
												assign node2505 = (inp[10]) ? 1'b0 : node2506;
													assign node2506 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2510 = (inp[10]) ? 1'b1 : node2511;
													assign node2511 = (inp[9]) ? 1'b0 : 1'b1;
						assign node2516 = (inp[2]) ? node2660 : node2517;
							assign node2517 = (inp[14]) ? node2587 : node2518;
								assign node2518 = (inp[12]) ? node2536 : node2519;
									assign node2519 = (inp[6]) ? node2521 : 1'b1;
										assign node2521 = (inp[5]) ? 1'b1 : node2522;
											assign node2522 = (inp[7]) ? node2530 : node2523;
												assign node2523 = (inp[3]) ? 1'b1 : node2524;
													assign node2524 = (inp[10]) ? 1'b0 : node2525;
														assign node2525 = (inp[9]) ? 1'b1 : 1'b0;
												assign node2530 = (inp[10]) ? 1'b0 : node2531;
													assign node2531 = (inp[9]) ? 1'b1 : 1'b0;
									assign node2536 = (inp[15]) ? node2572 : node2537;
										assign node2537 = (inp[6]) ? node2555 : node2538;
											assign node2538 = (inp[9]) ? node2544 : node2539;
												assign node2539 = (inp[7]) ? 1'b0 : node2540;
													assign node2540 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2544 = (inp[10]) ? node2550 : node2545;
													assign node2545 = (inp[3]) ? node2547 : 1'b1;
														assign node2547 = (inp[7]) ? 1'b1 : 1'b0;
													assign node2550 = (inp[7]) ? 1'b0 : node2551;
														assign node2551 = (inp[3]) ? 1'b1 : 1'b0;
											assign node2555 = (inp[5]) ? node2557 : 1'b1;
												assign node2557 = (inp[9]) ? node2563 : node2558;
													assign node2558 = (inp[3]) ? node2560 : 1'b0;
														assign node2560 = (inp[0]) ? 1'b1 : 1'b0;
													assign node2563 = (inp[10]) ? node2567 : node2564;
														assign node2564 = (inp[3]) ? 1'b0 : 1'b1;
														assign node2567 = (inp[3]) ? node2569 : 1'b0;
															assign node2569 = (inp[7]) ? 1'b0 : 1'b1;
										assign node2572 = (inp[6]) ? node2574 : 1'b1;
											assign node2574 = (inp[5]) ? 1'b1 : node2575;
												assign node2575 = (inp[3]) ? node2579 : node2576;
													assign node2576 = (inp[9]) ? 1'b1 : 1'b0;
													assign node2579 = (inp[7]) ? node2581 : 1'b1;
														assign node2581 = (inp[10]) ? 1'b0 : node2582;
															assign node2582 = (inp[9]) ? 1'b1 : 1'b0;
								assign node2587 = (inp[6]) ? node2609 : node2588;
									assign node2588 = (inp[15]) ? 1'b0 : node2589;
										assign node2589 = (inp[12]) ? node2591 : 1'b0;
											assign node2591 = (inp[3]) ? node2597 : node2592;
												assign node2592 = (inp[9]) ? node2594 : 1'b1;
													assign node2594 = (inp[10]) ? 1'b1 : 1'b0;
												assign node2597 = (inp[7]) ? node2603 : node2598;
													assign node2598 = (inp[9]) ? node2600 : 1'b0;
														assign node2600 = (inp[10]) ? 1'b0 : 1'b1;
													assign node2603 = (inp[10]) ? 1'b1 : node2604;
														assign node2604 = (inp[9]) ? 1'b0 : 1'b1;
									assign node2609 = (inp[5]) ? node2639 : node2610;
										assign node2610 = (inp[15]) ? node2624 : node2611;
											assign node2611 = (inp[12]) ? 1'b0 : node2612;
												assign node2612 = (inp[10]) ? node2618 : node2613;
													assign node2613 = (inp[9]) ? 1'b0 : node2614;
														assign node2614 = (inp[3]) ? 1'b0 : 1'b1;
													assign node2618 = (inp[3]) ? node2620 : 1'b1;
														assign node2620 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2624 = (inp[10]) ? node2634 : node2625;
												assign node2625 = (inp[9]) ? node2629 : node2626;
													assign node2626 = (inp[3]) ? 1'b0 : 1'b1;
													assign node2629 = (inp[3]) ? node2631 : 1'b0;
														assign node2631 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2634 = (inp[7]) ? 1'b1 : node2635;
													assign node2635 = (inp[3]) ? 1'b0 : 1'b1;
										assign node2639 = (inp[12]) ? node2641 : 1'b0;
											assign node2641 = (inp[15]) ? 1'b0 : node2642;
												assign node2642 = (inp[9]) ? node2648 : node2643;
													assign node2643 = (inp[7]) ? 1'b1 : node2644;
														assign node2644 = (inp[3]) ? 1'b0 : 1'b1;
													assign node2648 = (inp[7]) ? node2656 : node2649;
														assign node2649 = (inp[3]) ? node2653 : node2650;
															assign node2650 = (inp[10]) ? 1'b1 : 1'b0;
															assign node2653 = (inp[10]) ? 1'b0 : 1'b1;
														assign node2656 = (inp[3]) ? 1'b1 : 1'b0;
							assign node2660 = (inp[15]) ? node2716 : node2661;
								assign node2661 = (inp[12]) ? node2683 : node2662;
									assign node2662 = (inp[6]) ? node2664 : 1'b1;
										assign node2664 = (inp[5]) ? 1'b1 : node2665;
											assign node2665 = (inp[9]) ? node2671 : node2666;
												assign node2666 = (inp[7]) ? 1'b0 : node2667;
													assign node2667 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2671 = (inp[10]) ? node2677 : node2672;
													assign node2672 = (inp[3]) ? node2674 : 1'b1;
														assign node2674 = (inp[7]) ? 1'b1 : 1'b0;
													assign node2677 = (inp[3]) ? node2679 : 1'b0;
														assign node2679 = (inp[7]) ? 1'b0 : 1'b1;
									assign node2683 = (inp[5]) ? node2699 : node2684;
										assign node2684 = (inp[6]) ? 1'b1 : node2685;
											assign node2685 = (inp[3]) ? node2691 : node2686;
												assign node2686 = (inp[9]) ? node2688 : 1'b0;
													assign node2688 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2691 = (inp[10]) ? 1'b1 : node2692;
													assign node2692 = (inp[7]) ? node2694 : 1'b0;
														assign node2694 = (inp[9]) ? 1'b1 : 1'b0;
										assign node2699 = (inp[10]) ? node2711 : node2700;
											assign node2700 = (inp[9]) ? node2706 : node2701;
												assign node2701 = (inp[3]) ? node2703 : 1'b0;
													assign node2703 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2706 = (inp[3]) ? node2708 : 1'b1;
													assign node2708 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2711 = (inp[3]) ? node2713 : 1'b0;
												assign node2713 = (inp[7]) ? 1'b0 : 1'b1;
								assign node2716 = (inp[5]) ? 1'b1 : node2717;
									assign node2717 = (inp[6]) ? node2719 : 1'b1;
										assign node2719 = (inp[10]) ? node2731 : node2720;
											assign node2720 = (inp[9]) ? node2726 : node2721;
												assign node2721 = (inp[7]) ? 1'b0 : node2722;
													assign node2722 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2726 = (inp[3]) ? node2728 : 1'b1;
													assign node2728 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2731 = (inp[7]) ? 1'b0 : node2732;
												assign node2732 = (inp[3]) ? 1'b1 : 1'b0;
					assign node2737 = (inp[2]) ? node2901 : node2738;
						assign node2738 = (inp[14]) ? node2820 : node2739;
							assign node2739 = (inp[12]) ? node2761 : node2740;
								assign node2740 = (inp[5]) ? 1'b0 : node2741;
									assign node2741 = (inp[6]) ? node2743 : 1'b0;
										assign node2743 = (inp[9]) ? node2749 : node2744;
											assign node2744 = (inp[7]) ? 1'b1 : node2745;
												assign node2745 = (inp[3]) ? 1'b0 : 1'b1;
											assign node2749 = (inp[10]) ? node2755 : node2750;
												assign node2750 = (inp[7]) ? 1'b0 : node2751;
													assign node2751 = (inp[3]) ? 1'b1 : 1'b0;
												assign node2755 = (inp[3]) ? node2757 : 1'b1;
													assign node2757 = (inp[7]) ? 1'b1 : 1'b0;
								assign node2761 = (inp[15]) ? node2797 : node2762;
									assign node2762 = (inp[7]) ? node2784 : node2763;
										assign node2763 = (inp[3]) ? node2777 : node2764;
											assign node2764 = (inp[9]) ? node2770 : node2765;
												assign node2765 = (inp[5]) ? 1'b1 : node2766;
													assign node2766 = (inp[6]) ? 1'b0 : 1'b1;
												assign node2770 = (inp[10]) ? node2772 : 1'b0;
													assign node2772 = (inp[6]) ? node2774 : 1'b1;
														assign node2774 = (inp[5]) ? 1'b1 : 1'b0;
											assign node2777 = (inp[10]) ? 1'b0 : node2778;
												assign node2778 = (inp[9]) ? node2780 : 1'b0;
													assign node2780 = (inp[6]) ? 1'b0 : 1'b1;
										assign node2784 = (inp[9]) ? node2790 : node2785;
											assign node2785 = (inp[5]) ? 1'b1 : node2786;
												assign node2786 = (inp[6]) ? 1'b0 : 1'b1;
											assign node2790 = (inp[10]) ? node2792 : 1'b0;
												assign node2792 = (inp[6]) ? node2794 : 1'b1;
													assign node2794 = (inp[5]) ? 1'b1 : 1'b0;
									assign node2797 = (inp[6]) ? node2799 : 1'b0;
										assign node2799 = (inp[5]) ? 1'b0 : node2800;
											assign node2800 = (inp[9]) ? node2806 : node2801;
												assign node2801 = (inp[3]) ? node2803 : 1'b1;
													assign node2803 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2806 = (inp[13]) ? node2812 : node2807;
													assign node2807 = (inp[3]) ? 1'b1 : node2808;
														assign node2808 = (inp[7]) ? 1'b1 : 1'b0;
													assign node2812 = (inp[10]) ? node2814 : 1'b0;
														assign node2814 = (inp[7]) ? 1'b1 : node2815;
															assign node2815 = (inp[3]) ? 1'b0 : 1'b1;
							assign node2820 = (inp[15]) ? node2880 : node2821;
								assign node2821 = (inp[12]) ? node2843 : node2822;
									assign node2822 = (inp[5]) ? 1'b1 : node2823;
										assign node2823 = (inp[6]) ? node2825 : 1'b1;
											assign node2825 = (inp[9]) ? node2831 : node2826;
												assign node2826 = (inp[3]) ? node2828 : 1'b0;
													assign node2828 = (inp[7]) ? 1'b0 : 1'b1;
												assign node2831 = (inp[10]) ? node2837 : node2832;
													assign node2832 = (inp[3]) ? node2834 : 1'b1;
														assign node2834 = (inp[7]) ? 1'b1 : 1'b0;
													assign node2837 = (inp[7]) ? 1'b0 : node2838;
														assign node2838 = (inp[3]) ? 1'b1 : 1'b0;
									assign node2843 = (inp[5]) ? node2863 : node2844;
										assign node2844 = (inp[6]) ? 1'b1 : node2845;
											assign node2845 = (inp[7]) ? node2857 : node2846;
												assign node2846 = (inp[3]) ? node2852 : node2847;
													assign node2847 = (inp[10]) ? 1'b0 : node2848;
														assign node2848 = (inp[13]) ? 1'b0 : 1'b1;
													assign node2852 = (inp[9]) ? node2854 : 1'b1;
														assign node2854 = (inp[10]) ? 1'b1 : 1'b0;
												assign node2857 = (inp[9]) ? node2859 : 1'b0;
													assign node2859 = (inp[10]) ? 1'b0 : 1'b1;
										assign node2863 = (inp[9]) ? node2869 : node2864;
											assign node2864 = (inp[7]) ? 1'b0 : node2865;
												assign node2865 = (inp[3]) ? 1'b1 : 1'b0;
											assign node2869 = (inp[10]) ? node2875 : node2870;
												assign node2870 = (inp[3]) ? node2872 : 1'b1;
													assign node2872 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2875 = (inp[7]) ? 1'b0 : node2876;
													assign node2876 = (inp[3]) ? 1'b1 : 1'b0;
								assign node2880 = (inp[6]) ? node2882 : 1'b1;
									assign node2882 = (inp[5]) ? 1'b1 : node2883;
										assign node2883 = (inp[7]) ? node2895 : node2884;
											assign node2884 = (inp[3]) ? node2890 : node2885;
												assign node2885 = (inp[9]) ? node2887 : 1'b0;
													assign node2887 = (inp[10]) ? 1'b0 : 1'b1;
												assign node2890 = (inp[10]) ? 1'b1 : node2891;
													assign node2891 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2895 = (inp[9]) ? node2897 : 1'b0;
												assign node2897 = (inp[10]) ? 1'b0 : 1'b1;
						assign node2901 = (inp[5]) ? node2961 : node2902;
							assign node2902 = (inp[6]) ? node2924 : node2903;
								assign node2903 = (inp[15]) ? 1'b0 : node2904;
									assign node2904 = (inp[12]) ? node2906 : 1'b0;
										assign node2906 = (inp[10]) ? node2918 : node2907;
											assign node2907 = (inp[9]) ? node2913 : node2908;
												assign node2908 = (inp[3]) ? node2910 : 1'b1;
													assign node2910 = (inp[7]) ? 1'b1 : 1'b0;
												assign node2913 = (inp[7]) ? 1'b0 : node2914;
													assign node2914 = (inp[3]) ? 1'b1 : 1'b0;
											assign node2918 = (inp[3]) ? node2920 : 1'b1;
												assign node2920 = (inp[7]) ? 1'b1 : 1'b0;
								assign node2924 = (inp[15]) ? node2944 : node2925;
									assign node2925 = (inp[12]) ? 1'b0 : node2926;
										assign node2926 = (inp[7]) ? node2938 : node2927;
											assign node2927 = (inp[3]) ? node2933 : node2928;
												assign node2928 = (inp[10]) ? 1'b1 : node2929;
													assign node2929 = (inp[9]) ? 1'b0 : 1'b1;
												assign node2933 = (inp[10]) ? 1'b0 : node2934;
													assign node2934 = (inp[9]) ? 1'b1 : 1'b0;
											assign node2938 = (inp[9]) ? node2940 : 1'b1;
												assign node2940 = (inp[10]) ? 1'b1 : 1'b0;
									assign node2944 = (inp[10]) ? node2956 : node2945;
										assign node2945 = (inp[9]) ? node2951 : node2946;
											assign node2946 = (inp[3]) ? node2948 : 1'b1;
												assign node2948 = (inp[7]) ? 1'b1 : 1'b0;
											assign node2951 = (inp[7]) ? 1'b0 : node2952;
												assign node2952 = (inp[3]) ? 1'b1 : 1'b0;
										assign node2956 = (inp[7]) ? 1'b1 : node2957;
											assign node2957 = (inp[3]) ? 1'b0 : 1'b1;
							assign node2961 = (inp[12]) ? node2963 : 1'b0;
								assign node2963 = (inp[15]) ? 1'b0 : node2964;
									assign node2964 = (inp[7]) ? node2976 : node2965;
										assign node2965 = (inp[3]) ? node2971 : node2966;
											assign node2966 = (inp[10]) ? 1'b1 : node2967;
												assign node2967 = (inp[9]) ? 1'b0 : 1'b1;
											assign node2971 = (inp[10]) ? 1'b0 : node2972;
												assign node2972 = (inp[9]) ? 1'b1 : 1'b0;
										assign node2976 = (inp[10]) ? 1'b1 : node2977;
											assign node2977 = (inp[9]) ? 1'b0 : 1'b1;
				assign node2982 = (inp[12]) ? node3004 : node2983;
					assign node2983 = (inp[6]) ? node2985 : 1'b1;
						assign node2985 = (inp[5]) ? 1'b1 : node2986;
							assign node2986 = (inp[9]) ? node2992 : node2987;
								assign node2987 = (inp[3]) ? node2989 : 1'b0;
									assign node2989 = (inp[7]) ? 1'b0 : 1'b1;
								assign node2992 = (inp[10]) ? node2998 : node2993;
									assign node2993 = (inp[3]) ? node2995 : 1'b1;
										assign node2995 = (inp[7]) ? 1'b1 : 1'b0;
									assign node2998 = (inp[3]) ? node3000 : 1'b0;
										assign node3000 = (inp[7]) ? 1'b0 : 1'b1;
					assign node3004 = (inp[15]) ? node3042 : node3005;
						assign node3005 = (inp[6]) ? node3023 : node3006;
							assign node3006 = (inp[10]) ? node3018 : node3007;
								assign node3007 = (inp[9]) ? node3013 : node3008;
									assign node3008 = (inp[3]) ? node3010 : 1'b0;
										assign node3010 = (inp[7]) ? 1'b0 : 1'b1;
									assign node3013 = (inp[3]) ? node3015 : 1'b1;
										assign node3015 = (inp[7]) ? 1'b1 : 1'b0;
								assign node3018 = (inp[3]) ? node3020 : 1'b0;
									assign node3020 = (inp[7]) ? 1'b0 : 1'b1;
							assign node3023 = (inp[5]) ? node3025 : 1'b1;
								assign node3025 = (inp[10]) ? node3037 : node3026;
									assign node3026 = (inp[9]) ? node3032 : node3027;
										assign node3027 = (inp[7]) ? 1'b0 : node3028;
											assign node3028 = (inp[3]) ? 1'b1 : 1'b0;
										assign node3032 = (inp[7]) ? 1'b1 : node3033;
											assign node3033 = (inp[3]) ? 1'b0 : 1'b1;
									assign node3037 = (inp[3]) ? node3039 : 1'b0;
										assign node3039 = (inp[7]) ? 1'b0 : 1'b1;
						assign node3042 = (inp[6]) ? node3044 : 1'b1;
							assign node3044 = (inp[5]) ? 1'b1 : node3045;
								assign node3045 = (inp[9]) ? node3051 : node3046;
									assign node3046 = (inp[3]) ? node3048 : 1'b0;
										assign node3048 = (inp[7]) ? 1'b0 : 1'b1;
									assign node3051 = (inp[10]) ? node3057 : node3052;
										assign node3052 = (inp[3]) ? node3054 : 1'b1;
											assign node3054 = (inp[7]) ? 1'b1 : 1'b0;
										assign node3057 = (inp[3]) ? node3059 : 1'b0;
											assign node3059 = (inp[7]) ? 1'b0 : 1'b1;

endmodule