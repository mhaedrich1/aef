module dtc_split33_bm50 (
	input  wire [8-1:0] inp,
	output wire [2-1:0] outp
);

	wire [2-1:0] node1;
	wire [2-1:0] node2;
	wire [2-1:0] node3;
	wire [2-1:0] node4;
	wire [2-1:0] node5;
	wire [2-1:0] node8;
	wire [2-1:0] node10;
	wire [2-1:0] node13;
	wire [2-1:0] node15;
	wire [2-1:0] node16;
	wire [2-1:0] node19;
	wire [2-1:0] node22;
	wire [2-1:0] node23;
	wire [2-1:0] node24;
	wire [2-1:0] node26;
	wire [2-1:0] node30;
	wire [2-1:0] node31;
	wire [2-1:0] node32;
	wire [2-1:0] node33;
	wire [2-1:0] node38;
	wire [2-1:0] node41;
	wire [2-1:0] node42;
	wire [2-1:0] node43;
	wire [2-1:0] node44;
	wire [2-1:0] node45;
	wire [2-1:0] node48;
	wire [2-1:0] node52;
	wire [2-1:0] node53;
	wire [2-1:0] node57;
	wire [2-1:0] node58;
	wire [2-1:0] node59;
	wire [2-1:0] node61;
	wire [2-1:0] node63;
	wire [2-1:0] node66;
	wire [2-1:0] node69;
	wire [2-1:0] node70;
	wire [2-1:0] node73;
	wire [2-1:0] node75;
	wire [2-1:0] node76;
	wire [2-1:0] node79;
	wire [2-1:0] node82;
	wire [2-1:0] node83;
	wire [2-1:0] node84;
	wire [2-1:0] node85;
	wire [2-1:0] node87;
	wire [2-1:0] node91;
	wire [2-1:0] node92;
	wire [2-1:0] node94;
	wire [2-1:0] node97;
	wire [2-1:0] node99;
	wire [2-1:0] node101;
	wire [2-1:0] node104;
	wire [2-1:0] node105;
	wire [2-1:0] node106;
	wire [2-1:0] node108;
	wire [2-1:0] node111;
	wire [2-1:0] node113;
	wire [2-1:0] node116;
	wire [2-1:0] node117;
	wire [2-1:0] node118;
	wire [2-1:0] node122;
	wire [2-1:0] node124;

	assign outp = (inp[2]) ? node82 : node1;
		assign node1 = (inp[3]) ? node41 : node2;
			assign node2 = (inp[0]) ? node22 : node3;
				assign node3 = (inp[6]) ? node13 : node4;
					assign node4 = (inp[7]) ? node8 : node5;
						assign node5 = (inp[5]) ? 2'b01 : 2'b11;
						assign node8 = (inp[5]) ? node10 : 2'b10;
							assign node10 = (inp[1]) ? 2'b10 : 2'b00;
					assign node13 = (inp[4]) ? node15 : 2'b10;
						assign node15 = (inp[1]) ? node19 : node16;
							assign node16 = (inp[5]) ? 2'b00 : 2'b10;
							assign node19 = (inp[5]) ? 2'b10 : 2'b00;
				assign node22 = (inp[7]) ? node30 : node23;
					assign node23 = (inp[6]) ? 2'b11 : node24;
						assign node24 = (inp[5]) ? node26 : 2'b10;
							assign node26 = (inp[1]) ? 2'b10 : 2'b00;
					assign node30 = (inp[6]) ? node38 : node31;
						assign node31 = (inp[1]) ? 2'b01 : node32;
							assign node32 = (inp[4]) ? 2'b11 : node33;
								assign node33 = (inp[5]) ? 2'b01 : 2'b11;
						assign node38 = (inp[1]) ? 2'b00 : 2'b10;
			assign node41 = (inp[1]) ? node57 : node42;
				assign node42 = (inp[0]) ? node52 : node43;
					assign node43 = (inp[5]) ? 2'b11 : node44;
						assign node44 = (inp[4]) ? node48 : node45;
							assign node45 = (inp[6]) ? 2'b01 : 2'b11;
							assign node48 = (inp[7]) ? 2'b00 : 2'b01;
					assign node52 = (inp[6]) ? 2'b00 : node53;
						assign node53 = (inp[7]) ? 2'b01 : 2'b00;
				assign node57 = (inp[5]) ? node69 : node58;
					assign node58 = (inp[4]) ? node66 : node59;
						assign node59 = (inp[6]) ? node61 : 2'b00;
							assign node61 = (inp[0]) ? node63 : 2'b00;
								assign node63 = (inp[7]) ? 2'b10 : 2'b11;
						assign node66 = (inp[6]) ? 2'b10 : 2'b11;
					assign node69 = (inp[6]) ? node73 : node70;
						assign node70 = (inp[7]) ? 2'b00 : 2'b10;
						assign node73 = (inp[4]) ? node75 : 2'b01;
							assign node75 = (inp[7]) ? node79 : node76;
								assign node76 = (inp[0]) ? 2'b01 : 2'b00;
								assign node79 = (inp[0]) ? 2'b00 : 2'b01;
		assign node82 = (inp[0]) ? node104 : node83;
			assign node83 = (inp[7]) ? node91 : node84;
				assign node84 = (inp[3]) ? 2'b00 : node85;
					assign node85 = (inp[5]) ? node87 : 2'b10;
						assign node87 = (inp[1]) ? 2'b10 : 2'b00;
				assign node91 = (inp[6]) ? node97 : node92;
					assign node92 = (inp[4]) ? node94 : 2'b01;
						assign node94 = (inp[3]) ? 2'b11 : 2'b01;
					assign node97 = (inp[1]) ? node99 : 2'b11;
						assign node99 = (inp[5]) ? node101 : 2'b11;
							assign node101 = (inp[3]) ? 2'b01 : 2'b11;
			assign node104 = (inp[7]) ? node116 : node105;
				assign node105 = (inp[3]) ? node111 : node106;
					assign node106 = (inp[1]) ? node108 : 2'b01;
						assign node108 = (inp[4]) ? 2'b11 : 2'b01;
					assign node111 = (inp[1]) ? node113 : 2'b11;
						assign node113 = (inp[5]) ? 2'b01 : 2'b11;
				assign node116 = (inp[3]) ? node122 : node117;
					assign node117 = (inp[4]) ? 2'b00 : node118;
						assign node118 = (inp[5]) ? 2'b10 : 2'b00;
					assign node122 = (inp[1]) ? node124 : 2'b10;
						assign node124 = (inp[5]) ? 2'b00 : 2'b10;

endmodule