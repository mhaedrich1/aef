module dtc_split125_bm48 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node9;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node15;
	wire [14-1:0] node19;
	wire [14-1:0] node20;
	wire [14-1:0] node22;
	wire [14-1:0] node23;
	wire [14-1:0] node25;
	wire [14-1:0] node26;
	wire [14-1:0] node31;
	wire [14-1:0] node32;
	wire [14-1:0] node34;
	wire [14-1:0] node35;
	wire [14-1:0] node36;
	wire [14-1:0] node41;
	wire [14-1:0] node42;
	wire [14-1:0] node43;
	wire [14-1:0] node45;
	wire [14-1:0] node49;
	wire [14-1:0] node50;
	wire [14-1:0] node51;
	wire [14-1:0] node55;
	wire [14-1:0] node58;
	wire [14-1:0] node59;
	wire [14-1:0] node61;
	wire [14-1:0] node62;
	wire [14-1:0] node64;
	wire [14-1:0] node66;
	wire [14-1:0] node67;
	wire [14-1:0] node70;
	wire [14-1:0] node73;
	wire [14-1:0] node74;
	wire [14-1:0] node75;
	wire [14-1:0] node79;
	wire [14-1:0] node80;
	wire [14-1:0] node81;
	wire [14-1:0] node86;
	wire [14-1:0] node87;
	wire [14-1:0] node88;
	wire [14-1:0] node90;
	wire [14-1:0] node91;
	wire [14-1:0] node96;
	wire [14-1:0] node97;
	wire [14-1:0] node99;
	wire [14-1:0] node100;
	wire [14-1:0] node104;
	wire [14-1:0] node105;
	wire [14-1:0] node106;
	wire [14-1:0] node109;
	wire [14-1:0] node112;
	wire [14-1:0] node114;
	wire [14-1:0] node116;
	wire [14-1:0] node119;
	wire [14-1:0] node120;
	wire [14-1:0] node121;
	wire [14-1:0] node122;
	wire [14-1:0] node123;
	wire [14-1:0] node125;
	wire [14-1:0] node126;
	wire [14-1:0] node127;
	wire [14-1:0] node130;
	wire [14-1:0] node135;
	wire [14-1:0] node136;
	wire [14-1:0] node138;
	wire [14-1:0] node139;
	wire [14-1:0] node140;
	wire [14-1:0] node145;
	wire [14-1:0] node146;
	wire [14-1:0] node147;
	wire [14-1:0] node149;
	wire [14-1:0] node152;
	wire [14-1:0] node153;
	wire [14-1:0] node156;
	wire [14-1:0] node159;
	wire [14-1:0] node161;
	wire [14-1:0] node162;
	wire [14-1:0] node165;
	wire [14-1:0] node168;
	wire [14-1:0] node169;
	wire [14-1:0] node170;
	wire [14-1:0] node171;
	wire [14-1:0] node172;
	wire [14-1:0] node173;
	wire [14-1:0] node176;
	wire [14-1:0] node179;
	wire [14-1:0] node180;
	wire [14-1:0] node186;
	wire [14-1:0] node188;
	wire [14-1:0] node190;
	wire [14-1:0] node191;
	wire [14-1:0] node193;
	wire [14-1:0] node197;
	wire [14-1:0] node198;
	wire [14-1:0] node199;
	wire [14-1:0] node201;
	wire [14-1:0] node202;
	wire [14-1:0] node204;
	wire [14-1:0] node206;
	wire [14-1:0] node209;
	wire [14-1:0] node210;
	wire [14-1:0] node212;
	wire [14-1:0] node215;
	wire [14-1:0] node217;
	wire [14-1:0] node221;
	wire [14-1:0] node222;
	wire [14-1:0] node223;
	wire [14-1:0] node224;
	wire [14-1:0] node225;
	wire [14-1:0] node226;
	wire [14-1:0] node232;
	wire [14-1:0] node233;
	wire [14-1:0] node235;
	wire [14-1:0] node236;
	wire [14-1:0] node240;
	wire [14-1:0] node241;
	wire [14-1:0] node244;
	wire [14-1:0] node246;
	wire [14-1:0] node250;
	wire [14-1:0] node251;
	wire [14-1:0] node252;
	wire [14-1:0] node253;
	wire [14-1:0] node255;
	wire [14-1:0] node256;
	wire [14-1:0] node257;
	wire [14-1:0] node259;
	wire [14-1:0] node260;
	wire [14-1:0] node266;
	wire [14-1:0] node267;
	wire [14-1:0] node268;
	wire [14-1:0] node270;
	wire [14-1:0] node271;
	wire [14-1:0] node272;
	wire [14-1:0] node278;
	wire [14-1:0] node280;
	wire [14-1:0] node282;
	wire [14-1:0] node284;
	wire [14-1:0] node285;
	wire [14-1:0] node289;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node292;
	wire [14-1:0] node293;
	wire [14-1:0] node294;
	wire [14-1:0] node296;
	wire [14-1:0] node299;
	wire [14-1:0] node301;
	wire [14-1:0] node304;
	wire [14-1:0] node306;
	wire [14-1:0] node307;
	wire [14-1:0] node311;
	wire [14-1:0] node313;
	wire [14-1:0] node315;
	wire [14-1:0] node317;
	wire [14-1:0] node320;
	wire [14-1:0] node322;
	wire [14-1:0] node324;
	wire [14-1:0] node325;
	wire [14-1:0] node327;
	wire [14-1:0] node331;
	wire [14-1:0] node332;
	wire [14-1:0] node333;
	wire [14-1:0] node334;
	wire [14-1:0] node335;
	wire [14-1:0] node337;
	wire [14-1:0] node344;
	wire [14-1:0] node345;
	wire [14-1:0] node346;
	wire [14-1:0] node348;
	wire [14-1:0] node350;
	wire [14-1:0] node352;
	wire [14-1:0] node354;
	wire [14-1:0] node357;
	wire [14-1:0] node358;
	wire [14-1:0] node359;
	wire [14-1:0] node360;
	wire [14-1:0] node361;
	wire [14-1:0] node362;
	wire [14-1:0] node365;
	wire [14-1:0] node368;
	wire [14-1:0] node369;
	wire [14-1:0] node373;
	wire [14-1:0] node374;
	wire [14-1:0] node376;
	wire [14-1:0] node381;
	wire [14-1:0] node382;
	wire [14-1:0] node383;
	wire [14-1:0] node384;
	wire [14-1:0] node388;
	wire [14-1:0] node389;
	wire [14-1:0] node391;
	wire [14-1:0] node395;
	wire [14-1:0] node396;
	wire [14-1:0] node397;
	wire [14-1:0] node398;
	wire [14-1:0] node402;
	wire [14-1:0] node406;
	wire [14-1:0] node407;
	wire [14-1:0] node409;
	wire [14-1:0] node410;
	wire [14-1:0] node411;
	wire [14-1:0] node412;
	wire [14-1:0] node413;
	wire [14-1:0] node419;
	wire [14-1:0] node420;
	wire [14-1:0] node421;
	wire [14-1:0] node424;
	wire [14-1:0] node425;
	wire [14-1:0] node428;
	wire [14-1:0] node431;
	wire [14-1:0] node433;
	wire [14-1:0] node436;
	wire [14-1:0] node437;
	wire [14-1:0] node438;
	wire [14-1:0] node440;
	wire [14-1:0] node441;

	assign outp = (inp[10]) ? node250 : node1;
		assign node1 = (inp[13]) ? node119 : node2;
			assign node2 = (inp[11]) ? node58 : node3;
				assign node3 = (inp[12]) ? node19 : node4;
					assign node4 = (inp[8]) ? node6 : 14'b00000100000011;
						assign node6 = (inp[4]) ? 14'b00000000000000 : node7;
							assign node7 = (inp[1]) ? node9 : 14'b00000000000000;
								assign node9 = (inp[5]) ? node11 : 14'b00000000000000;
									assign node11 = (inp[3]) ? node15 : node12;
										assign node12 = (inp[0]) ? 14'b10000000011010 : 14'b00000000000000;
										assign node15 = (inp[2]) ? 14'b00000000000000 : 14'b10100100111000;
					assign node19 = (inp[6]) ? node31 : node20;
						assign node20 = (inp[9]) ? node22 : 14'b00000000000000;
							assign node22 = (inp[0]) ? 14'b00000000000000 : node23;
								assign node23 = (inp[1]) ? node25 : 14'b00000000000000;
									assign node25 = (inp[7]) ? 14'b00000000000000 : node26;
										assign node26 = (inp[3]) ? 14'b00001000000101 : 14'b00000000000000;
						assign node31 = (inp[8]) ? node41 : node32;
							assign node32 = (inp[4]) ? node34 : 14'b00000000000000;
								assign node34 = (inp[2]) ? 14'b00000000000000 : node35;
									assign node35 = (inp[7]) ? 14'b00000000000000 : node36;
										assign node36 = (inp[0]) ? 14'b00000000000000 : 14'b00100000000011;
							assign node41 = (inp[3]) ? node49 : node42;
								assign node42 = (inp[2]) ? 14'b00000000000000 : node43;
									assign node43 = (inp[1]) ? node45 : 14'b00000000000000;
										assign node45 = (inp[4]) ? 14'b10100100111111 : 14'b00000000000000;
								assign node49 = (inp[4]) ? node55 : node50;
									assign node50 = (inp[7]) ? 14'b00000000000000 : node51;
										assign node51 = (inp[9]) ? 14'b11110111110010 : 14'b00000000000000;
									assign node55 = (inp[1]) ? 14'b00000000000000 : 14'b11110111110010;
				assign node58 = (inp[12]) ? node86 : node59;
					assign node59 = (inp[1]) ? node61 : 14'b00000000000000;
						assign node61 = (inp[8]) ? node73 : node62;
							assign node62 = (inp[7]) ? node64 : 14'b00000000000000;
								assign node64 = (inp[9]) ? node66 : 14'b00000000000000;
									assign node66 = (inp[0]) ? node70 : node67;
										assign node67 = (inp[6]) ? 14'b00000000000000 : 14'b10010000001101;
										assign node70 = (inp[2]) ? 14'b01001000000100 : 14'b00000000000000;
							assign node73 = (inp[6]) ? node79 : node74;
								assign node74 = (inp[9]) ? 14'b00000000000000 : node75;
									assign node75 = (inp[3]) ? 14'b00000000000000 : 14'b01001000000100;
								assign node79 = (inp[5]) ? 14'b00000000000000 : node80;
									assign node80 = (inp[4]) ? 14'b00000000000000 : node81;
										assign node81 = (inp[9]) ? 14'b01100000001010 : 14'b00000000000000;
					assign node86 = (inp[6]) ? node96 : node87;
						assign node87 = (inp[3]) ? 14'b00000000000000 : node88;
							assign node88 = (inp[1]) ? node90 : 14'b00000000000000;
								assign node90 = (inp[9]) ? 14'b00000000000000 : node91;
									assign node91 = (inp[8]) ? 14'b00100100011111 : 14'b10000100011000;
						assign node96 = (inp[3]) ? node104 : node97;
							assign node97 = (inp[1]) ? node99 : 14'b00000000000000;
								assign node99 = (inp[9]) ? 14'b00000000000000 : node100;
									assign node100 = (inp[8]) ? 14'b01000100000100 : 14'b00000000000000;
							assign node104 = (inp[1]) ? node112 : node105;
								assign node105 = (inp[9]) ? node109 : node106;
									assign node106 = (inp[8]) ? 14'b00000000000000 : 14'b01100000001010;
									assign node109 = (inp[8]) ? 14'b10100010001100 : 14'b00000000000000;
								assign node112 = (inp[5]) ? node114 : 14'b00000000000000;
									assign node114 = (inp[9]) ? node116 : 14'b00000000000000;
										assign node116 = (inp[7]) ? 14'b00000000000000 : 14'b01001000001100;
			assign node119 = (inp[8]) ? node197 : node120;
				assign node120 = (inp[2]) ? node168 : node121;
					assign node121 = (inp[3]) ? node135 : node122;
						assign node122 = (inp[9]) ? 14'b00000000000000 : node123;
							assign node123 = (inp[1]) ? node125 : 14'b00000000000000;
								assign node125 = (inp[6]) ? 14'b00000000000000 : node126;
									assign node126 = (inp[11]) ? node130 : node127;
										assign node127 = (inp[12]) ? 14'b00000000000000 : 14'b11000000000100;
										assign node130 = (inp[0]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node135 = (inp[7]) ? node145 : node136;
							assign node136 = (inp[6]) ? node138 : 14'b00000000000000;
								assign node138 = (inp[11]) ? 14'b00000000000000 : node139;
									assign node139 = (inp[9]) ? 14'b00000000000000 : node140;
										assign node140 = (inp[1]) ? 14'b00000000000000 : 14'b11000000000100;
							assign node145 = (inp[6]) ? node159 : node146;
								assign node146 = (inp[9]) ? node152 : node147;
									assign node147 = (inp[1]) ? node149 : 14'b00000000000000;
										assign node149 = (inp[0]) ? 14'b00000000000000 : 14'b10000100111010;
									assign node152 = (inp[11]) ? node156 : node153;
										assign node153 = (inp[12]) ? 14'b11110111110010 : 14'b00000000000000;
										assign node156 = (inp[0]) ? 14'b00000000000000 : 14'b10100010001100;
								assign node159 = (inp[4]) ? node161 : 14'b00000000000000;
									assign node161 = (inp[0]) ? node165 : node162;
										assign node162 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
										assign node165 = (inp[12]) ? 14'b00000000000000 : 14'b01000000000100;
					assign node168 = (inp[12]) ? node186 : node169;
						assign node169 = (inp[11]) ? 14'b00000000000000 : node170;
							assign node170 = (inp[9]) ? 14'b00000000000000 : node171;
								assign node171 = (inp[7]) ? node179 : node172;
									assign node172 = (inp[4]) ? node176 : node173;
										assign node173 = (inp[1]) ? 14'b11000000000100 : 14'b00000000000000;
										assign node176 = (inp[1]) ? 14'b00000000000000 : 14'b00000000000000;
									assign node179 = (inp[6]) ? 14'b00000000000000 : node180;
										assign node180 = (inp[3]) ? 14'b00000000000000 : 14'b11000000000100;
						assign node186 = (inp[0]) ? node188 : 14'b00000000000000;
							assign node188 = (inp[7]) ? node190 : 14'b00000000000000;
								assign node190 = (inp[1]) ? 14'b00000000000000 : node191;
									assign node191 = (inp[3]) ? node193 : 14'b00000000000000;
										assign node193 = (inp[5]) ? 14'b00000000000000 : 14'b00100100001101;
				assign node197 = (inp[12]) ? node221 : node198;
					assign node198 = (inp[0]) ? 14'b00000000000000 : node199;
						assign node199 = (inp[1]) ? node201 : 14'b00000000000000;
							assign node201 = (inp[11]) ? node209 : node202;
								assign node202 = (inp[9]) ? node204 : 14'b00000000000000;
									assign node204 = (inp[3]) ? node206 : 14'b00000000000000;
										assign node206 = (inp[5]) ? 14'b00000000000000 : 14'b00000000011100;
								assign node209 = (inp[9]) ? node215 : node210;
									assign node210 = (inp[3]) ? node212 : 14'b00000000011100;
										assign node212 = (inp[2]) ? 14'b00000000000000 : 14'b00000000011100;
									assign node215 = (inp[3]) ? node217 : 14'b00000000000000;
										assign node217 = (inp[7]) ? 14'b10100010001100 : 14'b00000000000000;
					assign node221 = (inp[11]) ? 14'b01000000010100 : node222;
						assign node222 = (inp[6]) ? node232 : node223;
							assign node223 = (inp[2]) ? 14'b00000000000000 : node224;
								assign node224 = (inp[3]) ? 14'b00000000000000 : node225;
									assign node225 = (inp[0]) ? 14'b00000000000000 : node226;
										assign node226 = (inp[4]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node232 = (inp[9]) ? node240 : node233;
								assign node233 = (inp[1]) ? node235 : 14'b00000000000000;
									assign node235 = (inp[3]) ? 14'b00000000000000 : node236;
										assign node236 = (inp[7]) ? 14'b11100100010100 : 14'b10010100011100;
								assign node240 = (inp[1]) ? node244 : node241;
									assign node241 = (inp[3]) ? 14'b01001000000100 : 14'b00000000000000;
									assign node244 = (inp[7]) ? node246 : 14'b00000000000000;
										assign node246 = (inp[5]) ? 14'b01001000001001 : 14'b00000000000000;
		assign node250 = (inp[13]) ? node344 : node251;
			assign node251 = (inp[12]) ? node289 : node252;
				assign node252 = (inp[11]) ? node266 : node253;
					assign node253 = (inp[8]) ? node255 : 14'b10000100001000;
						assign node255 = (inp[3]) ? 14'b00000000000000 : node256;
							assign node256 = (inp[0]) ? 14'b00000000000000 : node257;
								assign node257 = (inp[2]) ? node259 : 14'b00000000000000;
									assign node259 = (inp[9]) ? 14'b00000000000000 : node260;
										assign node260 = (inp[5]) ? 14'b00000000000000 : 14'b00100000000011;
					assign node266 = (inp[4]) ? node278 : node267;
						assign node267 = (inp[2]) ? 14'b00000000000000 : node268;
							assign node268 = (inp[1]) ? node270 : 14'b00000000000000;
								assign node270 = (inp[6]) ? 14'b00000000000000 : node271;
									assign node271 = (inp[7]) ? 14'b10100000001101 : node272;
										assign node272 = (inp[0]) ? 14'b00000000000000 : 14'b00100000000011;
						assign node278 = (inp[1]) ? node280 : 14'b00000000000000;
							assign node280 = (inp[8]) ? node282 : 14'b00000000000000;
								assign node282 = (inp[3]) ? node284 : 14'b00000000000000;
									assign node284 = (inp[5]) ? 14'b00000000000000 : node285;
										assign node285 = (inp[6]) ? 14'b01001000000100 : 14'b00000000000000;
				assign node289 = (inp[11]) ? node331 : node290;
					assign node290 = (inp[2]) ? node320 : node291;
						assign node291 = (inp[0]) ? node311 : node292;
							assign node292 = (inp[7]) ? node304 : node293;
								assign node293 = (inp[3]) ? node299 : node294;
									assign node294 = (inp[4]) ? node296 : 14'b00000000000000;
										assign node296 = (inp[8]) ? 14'b00000000000000 : 14'b00000000000000;
									assign node299 = (inp[1]) ? node301 : 14'b10100100101000;
										assign node301 = (inp[8]) ? 14'b00000000011100 : 14'b00000000000000;
								assign node304 = (inp[1]) ? node306 : 14'b00000000000000;
									assign node306 = (inp[3]) ? 14'b00000000000000 : node307;
										assign node307 = (inp[9]) ? 14'b00000000000000 : 14'b10100100111000;
							assign node311 = (inp[8]) ? node313 : 14'b00000000000000;
								assign node313 = (inp[6]) ? node315 : 14'b00000000000000;
									assign node315 = (inp[3]) ? node317 : 14'b00000000000000;
										assign node317 = (inp[9]) ? 14'b01100000001010 : 14'b00000000000000;
						assign node320 = (inp[9]) ? node322 : 14'b00000000000000;
							assign node322 = (inp[7]) ? node324 : 14'b00000000000000;
								assign node324 = (inp[4]) ? 14'b00000000000000 : node325;
									assign node325 = (inp[8]) ? node327 : 14'b00000000000000;
										assign node327 = (inp[3]) ? 14'b01100000000010 : 14'b00000000000000;
					assign node331 = (inp[2]) ? 14'b00000000000000 : node332;
						assign node332 = (inp[5]) ? 14'b00000000000000 : node333;
							assign node333 = (inp[7]) ? 14'b00000000000000 : node334;
								assign node334 = (inp[0]) ? 14'b00000000000000 : node335;
									assign node335 = (inp[4]) ? node337 : 14'b00000000000000;
										assign node337 = (inp[8]) ? 14'b00000000000000 : 14'b00000000000000;
			assign node344 = (inp[11]) ? node406 : node345;
				assign node345 = (inp[1]) ? node357 : node346;
					assign node346 = (inp[6]) ? node348 : 14'b00000000000000;
						assign node348 = (inp[3]) ? node350 : 14'b00000000000000;
							assign node350 = (inp[9]) ? node352 : 14'b00000000000000;
								assign node352 = (inp[8]) ? node354 : 14'b00000000000000;
									assign node354 = (inp[7]) ? 14'b00100100001101 : 14'b00000000000000;
					assign node357 = (inp[12]) ? node381 : node358;
						assign node358 = (inp[2]) ? 14'b00000000000000 : node359;
							assign node359 = (inp[5]) ? node373 : node360;
								assign node360 = (inp[6]) ? node368 : node361;
									assign node361 = (inp[9]) ? node365 : node362;
										assign node362 = (inp[0]) ? 14'b00000000000000 : 14'b00000000000000;
										assign node365 = (inp[0]) ? 14'b00000000000000 : 14'b00001000000000;
									assign node368 = (inp[0]) ? 14'b00000000000000 : node369;
										assign node369 = (inp[7]) ? 14'b00000000011101 : 14'b00000000000000;
								assign node373 = (inp[7]) ? 14'b00000000000000 : node374;
									assign node374 = (inp[9]) ? node376 : 14'b00000000000000;
										assign node376 = (inp[8]) ? 14'b00000000000000 : 14'b00000000000000;
						assign node381 = (inp[7]) ? node395 : node382;
							assign node382 = (inp[9]) ? node388 : node383;
								assign node383 = (inp[3]) ? 14'b00000000000000 : node384;
									assign node384 = (inp[8]) ? 14'b00000100001110 : 14'b00000000000000;
								assign node388 = (inp[8]) ? 14'b00000000000000 : node389;
									assign node389 = (inp[3]) ? node391 : 14'b00000000000000;
										assign node391 = (inp[2]) ? 14'b00000000000000 : 14'b10100000001000;
							assign node395 = (inp[0]) ? 14'b00000000000000 : node396;
								assign node396 = (inp[9]) ? node402 : node397;
									assign node397 = (inp[3]) ? 14'b00000000000000 : node398;
										assign node398 = (inp[8]) ? 14'b10000000101000 : 14'b00000000011101;
									assign node402 = (inp[2]) ? 14'b00000000011100 : 14'b00000000000000;
				assign node406 = (inp[12]) ? node436 : node407;
					assign node407 = (inp[1]) ? node409 : 14'b00000000000000;
						assign node409 = (inp[3]) ? node419 : node410;
							assign node410 = (inp[6]) ? 14'b00000000000000 : node411;
								assign node411 = (inp[9]) ? 14'b00000000000000 : node412;
									assign node412 = (inp[8]) ? 14'b10100100011000 : node413;
										assign node413 = (inp[5]) ? 14'b00000000011100 : 14'b00000000000000;
							assign node419 = (inp[8]) ? node431 : node420;
								assign node420 = (inp[9]) ? node424 : node421;
									assign node421 = (inp[2]) ? 14'b00000000000000 : 14'b00100000000011;
									assign node424 = (inp[5]) ? node428 : node425;
										assign node425 = (inp[7]) ? 14'b01000100000010 : 14'b00000000000000;
										assign node428 = (inp[6]) ? 14'b10100101111111 : 14'b00100000000011;
								assign node431 = (inp[7]) ? node433 : 14'b00000000000000;
									assign node433 = (inp[6]) ? 14'b00100100001101 : 14'b00000000000000;
					assign node436 = (inp[8]) ? 14'b10000100001000 : node437;
						assign node437 = (inp[1]) ? 14'b00000000000000 : node438;
							assign node438 = (inp[6]) ? node440 : 14'b00000000000000;
								assign node440 = (inp[9]) ? 14'b00000000000000 : node441;
									assign node441 = (inp[3]) ? 14'b10010101111110 : 14'b00000000000000;

endmodule