module dtc_split125_bm68 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node98;
	wire [3-1:0] node100;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node123;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node232;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node250;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node269;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node278;
	wire [3-1:0] node280;

	assign outp = (inp[9]) ? node192 : node1;
		assign node1 = (inp[6]) ? node87 : node2;
			assign node2 = (inp[10]) ? node42 : node3;
				assign node3 = (inp[7]) ? node11 : node4;
					assign node4 = (inp[8]) ? node6 : 3'b111;
						assign node6 = (inp[11]) ? node8 : 3'b111;
							assign node8 = (inp[5]) ? 3'b011 : 3'b111;
					assign node11 = (inp[11]) ? node21 : node12;
						assign node12 = (inp[1]) ? node14 : 3'b111;
							assign node14 = (inp[4]) ? 3'b011 : node15;
								assign node15 = (inp[8]) ? node17 : 3'b111;
									assign node17 = (inp[0]) ? 3'b011 : 3'b111;
						assign node21 = (inp[3]) ? node33 : node22;
							assign node22 = (inp[0]) ? node28 : node23;
								assign node23 = (inp[4]) ? 3'b011 : node24;
									assign node24 = (inp[8]) ? 3'b011 : 3'b111;
								assign node28 = (inp[5]) ? 3'b101 : node29;
									assign node29 = (inp[1]) ? 3'b011 : 3'b111;
							assign node33 = (inp[0]) ? node37 : node34;
								assign node34 = (inp[8]) ? 3'b101 : 3'b011;
								assign node37 = (inp[5]) ? node39 : 3'b101;
									assign node39 = (inp[8]) ? 3'b001 : 3'b101;
				assign node42 = (inp[11]) ? node64 : node43;
					assign node43 = (inp[7]) ? node51 : node44;
						assign node44 = (inp[0]) ? node46 : 3'b011;
							assign node46 = (inp[2]) ? node48 : 3'b011;
								assign node48 = (inp[8]) ? 3'b101 : 3'b111;
						assign node51 = (inp[4]) ? node59 : node52;
							assign node52 = (inp[2]) ? 3'b101 : node53;
								assign node53 = (inp[1]) ? 3'b101 : node54;
									assign node54 = (inp[3]) ? 3'b001 : 3'b011;
							assign node59 = (inp[8]) ? 3'b001 : node60;
								assign node60 = (inp[2]) ? 3'b001 : 3'b101;
					assign node64 = (inp[7]) ? node76 : node65;
						assign node65 = (inp[0]) ? node71 : node66;
							assign node66 = (inp[2]) ? node68 : 3'b101;
								assign node68 = (inp[4]) ? 3'b011 : 3'b101;
							assign node71 = (inp[2]) ? 3'b101 : node72;
								assign node72 = (inp[3]) ? 3'b001 : 3'b011;
						assign node76 = (inp[8]) ? node82 : node77;
							assign node77 = (inp[0]) ? node79 : 3'b001;
								assign node79 = (inp[4]) ? 3'b110 : 3'b001;
							assign node82 = (inp[3]) ? 3'b110 : node83;
								assign node83 = (inp[2]) ? 3'b001 : 3'b110;
			assign node87 = (inp[10]) ? node147 : node88;
				assign node88 = (inp[11]) ? node116 : node89;
					assign node89 = (inp[7]) ? node103 : node90;
						assign node90 = (inp[3]) ? node98 : node91;
							assign node91 = (inp[8]) ? node93 : 3'b011;
								assign node93 = (inp[2]) ? 3'b101 : node94;
									assign node94 = (inp[5]) ? 3'b101 : 3'b011;
							assign node98 = (inp[8]) ? node100 : 3'b101;
								assign node100 = (inp[0]) ? 3'b001 : 3'b101;
						assign node103 = (inp[4]) ? node109 : node104;
							assign node104 = (inp[1]) ? 3'b001 : node105;
								assign node105 = (inp[8]) ? 3'b001 : 3'b101;
							assign node109 = (inp[5]) ? 3'b110 : node110;
								assign node110 = (inp[0]) ? node112 : 3'b001;
									assign node112 = (inp[8]) ? 3'b110 : 3'b001;
					assign node116 = (inp[7]) ? node128 : node117;
						assign node117 = (inp[8]) ? node121 : node118;
							assign node118 = (inp[2]) ? 3'b001 : 3'b101;
							assign node121 = (inp[3]) ? node123 : 3'b001;
								assign node123 = (inp[1]) ? node125 : 3'b110;
									assign node125 = (inp[4]) ? 3'b110 : 3'b001;
						assign node128 = (inp[0]) ? node138 : node129;
							assign node129 = (inp[3]) ? node135 : node130;
								assign node130 = (inp[2]) ? 3'b110 : node131;
									assign node131 = (inp[8]) ? 3'b110 : 3'b001;
								assign node135 = (inp[5]) ? 3'b010 : 3'b110;
							assign node138 = (inp[1]) ? node144 : node139;
								assign node139 = (inp[8]) ? node141 : 3'b110;
									assign node141 = (inp[4]) ? 3'b100 : 3'b110;
								assign node144 = (inp[4]) ? 3'b010 : 3'b110;
				assign node147 = (inp[7]) ? node171 : node148;
					assign node148 = (inp[8]) ? node156 : node149;
						assign node149 = (inp[11]) ? node153 : node150;
							assign node150 = (inp[3]) ? 3'b110 : 3'b001;
							assign node153 = (inp[3]) ? 3'b010 : 3'b110;
						assign node156 = (inp[4]) ? node168 : node157;
							assign node157 = (inp[0]) ? node163 : node158;
								assign node158 = (inp[11]) ? 3'b010 : node159;
									assign node159 = (inp[5]) ? 3'b010 : 3'b110;
								assign node163 = (inp[1]) ? node165 : 3'b100;
									assign node165 = (inp[3]) ? 3'b010 : 3'b110;
							assign node168 = (inp[3]) ? 3'b100 : 3'b110;
					assign node171 = (inp[11]) ? node187 : node172;
						assign node172 = (inp[8]) ? node182 : node173;
							assign node173 = (inp[4]) ? node177 : node174;
								assign node174 = (inp[5]) ? 3'b010 : 3'b110;
								assign node177 = (inp[1]) ? node179 : 3'b010;
									assign node179 = (inp[3]) ? 3'b100 : 3'b010;
							assign node182 = (inp[3]) ? 3'b100 : node183;
								assign node183 = (inp[4]) ? 3'b100 : 3'b010;
						assign node187 = (inp[8]) ? node189 : 3'b100;
							assign node189 = (inp[4]) ? 3'b000 : 3'b100;
		assign node192 = (inp[6]) ? node264 : node193;
			assign node193 = (inp[10]) ? node237 : node194;
				assign node194 = (inp[7]) ? node214 : node195;
					assign node195 = (inp[11]) ? node203 : node196;
						assign node196 = (inp[3]) ? node200 : node197;
							assign node197 = (inp[8]) ? 3'b001 : 3'b101;
							assign node200 = (inp[8]) ? 3'b110 : 3'b001;
						assign node203 = (inp[8]) ? node211 : node204;
							assign node204 = (inp[3]) ? 3'b110 : node205;
								assign node205 = (inp[1]) ? node207 : 3'b001;
									assign node207 = (inp[4]) ? 3'b110 : 3'b001;
							assign node211 = (inp[3]) ? 3'b010 : 3'b110;
					assign node214 = (inp[11]) ? node224 : node215;
						assign node215 = (inp[8]) ? 3'b010 : node216;
							assign node216 = (inp[3]) ? node218 : 3'b110;
								assign node218 = (inp[2]) ? 3'b010 : node219;
									assign node219 = (inp[5]) ? 3'b010 : 3'b110;
						assign node224 = (inp[1]) ? node230 : node225;
							assign node225 = (inp[4]) ? node227 : 3'b010;
								assign node227 = (inp[2]) ? 3'b100 : 3'b010;
							assign node230 = (inp[8]) ? node232 : 3'b010;
								assign node232 = (inp[3]) ? node234 : 3'b100;
									assign node234 = (inp[2]) ? 3'b000 : 3'b100;
				assign node237 = (inp[7]) ? node255 : node238;
					assign node238 = (inp[11]) ? node246 : node239;
						assign node239 = (inp[5]) ? node241 : 3'b010;
							assign node241 = (inp[2]) ? 3'b010 : node242;
								assign node242 = (inp[4]) ? 3'b010 : 3'b110;
						assign node246 = (inp[4]) ? 3'b100 : node247;
							assign node247 = (inp[2]) ? 3'b010 : node248;
								assign node248 = (inp[5]) ? node250 : 3'b100;
									assign node250 = (inp[8]) ? 3'b000 : 3'b010;
					assign node255 = (inp[11]) ? 3'b000 : node256;
						assign node256 = (inp[8]) ? 3'b000 : node257;
							assign node257 = (inp[3]) ? node259 : 3'b100;
								assign node259 = (inp[1]) ? 3'b100 : 3'b000;
			assign node264 = (inp[7]) ? 3'b000 : node265;
				assign node265 = (inp[10]) ? 3'b000 : node266;
					assign node266 = (inp[11]) ? node276 : node267;
						assign node267 = (inp[3]) ? node273 : node268;
							assign node268 = (inp[8]) ? 3'b100 : node269;
								assign node269 = (inp[5]) ? 3'b100 : 3'b010;
							assign node273 = (inp[8]) ? 3'b000 : 3'b100;
						assign node276 = (inp[8]) ? 3'b000 : node277;
							assign node277 = (inp[3]) ? 3'b000 : node278;
								assign node278 = (inp[5]) ? node280 : 3'b100;
									assign node280 = (inp[2]) ? 3'b100 : 3'b000;

endmodule