module dtc_split33_bm83 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node16;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node33;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node103;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node235;
	wire [3-1:0] node238;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node275;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node293;
	wire [3-1:0] node294;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node327;
	wire [3-1:0] node329;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node432;
	wire [3-1:0] node435;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node443;
	wire [3-1:0] node444;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node462;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node475;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node485;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node492;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node502;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node510;
	wire [3-1:0] node511;
	wire [3-1:0] node515;
	wire [3-1:0] node516;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node526;
	wire [3-1:0] node527;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node538;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node559;
	wire [3-1:0] node563;
	wire [3-1:0] node565;
	wire [3-1:0] node568;
	wire [3-1:0] node569;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node581;
	wire [3-1:0] node584;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node591;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node601;
	wire [3-1:0] node604;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node623;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node638;
	wire [3-1:0] node639;
	wire [3-1:0] node640;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node645;
	wire [3-1:0] node649;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node658;
	wire [3-1:0] node659;
	wire [3-1:0] node660;
	wire [3-1:0] node662;
	wire [3-1:0] node665;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node673;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node679;
	wire [3-1:0] node680;
	wire [3-1:0] node682;
	wire [3-1:0] node685;
	wire [3-1:0] node686;
	wire [3-1:0] node689;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node728;
	wire [3-1:0] node729;
	wire [3-1:0] node731;
	wire [3-1:0] node732;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node760;
	wire [3-1:0] node763;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node772;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node775;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node782;
	wire [3-1:0] node784;
	wire [3-1:0] node787;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node796;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node802;
	wire [3-1:0] node806;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node812;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node822;
	wire [3-1:0] node826;
	wire [3-1:0] node827;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node850;
	wire [3-1:0] node853;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node859;
	wire [3-1:0] node860;
	wire [3-1:0] node863;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node877;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node884;
	wire [3-1:0] node887;
	wire [3-1:0] node889;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node899;
	wire [3-1:0] node901;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node909;
	wire [3-1:0] node910;
	wire [3-1:0] node911;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node923;
	wire [3-1:0] node926;
	wire [3-1:0] node927;
	wire [3-1:0] node928;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node935;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node941;
	wire [3-1:0] node943;
	wire [3-1:0] node946;
	wire [3-1:0] node947;
	wire [3-1:0] node950;
	wire [3-1:0] node953;
	wire [3-1:0] node954;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node964;
	wire [3-1:0] node965;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node984;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node992;
	wire [3-1:0] node993;
	wire [3-1:0] node994;
	wire [3-1:0] node997;
	wire [3-1:0] node1000;
	wire [3-1:0] node1001;
	wire [3-1:0] node1005;
	wire [3-1:0] node1006;
	wire [3-1:0] node1007;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1012;
	wire [3-1:0] node1013;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1025;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1039;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1057;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1069;
	wire [3-1:0] node1071;
	wire [3-1:0] node1074;
	wire [3-1:0] node1075;
	wire [3-1:0] node1077;
	wire [3-1:0] node1079;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1086;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1093;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1100;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1116;
	wire [3-1:0] node1118;
	wire [3-1:0] node1120;

	assign outp = (inp[3]) ? node636 : node1;
		assign node1 = (inp[4]) ? node261 : node2;
			assign node2 = (inp[9]) ? node112 : node3;
				assign node3 = (inp[5]) ? node53 : node4;
					assign node4 = (inp[7]) ? node44 : node5;
						assign node5 = (inp[0]) ? node29 : node6;
							assign node6 = (inp[11]) ? node16 : node7;
								assign node7 = (inp[1]) ? node11 : node8;
									assign node8 = (inp[6]) ? 3'b111 : 3'b001;
									assign node11 = (inp[10]) ? 3'b011 : node12;
										assign node12 = (inp[8]) ? 3'b001 : 3'b001;
								assign node16 = (inp[1]) ? node22 : node17;
									assign node17 = (inp[6]) ? 3'b011 : node18;
										assign node18 = (inp[8]) ? 3'b001 : 3'b101;
									assign node22 = (inp[8]) ? node26 : node23;
										assign node23 = (inp[6]) ? 3'b101 : 3'b101;
										assign node26 = (inp[10]) ? 3'b111 : 3'b101;
							assign node29 = (inp[8]) ? node37 : node30;
								assign node30 = (inp[2]) ? 3'b111 : node31;
									assign node31 = (inp[1]) ? node33 : 3'b011;
										assign node33 = (inp[6]) ? 3'b111 : 3'b011;
								assign node37 = (inp[11]) ? 3'b111 : node38;
									assign node38 = (inp[2]) ? node40 : 3'b111;
										assign node40 = (inp[6]) ? 3'b111 : 3'b011;
						assign node44 = (inp[8]) ? node46 : 3'b111;
							assign node46 = (inp[0]) ? 3'b111 : node47;
								assign node47 = (inp[2]) ? node49 : 3'b111;
									assign node49 = (inp[11]) ? 3'b111 : 3'b101;
					assign node53 = (inp[7]) ? node89 : node54;
						assign node54 = (inp[1]) ? node74 : node55;
							assign node55 = (inp[0]) ? node67 : node56;
								assign node56 = (inp[6]) ? node62 : node57;
									assign node57 = (inp[2]) ? node59 : 3'b110;
										assign node59 = (inp[8]) ? 3'b101 : 3'b001;
									assign node62 = (inp[11]) ? 3'b011 : node63;
										assign node63 = (inp[2]) ? 3'b011 : 3'b011;
								assign node67 = (inp[8]) ? node71 : node68;
									assign node68 = (inp[2]) ? 3'b101 : 3'b001;
									assign node71 = (inp[2]) ? 3'b001 : 3'b101;
							assign node74 = (inp[0]) ? node84 : node75;
								assign node75 = (inp[11]) ? node81 : node76;
									assign node76 = (inp[8]) ? node78 : 3'b011;
										assign node78 = (inp[2]) ? 3'b111 : 3'b101;
									assign node81 = (inp[6]) ? 3'b011 : 3'b001;
								assign node84 = (inp[6]) ? 3'b111 : node85;
									assign node85 = (inp[10]) ? 3'b011 : 3'b111;
						assign node89 = (inp[0]) ? node103 : node90;
							assign node90 = (inp[6]) ? node98 : node91;
								assign node91 = (inp[1]) ? node93 : 3'b111;
									assign node93 = (inp[8]) ? node95 : 3'b011;
										assign node95 = (inp[11]) ? 3'b011 : 3'b111;
								assign node98 = (inp[2]) ? 3'b111 : node99;
									assign node99 = (inp[10]) ? 3'b101 : 3'b111;
							assign node103 = (inp[1]) ? node105 : 3'b011;
								assign node105 = (inp[6]) ? 3'b111 : node106;
									assign node106 = (inp[11]) ? 3'b011 : node107;
										assign node107 = (inp[8]) ? 3'b111 : 3'b011;
				assign node112 = (inp[6]) ? node192 : node113;
					assign node113 = (inp[0]) ? node153 : node114;
						assign node114 = (inp[5]) ? node138 : node115;
							assign node115 = (inp[1]) ? node125 : node116;
								assign node116 = (inp[10]) ? node120 : node117;
									assign node117 = (inp[7]) ? 3'b001 : 3'b110;
									assign node120 = (inp[2]) ? 3'b110 : node121;
										assign node121 = (inp[7]) ? 3'b110 : 3'b010;
								assign node125 = (inp[10]) ? node131 : node126;
									assign node126 = (inp[8]) ? 3'b101 : node127;
										assign node127 = (inp[2]) ? 3'b101 : 3'b001;
									assign node131 = (inp[11]) ? node135 : node132;
										assign node132 = (inp[2]) ? 3'b001 : 3'b001;
										assign node135 = (inp[8]) ? 3'b000 : 3'b110;
							assign node138 = (inp[11]) ? node146 : node139;
								assign node139 = (inp[10]) ? node141 : 3'b001;
									assign node141 = (inp[7]) ? 3'b110 : node142;
										assign node142 = (inp[2]) ? 3'b010 : 3'b100;
								assign node146 = (inp[1]) ? node148 : 3'b010;
									assign node148 = (inp[10]) ? node150 : 3'b110;
										assign node150 = (inp[7]) ? 3'b110 : 3'b010;
						assign node153 = (inp[10]) ? node173 : node154;
							assign node154 = (inp[1]) ? node166 : node155;
								assign node155 = (inp[7]) ? node163 : node156;
									assign node156 = (inp[5]) ? node160 : node157;
										assign node157 = (inp[8]) ? 3'b101 : 3'b101;
										assign node160 = (inp[8]) ? 3'b001 : 3'b001;
									assign node163 = (inp[11]) ? 3'b011 : 3'b101;
								assign node166 = (inp[2]) ? 3'b011 : node167;
									assign node167 = (inp[5]) ? 3'b101 : node168;
										assign node168 = (inp[7]) ? 3'b111 : 3'b011;
							assign node173 = (inp[5]) ? node181 : node174;
								assign node174 = (inp[7]) ? 3'b101 : node175;
									assign node175 = (inp[1]) ? 3'b101 : node176;
										assign node176 = (inp[2]) ? 3'b001 : 3'b001;
								assign node181 = (inp[1]) ? node187 : node182;
									assign node182 = (inp[7]) ? node184 : 3'b110;
										assign node184 = (inp[8]) ? 3'b001 : 3'b110;
									assign node187 = (inp[2]) ? 3'b001 : node188;
										assign node188 = (inp[8]) ? 3'b110 : 3'b001;
					assign node192 = (inp[0]) ? node230 : node193;
						assign node193 = (inp[7]) ? node217 : node194;
							assign node194 = (inp[10]) ? node206 : node195;
								assign node195 = (inp[11]) ? node201 : node196;
									assign node196 = (inp[8]) ? node198 : 3'b101;
										assign node198 = (inp[2]) ? 3'b111 : 3'b011;
									assign node201 = (inp[1]) ? 3'b101 : node202;
										assign node202 = (inp[5]) ? 3'b001 : 3'b101;
								assign node206 = (inp[8]) ? node214 : node207;
									assign node207 = (inp[2]) ? node211 : node208;
										assign node208 = (inp[1]) ? 3'b110 : 3'b010;
										assign node211 = (inp[1]) ? 3'b001 : 3'b110;
									assign node214 = (inp[1]) ? 3'b101 : 3'b001;
							assign node217 = (inp[5]) ? node227 : node218;
								assign node218 = (inp[8]) ? node220 : 3'b101;
									assign node220 = (inp[1]) ? node224 : node221;
										assign node221 = (inp[2]) ? 3'b011 : 3'b101;
										assign node224 = (inp[10]) ? 3'b011 : 3'b001;
								assign node227 = (inp[1]) ? 3'b101 : 3'b001;
						assign node230 = (inp[10]) ? node242 : node231;
							assign node231 = (inp[11]) ? node233 : 3'b111;
								assign node233 = (inp[1]) ? 3'b111 : node234;
									assign node234 = (inp[5]) ? node238 : node235;
										assign node235 = (inp[7]) ? 3'b111 : 3'b011;
										assign node238 = (inp[7]) ? 3'b011 : 3'b001;
							assign node242 = (inp[5]) ? node250 : node243;
								assign node243 = (inp[8]) ? 3'b111 : node244;
									assign node244 = (inp[2]) ? 3'b011 : node245;
										assign node245 = (inp[1]) ? 3'b011 : 3'b101;
								assign node250 = (inp[11]) ? node256 : node251;
									assign node251 = (inp[8]) ? 3'b011 : node252;
										assign node252 = (inp[7]) ? 3'b011 : 3'b101;
									assign node256 = (inp[7]) ? node258 : 3'b101;
										assign node258 = (inp[1]) ? 3'b011 : 3'b101;
			assign node261 = (inp[9]) ? node461 : node262;
				assign node262 = (inp[0]) ? node360 : node263;
					assign node263 = (inp[11]) ? node311 : node264;
						assign node264 = (inp[7]) ? node286 : node265;
							assign node265 = (inp[6]) ? node275 : node266;
								assign node266 = (inp[5]) ? node270 : node267;
									assign node267 = (inp[2]) ? 3'b110 : 3'b101;
									assign node270 = (inp[2]) ? 3'b110 : node271;
										assign node271 = (inp[8]) ? 3'b010 : 3'b010;
								assign node275 = (inp[5]) ? node281 : node276;
									assign node276 = (inp[10]) ? node278 : 3'b101;
										assign node278 = (inp[1]) ? 3'b001 : 3'b001;
									assign node281 = (inp[1]) ? 3'b010 : node282;
										assign node282 = (inp[10]) ? 3'b110 : 3'b101;
							assign node286 = (inp[1]) ? node298 : node287;
								assign node287 = (inp[6]) ? node293 : node288;
									assign node288 = (inp[8]) ? 3'b001 : node289;
										assign node289 = (inp[2]) ? 3'b001 : 3'b101;
									assign node293 = (inp[2]) ? 3'b101 : node294;
										assign node294 = (inp[5]) ? 3'b101 : 3'b001;
								assign node298 = (inp[5]) ? node306 : node299;
									assign node299 = (inp[6]) ? node303 : node300;
										assign node300 = (inp[10]) ? 3'b001 : 3'b100;
										assign node303 = (inp[10]) ? 3'b010 : 3'b000;
									assign node306 = (inp[10]) ? 3'b101 : node307;
										assign node307 = (inp[8]) ? 3'b111 : 3'b011;
						assign node311 = (inp[6]) ? node333 : node312;
							assign node312 = (inp[10]) ? node326 : node313;
								assign node313 = (inp[1]) ? node319 : node314;
									assign node314 = (inp[8]) ? 3'b110 : node315;
										assign node315 = (inp[7]) ? 3'b110 : 3'b010;
									assign node319 = (inp[7]) ? node323 : node320;
										assign node320 = (inp[5]) ? 3'b010 : 3'b110;
										assign node323 = (inp[5]) ? 3'b000 : 3'b101;
								assign node326 = (inp[7]) ? 3'b110 : node327;
									assign node327 = (inp[8]) ? node329 : 3'b100;
										assign node329 = (inp[5]) ? 3'b010 : 3'b110;
							assign node333 = (inp[8]) ? node347 : node334;
								assign node334 = (inp[5]) ? node342 : node335;
									assign node335 = (inp[10]) ? node339 : node336;
										assign node336 = (inp[1]) ? 3'b010 : 3'b101;
										assign node339 = (inp[2]) ? 3'b001 : 3'b000;
									assign node342 = (inp[10]) ? node344 : 3'b000;
										assign node344 = (inp[1]) ? 3'b010 : 3'b110;
								assign node347 = (inp[10]) ? node353 : node348;
									assign node348 = (inp[7]) ? 3'b110 : node349;
										assign node349 = (inp[1]) ? 3'b010 : 3'b011;
									assign node353 = (inp[7]) ? node357 : node354;
										assign node354 = (inp[2]) ? 3'b100 : 3'b110;
										assign node357 = (inp[1]) ? 3'b001 : 3'b110;
					assign node360 = (inp[8]) ? node414 : node361;
						assign node361 = (inp[6]) ? node385 : node362;
							assign node362 = (inp[2]) ? node372 : node363;
								assign node363 = (inp[10]) ? 3'b001 : node364;
									assign node364 = (inp[7]) ? node368 : node365;
										assign node365 = (inp[11]) ? 3'b001 : 3'b000;
										assign node368 = (inp[11]) ? 3'b010 : 3'b001;
								assign node372 = (inp[11]) ? node378 : node373;
									assign node373 = (inp[10]) ? 3'b101 : node374;
										assign node374 = (inp[5]) ? 3'b001 : 3'b101;
									assign node378 = (inp[10]) ? node382 : node379;
										assign node379 = (inp[5]) ? 3'b101 : 3'b011;
										assign node382 = (inp[7]) ? 3'b001 : 3'b001;
							assign node385 = (inp[1]) ? node401 : node386;
								assign node386 = (inp[10]) ? node394 : node387;
									assign node387 = (inp[7]) ? node391 : node388;
										assign node388 = (inp[2]) ? 3'b011 : 3'b001;
										assign node391 = (inp[5]) ? 3'b001 : 3'b111;
									assign node394 = (inp[5]) ? node398 : node395;
										assign node395 = (inp[11]) ? 3'b000 : 3'b000;
										assign node398 = (inp[2]) ? 3'b011 : 3'b000;
								assign node401 = (inp[10]) ? node407 : node402;
									assign node402 = (inp[5]) ? 3'b111 : node403;
										assign node403 = (inp[7]) ? 3'b101 : 3'b001;
									assign node407 = (inp[5]) ? node411 : node408;
										assign node408 = (inp[2]) ? 3'b011 : 3'b111;
										assign node411 = (inp[7]) ? 3'b001 : 3'b101;
						assign node414 = (inp[7]) ? node438 : node415;
							assign node415 = (inp[1]) ? node429 : node416;
								assign node416 = (inp[6]) ? node424 : node417;
									assign node417 = (inp[5]) ? node421 : node418;
										assign node418 = (inp[2]) ? 3'b010 : 3'b001;
										assign node421 = (inp[2]) ? 3'b000 : 3'b110;
									assign node424 = (inp[11]) ? 3'b101 : node425;
										assign node425 = (inp[5]) ? 3'b001 : 3'b110;
								assign node429 = (inp[11]) ? node431 : 3'b011;
									assign node431 = (inp[10]) ? node435 : node432;
										assign node432 = (inp[5]) ? 3'b101 : 3'b001;
										assign node435 = (inp[5]) ? 3'b011 : 3'b101;
							assign node438 = (inp[2]) ? node450 : node439;
								assign node439 = (inp[5]) ? node443 : node440;
									assign node440 = (inp[10]) ? 3'b111 : 3'b011;
									assign node443 = (inp[1]) ? node447 : node444;
										assign node444 = (inp[10]) ? 3'b001 : 3'b101;
										assign node447 = (inp[6]) ? 3'b011 : 3'b111;
								assign node450 = (inp[5]) ? node456 : node451;
									assign node451 = (inp[6]) ? node453 : 3'b011;
										assign node453 = (inp[11]) ? 3'b001 : 3'b001;
									assign node456 = (inp[11]) ? node458 : 3'b011;
										assign node458 = (inp[1]) ? 3'b011 : 3'b001;
				assign node461 = (inp[0]) ? node543 : node462;
					assign node462 = (inp[6]) ? node502 : node463;
						assign node463 = (inp[1]) ? node483 : node464;
							assign node464 = (inp[8]) ? node472 : node465;
								assign node465 = (inp[5]) ? 3'b000 : node466;
									assign node466 = (inp[2]) ? 3'b010 : node467;
										assign node467 = (inp[11]) ? 3'b100 : 3'b000;
								assign node472 = (inp[7]) ? node478 : node473;
									assign node473 = (inp[5]) ? node475 : 3'b010;
										assign node475 = (inp[10]) ? 3'b000 : 3'b100;
									assign node478 = (inp[10]) ? 3'b010 : node479;
										assign node479 = (inp[5]) ? 3'b010 : 3'b100;
							assign node483 = (inp[10]) ? node495 : node484;
								assign node484 = (inp[5]) ? node490 : node485;
									assign node485 = (inp[7]) ? node487 : 3'b010;
										assign node487 = (inp[11]) ? 3'b110 : 3'b010;
									assign node490 = (inp[7]) ? node492 : 3'b100;
										assign node492 = (inp[11]) ? 3'b010 : 3'b100;
								assign node495 = (inp[2]) ? 3'b100 : node496;
									assign node496 = (inp[11]) ? 3'b100 : node497;
										assign node497 = (inp[8]) ? 3'b010 : 3'b100;
						assign node502 = (inp[5]) ? node526 : node503;
							assign node503 = (inp[8]) ? node515 : node504;
								assign node504 = (inp[10]) ? node510 : node505;
									assign node505 = (inp[7]) ? 3'b011 : node506;
										assign node506 = (inp[1]) ? 3'b111 : 3'b110;
									assign node510 = (inp[1]) ? 3'b110 : node511;
										assign node511 = (inp[2]) ? 3'b010 : 3'b010;
								assign node515 = (inp[10]) ? node521 : node516;
									assign node516 = (inp[1]) ? node518 : 3'b001;
										assign node518 = (inp[7]) ? 3'b101 : 3'b001;
									assign node521 = (inp[11]) ? 3'b110 : node522;
										assign node522 = (inp[7]) ? 3'b001 : 3'b110;
							assign node526 = (inp[7]) ? node536 : node527;
								assign node527 = (inp[1]) ? node529 : 3'b010;
									assign node529 = (inp[8]) ? node533 : node530;
										assign node530 = (inp[10]) ? 3'b100 : 3'b110;
										assign node533 = (inp[2]) ? 3'b000 : 3'b100;
								assign node536 = (inp[10]) ? node538 : 3'b110;
									assign node538 = (inp[8]) ? node540 : 3'b010;
										assign node540 = (inp[11]) ? 3'b010 : 3'b110;
					assign node543 = (inp[6]) ? node587 : node544;
						assign node544 = (inp[10]) ? node568 : node545;
							assign node545 = (inp[7]) ? node557 : node546;
								assign node546 = (inp[5]) ? node552 : node547;
									assign node547 = (inp[11]) ? 3'b110 : node548;
										assign node548 = (inp[2]) ? 3'b001 : 3'b110;
									assign node552 = (inp[11]) ? 3'b010 : node553;
										assign node553 = (inp[1]) ? 3'b110 : 3'b010;
								assign node557 = (inp[11]) ? node563 : node558;
									assign node558 = (inp[8]) ? 3'b001 : node559;
										assign node559 = (inp[1]) ? 3'b101 : 3'b001;
									assign node563 = (inp[1]) ? node565 : 3'b110;
										assign node565 = (inp[8]) ? 3'b001 : 3'b101;
							assign node568 = (inp[1]) ? node578 : node569;
								assign node569 = (inp[7]) ? node575 : node570;
									assign node570 = (inp[5]) ? 3'b100 : node571;
										assign node571 = (inp[8]) ? 3'b010 : 3'b000;
									assign node575 = (inp[5]) ? 3'b010 : 3'b110;
								assign node578 = (inp[8]) ? node584 : node579;
									assign node579 = (inp[7]) ? node581 : 3'b010;
										assign node581 = (inp[5]) ? 3'b010 : 3'b110;
									assign node584 = (inp[7]) ? 3'b001 : 3'b110;
						assign node587 = (inp[1]) ? node617 : node588;
							assign node588 = (inp[5]) ? node604 : node589;
								assign node589 = (inp[11]) ? node597 : node590;
									assign node590 = (inp[2]) ? node594 : node591;
										assign node591 = (inp[7]) ? 3'b001 : 3'b001;
										assign node594 = (inp[7]) ? 3'b101 : 3'b101;
									assign node597 = (inp[7]) ? node601 : node598;
										assign node598 = (inp[10]) ? 3'b110 : 3'b101;
										assign node601 = (inp[10]) ? 3'b101 : 3'b001;
								assign node604 = (inp[10]) ? node610 : node605;
									assign node605 = (inp[7]) ? 3'b001 : node606;
										assign node606 = (inp[2]) ? 3'b111 : 3'b110;
									assign node610 = (inp[11]) ? node614 : node611;
										assign node611 = (inp[7]) ? 3'b000 : 3'b010;
										assign node614 = (inp[7]) ? 3'b110 : 3'b010;
							assign node617 = (inp[2]) ? node627 : node618;
								assign node618 = (inp[11]) ? node622 : node619;
									assign node619 = (inp[8]) ? 3'b001 : 3'b101;
									assign node622 = (inp[5]) ? 3'b110 : node623;
										assign node623 = (inp[8]) ? 3'b101 : 3'b001;
								assign node627 = (inp[7]) ? node633 : node628;
									assign node628 = (inp[5]) ? node630 : 3'b001;
										assign node630 = (inp[8]) ? 3'b101 : 3'b001;
									assign node633 = (inp[11]) ? 3'b101 : 3'b011;
		assign node636 = (inp[4]) ? node958 : node637;
			assign node637 = (inp[9]) ? node815 : node638;
				assign node638 = (inp[6]) ? node726 : node639;
					assign node639 = (inp[0]) ? node677 : node640;
						assign node640 = (inp[7]) ? node658 : node641;
							assign node641 = (inp[5]) ? node649 : node642;
								assign node642 = (inp[8]) ? 3'b100 : node643;
									assign node643 = (inp[1]) ? node645 : 3'b000;
										assign node645 = (inp[10]) ? 3'b100 : 3'b000;
								assign node649 = (inp[10]) ? 3'b000 : node650;
									assign node650 = (inp[8]) ? node654 : node651;
										assign node651 = (inp[2]) ? 3'b100 : 3'b000;
										assign node654 = (inp[2]) ? 3'b000 : 3'b100;
							assign node658 = (inp[11]) ? node668 : node659;
								assign node659 = (inp[8]) ? node665 : node660;
									assign node660 = (inp[1]) ? node662 : 3'b100;
										assign node662 = (inp[2]) ? 3'b010 : 3'b110;
									assign node665 = (inp[5]) ? 3'b110 : 3'b010;
								assign node668 = (inp[5]) ? 3'b000 : node669;
									assign node669 = (inp[1]) ? node673 : node670;
										assign node670 = (inp[10]) ? 3'b100 : 3'b110;
										assign node673 = (inp[8]) ? 3'b000 : 3'b100;
						assign node677 = (inp[11]) ? node703 : node678;
							assign node678 = (inp[1]) ? node692 : node679;
								assign node679 = (inp[2]) ? node685 : node680;
									assign node680 = (inp[10]) ? node682 : 3'b010;
										assign node682 = (inp[5]) ? 3'b000 : 3'b010;
									assign node685 = (inp[7]) ? node689 : node686;
										assign node686 = (inp[10]) ? 3'b000 : 3'b000;
										assign node689 = (inp[10]) ? 3'b110 : 3'b100;
								assign node692 = (inp[7]) ? node696 : node693;
									assign node693 = (inp[5]) ? 3'b010 : 3'b110;
									assign node696 = (inp[8]) ? node700 : node697;
										assign node697 = (inp[10]) ? 3'b010 : 3'b001;
										assign node700 = (inp[10]) ? 3'b001 : 3'b001;
							assign node703 = (inp[10]) ? node715 : node704;
								assign node704 = (inp[5]) ? node712 : node705;
									assign node705 = (inp[1]) ? node709 : node706;
										assign node706 = (inp[7]) ? 3'b100 : 3'b110;
										assign node709 = (inp[7]) ? 3'b011 : 3'b110;
									assign node712 = (inp[1]) ? 3'b110 : 3'b010;
								assign node715 = (inp[7]) ? node721 : node716;
									assign node716 = (inp[8]) ? node718 : 3'b100;
										assign node718 = (inp[1]) ? 3'b010 : 3'b100;
									assign node721 = (inp[8]) ? node723 : 3'b110;
										assign node723 = (inp[1]) ? 3'b000 : 3'b100;
					assign node726 = (inp[0]) ? node772 : node727;
						assign node727 = (inp[7]) ? node749 : node728;
							assign node728 = (inp[1]) ? node736 : node729;
								assign node729 = (inp[2]) ? node731 : 3'b000;
									assign node731 = (inp[10]) ? 3'b100 : node732;
										assign node732 = (inp[5]) ? 3'b000 : 3'b100;
								assign node736 = (inp[2]) ? node742 : node737;
									assign node737 = (inp[11]) ? node739 : 3'b110;
										assign node739 = (inp[5]) ? 3'b100 : 3'b110;
									assign node742 = (inp[8]) ? node746 : node743;
										assign node743 = (inp[10]) ? 3'b010 : 3'b000;
										assign node746 = (inp[5]) ? 3'b110 : 3'b110;
							assign node749 = (inp[10]) ? node763 : node750;
								assign node750 = (inp[11]) ? node756 : node751;
									assign node751 = (inp[1]) ? 3'b001 : node752;
										assign node752 = (inp[2]) ? 3'b010 : 3'b000;
									assign node756 = (inp[5]) ? node760 : node757;
										assign node757 = (inp[8]) ? 3'b101 : 3'b100;
										assign node760 = (inp[1]) ? 3'b001 : 3'b110;
								assign node763 = (inp[2]) ? node765 : 3'b110;
									assign node765 = (inp[5]) ? node769 : node766;
										assign node766 = (inp[1]) ? 3'b011 : 3'b001;
										assign node769 = (inp[11]) ? 3'b010 : 3'b110;
						assign node772 = (inp[1]) ? node796 : node773;
							assign node773 = (inp[7]) ? node787 : node774;
								assign node774 = (inp[10]) ? node782 : node775;
									assign node775 = (inp[8]) ? node779 : node776;
										assign node776 = (inp[2]) ? 3'b011 : 3'b110;
										assign node779 = (inp[5]) ? 3'b001 : 3'b100;
									assign node782 = (inp[8]) ? node784 : 3'b010;
										assign node784 = (inp[11]) ? 3'b010 : 3'b110;
								assign node787 = (inp[8]) ? node791 : node788;
									assign node788 = (inp[5]) ? 3'b001 : 3'b101;
									assign node791 = (inp[5]) ? 3'b110 : node792;
										assign node792 = (inp[10]) ? 3'b001 : 3'b010;
							assign node796 = (inp[5]) ? node806 : node797;
								assign node797 = (inp[10]) ? 3'b101 : node798;
									assign node798 = (inp[8]) ? node802 : node799;
										assign node799 = (inp[11]) ? 3'b101 : 3'b111;
										assign node802 = (inp[2]) ? 3'b011 : 3'b011;
								assign node806 = (inp[10]) ? node812 : node807;
									assign node807 = (inp[8]) ? 3'b101 : node808;
										assign node808 = (inp[11]) ? 3'b001 : 3'b101;
									assign node812 = (inp[2]) ? 3'b001 : 3'b101;
				assign node815 = (inp[6]) ? node871 : node816;
					assign node816 = (inp[0]) ? node832 : node817;
						assign node817 = (inp[1]) ? node819 : 3'b000;
							assign node819 = (inp[10]) ? 3'b000 : node820;
								assign node820 = (inp[5]) ? node826 : node821;
									assign node821 = (inp[7]) ? 3'b010 : node822;
										assign node822 = (inp[8]) ? 3'b100 : 3'b000;
									assign node826 = (inp[8]) ? 3'b000 : node827;
										assign node827 = (inp[7]) ? 3'b100 : 3'b000;
						assign node832 = (inp[7]) ? node846 : node833;
							assign node833 = (inp[1]) ? node835 : 3'b000;
								assign node835 = (inp[11]) ? node841 : node836;
									assign node836 = (inp[2]) ? 3'b100 : node837;
										assign node837 = (inp[5]) ? 3'b000 : 3'b100;
									assign node841 = (inp[10]) ? 3'b000 : node842;
										assign node842 = (inp[2]) ? 3'b010 : 3'b000;
							assign node846 = (inp[1]) ? node858 : node847;
								assign node847 = (inp[2]) ? node853 : node848;
									assign node848 = (inp[11]) ? node850 : 3'b100;
										assign node850 = (inp[10]) ? 3'b000 : 3'b100;
									assign node853 = (inp[8]) ? node855 : 3'b000;
										assign node855 = (inp[11]) ? 3'b100 : 3'b000;
								assign node858 = (inp[2]) ? node866 : node859;
									assign node859 = (inp[10]) ? node863 : node860;
										assign node860 = (inp[8]) ? 3'b110 : 3'b100;
										assign node863 = (inp[5]) ? 3'b000 : 3'b100;
									assign node866 = (inp[5]) ? 3'b010 : node867;
										assign node867 = (inp[10]) ? 3'b010 : 3'b110;
					assign node871 = (inp[0]) ? node909 : node872;
						assign node872 = (inp[11]) ? node892 : node873;
							assign node873 = (inp[8]) ? node881 : node874;
								assign node874 = (inp[10]) ? 3'b100 : node875;
									assign node875 = (inp[2]) ? node877 : 3'b000;
										assign node877 = (inp[1]) ? 3'b100 : 3'b000;
								assign node881 = (inp[10]) ? node887 : node882;
									assign node882 = (inp[5]) ? node884 : 3'b100;
										assign node884 = (inp[7]) ? 3'b000 : 3'b100;
									assign node887 = (inp[1]) ? node889 : 3'b000;
										assign node889 = (inp[5]) ? 3'b000 : 3'b000;
							assign node892 = (inp[10]) ? node904 : node893;
								assign node893 = (inp[7]) ? node899 : node894;
									assign node894 = (inp[5]) ? 3'b000 : node895;
										assign node895 = (inp[8]) ? 3'b110 : 3'b100;
									assign node899 = (inp[5]) ? node901 : 3'b010;
										assign node901 = (inp[8]) ? 3'b010 : 3'b100;
								assign node904 = (inp[5]) ? 3'b000 : node905;
									assign node905 = (inp[7]) ? 3'b100 : 3'b000;
						assign node909 = (inp[1]) ? node939 : node910;
							assign node910 = (inp[10]) ? node926 : node911;
								assign node911 = (inp[11]) ? node919 : node912;
									assign node912 = (inp[8]) ? node916 : node913;
										assign node913 = (inp[5]) ? 3'b010 : 3'b110;
										assign node916 = (inp[5]) ? 3'b110 : 3'b001;
									assign node919 = (inp[8]) ? node923 : node920;
										assign node920 = (inp[2]) ? 3'b110 : 3'b100;
										assign node923 = (inp[7]) ? 3'b110 : 3'b010;
								assign node926 = (inp[7]) ? node934 : node927;
									assign node927 = (inp[5]) ? node931 : node928;
										assign node928 = (inp[2]) ? 3'b010 : 3'b100;
										assign node931 = (inp[11]) ? 3'b000 : 3'b000;
									assign node934 = (inp[11]) ? 3'b010 : node935;
										assign node935 = (inp[5]) ? 3'b010 : 3'b110;
							assign node939 = (inp[10]) ? node953 : node940;
								assign node940 = (inp[5]) ? node946 : node941;
									assign node941 = (inp[2]) ? node943 : 3'b001;
										assign node943 = (inp[8]) ? 3'b001 : 3'b001;
									assign node946 = (inp[7]) ? node950 : node947;
										assign node947 = (inp[8]) ? 3'b110 : 3'b010;
										assign node950 = (inp[2]) ? 3'b001 : 3'b000;
								assign node953 = (inp[5]) ? 3'b100 : node954;
									assign node954 = (inp[7]) ? 3'b110 : 3'b010;
			assign node958 = (inp[9]) ? node1074 : node959;
				assign node959 = (inp[6]) ? node1005 : node960;
					assign node960 = (inp[1]) ? node974 : node961;
						assign node961 = (inp[5]) ? 3'b000 : node962;
							assign node962 = (inp[0]) ? node964 : 3'b000;
								assign node964 = (inp[11]) ? node968 : node965;
									assign node965 = (inp[7]) ? 3'b001 : 3'b000;
									assign node968 = (inp[10]) ? 3'b000 : node969;
										assign node969 = (inp[7]) ? 3'b100 : 3'b000;
						assign node974 = (inp[0]) ? node980 : node975;
							assign node975 = (inp[2]) ? node977 : 3'b000;
								assign node977 = (inp[7]) ? 3'b100 : 3'b000;
							assign node980 = (inp[2]) ? node992 : node981;
								assign node981 = (inp[10]) ? node987 : node982;
									assign node982 = (inp[7]) ? node984 : 3'b100;
										assign node984 = (inp[5]) ? 3'b100 : 3'b110;
									assign node987 = (inp[8]) ? 3'b100 : node988;
										assign node988 = (inp[5]) ? 3'b000 : 3'b000;
								assign node992 = (inp[7]) ? node1000 : node993;
									assign node993 = (inp[8]) ? node997 : node994;
										assign node994 = (inp[10]) ? 3'b000 : 3'b001;
										assign node997 = (inp[11]) ? 3'b000 : 3'b000;
									assign node1000 = (inp[11]) ? 3'b100 : node1001;
										assign node1001 = (inp[10]) ? 3'b010 : 3'b000;
					assign node1005 = (inp[0]) ? node1035 : node1006;
						assign node1006 = (inp[10]) ? node1028 : node1007;
							assign node1007 = (inp[8]) ? node1017 : node1008;
								assign node1008 = (inp[5]) ? node1012 : node1009;
									assign node1009 = (inp[2]) ? 3'b110 : 3'b100;
									assign node1012 = (inp[11]) ? 3'b100 : node1013;
										assign node1013 = (inp[7]) ? 3'b000 : 3'b100;
								assign node1017 = (inp[1]) ? node1021 : node1018;
									assign node1018 = (inp[11]) ? 3'b100 : 3'b000;
									assign node1021 = (inp[11]) ? node1025 : node1022;
										assign node1022 = (inp[7]) ? 3'b010 : 3'b100;
										assign node1025 = (inp[5]) ? 3'b100 : 3'b000;
							assign node1028 = (inp[5]) ? 3'b000 : node1029;
								assign node1029 = (inp[7]) ? 3'b010 : node1030;
									assign node1030 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1035 = (inp[10]) ? node1051 : node1036;
							assign node1036 = (inp[5]) ? node1044 : node1037;
								assign node1037 = (inp[11]) ? node1039 : 3'b001;
									assign node1039 = (inp[1]) ? node1041 : 3'b110;
										assign node1041 = (inp[7]) ? 3'b001 : 3'b010;
								assign node1044 = (inp[11]) ? node1046 : 3'b110;
									assign node1046 = (inp[8]) ? 3'b010 : node1047;
										assign node1047 = (inp[1]) ? 3'b010 : 3'b100;
							assign node1051 = (inp[7]) ? node1067 : node1052;
								assign node1052 = (inp[5]) ? node1060 : node1053;
									assign node1053 = (inp[11]) ? node1057 : node1054;
										assign node1054 = (inp[8]) ? 3'b010 : 3'b110;
										assign node1057 = (inp[1]) ? 3'b010 : 3'b000;
									assign node1060 = (inp[1]) ? node1064 : node1061;
										assign node1061 = (inp[2]) ? 3'b100 : 3'b000;
										assign node1064 = (inp[11]) ? 3'b100 : 3'b000;
								assign node1067 = (inp[8]) ? node1069 : 3'b010;
									assign node1069 = (inp[5]) ? node1071 : 3'b110;
										assign node1071 = (inp[11]) ? 3'b000 : 3'b010;
				assign node1074 = (inp[0]) ? node1086 : node1075;
					assign node1075 = (inp[1]) ? node1077 : 3'b000;
						assign node1077 = (inp[11]) ? node1079 : 3'b000;
							assign node1079 = (inp[5]) ? 3'b000 : node1080;
								assign node1080 = (inp[10]) ? 3'b000 : node1081;
									assign node1081 = (inp[7]) ? 3'b100 : 3'b000;
					assign node1086 = (inp[7]) ? node1098 : node1087;
						assign node1087 = (inp[5]) ? 3'b000 : node1088;
							assign node1088 = (inp[1]) ? node1090 : 3'b000;
								assign node1090 = (inp[10]) ? 3'b000 : node1091;
									assign node1091 = (inp[6]) ? node1093 : 3'b000;
										assign node1093 = (inp[8]) ? 3'b000 : 3'b100;
						assign node1098 = (inp[10]) ? node1116 : node1099;
							assign node1099 = (inp[1]) ? node1105 : node1100;
								assign node1100 = (inp[11]) ? node1102 : 3'b010;
									assign node1102 = (inp[8]) ? 3'b000 : 3'b100;
								assign node1105 = (inp[11]) ? node1113 : node1106;
									assign node1106 = (inp[5]) ? node1110 : node1107;
										assign node1107 = (inp[6]) ? 3'b110 : 3'b100;
										assign node1110 = (inp[2]) ? 3'b000 : 3'b100;
									assign node1113 = (inp[6]) ? 3'b100 : 3'b000;
							assign node1116 = (inp[1]) ? node1118 : 3'b000;
								assign node1118 = (inp[11]) ? node1120 : 3'b000;
									assign node1120 = (inp[8]) ? 3'b100 : 3'b000;

endmodule