module dtc_split75_bm98 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node19;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node48;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node147;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node164;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node202;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node235;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node244;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node256;
	wire [3-1:0] node258;
	wire [3-1:0] node260;
	wire [3-1:0] node263;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node302;
	wire [3-1:0] node304;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node330;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node341;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node350;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node358;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node383;
	wire [3-1:0] node384;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node392;
	wire [3-1:0] node395;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node402;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node413;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node418;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node436;
	wire [3-1:0] node439;
	wire [3-1:0] node441;
	wire [3-1:0] node444;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node456;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node461;
	wire [3-1:0] node465;
	wire [3-1:0] node467;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node474;
	wire [3-1:0] node477;
	wire [3-1:0] node478;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node486;
	wire [3-1:0] node487;
	wire [3-1:0] node488;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node509;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node518;
	wire [3-1:0] node519;
	wire [3-1:0] node522;
	wire [3-1:0] node524;
	wire [3-1:0] node526;
	wire [3-1:0] node529;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node538;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node542;
	wire [3-1:0] node545;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node552;
	wire [3-1:0] node554;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node564;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node578;
	wire [3-1:0] node581;
	wire [3-1:0] node582;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node588;
	wire [3-1:0] node591;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node597;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node604;
	wire [3-1:0] node607;
	wire [3-1:0] node610;
	wire [3-1:0] node611;
	wire [3-1:0] node613;
	wire [3-1:0] node616;
	wire [3-1:0] node618;
	wire [3-1:0] node619;
	wire [3-1:0] node622;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node631;
	wire [3-1:0] node632;
	wire [3-1:0] node633;
	wire [3-1:0] node634;
	wire [3-1:0] node636;
	wire [3-1:0] node640;
	wire [3-1:0] node642;
	wire [3-1:0] node643;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node650;
	wire [3-1:0] node653;
	wire [3-1:0] node654;
	wire [3-1:0] node657;
	wire [3-1:0] node660;
	wire [3-1:0] node661;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node680;
	wire [3-1:0] node683;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node689;
	wire [3-1:0] node691;
	wire [3-1:0] node695;
	wire [3-1:0] node696;
	wire [3-1:0] node697;
	wire [3-1:0] node699;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node710;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node719;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node725;
	wire [3-1:0] node728;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node735;
	wire [3-1:0] node736;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node744;
	wire [3-1:0] node745;
	wire [3-1:0] node748;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node763;
	wire [3-1:0] node766;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node772;
	wire [3-1:0] node775;
	wire [3-1:0] node777;
	wire [3-1:0] node778;
	wire [3-1:0] node782;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node797;
	wire [3-1:0] node798;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node808;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node814;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node834;

	assign outp = (inp[0]) ? node312 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b111;
			assign node3 = (inp[9]) ? node101 : node4;
				assign node4 = (inp[3]) ? node70 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b100;
						assign node7 = (inp[1]) ? node43 : node8;
							assign node8 = (inp[7]) ? node10 : 3'b100;
								assign node10 = (inp[5]) ? node22 : node11;
									assign node11 = (inp[2]) ? node17 : node12;
										assign node12 = (inp[11]) ? node14 : 3'b000;
											assign node14 = (inp[10]) ? 3'b100 : 3'b000;
										assign node17 = (inp[10]) ? node19 : 3'b100;
											assign node19 = (inp[11]) ? 3'b000 : 3'b100;
									assign node22 = (inp[2]) ? node28 : node23;
										assign node23 = (inp[10]) ? node25 : 3'b100;
											assign node25 = (inp[11]) ? 3'b000 : 3'b100;
										assign node28 = (inp[8]) ? node36 : node29;
											assign node29 = (inp[11]) ? node33 : node30;
												assign node30 = (inp[10]) ? 3'b000 : 3'b100;
												assign node33 = (inp[10]) ? 3'b100 : 3'b000;
											assign node36 = (inp[10]) ? node40 : node37;
												assign node37 = (inp[11]) ? 3'b000 : 3'b100;
												assign node40 = (inp[11]) ? 3'b100 : 3'b000;
							assign node43 = (inp[7]) ? node45 : 3'b000;
								assign node45 = (inp[2]) ? node57 : node46;
									assign node46 = (inp[10]) ? node48 : 3'b101;
										assign node48 = (inp[8]) ? node50 : 3'b101;
											assign node50 = (inp[11]) ? node54 : node51;
												assign node51 = (inp[5]) ? 3'b100 : 3'b101;
												assign node54 = (inp[5]) ? 3'b101 : 3'b100;
									assign node57 = (inp[10]) ? node63 : node58;
										assign node58 = (inp[11]) ? node60 : 3'b100;
											assign node60 = (inp[8]) ? 3'b101 : 3'b100;
										assign node63 = (inp[5]) ? node67 : node64;
											assign node64 = (inp[11]) ? 3'b101 : 3'b100;
											assign node67 = (inp[11]) ? 3'b100 : 3'b101;
					assign node70 = (inp[1]) ? node72 : 3'b010;
						assign node72 = (inp[7]) ? node74 : 3'b010;
							assign node74 = (inp[4]) ? node76 : 3'b010;
								assign node76 = (inp[5]) ? node88 : node77;
									assign node77 = (inp[2]) ? node83 : node78;
										assign node78 = (inp[11]) ? node80 : 3'b110;
											assign node80 = (inp[10]) ? 3'b010 : 3'b110;
										assign node83 = (inp[11]) ? node85 : 3'b010;
											assign node85 = (inp[10]) ? 3'b110 : 3'b010;
									assign node88 = (inp[11]) ? node96 : node89;
										assign node89 = (inp[10]) ? node93 : node90;
											assign node90 = (inp[2]) ? 3'b010 : 3'b110;
											assign node93 = (inp[2]) ? 3'b110 : 3'b010;
										assign node96 = (inp[10]) ? node98 : 3'b110;
											assign node98 = (inp[2]) ? 3'b010 : 3'b110;
				assign node101 = (inp[3]) ? node263 : node102;
					assign node102 = (inp[1]) ? node176 : node103;
						assign node103 = (inp[4]) ? node123 : node104;
							assign node104 = (inp[2]) ? node114 : node105;
								assign node105 = (inp[7]) ? 3'b001 : node106;
									assign node106 = (inp[11]) ? node110 : node107;
										assign node107 = (inp[5]) ? 3'b101 : 3'b001;
										assign node110 = (inp[5]) ? 3'b001 : 3'b101;
								assign node114 = (inp[7]) ? 3'b101 : node115;
									assign node115 = (inp[5]) ? node119 : node116;
										assign node116 = (inp[11]) ? 3'b101 : 3'b001;
										assign node119 = (inp[11]) ? 3'b001 : 3'b101;
							assign node123 = (inp[2]) ? node139 : node124;
								assign node124 = (inp[7]) ? node132 : node125;
									assign node125 = (inp[11]) ? 3'b101 : node126;
										assign node126 = (inp[8]) ? node128 : 3'b111;
											assign node128 = (inp[5]) ? 3'b111 : 3'b101;
									assign node132 = (inp[11]) ? node136 : node133;
										assign node133 = (inp[5]) ? 3'b111 : 3'b011;
										assign node136 = (inp[5]) ? 3'b011 : 3'b111;
								assign node139 = (inp[7]) ? node161 : node140;
									assign node140 = (inp[10]) ? node150 : node141;
										assign node141 = (inp[8]) ? node145 : node142;
											assign node142 = (inp[5]) ? 3'b011 : 3'b001;
											assign node145 = (inp[11]) ? node147 : 3'b111;
												assign node147 = (inp[5]) ? 3'b101 : 3'b111;
										assign node150 = (inp[8]) ? node154 : node151;
											assign node151 = (inp[11]) ? 3'b111 : 3'b101;
											assign node154 = (inp[11]) ? node158 : node155;
												assign node155 = (inp[5]) ? 3'b001 : 3'b011;
												assign node158 = (inp[5]) ? 3'b011 : 3'b001;
									assign node161 = (inp[11]) ? node169 : node162;
										assign node162 = (inp[8]) ? node164 : 3'b001;
											assign node164 = (inp[5]) ? node166 : 3'b101;
												assign node166 = (inp[10]) ? 3'b001 : 3'b101;
										assign node169 = (inp[8]) ? node171 : 3'b101;
											assign node171 = (inp[5]) ? node173 : 3'b001;
												assign node173 = (inp[10]) ? 3'b101 : 3'b001;
						assign node176 = (inp[4]) ? node202 : node177;
							assign node177 = (inp[2]) ? node193 : node178;
								assign node178 = (inp[7]) ? 3'b001 : node179;
									assign node179 = (inp[10]) ? node185 : node180;
										assign node180 = (inp[11]) ? node182 : 3'b001;
											assign node182 = (inp[5]) ? 3'b001 : 3'b100;
										assign node185 = (inp[11]) ? node189 : node186;
											assign node186 = (inp[5]) ? 3'b100 : 3'b001;
											assign node189 = (inp[5]) ? 3'b001 : 3'b100;
								assign node193 = (inp[7]) ? 3'b100 : node194;
									assign node194 = (inp[5]) ? node198 : node195;
										assign node195 = (inp[11]) ? 3'b100 : 3'b001;
										assign node198 = (inp[11]) ? 3'b001 : 3'b100;
							assign node202 = (inp[7]) ? node240 : node203;
								assign node203 = (inp[2]) ? node219 : node204;
									assign node204 = (inp[11]) ? node212 : node205;
										assign node205 = (inp[8]) ? node207 : 3'b110;
											assign node207 = (inp[10]) ? node209 : 3'b100;
												assign node209 = (inp[5]) ? 3'b110 : 3'b100;
										assign node212 = (inp[8]) ? node214 : 3'b100;
											assign node214 = (inp[5]) ? 3'b100 : node215;
												assign node215 = (inp[10]) ? 3'b110 : 3'b100;
									assign node219 = (inp[11]) ? node229 : node220;
										assign node220 = (inp[8]) ? node224 : node221;
											assign node221 = (inp[10]) ? 3'b100 : 3'b001;
											assign node224 = (inp[10]) ? node226 : 3'b110;
												assign node226 = (inp[5]) ? 3'b001 : 3'b011;
										assign node229 = (inp[5]) ? node235 : node230;
											assign node230 = (inp[10]) ? 3'b110 : node231;
												assign node231 = (inp[8]) ? 3'b110 : 3'b011;
											assign node235 = (inp[10]) ? node237 : 3'b100;
												assign node237 = (inp[8]) ? 3'b011 : 3'b110;
								assign node240 = (inp[11]) ? node250 : node241;
									assign node241 = (inp[5]) ? node247 : node242;
										assign node242 = (inp[8]) ? node244 : 3'b001;
											assign node244 = (inp[2]) ? 3'b110 : 3'b001;
										assign node247 = (inp[2]) ? 3'b001 : 3'b110;
									assign node250 = (inp[5]) ? node256 : node251;
										assign node251 = (inp[10]) ? node253 : 3'b110;
											assign node253 = (inp[2]) ? 3'b001 : 3'b110;
										assign node256 = (inp[2]) ? node258 : 3'b001;
											assign node258 = (inp[8]) ? node260 : 3'b110;
												assign node260 = (inp[10]) ? 3'b110 : 3'b001;
					assign node263 = (inp[1]) ? node265 : 3'b111;
						assign node265 = (inp[7]) ? node283 : node266;
							assign node266 = (inp[4]) ? node274 : node267;
								assign node267 = (inp[5]) ? node271 : node268;
									assign node268 = (inp[11]) ? 3'b011 : 3'b111;
									assign node271 = (inp[11]) ? 3'b111 : 3'b011;
								assign node274 = (inp[2]) ? node276 : 3'b001;
									assign node276 = (inp[8]) ? node280 : node277;
										assign node277 = (inp[10]) ? 3'b001 : 3'b111;
										assign node280 = (inp[10]) ? 3'b111 : 3'b011;
							assign node283 = (inp[4]) ? node287 : node284;
								assign node284 = (inp[2]) ? 3'b001 : 3'b101;
								assign node287 = (inp[2]) ? node301 : node288;
									assign node288 = (inp[10]) ? node294 : node289;
										assign node289 = (inp[11]) ? 3'b011 : node290;
											assign node290 = (inp[5]) ? 3'b011 : 3'b111;
										assign node294 = (inp[5]) ? node298 : node295;
											assign node295 = (inp[11]) ? 3'b011 : 3'b111;
											assign node298 = (inp[11]) ? 3'b111 : 3'b011;
									assign node301 = (inp[11]) ? node307 : node302;
										assign node302 = (inp[8]) ? node304 : 3'b101;
											assign node304 = (inp[5]) ? 3'b101 : 3'b001;
										assign node307 = (inp[10]) ? 3'b011 : node308;
											assign node308 = (inp[5]) ? 3'b101 : 3'b001;
		assign node312 = (inp[3]) ? node506 : node313;
			assign node313 = (inp[6]) ? node465 : node314;
				assign node314 = (inp[9]) ? node358 : node315;
					assign node315 = (inp[4]) ? node317 : 3'b010;
						assign node317 = (inp[1]) ? node355 : node318;
							assign node318 = (inp[7]) ? node320 : 3'b010;
								assign node320 = (inp[2]) ? node338 : node321;
									assign node321 = (inp[10]) ? node327 : node322;
										assign node322 = (inp[11]) ? node324 : 3'b000;
											assign node324 = (inp[5]) ? 3'b010 : 3'b000;
										assign node327 = (inp[8]) ? node333 : node328;
											assign node328 = (inp[5]) ? node330 : 3'b010;
												assign node330 = (inp[11]) ? 3'b000 : 3'b010;
											assign node333 = (inp[5]) ? 3'b010 : node334;
												assign node334 = (inp[11]) ? 3'b010 : 3'b000;
									assign node338 = (inp[5]) ? node344 : node339;
										assign node339 = (inp[11]) ? node341 : 3'b010;
											assign node341 = (inp[10]) ? 3'b000 : 3'b010;
										assign node344 = (inp[8]) ? node350 : node345;
											assign node345 = (inp[11]) ? 3'b010 : node346;
												assign node346 = (inp[10]) ? 3'b000 : 3'b010;
											assign node350 = (inp[10]) ? node352 : 3'b000;
												assign node352 = (inp[11]) ? 3'b010 : 3'b000;
							assign node355 = (inp[7]) ? 3'b010 : 3'b000;
					assign node358 = (inp[4]) ? node406 : node359;
						assign node359 = (inp[2]) ? node383 : node360;
							assign node360 = (inp[7]) ? 3'b000 : node361;
								assign node361 = (inp[10]) ? node375 : node362;
									assign node362 = (inp[8]) ? node368 : node363;
										assign node363 = (inp[5]) ? 3'b000 : node364;
											assign node364 = (inp[11]) ? 3'b010 : 3'b000;
										assign node368 = (inp[5]) ? node372 : node369;
											assign node369 = (inp[11]) ? 3'b010 : 3'b000;
											assign node372 = (inp[11]) ? 3'b000 : 3'b010;
									assign node375 = (inp[11]) ? node379 : node376;
										assign node376 = (inp[5]) ? 3'b010 : 3'b000;
										assign node379 = (inp[5]) ? 3'b000 : 3'b010;
							assign node383 = (inp[7]) ? 3'b010 : node384;
								assign node384 = (inp[10]) ? node398 : node385;
									assign node385 = (inp[1]) ? node391 : node386;
										assign node386 = (inp[11]) ? node388 : 3'b010;
											assign node388 = (inp[5]) ? 3'b000 : 3'b010;
										assign node391 = (inp[5]) ? node395 : node392;
											assign node392 = (inp[11]) ? 3'b010 : 3'b000;
											assign node395 = (inp[11]) ? 3'b000 : 3'b010;
									assign node398 = (inp[5]) ? node402 : node399;
										assign node399 = (inp[11]) ? 3'b010 : 3'b000;
										assign node402 = (inp[11]) ? 3'b000 : 3'b010;
						assign node406 = (inp[2]) ? node416 : node407;
							assign node407 = (inp[7]) ? node409 : 3'b010;
								assign node409 = (inp[5]) ? node413 : node410;
									assign node410 = (inp[11]) ? 3'b010 : 3'b000;
									assign node413 = (inp[11]) ? 3'b000 : 3'b010;
							assign node416 = (inp[1]) ? node444 : node417;
								assign node417 = (inp[11]) ? node429 : node418;
									assign node418 = (inp[8]) ? node424 : node419;
										assign node419 = (inp[10]) ? node421 : 3'b000;
											assign node421 = (inp[7]) ? 3'b000 : 3'b010;
										assign node424 = (inp[10]) ? node426 : 3'b010;
											assign node426 = (inp[7]) ? 3'b010 : 3'b000;
									assign node429 = (inp[10]) ? node439 : node430;
										assign node430 = (inp[8]) ? node434 : node431;
											assign node431 = (inp[7]) ? 3'b010 : 3'b000;
											assign node434 = (inp[7]) ? node436 : 3'b010;
												assign node436 = (inp[5]) ? 3'b000 : 3'b010;
										assign node439 = (inp[8]) ? node441 : 3'b010;
											assign node441 = (inp[5]) ? 3'b010 : 3'b000;
								assign node444 = (inp[7]) ? node452 : node445;
									assign node445 = (inp[8]) ? node449 : node446;
										assign node446 = (inp[10]) ? 3'b010 : 3'b000;
										assign node449 = (inp[10]) ? 3'b000 : 3'b010;
									assign node452 = (inp[8]) ? node456 : node453;
										assign node453 = (inp[11]) ? 3'b110 : 3'b100;
										assign node456 = (inp[10]) ? 3'b010 : node457;
											assign node457 = (inp[11]) ? node461 : node458;
												assign node458 = (inp[5]) ? 3'b110 : 3'b010;
												assign node461 = (inp[5]) ? 3'b000 : 3'b110;
				assign node465 = (inp[9]) ? node467 : 3'b000;
					assign node467 = (inp[4]) ? node469 : 3'b000;
						assign node469 = (inp[1]) ? node503 : node470;
							assign node470 = (inp[11]) ? node486 : node471;
								assign node471 = (inp[5]) ? node477 : node472;
									assign node472 = (inp[8]) ? node474 : 3'b010;
										assign node474 = (inp[2]) ? 3'b110 : 3'b010;
									assign node477 = (inp[2]) ? node481 : node478;
										assign node478 = (inp[10]) ? 3'b100 : 3'b110;
										assign node481 = (inp[10]) ? 3'b010 : node482;
											assign node482 = (inp[8]) ? 3'b110 : 3'b010;
								assign node486 = (inp[2]) ? node494 : node487;
									assign node487 = (inp[5]) ? node491 : node488;
										assign node488 = (inp[10]) ? 3'b100 : 3'b110;
										assign node491 = (inp[10]) ? 3'b010 : 3'b000;
									assign node494 = (inp[8]) ? node496 : 3'b100;
										assign node496 = (inp[10]) ? node500 : node497;
											assign node497 = (inp[5]) ? 3'b000 : 3'b100;
											assign node500 = (inp[5]) ? 3'b100 : 3'b000;
							assign node503 = (inp[7]) ? 3'b000 : 3'b100;
			assign node506 = (inp[9]) ? node626 : node507;
				assign node507 = (inp[1]) ? node569 : node508;
					assign node508 = (inp[6]) ? node532 : node509;
						assign node509 = (inp[4]) ? node511 : 3'b001;
							assign node511 = (inp[7]) ? node529 : node512;
								assign node512 = (inp[2]) ? node518 : node513;
									assign node513 = (inp[8]) ? 3'b011 : node514;
										assign node514 = (inp[11]) ? 3'b011 : 3'b111;
									assign node518 = (inp[11]) ? node522 : node519;
										assign node519 = (inp[8]) ? 3'b101 : 3'b011;
										assign node522 = (inp[8]) ? node524 : 3'b101;
											assign node524 = (inp[10]) ? node526 : 3'b011;
												assign node526 = (inp[5]) ? 3'b101 : 3'b011;
								assign node529 = (inp[2]) ? 3'b001 : 3'b101;
						assign node532 = (inp[7]) ? node536 : node533;
							assign node533 = (inp[4]) ? 3'b001 : 3'b000;
							assign node536 = (inp[4]) ? node538 : 3'b000;
								assign node538 = (inp[11]) ? node550 : node539;
									assign node539 = (inp[2]) ? node545 : node540;
										assign node540 = (inp[5]) ? node542 : 3'b100;
											assign node542 = (inp[10]) ? 3'b010 : 3'b100;
										assign node545 = (inp[10]) ? node547 : 3'b000;
											assign node547 = (inp[5]) ? 3'b100 : 3'b000;
									assign node550 = (inp[2]) ? node564 : node551;
										assign node551 = (inp[8]) ? node557 : node552;
											assign node552 = (inp[10]) ? node554 : 3'b100;
												assign node554 = (inp[5]) ? 3'b100 : 3'b010;
											assign node557 = (inp[10]) ? node561 : node558;
												assign node558 = (inp[5]) ? 3'b010 : 3'b100;
												assign node561 = (inp[5]) ? 3'b100 : 3'b010;
										assign node564 = (inp[10]) ? node566 : 3'b110;
											assign node566 = (inp[5]) ? 3'b010 : 3'b110;
					assign node569 = (inp[4]) ? node571 : 3'b000;
						assign node571 = (inp[7]) ? node601 : node572;
							assign node572 = (inp[6]) ? 3'b100 : node573;
								assign node573 = (inp[2]) ? node581 : node574;
									assign node574 = (inp[11]) ? node578 : node575;
										assign node575 = (inp[8]) ? 3'b001 : 3'b101;
										assign node578 = (inp[8]) ? 3'b101 : 3'b001;
									assign node581 = (inp[10]) ? node591 : node582;
										assign node582 = (inp[5]) ? node584 : 3'b110;
											assign node584 = (inp[8]) ? node588 : node585;
												assign node585 = (inp[11]) ? 3'b110 : 3'b001;
												assign node588 = (inp[11]) ? 3'b001 : 3'b110;
										assign node591 = (inp[8]) ? node593 : 3'b001;
											assign node593 = (inp[5]) ? node597 : node594;
												assign node594 = (inp[11]) ? 3'b001 : 3'b110;
												assign node597 = (inp[11]) ? 3'b110 : 3'b001;
							assign node601 = (inp[6]) ? 3'b000 : node602;
								assign node602 = (inp[2]) ? node610 : node603;
									assign node603 = (inp[11]) ? node607 : node604;
										assign node604 = (inp[5]) ? 3'b110 : 3'b010;
										assign node607 = (inp[5]) ? 3'b010 : 3'b110;
									assign node610 = (inp[11]) ? node616 : node611;
										assign node611 = (inp[8]) ? node613 : 3'b010;
											assign node613 = (inp[5]) ? 3'b010 : 3'b100;
										assign node616 = (inp[8]) ? node618 : 3'b100;
											assign node618 = (inp[10]) ? node622 : node619;
												assign node619 = (inp[5]) ? 3'b010 : 3'b100;
												assign node622 = (inp[5]) ? 3'b100 : 3'b010;
				assign node626 = (inp[6]) ? node732 : node627;
					assign node627 = (inp[1]) ? node629 : 3'b111;
						assign node629 = (inp[4]) ? node695 : node630;
							assign node630 = (inp[11]) ? node660 : node631;
								assign node631 = (inp[8]) ? node647 : node632;
									assign node632 = (inp[5]) ? node640 : node633;
										assign node633 = (inp[7]) ? 3'b110 : node634;
											assign node634 = (inp[2]) ? node636 : 3'b010;
												assign node636 = (inp[10]) ? 3'b010 : 3'b110;
										assign node640 = (inp[2]) ? node642 : 3'b010;
											assign node642 = (inp[7]) ? 3'b110 : node643;
												assign node643 = (inp[10]) ? 3'b010 : 3'b110;
									assign node647 = (inp[10]) ? node653 : node648;
										assign node648 = (inp[7]) ? node650 : 3'b001;
											assign node650 = (inp[2]) ? 3'b001 : 3'b101;
										assign node653 = (inp[5]) ? node657 : node654;
											assign node654 = (inp[7]) ? 3'b101 : 3'b001;
											assign node657 = (inp[2]) ? 3'b110 : 3'b010;
								assign node660 = (inp[8]) ? node676 : node661;
									assign node661 = (inp[10]) ? node671 : node662;
										assign node662 = (inp[5]) ? node666 : node663;
											assign node663 = (inp[7]) ? 3'b001 : 3'b101;
											assign node666 = (inp[2]) ? 3'b101 : node667;
												assign node667 = (inp[7]) ? 3'b101 : 3'b001;
										assign node671 = (inp[2]) ? 3'b001 : node672;
											assign node672 = (inp[7]) ? 3'b101 : 3'b001;
									assign node676 = (inp[7]) ? node688 : node677;
										assign node677 = (inp[2]) ? node683 : node678;
											assign node678 = (inp[5]) ? node680 : 3'b001;
												assign node680 = (inp[10]) ? 3'b001 : 3'b010;
											assign node683 = (inp[10]) ? node685 : 3'b001;
												assign node685 = (inp[5]) ? 3'b101 : 3'b110;
										assign node688 = (inp[5]) ? 3'b110 : node689;
											assign node689 = (inp[10]) ? node691 : 3'b001;
												assign node691 = (inp[2]) ? 3'b110 : 3'b010;
							assign node695 = (inp[7]) ? node713 : node696;
								assign node696 = (inp[11]) ? node704 : node697;
									assign node697 = (inp[8]) ? node699 : 3'b011;
										assign node699 = (inp[10]) ? node701 : 3'b111;
											assign node701 = (inp[5]) ? 3'b011 : 3'b111;
									assign node704 = (inp[8]) ? node706 : 3'b111;
										assign node706 = (inp[5]) ? node710 : node707;
											assign node707 = (inp[10]) ? 3'b011 : 3'b111;
											assign node710 = (inp[10]) ? 3'b111 : 3'b011;
								assign node713 = (inp[2]) ? node723 : node714;
									assign node714 = (inp[8]) ? 3'b001 : node715;
										assign node715 = (inp[11]) ? node719 : node716;
											assign node716 = (inp[5]) ? 3'b001 : 3'b011;
											assign node719 = (inp[5]) ? 3'b011 : 3'b001;
									assign node723 = (inp[8]) ? 3'b101 : node724;
										assign node724 = (inp[11]) ? node728 : node725;
											assign node725 = (inp[5]) ? 3'b101 : 3'b011;
											assign node728 = (inp[5]) ? 3'b011 : 3'b101;
					assign node732 = (inp[1]) ? node782 : node733;
						assign node733 = (inp[7]) ? node751 : node734;
							assign node734 = (inp[4]) ? node742 : node735;
								assign node735 = (inp[5]) ? node739 : node736;
									assign node736 = (inp[11]) ? 3'b001 : 3'b101;
									assign node739 = (inp[11]) ? 3'b101 : 3'b001;
								assign node742 = (inp[2]) ? node744 : 3'b010;
									assign node744 = (inp[10]) ? node748 : node745;
										assign node745 = (inp[8]) ? 3'b001 : 3'b101;
										assign node748 = (inp[8]) ? 3'b101 : 3'b010;
							assign node751 = (inp[4]) ? node755 : node752;
								assign node752 = (inp[2]) ? 3'b010 : 3'b110;
								assign node755 = (inp[2]) ? node769 : node756;
									assign node756 = (inp[10]) ? node762 : node757;
										assign node757 = (inp[5]) ? node759 : 3'b001;
											assign node759 = (inp[11]) ? 3'b101 : 3'b001;
										assign node762 = (inp[11]) ? node766 : node763;
											assign node763 = (inp[5]) ? 3'b001 : 3'b101;
											assign node766 = (inp[5]) ? 3'b101 : 3'b001;
									assign node769 = (inp[11]) ? node775 : node770;
										assign node770 = (inp[10]) ? node772 : 3'b010;
											assign node772 = (inp[5]) ? 3'b110 : 3'b010;
										assign node775 = (inp[8]) ? node777 : 3'b001;
											assign node777 = (inp[5]) ? 3'b001 : node778;
												assign node778 = (inp[10]) ? 3'b110 : 3'b010;
						assign node782 = (inp[7]) ? node804 : node783;
							assign node783 = (inp[4]) ? node791 : node784;
								assign node784 = (inp[11]) ? node788 : node785;
									assign node785 = (inp[5]) ? 3'b010 : 3'b110;
									assign node788 = (inp[5]) ? 3'b110 : 3'b010;
								assign node791 = (inp[2]) ? node797 : node792;
									assign node792 = (inp[8]) ? 3'b000 : node793;
										assign node793 = (inp[10]) ? 3'b001 : 3'b000;
									assign node797 = (inp[10]) ? node801 : node798;
										assign node798 = (inp[8]) ? 3'b010 : 3'b110;
										assign node801 = (inp[8]) ? 3'b110 : 3'b001;
							assign node804 = (inp[4]) ? node808 : node805;
								assign node805 = (inp[2]) ? 3'b000 : 3'b100;
								assign node808 = (inp[2]) ? node822 : node809;
									assign node809 = (inp[10]) ? node817 : node810;
										assign node810 = (inp[11]) ? node814 : node811;
											assign node811 = (inp[5]) ? 3'b010 : 3'b110;
											assign node814 = (inp[5]) ? 3'b110 : 3'b010;
										assign node817 = (inp[11]) ? node819 : 3'b110;
											assign node819 = (inp[5]) ? 3'b110 : 3'b010;
									assign node822 = (inp[11]) ? node828 : node823;
										assign node823 = (inp[8]) ? node825 : 3'b100;
											assign node825 = (inp[10]) ? 3'b100 : 3'b000;
										assign node828 = (inp[8]) ? node830 : 3'b010;
											assign node830 = (inp[5]) ? node834 : node831;
												assign node831 = (inp[10]) ? 3'b100 : 3'b000;
												assign node834 = (inp[10]) ? 3'b010 : 3'b100;

endmodule