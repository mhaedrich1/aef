module dtc_split875_bm11 (
	input  wire [7-1:0] inp,
	output wire [1-1:0] outp
);

	wire [1-1:0] node1;
	wire [1-1:0] node2;
	wire [1-1:0] node4;
	wire [1-1:0] node5;
	wire [1-1:0] node7;
	wire [1-1:0] node9;
	wire [1-1:0] node12;
	wire [1-1:0] node13;
	wire [1-1:0] node15;
	wire [1-1:0] node18;
	wire [1-1:0] node19;
	wire [1-1:0] node23;
	wire [1-1:0] node24;
	wire [1-1:0] node26;
	wire [1-1:0] node27;
	wire [1-1:0] node29;
	wire [1-1:0] node33;
	wire [1-1:0] node34;
	wire [1-1:0] node35;
	wire [1-1:0] node37;
	wire [1-1:0] node40;
	wire [1-1:0] node41;
	wire [1-1:0] node45;
	wire [1-1:0] node46;
	wire [1-1:0] node47;
	wire [1-1:0] node52;
	wire [1-1:0] node53;
	wire [1-1:0] node54;
	wire [1-1:0] node55;
	wire [1-1:0] node57;
	wire [1-1:0] node59;
	wire [1-1:0] node62;
	wire [1-1:0] node63;
	wire [1-1:0] node65;
	wire [1-1:0] node69;
	wire [1-1:0] node70;
	wire [1-1:0] node71;
	wire [1-1:0] node73;
	wire [1-1:0] node76;
	wire [1-1:0] node77;
	wire [1-1:0] node81;
	wire [1-1:0] node82;
	wire [1-1:0] node83;
	wire [1-1:0] node88;
	wire [1-1:0] node89;
	wire [1-1:0] node90;
	wire [1-1:0] node92;
	wire [1-1:0] node93;

	assign outp = (inp[1]) ? node52 : node1;
		assign node1 = (inp[6]) ? node23 : node2;
			assign node2 = (inp[3]) ? node4 : 1'b1;
				assign node4 = (inp[0]) ? node12 : node5;
					assign node5 = (inp[4]) ? node7 : 1'b1;
						assign node7 = (inp[5]) ? node9 : 1'b1;
							assign node9 = (inp[2]) ? 1'b0 : 1'b1;
					assign node12 = (inp[4]) ? node18 : node13;
						assign node13 = (inp[2]) ? node15 : 1'b1;
							assign node15 = (inp[5]) ? 1'b0 : 1'b1;
						assign node18 = (inp[5]) ? 1'b0 : node19;
							assign node19 = (inp[2]) ? 1'b0 : 1'b1;
			assign node23 = (inp[2]) ? node33 : node24;
				assign node24 = (inp[4]) ? node26 : 1'b1;
					assign node26 = (inp[5]) ? 1'b0 : node27;
						assign node27 = (inp[0]) ? node29 : 1'b1;
							assign node29 = (inp[3]) ? 1'b0 : 1'b1;
				assign node33 = (inp[0]) ? node45 : node34;
					assign node34 = (inp[3]) ? node40 : node35;
						assign node35 = (inp[4]) ? node37 : 1'b1;
							assign node37 = (inp[5]) ? 1'b0 : 1'b1;
						assign node40 = (inp[5]) ? 1'b0 : node41;
							assign node41 = (inp[4]) ? 1'b0 : 1'b1;
					assign node45 = (inp[4]) ? 1'b0 : node46;
						assign node46 = (inp[5]) ? 1'b0 : node47;
							assign node47 = (inp[3]) ? 1'b0 : 1'b1;
		assign node52 = (inp[2]) ? node88 : node53;
			assign node53 = (inp[4]) ? node69 : node54;
				assign node54 = (inp[5]) ? node62 : node55;
					assign node55 = (inp[3]) ? node57 : 1'b1;
						assign node57 = (inp[0]) ? node59 : 1'b1;
							assign node59 = (inp[6]) ? 1'b0 : 1'b1;
					assign node62 = (inp[3]) ? 1'b0 : node63;
						assign node63 = (inp[6]) ? node65 : 1'b1;
							assign node65 = (inp[0]) ? 1'b0 : 1'b1;
				assign node69 = (inp[6]) ? node81 : node70;
					assign node70 = (inp[0]) ? node76 : node71;
						assign node71 = (inp[3]) ? node73 : 1'b1;
							assign node73 = (inp[5]) ? 1'b0 : 1'b1;
						assign node76 = (inp[5]) ? 1'b0 : node77;
							assign node77 = (inp[3]) ? 1'b0 : 1'b1;
					assign node81 = (inp[3]) ? 1'b0 : node82;
						assign node82 = (inp[0]) ? 1'b0 : node83;
							assign node83 = (inp[5]) ? 1'b0 : 1'b1;
			assign node88 = (inp[4]) ? 1'b0 : node89;
				assign node89 = (inp[0]) ? 1'b0 : node90;
					assign node90 = (inp[3]) ? node92 : 1'b1;
						assign node92 = (inp[5]) ? 1'b0 : node93;
							assign node93 = (inp[6]) ? 1'b0 : 1'b1;

endmodule