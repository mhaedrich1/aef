module dtc_split75_bm87 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node73;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node117;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node163;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node228;
	wire [3-1:0] node232;
	wire [3-1:0] node233;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node261;
	wire [3-1:0] node266;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node277;
	wire [3-1:0] node279;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node296;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node312;
	wire [3-1:0] node315;
	wire [3-1:0] node317;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node326;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node334;
	wire [3-1:0] node335;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node349;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node355;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node366;
	wire [3-1:0] node368;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node376;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node383;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node389;
	wire [3-1:0] node392;
	wire [3-1:0] node393;
	wire [3-1:0] node394;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node403;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node423;
	wire [3-1:0] node427;
	wire [3-1:0] node428;
	wire [3-1:0] node429;
	wire [3-1:0] node431;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node446;
	wire [3-1:0] node447;
	wire [3-1:0] node448;
	wire [3-1:0] node449;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node464;
	wire [3-1:0] node465;
	wire [3-1:0] node467;
	wire [3-1:0] node471;
	wire [3-1:0] node472;
	wire [3-1:0] node473;
	wire [3-1:0] node474;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node478;
	wire [3-1:0] node479;
	wire [3-1:0] node483;
	wire [3-1:0] node485;
	wire [3-1:0] node486;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node496;
	wire [3-1:0] node498;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node504;
	wire [3-1:0] node505;
	wire [3-1:0] node507;
	wire [3-1:0] node508;
	wire [3-1:0] node512;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node519;
	wire [3-1:0] node520;
	wire [3-1:0] node521;
	wire [3-1:0] node525;
	wire [3-1:0] node526;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node535;
	wire [3-1:0] node536;
	wire [3-1:0] node540;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node545;
	wire [3-1:0] node547;
	wire [3-1:0] node550;
	wire [3-1:0] node552;
	wire [3-1:0] node553;
	wire [3-1:0] node557;
	wire [3-1:0] node558;
	wire [3-1:0] node560;
	wire [3-1:0] node561;
	wire [3-1:0] node565;
	wire [3-1:0] node567;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node572;
	wire [3-1:0] node573;
	wire [3-1:0] node575;
	wire [3-1:0] node579;
	wire [3-1:0] node580;
	wire [3-1:0] node584;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node592;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node598;
	wire [3-1:0] node599;
	wire [3-1:0] node600;
	wire [3-1:0] node601;
	wire [3-1:0] node605;
	wire [3-1:0] node606;
	wire [3-1:0] node607;
	wire [3-1:0] node612;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node623;
	wire [3-1:0] node625;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node652;
	wire [3-1:0] node653;
	wire [3-1:0] node657;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node666;
	wire [3-1:0] node669;
	wire [3-1:0] node671;
	wire [3-1:0] node674;
	wire [3-1:0] node675;
	wire [3-1:0] node677;
	wire [3-1:0] node680;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node693;
	wire [3-1:0] node694;
	wire [3-1:0] node698;
	wire [3-1:0] node700;
	wire [3-1:0] node703;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node710;
	wire [3-1:0] node711;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node716;
	wire [3-1:0] node717;
	wire [3-1:0] node719;
	wire [3-1:0] node723;
	wire [3-1:0] node724;
	wire [3-1:0] node727;
	wire [3-1:0] node729;
	wire [3-1:0] node732;
	wire [3-1:0] node733;
	wire [3-1:0] node735;
	wire [3-1:0] node737;
	wire [3-1:0] node739;
	wire [3-1:0] node742;
	wire [3-1:0] node743;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node749;
	wire [3-1:0] node750;
	wire [3-1:0] node752;
	wire [3-1:0] node756;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node763;
	wire [3-1:0] node764;
	wire [3-1:0] node765;
	wire [3-1:0] node767;
	wire [3-1:0] node769;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node778;
	wire [3-1:0] node779;
	wire [3-1:0] node780;
	wire [3-1:0] node781;
	wire [3-1:0] node784;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node793;
	wire [3-1:0] node795;
	wire [3-1:0] node796;
	wire [3-1:0] node799;
	wire [3-1:0] node802;
	wire [3-1:0] node803;
	wire [3-1:0] node806;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node813;
	wire [3-1:0] node816;
	wire [3-1:0] node817;
	wire [3-1:0] node819;
	wire [3-1:0] node820;
	wire [3-1:0] node821;
	wire [3-1:0] node823;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node834;
	wire [3-1:0] node835;
	wire [3-1:0] node837;
	wire [3-1:0] node841;
	wire [3-1:0] node842;
	wire [3-1:0] node844;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node850;
	wire [3-1:0] node852;
	wire [3-1:0] node857;
	wire [3-1:0] node858;
	wire [3-1:0] node860;
	wire [3-1:0] node861;
	wire [3-1:0] node865;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node872;
	wire [3-1:0] node873;
	wire [3-1:0] node874;
	wire [3-1:0] node875;
	wire [3-1:0] node881;
	wire [3-1:0] node882;
	wire [3-1:0] node884;
	wire [3-1:0] node888;
	wire [3-1:0] node889;
	wire [3-1:0] node890;
	wire [3-1:0] node892;
	wire [3-1:0] node895;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node903;
	wire [3-1:0] node904;
	wire [3-1:0] node905;
	wire [3-1:0] node906;
	wire [3-1:0] node909;
	wire [3-1:0] node912;
	wire [3-1:0] node913;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node924;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node931;
	wire [3-1:0] node935;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node939;
	wire [3-1:0] node942;
	wire [3-1:0] node944;
	wire [3-1:0] node947;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node959;
	wire [3-1:0] node960;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node964;
	wire [3-1:0] node968;
	wire [3-1:0] node970;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node975;
	wire [3-1:0] node981;
	wire [3-1:0] node982;
	wire [3-1:0] node983;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node988;
	wire [3-1:0] node991;
	wire [3-1:0] node992;
	wire [3-1:0] node994;
	wire [3-1:0] node998;
	wire [3-1:0] node999;
	wire [3-1:0] node1001;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1009;
	wire [3-1:0] node1010;
	wire [3-1:0] node1011;
	wire [3-1:0] node1014;
	wire [3-1:0] node1017;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1024;
	wire [3-1:0] node1026;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1031;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1039;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1043;
	wire [3-1:0] node1047;
	wire [3-1:0] node1048;

	assign outp = (inp[6]) ? node220 : node1;
		assign node1 = (inp[7]) ? node33 : node2;
			assign node2 = (inp[1]) ? 3'b000 : node3;
				assign node3 = (inp[0]) ? node5 : 3'b000;
					assign node5 = (inp[8]) ? node7 : 3'b000;
						assign node7 = (inp[10]) ? 3'b000 : node8;
							assign node8 = (inp[9]) ? 3'b000 : node9;
								assign node9 = (inp[4]) ? node17 : node10;
									assign node10 = (inp[11]) ? node14 : node11;
										assign node11 = (inp[2]) ? 3'b000 : 3'b100;
										assign node14 = (inp[2]) ? 3'b100 : 3'b000;
									assign node17 = (inp[3]) ? node23 : node18;
										assign node18 = (inp[11]) ? node20 : 3'b100;
											assign node20 = (inp[2]) ? 3'b100 : 3'b000;
										assign node23 = (inp[11]) ? node27 : node24;
											assign node24 = (inp[2]) ? 3'b000 : 3'b100;
											assign node27 = (inp[2]) ? 3'b100 : 3'b000;
			assign node33 = (inp[9]) ? node191 : node34;
				assign node34 = (inp[0]) ? node106 : node35;
					assign node35 = (inp[10]) ? node77 : node36;
						assign node36 = (inp[1]) ? node40 : node37;
							assign node37 = (inp[11]) ? 3'b001 : 3'b101;
							assign node40 = (inp[8]) ? node56 : node41;
								assign node41 = (inp[11]) ? node49 : node42;
									assign node42 = (inp[2]) ? node44 : 3'b110;
										assign node44 = (inp[4]) ? 3'b010 : node45;
											assign node45 = (inp[3]) ? 3'b010 : 3'b110;
									assign node49 = (inp[2]) ? node51 : 3'b010;
										assign node51 = (inp[4]) ? 3'b110 : node52;
											assign node52 = (inp[3]) ? 3'b110 : 3'b010;
								assign node56 = (inp[11]) ? node70 : node57;
									assign node57 = (inp[4]) ? 3'b001 : node58;
										assign node58 = (inp[2]) ? node64 : node59;
											assign node59 = (inp[5]) ? 3'b001 : node60;
												assign node60 = (inp[3]) ? 3'b001 : 3'b101;
											assign node64 = (inp[3]) ? 3'b110 : node65;
												assign node65 = (inp[5]) ? 3'b110 : 3'b001;
									assign node70 = (inp[5]) ? node72 : 3'b110;
										assign node72 = (inp[4]) ? 3'b110 : node73;
											assign node73 = (inp[2]) ? 3'b010 : 3'b110;
						assign node77 = (inp[1]) ? node79 : 3'b110;
							assign node79 = (inp[8]) ? node83 : node80;
								assign node80 = (inp[11]) ? 3'b000 : 3'b100;
								assign node83 = (inp[3]) ? node97 : node84;
									assign node84 = (inp[11]) ? node94 : node85;
										assign node85 = (inp[4]) ? 3'b010 : node86;
											assign node86 = (inp[5]) ? node90 : node87;
												assign node87 = (inp[2]) ? 3'b010 : 3'b110;
												assign node90 = (inp[2]) ? 3'b110 : 3'b010;
										assign node94 = (inp[4]) ? 3'b100 : 3'b010;
									assign node97 = (inp[4]) ? 3'b100 : node98;
										assign node98 = (inp[5]) ? node102 : node99;
											assign node99 = (inp[11]) ? 3'b110 : 3'b010;
											assign node102 = (inp[2]) ? 3'b000 : 3'b100;
					assign node106 = (inp[10]) ? node178 : node107;
						assign node107 = (inp[1]) ? node147 : node108;
							assign node108 = (inp[11]) ? node124 : node109;
								assign node109 = (inp[8]) ? node117 : node110;
									assign node110 = (inp[2]) ? node112 : 3'b010;
										assign node112 = (inp[4]) ? 3'b100 : node113;
											assign node113 = (inp[3]) ? 3'b100 : 3'b010;
									assign node117 = (inp[2]) ? node119 : 3'b110;
										assign node119 = (inp[4]) ? 3'b010 : node120;
											assign node120 = (inp[3]) ? 3'b010 : 3'b110;
								assign node124 = (inp[5]) ? node138 : node125;
									assign node125 = (inp[8]) ? node133 : node126;
										assign node126 = (inp[2]) ? node128 : 3'b100;
											assign node128 = (inp[4]) ? 3'b010 : node129;
												assign node129 = (inp[3]) ? 3'b010 : 3'b100;
										assign node133 = (inp[2]) ? node135 : 3'b010;
											assign node135 = (inp[4]) ? 3'b100 : 3'b010;
									assign node138 = (inp[8]) ? node144 : node139;
										assign node139 = (inp[2]) ? node141 : 3'b100;
											assign node141 = (inp[4]) ? 3'b010 : 3'b100;
										assign node144 = (inp[2]) ? 3'b100 : 3'b010;
							assign node147 = (inp[8]) ? node155 : node148;
								assign node148 = (inp[2]) ? 3'b000 : node149;
									assign node149 = (inp[11]) ? 3'b000 : node150;
										assign node150 = (inp[3]) ? 3'b000 : 3'b100;
								assign node155 = (inp[11]) ? node167 : node156;
									assign node156 = (inp[2]) ? 3'b100 : node157;
										assign node157 = (inp[3]) ? node163 : node158;
											assign node158 = (inp[4]) ? 3'b010 : node159;
												assign node159 = (inp[5]) ? 3'b100 : 3'b010;
											assign node163 = (inp[4]) ? 3'b100 : 3'b010;
									assign node167 = (inp[2]) ? node173 : node168;
										assign node168 = (inp[3]) ? node170 : 3'b100;
											assign node170 = (inp[4]) ? 3'b000 : 3'b100;
										assign node173 = (inp[4]) ? 3'b000 : node174;
											assign node174 = (inp[5]) ? 3'b100 : 3'b000;
						assign node178 = (inp[8]) ? node180 : 3'b000;
							assign node180 = (inp[11]) ? 3'b000 : node181;
								assign node181 = (inp[1]) ? 3'b000 : node182;
									assign node182 = (inp[2]) ? node184 : 3'b100;
										assign node184 = (inp[4]) ? 3'b000 : node185;
											assign node185 = (inp[3]) ? 3'b000 : 3'b100;
				assign node191 = (inp[10]) ? 3'b000 : node192;
					assign node192 = (inp[0]) ? 3'b000 : node193;
						assign node193 = (inp[1]) ? node201 : node194;
							assign node194 = (inp[2]) ? node198 : node195;
								assign node195 = (inp[11]) ? 3'b110 : 3'b010;
								assign node198 = (inp[11]) ? 3'b000 : 3'b100;
							assign node201 = (inp[8]) ? node203 : 3'b000;
								assign node203 = (inp[11]) ? node213 : node204;
									assign node204 = (inp[3]) ? node208 : node205;
										assign node205 = (inp[2]) ? 3'b000 : 3'b100;
										assign node208 = (inp[4]) ? node210 : 3'b000;
											assign node210 = (inp[2]) ? 3'b100 : 3'b000;
									assign node213 = (inp[3]) ? 3'b100 : node214;
										assign node214 = (inp[4]) ? 3'b000 : 3'b100;
		assign node220 = (inp[9]) ? node710 : node221;
			assign node221 = (inp[0]) ? node471 : node222;
				assign node222 = (inp[7]) ? node392 : node223;
					assign node223 = (inp[10]) ? node305 : node224;
						assign node224 = (inp[1]) ? node256 : node225;
							assign node225 = (inp[11]) ? node241 : node226;
								assign node226 = (inp[8]) ? node232 : node227;
									assign node227 = (inp[2]) ? 3'b011 : node228;
										assign node228 = (inp[3]) ? 3'b011 : 3'b111;
									assign node232 = (inp[2]) ? 3'b111 : node233;
										assign node233 = (inp[3]) ? node235 : 3'b011;
											assign node235 = (inp[5]) ? 3'b111 : node236;
												assign node236 = (inp[4]) ? 3'b111 : 3'b011;
								assign node241 = (inp[8]) ? node247 : node242;
									assign node242 = (inp[2]) ? 3'b101 : node243;
										assign node243 = (inp[3]) ? 3'b101 : 3'b001;
									assign node247 = (inp[2]) ? 3'b011 : node248;
										assign node248 = (inp[3]) ? node250 : 3'b111;
											assign node250 = (inp[5]) ? 3'b011 : node251;
												assign node251 = (inp[4]) ? 3'b011 : 3'b111;
							assign node256 = (inp[11]) ? node282 : node257;
								assign node257 = (inp[8]) ? node271 : node258;
									assign node258 = (inp[3]) ? node266 : node259;
										assign node259 = (inp[4]) ? 3'b101 : node260;
											assign node260 = (inp[2]) ? 3'b101 : node261;
												assign node261 = (inp[5]) ? 3'b110 : 3'b010;
										assign node266 = (inp[2]) ? node268 : 3'b101;
											assign node268 = (inp[5]) ? 3'b001 : 3'b101;
									assign node271 = (inp[3]) ? node277 : node272;
										assign node272 = (inp[2]) ? 3'b011 : node273;
											assign node273 = (inp[4]) ? 3'b011 : 3'b101;
										assign node277 = (inp[2]) ? node279 : 3'b011;
											assign node279 = (inp[4]) ? 3'b101 : 3'b011;
								assign node282 = (inp[8]) ? node294 : node283;
									assign node283 = (inp[3]) ? node289 : node284;
										assign node284 = (inp[2]) ? 3'b001 : node285;
											assign node285 = (inp[5]) ? 3'b001 : 3'b101;
										assign node289 = (inp[5]) ? node291 : 3'b001;
											assign node291 = (inp[2]) ? 3'b110 : 3'b001;
									assign node294 = (inp[2]) ? node300 : node295;
										assign node295 = (inp[3]) ? 3'b101 : node296;
											assign node296 = (inp[4]) ? 3'b101 : 3'b011;
										assign node300 = (inp[3]) ? node302 : 3'b101;
											assign node302 = (inp[4]) ? 3'b001 : 3'b101;
						assign node305 = (inp[1]) ? node347 : node306;
							assign node306 = (inp[8]) ? node334 : node307;
								assign node307 = (inp[11]) ? node321 : node308;
									assign node308 = (inp[2]) ? 3'b001 : node309;
										assign node309 = (inp[5]) ? node315 : node310;
											assign node310 = (inp[3]) ? node312 : 3'b101;
												assign node312 = (inp[4]) ? 3'b001 : 3'b101;
											assign node315 = (inp[4]) ? node317 : 3'b001;
												assign node317 = (inp[3]) ? 3'b001 : 3'b101;
									assign node321 = (inp[5]) ? node325 : node322;
										assign node322 = (inp[2]) ? 3'b101 : 3'b001;
										assign node325 = (inp[2]) ? node331 : node326;
											assign node326 = (inp[3]) ? node328 : 3'b001;
												assign node328 = (inp[4]) ? 3'b110 : 3'b000;
											assign node331 = (inp[4]) ? 3'b110 : 3'b010;
								assign node334 = (inp[2]) ? node340 : node335;
									assign node335 = (inp[11]) ? node337 : 3'b011;
										assign node337 = (inp[3]) ? 3'b001 : 3'b101;
									assign node340 = (inp[11]) ? node342 : 3'b101;
										assign node342 = (inp[4]) ? node344 : 3'b001;
											assign node344 = (inp[5]) ? 3'b001 : 3'b011;
							assign node347 = (inp[8]) ? node371 : node348;
								assign node348 = (inp[11]) ? node360 : node349;
									assign node349 = (inp[2]) ? node355 : node350;
										assign node350 = (inp[4]) ? 3'b110 : node351;
											assign node351 = (inp[3]) ? 3'b110 : 3'b001;
										assign node355 = (inp[4]) ? node357 : 3'b110;
											assign node357 = (inp[3]) ? 3'b010 : 3'b110;
									assign node360 = (inp[4]) ? node366 : node361;
										assign node361 = (inp[2]) ? 3'b010 : node362;
											assign node362 = (inp[3]) ? 3'b010 : 3'b110;
										assign node366 = (inp[2]) ? node368 : 3'b010;
											assign node368 = (inp[3]) ? 3'b100 : 3'b010;
								assign node371 = (inp[11]) ? node379 : node372;
									assign node372 = (inp[3]) ? node374 : 3'b001;
										assign node374 = (inp[2]) ? node376 : 3'b001;
											assign node376 = (inp[4]) ? 3'b110 : 3'b001;
									assign node379 = (inp[4]) ? node383 : node380;
										assign node380 = (inp[2]) ? 3'b110 : 3'b010;
										assign node383 = (inp[3]) ? node385 : 3'b001;
											assign node385 = (inp[5]) ? node389 : node386;
												assign node386 = (inp[2]) ? 3'b001 : 3'b101;
												assign node389 = (inp[2]) ? 3'b010 : 3'b110;
					assign node392 = (inp[10]) ? node414 : node393;
						assign node393 = (inp[8]) ? 3'b111 : node394;
							assign node394 = (inp[1]) ? node396 : 3'b111;
								assign node396 = (inp[11]) ? node406 : node397;
									assign node397 = (inp[5]) ? node403 : node398;
										assign node398 = (inp[4]) ? 3'b111 : node399;
											assign node399 = (inp[2]) ? 3'b111 : 3'b011;
										assign node403 = (inp[4]) ? 3'b011 : 3'b111;
									assign node406 = (inp[2]) ? 3'b011 : node407;
										assign node407 = (inp[3]) ? 3'b011 : node408;
											assign node408 = (inp[4]) ? 3'b011 : 3'b111;
						assign node414 = (inp[1]) ? node446 : node415;
							assign node415 = (inp[2]) ? node427 : node416;
								assign node416 = (inp[8]) ? 3'b111 : node417;
									assign node417 = (inp[11]) ? node419 : 3'b111;
										assign node419 = (inp[5]) ? node421 : 3'b011;
											assign node421 = (inp[3]) ? node423 : 3'b011;
												assign node423 = (inp[4]) ? 3'b101 : 3'b001;
								assign node427 = (inp[4]) ? node437 : node428;
									assign node428 = (inp[8]) ? node434 : node429;
										assign node429 = (inp[11]) ? node431 : 3'b011;
											assign node431 = (inp[5]) ? 3'b001 : 3'b011;
										assign node434 = (inp[11]) ? 3'b011 : 3'b111;
									assign node437 = (inp[11]) ? node441 : node438;
										assign node438 = (inp[8]) ? 3'b111 : 3'b011;
										assign node441 = (inp[8]) ? 3'b011 : node442;
											assign node442 = (inp[5]) ? 3'b101 : 3'b111;
							assign node446 = (inp[11]) ? node458 : node447;
								assign node447 = (inp[8]) ? node453 : node448;
									assign node448 = (inp[3]) ? 3'b101 : node449;
										assign node449 = (inp[2]) ? 3'b101 : 3'b011;
									assign node453 = (inp[2]) ? 3'b011 : node454;
										assign node454 = (inp[3]) ? 3'b011 : 3'b111;
								assign node458 = (inp[8]) ? node464 : node459;
									assign node459 = (inp[2]) ? 3'b001 : node460;
										assign node460 = (inp[3]) ? 3'b001 : 3'b101;
									assign node464 = (inp[2]) ? 3'b101 : node465;
										assign node465 = (inp[3]) ? node467 : 3'b001;
											assign node467 = (inp[4]) ? 3'b101 : 3'b001;
				assign node471 = (inp[7]) ? node595 : node472;
					assign node472 = (inp[10]) ? node540 : node473;
						assign node473 = (inp[8]) ? node503 : node474;
							assign node474 = (inp[1]) ? node490 : node475;
								assign node475 = (inp[11]) ? node483 : node476;
									assign node476 = (inp[2]) ? node478 : 3'b001;
										assign node478 = (inp[4]) ? 3'b110 : node479;
											assign node479 = (inp[3]) ? 3'b110 : 3'b001;
									assign node483 = (inp[2]) ? node485 : 3'b110;
										assign node485 = (inp[4]) ? 3'b010 : node486;
											assign node486 = (inp[3]) ? 3'b010 : 3'b110;
								assign node490 = (inp[11]) ? node496 : node491;
									assign node491 = (inp[2]) ? 3'b010 : node492;
										assign node492 = (inp[4]) ? 3'b010 : 3'b110;
									assign node496 = (inp[2]) ? node498 : 3'b010;
										assign node498 = (inp[4]) ? node500 : 3'b100;
											assign node500 = (inp[5]) ? 3'b100 : 3'b010;
							assign node503 = (inp[1]) ? node519 : node504;
								assign node504 = (inp[11]) ? node512 : node505;
									assign node505 = (inp[2]) ? node507 : 3'b101;
										assign node507 = (inp[4]) ? 3'b001 : node508;
											assign node508 = (inp[3]) ? 3'b001 : 3'b101;
									assign node512 = (inp[2]) ? node514 : 3'b001;
										assign node514 = (inp[3]) ? 3'b110 : node515;
											assign node515 = (inp[4]) ? 3'b101 : 3'b001;
								assign node519 = (inp[4]) ? node525 : node520;
									assign node520 = (inp[11]) ? 3'b110 : node521;
										assign node521 = (inp[2]) ? 3'b110 : 3'b001;
									assign node525 = (inp[5]) ? node529 : node526;
										assign node526 = (inp[11]) ? 3'b001 : 3'b110;
										assign node529 = (inp[11]) ? node535 : node530;
											assign node530 = (inp[3]) ? 3'b110 : node531;
												assign node531 = (inp[2]) ? 3'b110 : 3'b001;
											assign node535 = (inp[2]) ? 3'b010 : node536;
												assign node536 = (inp[3]) ? 3'b010 : 3'b110;
						assign node540 = (inp[11]) ? node570 : node541;
							assign node541 = (inp[8]) ? node557 : node542;
								assign node542 = (inp[1]) ? node550 : node543;
									assign node543 = (inp[2]) ? node545 : 3'b010;
										assign node545 = (inp[5]) ? node547 : 3'b100;
											assign node547 = (inp[4]) ? 3'b100 : 3'b010;
									assign node550 = (inp[4]) ? node552 : 3'b100;
										assign node552 = (inp[2]) ? 3'b000 : node553;
											assign node553 = (inp[3]) ? 3'b000 : 3'b100;
								assign node557 = (inp[1]) ? node565 : node558;
									assign node558 = (inp[2]) ? node560 : 3'b110;
										assign node560 = (inp[3]) ? 3'b010 : node561;
											assign node561 = (inp[4]) ? 3'b010 : 3'b110;
									assign node565 = (inp[2]) ? node567 : 3'b010;
										assign node567 = (inp[3]) ? 3'b100 : 3'b110;
							assign node570 = (inp[8]) ? node584 : node571;
								assign node571 = (inp[4]) ? node579 : node572;
									assign node572 = (inp[1]) ? 3'b100 : node573;
										assign node573 = (inp[3]) ? node575 : 3'b000;
											assign node575 = (inp[2]) ? 3'b000 : 3'b100;
									assign node579 = (inp[1]) ? 3'b000 : node580;
										assign node580 = (inp[2]) ? 3'b000 : 3'b100;
								assign node584 = (inp[2]) ? node592 : node585;
									assign node585 = (inp[1]) ? 3'b100 : node586;
										assign node586 = (inp[3]) ? 3'b010 : node587;
											assign node587 = (inp[4]) ? 3'b010 : 3'b110;
									assign node592 = (inp[1]) ? 3'b000 : 3'b100;
					assign node595 = (inp[10]) ? node643 : node596;
						assign node596 = (inp[1]) ? node628 : node597;
							assign node597 = (inp[8]) ? node619 : node598;
								assign node598 = (inp[11]) ? node612 : node599;
									assign node599 = (inp[2]) ? node605 : node600;
										assign node600 = (inp[4]) ? 3'b011 : node601;
											assign node601 = (inp[5]) ? 3'b001 : 3'b101;
										assign node605 = (inp[3]) ? 3'b101 : node606;
											assign node606 = (inp[4]) ? 3'b101 : node607;
												assign node607 = (inp[5]) ? 3'b111 : 3'b011;
									assign node612 = (inp[2]) ? node614 : 3'b101;
										assign node614 = (inp[4]) ? 3'b001 : node615;
											assign node615 = (inp[5]) ? 3'b001 : 3'b101;
								assign node619 = (inp[2]) ? node623 : node620;
									assign node620 = (inp[11]) ? 3'b011 : 3'b111;
									assign node623 = (inp[11]) ? node625 : 3'b011;
										assign node625 = (inp[4]) ? 3'b101 : 3'b011;
							assign node628 = (inp[8]) ? node636 : node629;
								assign node629 = (inp[2]) ? node633 : node630;
									assign node630 = (inp[11]) ? 3'b001 : 3'b101;
									assign node633 = (inp[11]) ? 3'b111 : 3'b001;
								assign node636 = (inp[2]) ? node640 : node637;
									assign node637 = (inp[11]) ? 3'b101 : 3'b011;
									assign node640 = (inp[11]) ? 3'b001 : 3'b101;
						assign node643 = (inp[1]) ? node683 : node644;
							assign node644 = (inp[4]) ? node662 : node645;
								assign node645 = (inp[8]) ? node657 : node646;
									assign node646 = (inp[11]) ? node652 : node647;
										assign node647 = (inp[3]) ? 3'b001 : node648;
											assign node648 = (inp[2]) ? 3'b001 : 3'b101;
										assign node652 = (inp[2]) ? 3'b101 : node653;
											assign node653 = (inp[3]) ? 3'b101 : 3'b001;
									assign node657 = (inp[11]) ? node659 : 3'b101;
										assign node659 = (inp[2]) ? 3'b010 : 3'b001;
								assign node662 = (inp[2]) ? node674 : node663;
									assign node663 = (inp[8]) ? node669 : node664;
										assign node664 = (inp[11]) ? node666 : 3'b001;
											assign node666 = (inp[5]) ? 3'b110 : 3'b101;
										assign node669 = (inp[3]) ? node671 : 3'b101;
											assign node671 = (inp[11]) ? 3'b001 : 3'b101;
									assign node674 = (inp[11]) ? node680 : node675;
										assign node675 = (inp[8]) ? node677 : 3'b110;
											assign node677 = (inp[3]) ? 3'b001 : 3'b101;
										assign node680 = (inp[8]) ? 3'b110 : 3'b010;
							assign node683 = (inp[8]) ? node691 : node684;
								assign node684 = (inp[2]) ? node688 : node685;
									assign node685 = (inp[11]) ? 3'b010 : 3'b110;
									assign node688 = (inp[11]) ? 3'b100 : 3'b010;
								assign node691 = (inp[11]) ? node703 : node692;
									assign node692 = (inp[2]) ? node698 : node693;
										assign node693 = (inp[4]) ? 3'b001 : node694;
											assign node694 = (inp[3]) ? 3'b001 : 3'b000;
										assign node698 = (inp[3]) ? node700 : 3'b111;
											assign node700 = (inp[4]) ? 3'b110 : 3'b111;
									assign node703 = (inp[2]) ? 3'b010 : node704;
										assign node704 = (inp[3]) ? 3'b110 : node705;
											assign node705 = (inp[4]) ? 3'b110 : 3'b111;
			assign node710 = (inp[0]) ? node954 : node711;
				assign node711 = (inp[7]) ? node829 : node712;
					assign node712 = (inp[10]) ? node778 : node713;
						assign node713 = (inp[11]) ? node747 : node714;
							assign node714 = (inp[1]) ? node732 : node715;
								assign node715 = (inp[8]) ? node723 : node716;
									assign node716 = (inp[2]) ? 3'b010 : node717;
										assign node717 = (inp[4]) ? node719 : 3'b110;
											assign node719 = (inp[3]) ? 3'b010 : 3'b110;
									assign node723 = (inp[2]) ? node727 : node724;
										assign node724 = (inp[4]) ? 3'b110 : 3'b001;
										assign node727 = (inp[4]) ? node729 : 3'b110;
											assign node729 = (inp[5]) ? 3'b110 : 3'b010;
								assign node732 = (inp[8]) ? node742 : node733;
									assign node733 = (inp[4]) ? node735 : 3'b100;
										assign node735 = (inp[5]) ? node737 : 3'b000;
											assign node737 = (inp[2]) ? node739 : 3'b100;
												assign node739 = (inp[3]) ? 3'b000 : 3'b100;
									assign node742 = (inp[2]) ? 3'b010 : node743;
										assign node743 = (inp[3]) ? 3'b010 : 3'b110;
							assign node747 = (inp[8]) ? node763 : node748;
								assign node748 = (inp[1]) ? node756 : node749;
									assign node749 = (inp[2]) ? 3'b100 : node750;
										assign node750 = (inp[4]) ? node752 : 3'b000;
											assign node752 = (inp[3]) ? 3'b100 : 3'b000;
									assign node756 = (inp[2]) ? 3'b000 : node757;
										assign node757 = (inp[5]) ? 3'b000 : node758;
											assign node758 = (inp[3]) ? 3'b000 : 3'b100;
								assign node763 = (inp[1]) ? node773 : node764;
									assign node764 = (inp[2]) ? 3'b010 : node765;
										assign node765 = (inp[4]) ? node767 : 3'b101;
											assign node767 = (inp[5]) ? node769 : 3'b110;
												assign node769 = (inp[3]) ? 3'b010 : 3'b110;
									assign node773 = (inp[2]) ? 3'b100 : node774;
										assign node774 = (inp[3]) ? 3'b100 : 3'b010;
						assign node778 = (inp[1]) ? node816 : node779;
							assign node779 = (inp[11]) ? node791 : node780;
								assign node780 = (inp[8]) ? node784 : node781;
									assign node781 = (inp[2]) ? 3'b000 : 3'b100;
									assign node784 = (inp[2]) ? node786 : 3'b010;
										assign node786 = (inp[3]) ? 3'b100 : node787;
											assign node787 = (inp[4]) ? 3'b100 : 3'b110;
								assign node791 = (inp[5]) ? node809 : node792;
									assign node792 = (inp[3]) ? node802 : node793;
										assign node793 = (inp[4]) ? node795 : 3'b100;
											assign node795 = (inp[2]) ? node799 : node796;
												assign node796 = (inp[8]) ? 3'b100 : 3'b000;
												assign node799 = (inp[8]) ? 3'b000 : 3'b100;
										assign node802 = (inp[2]) ? node806 : node803;
											assign node803 = (inp[8]) ? 3'b100 : 3'b000;
											assign node806 = (inp[8]) ? 3'b000 : 3'b100;
									assign node809 = (inp[8]) ? node813 : node810;
										assign node810 = (inp[2]) ? 3'b100 : 3'b000;
										assign node813 = (inp[2]) ? 3'b000 : 3'b100;
							assign node816 = (inp[2]) ? 3'b000 : node817;
								assign node817 = (inp[4]) ? node819 : 3'b000;
									assign node819 = (inp[3]) ? 3'b000 : node820;
										assign node820 = (inp[5]) ? 3'b100 : node821;
											assign node821 = (inp[8]) ? node823 : 3'b000;
												assign node823 = (inp[11]) ? 3'b000 : 3'b100;
					assign node829 = (inp[10]) ? node903 : node830;
						assign node830 = (inp[1]) ? node870 : node831;
							assign node831 = (inp[8]) ? node857 : node832;
								assign node832 = (inp[2]) ? node848 : node833;
									assign node833 = (inp[5]) ? node841 : node834;
										assign node834 = (inp[4]) ? 3'b101 : node835;
											assign node835 = (inp[3]) ? node837 : 3'b101;
												assign node837 = (inp[11]) ? 3'b001 : 3'b101;
										assign node841 = (inp[4]) ? 3'b001 : node842;
											assign node842 = (inp[11]) ? node844 : 3'b101;
												assign node844 = (inp[3]) ? 3'b001 : 3'b101;
									assign node848 = (inp[11]) ? 3'b110 : node849;
										assign node849 = (inp[3]) ? 3'b001 : node850;
											assign node850 = (inp[5]) ? node852 : 3'b101;
												assign node852 = (inp[4]) ? 3'b001 : 3'b101;
								assign node857 = (inp[11]) ? node865 : node858;
									assign node858 = (inp[2]) ? node860 : 3'b011;
										assign node860 = (inp[3]) ? 3'b101 : node861;
											assign node861 = (inp[4]) ? 3'b101 : 3'b011;
									assign node865 = (inp[3]) ? node867 : 3'b001;
										assign node867 = (inp[2]) ? 3'b001 : 3'b101;
							assign node870 = (inp[11]) ? node888 : node871;
								assign node871 = (inp[8]) ? node881 : node872;
									assign node872 = (inp[2]) ? 3'b110 : node873;
										assign node873 = (inp[3]) ? 3'b110 : node874;
											assign node874 = (inp[4]) ? 3'b001 : node875;
												assign node875 = (inp[5]) ? 3'b110 : 3'b001;
									assign node881 = (inp[2]) ? 3'b001 : node882;
										assign node882 = (inp[3]) ? node884 : 3'b101;
											assign node884 = (inp[4]) ? 3'b001 : 3'b101;
								assign node888 = (inp[8]) ? node898 : node889;
									assign node889 = (inp[2]) ? node895 : node890;
										assign node890 = (inp[4]) ? node892 : 3'b110;
											assign node892 = (inp[3]) ? 3'b010 : 3'b110;
										assign node895 = (inp[4]) ? 3'b010 : 3'b001;
									assign node898 = (inp[2]) ? 3'b110 : node899;
										assign node899 = (inp[4]) ? 3'b110 : 3'b010;
						assign node903 = (inp[1]) ? node919 : node904;
							assign node904 = (inp[8]) ? node912 : node905;
								assign node905 = (inp[2]) ? node909 : node906;
									assign node906 = (inp[11]) ? 3'b010 : 3'b110;
									assign node909 = (inp[11]) ? 3'b100 : 3'b010;
								assign node912 = (inp[11]) ? node916 : node913;
									assign node913 = (inp[2]) ? 3'b110 : 3'b001;
									assign node916 = (inp[2]) ? 3'b010 : 3'b110;
							assign node919 = (inp[8]) ? node935 : node920;
								assign node920 = (inp[11]) ? node928 : node921;
									assign node921 = (inp[2]) ? 3'b100 : node922;
										assign node922 = (inp[3]) ? node924 : 3'b010;
											assign node924 = (inp[4]) ? 3'b100 : 3'b000;
									assign node928 = (inp[2]) ? 3'b000 : node929;
										assign node929 = (inp[3]) ? node931 : 3'b100;
											assign node931 = (inp[5]) ? 3'b000 : 3'b100;
								assign node935 = (inp[2]) ? node947 : node936;
									assign node936 = (inp[11]) ? node942 : node937;
										assign node937 = (inp[4]) ? node939 : 3'b100;
											assign node939 = (inp[3]) ? 3'b010 : 3'b110;
										assign node942 = (inp[5]) ? node944 : 3'b010;
											assign node944 = (inp[4]) ? 3'b100 : 3'b010;
									assign node947 = (inp[11]) ? 3'b100 : node948;
										assign node948 = (inp[5]) ? 3'b010 : node949;
											assign node949 = (inp[4]) ? 3'b100 : 3'b010;
				assign node954 = (inp[10]) ? node1036 : node955;
					assign node955 = (inp[7]) ? node981 : node956;
						assign node956 = (inp[1]) ? 3'b000 : node957;
							assign node957 = (inp[8]) ? node959 : 3'b000;
								assign node959 = (inp[11]) ? node973 : node960;
									assign node960 = (inp[5]) ? node962 : 3'b100;
										assign node962 = (inp[3]) ? node968 : node963;
											assign node963 = (inp[2]) ? 3'b100 : node964;
												assign node964 = (inp[4]) ? 3'b100 : 3'b010;
											assign node968 = (inp[4]) ? node970 : 3'b100;
												assign node970 = (inp[2]) ? 3'b000 : 3'b100;
									assign node973 = (inp[4]) ? 3'b000 : node974;
										assign node974 = (inp[2]) ? 3'b010 : node975;
											assign node975 = (inp[3]) ? 3'b010 : 3'b100;
						assign node981 = (inp[1]) ? node1009 : node982;
							assign node982 = (inp[8]) ? node998 : node983;
								assign node983 = (inp[4]) ? node985 : 3'b010;
									assign node985 = (inp[2]) ? node991 : node986;
										assign node986 = (inp[11]) ? node988 : 3'b010;
											assign node988 = (inp[5]) ? 3'b100 : 3'b010;
										assign node991 = (inp[3]) ? 3'b000 : node992;
											assign node992 = (inp[11]) ? node994 : 3'b100;
												assign node994 = (inp[5]) ? 3'b000 : 3'b100;
								assign node998 = (inp[2]) ? node1004 : node999;
									assign node999 = (inp[11]) ? node1001 : 3'b110;
										assign node1001 = (inp[4]) ? 3'b010 : 3'b110;
									assign node1004 = (inp[11]) ? 3'b100 : node1005;
										assign node1005 = (inp[4]) ? 3'b010 : 3'b110;
							assign node1009 = (inp[8]) ? node1017 : node1010;
								assign node1010 = (inp[2]) ? node1014 : node1011;
									assign node1011 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1014 = (inp[11]) ? 3'b100 : 3'b000;
								assign node1017 = (inp[11]) ? node1029 : node1018;
									assign node1018 = (inp[2]) ? node1024 : node1019;
										assign node1019 = (inp[3]) ? 3'b010 : node1020;
											assign node1020 = (inp[4]) ? 3'b010 : 3'b000;
										assign node1024 = (inp[4]) ? node1026 : 3'b110;
											assign node1026 = (inp[3]) ? 3'b100 : 3'b110;
									assign node1029 = (inp[2]) ? 3'b000 : node1030;
										assign node1030 = (inp[4]) ? 3'b100 : node1031;
											assign node1031 = (inp[3]) ? 3'b100 : 3'b110;
					assign node1036 = (inp[1]) ? 3'b000 : node1037;
						assign node1037 = (inp[8]) ? node1039 : 3'b000;
							assign node1039 = (inp[7]) ? node1041 : 3'b000;
								assign node1041 = (inp[11]) ? node1047 : node1042;
									assign node1042 = (inp[3]) ? 3'b100 : node1043;
										assign node1043 = (inp[2]) ? 3'b100 : 3'b010;
									assign node1047 = (inp[2]) ? 3'b000 : node1048;
										assign node1048 = (inp[3]) ? 3'b000 : 3'b100;

endmodule