module dtc_split33_bm20 (
	input  wire [9-1:0] inp,
	output wire [9-1:0] outp
);

	wire [9-1:0] node1;
	wire [9-1:0] node2;
	wire [9-1:0] node3;
	wire [9-1:0] node4;
	wire [9-1:0] node5;
	wire [9-1:0] node7;
	wire [9-1:0] node10;
	wire [9-1:0] node11;
	wire [9-1:0] node14;
	wire [9-1:0] node17;
	wire [9-1:0] node18;
	wire [9-1:0] node21;
	wire [9-1:0] node22;
	wire [9-1:0] node25;
	wire [9-1:0] node28;
	wire [9-1:0] node29;
	wire [9-1:0] node30;
	wire [9-1:0] node31;
	wire [9-1:0] node34;
	wire [9-1:0] node37;
	wire [9-1:0] node38;
	wire [9-1:0] node39;
	wire [9-1:0] node43;
	wire [9-1:0] node46;
	wire [9-1:0] node49;
	wire [9-1:0] node50;
	wire [9-1:0] node51;
	wire [9-1:0] node52;
	wire [9-1:0] node54;
	wire [9-1:0] node55;
	wire [9-1:0] node56;
	wire [9-1:0] node61;
	wire [9-1:0] node64;
	wire [9-1:0] node65;
	wire [9-1:0] node66;
	wire [9-1:0] node68;
	wire [9-1:0] node71;
	wire [9-1:0] node74;
	wire [9-1:0] node75;
	wire [9-1:0] node76;
	wire [9-1:0] node81;
	wire [9-1:0] node82;
	wire [9-1:0] node83;
	wire [9-1:0] node85;
	wire [9-1:0] node87;
	wire [9-1:0] node90;
	wire [9-1:0] node91;
	wire [9-1:0] node92;
	wire [9-1:0] node94;
	wire [9-1:0] node98;
	wire [9-1:0] node101;
	wire [9-1:0] node102;
	wire [9-1:0] node104;
	wire [9-1:0] node107;
	wire [9-1:0] node108;
	wire [9-1:0] node109;
	wire [9-1:0] node113;
	wire [9-1:0] node115;
	wire [9-1:0] node116;
	wire [9-1:0] node120;
	wire [9-1:0] node121;
	wire [9-1:0] node122;
	wire [9-1:0] node123;
	wire [9-1:0] node124;
	wire [9-1:0] node126;
	wire [9-1:0] node129;
	wire [9-1:0] node130;
	wire [9-1:0] node131;
	wire [9-1:0] node136;
	wire [9-1:0] node138;
	wire [9-1:0] node139;
	wire [9-1:0] node142;
	wire [9-1:0] node143;
	wire [9-1:0] node147;
	wire [9-1:0] node148;
	wire [9-1:0] node149;
	wire [9-1:0] node151;
	wire [9-1:0] node154;
	wire [9-1:0] node155;
	wire [9-1:0] node157;
	wire [9-1:0] node159;
	wire [9-1:0] node162;
	wire [9-1:0] node163;
	wire [9-1:0] node165;
	wire [9-1:0] node169;
	wire [9-1:0] node170;
	wire [9-1:0] node172;
	wire [9-1:0] node173;
	wire [9-1:0] node177;
	wire [9-1:0] node178;
	wire [9-1:0] node180;
	wire [9-1:0] node184;
	wire [9-1:0] node185;
	wire [9-1:0] node186;
	wire [9-1:0] node187;
	wire [9-1:0] node188;
	wire [9-1:0] node192;
	wire [9-1:0] node194;
	wire [9-1:0] node195;
	wire [9-1:0] node197;
	wire [9-1:0] node201;
	wire [9-1:0] node202;
	wire [9-1:0] node204;
	wire [9-1:0] node206;
	wire [9-1:0] node208;
	wire [9-1:0] node211;
	wire [9-1:0] node213;
	wire [9-1:0] node214;
	wire [9-1:0] node218;
	wire [9-1:0] node219;
	wire [9-1:0] node221;
	wire [9-1:0] node223;
	wire [9-1:0] node225;
	wire [9-1:0] node226;
	wire [9-1:0] node230;
	wire [9-1:0] node231;
	wire [9-1:0] node233;
	wire [9-1:0] node236;
	wire [9-1:0] node238;
	wire [9-1:0] node239;
	wire [9-1:0] node241;
	wire [9-1:0] node244;
	wire [9-1:0] node246;

	assign outp = (inp[7]) ? node120 : node1;
		assign node1 = (inp[1]) ? node49 : node2;
			assign node2 = (inp[8]) ? node28 : node3;
				assign node3 = (inp[3]) ? node17 : node4;
					assign node4 = (inp[0]) ? node10 : node5;
						assign node5 = (inp[5]) ? node7 : 9'b011111111;
							assign node7 = (inp[4]) ? 9'b000111111 : 9'b001111111;
						assign node10 = (inp[4]) ? node14 : node11;
							assign node11 = (inp[6]) ? 9'b001111111 : 9'b000111111;
							assign node14 = (inp[2]) ? 9'b000011111 : 9'b000111111;
					assign node17 = (inp[5]) ? node21 : node18;
						assign node18 = (inp[6]) ? 9'b000111111 : 9'b001111111;
						assign node21 = (inp[6]) ? node25 : node22;
							assign node22 = (inp[0]) ? 9'b000011111 : 9'b000111111;
							assign node25 = (inp[2]) ? 9'b000001111 : 9'b000011111;
				assign node28 = (inp[6]) ? node46 : node29;
					assign node29 = (inp[3]) ? node37 : node30;
						assign node30 = (inp[5]) ? node34 : node31;
							assign node31 = (inp[4]) ? 9'b000111111 : 9'b001111111;
							assign node34 = (inp[0]) ? 9'b000011111 : 9'b000111111;
						assign node37 = (inp[4]) ? node43 : node38;
							assign node38 = (inp[5]) ? 9'b000011111 : node39;
								assign node39 = (inp[2]) ? 9'b000011111 : 9'b000111111;
							assign node43 = (inp[5]) ? 9'b000001111 : 9'b000011111;
					assign node46 = (inp[0]) ? 9'b000001111 : 9'b000011111;
			assign node49 = (inp[2]) ? node81 : node50;
				assign node50 = (inp[4]) ? node64 : node51;
					assign node51 = (inp[8]) ? node61 : node52;
						assign node52 = (inp[0]) ? node54 : 9'b001111111;
							assign node54 = (inp[3]) ? 9'b000011111 : node55;
								assign node55 = (inp[5]) ? 9'b000111111 : node56;
									assign node56 = (inp[6]) ? 9'b000111111 : 9'b001111111;
						assign node61 = (inp[0]) ? 9'b000011111 : 9'b000111111;
					assign node64 = (inp[5]) ? node74 : node65;
						assign node65 = (inp[8]) ? node71 : node66;
							assign node66 = (inp[3]) ? node68 : 9'b000111111;
								assign node68 = (inp[6]) ? 9'b000011111 : 9'b000111111;
							assign node71 = (inp[6]) ? 9'b000001111 : 9'b000011111;
						assign node74 = (inp[3]) ? 9'b000001111 : node75;
							assign node75 = (inp[8]) ? 9'b000001111 : node76;
								assign node76 = (inp[0]) ? 9'b000001111 : 9'b000011111;
				assign node81 = (inp[6]) ? node101 : node82;
					assign node82 = (inp[8]) ? node90 : node83;
						assign node83 = (inp[0]) ? node85 : 9'b000111111;
							assign node85 = (inp[5]) ? node87 : 9'b000011111;
								assign node87 = (inp[4]) ? 9'b000001111 : 9'b000011111;
						assign node90 = (inp[0]) ? node98 : node91;
							assign node91 = (inp[3]) ? 9'b000001111 : node92;
								assign node92 = (inp[5]) ? node94 : 9'b000011111;
									assign node94 = (inp[4]) ? 9'b000001111 : 9'b000011111;
							assign node98 = (inp[3]) ? 9'b000000111 : 9'b000001111;
					assign node101 = (inp[3]) ? node107 : node102;
						assign node102 = (inp[0]) ? node104 : 9'b000001111;
							assign node104 = (inp[8]) ? 9'b000000111 : 9'b000001111;
						assign node107 = (inp[0]) ? node113 : node108;
							assign node108 = (inp[8]) ? 9'b000000111 : node109;
								assign node109 = (inp[4]) ? 9'b000000111 : 9'b000001111;
							assign node113 = (inp[8]) ? node115 : 9'b000000111;
								assign node115 = (inp[4]) ? 9'b000000011 : node116;
									assign node116 = (inp[5]) ? 9'b000000011 : 9'b000000111;
		assign node120 = (inp[3]) ? node184 : node121;
			assign node121 = (inp[5]) ? node147 : node122;
				assign node122 = (inp[2]) ? node136 : node123;
					assign node123 = (inp[1]) ? node129 : node124;
						assign node124 = (inp[0]) ? node126 : 9'b000111111;
							assign node126 = (inp[6]) ? 9'b000011111 : 9'b000111111;
						assign node129 = (inp[4]) ? 9'b000001111 : node130;
							assign node130 = (inp[0]) ? 9'b000011111 : node131;
								assign node131 = (inp[6]) ? 9'b000011111 : 9'b000111111;
					assign node136 = (inp[0]) ? node138 : 9'b000011111;
						assign node138 = (inp[1]) ? node142 : node139;
							assign node139 = (inp[8]) ? 9'b000001111 : 9'b000111111;
							assign node142 = (inp[8]) ? 9'b000000111 : node143;
								assign node143 = (inp[6]) ? 9'b000000111 : 9'b000001111;
				assign node147 = (inp[2]) ? node169 : node148;
					assign node148 = (inp[1]) ? node154 : node149;
						assign node149 = (inp[6]) ? node151 : 9'b000011111;
							assign node151 = (inp[0]) ? 9'b000000111 : 9'b000011111;
						assign node154 = (inp[0]) ? node162 : node155;
							assign node155 = (inp[8]) ? node157 : 9'b000011111;
								assign node157 = (inp[4]) ? node159 : 9'b000001111;
									assign node159 = (inp[6]) ? 9'b000000111 : 9'b000001111;
							assign node162 = (inp[6]) ? 9'b000000111 : node163;
								assign node163 = (inp[4]) ? node165 : 9'b000001111;
									assign node165 = (inp[8]) ? 9'b000000111 : 9'b000001111;
					assign node169 = (inp[4]) ? node177 : node170;
						assign node170 = (inp[0]) ? node172 : 9'b000001111;
							assign node172 = (inp[6]) ? 9'b000000111 : node173;
								assign node173 = (inp[8]) ? 9'b000000111 : 9'b000001111;
						assign node177 = (inp[6]) ? 9'b000000011 : node178;
							assign node178 = (inp[8]) ? node180 : 9'b000001111;
								assign node180 = (inp[0]) ? 9'b000000011 : 9'b000000111;
			assign node184 = (inp[5]) ? node218 : node185;
				assign node185 = (inp[4]) ? node201 : node186;
					assign node186 = (inp[6]) ? node192 : node187;
						assign node187 = (inp[2]) ? 9'b000001111 : node188;
							assign node188 = (inp[8]) ? 9'b000011111 : 9'b000111111;
						assign node192 = (inp[2]) ? node194 : 9'b000001111;
							assign node194 = (inp[1]) ? 9'b000000111 : node195;
								assign node195 = (inp[0]) ? node197 : 9'b000001111;
									assign node197 = (inp[8]) ? 9'b000000111 : 9'b000001111;
					assign node201 = (inp[0]) ? node211 : node202;
						assign node202 = (inp[2]) ? node204 : 9'b000001111;
							assign node204 = (inp[8]) ? node206 : 9'b000001111;
								assign node206 = (inp[1]) ? node208 : 9'b000000111;
									assign node208 = (inp[6]) ? 9'b000000011 : 9'b000000111;
						assign node211 = (inp[2]) ? node213 : 9'b000000111;
							assign node213 = (inp[1]) ? 9'b000000011 : node214;
								assign node214 = (inp[6]) ? 9'b000000011 : 9'b000000111;
				assign node218 = (inp[6]) ? node230 : node219;
					assign node219 = (inp[4]) ? node221 : 9'b000001111;
						assign node221 = (inp[1]) ? node223 : 9'b000001111;
							assign node223 = (inp[8]) ? node225 : 9'b000000111;
								assign node225 = (inp[2]) ? 9'b000000011 : node226;
									assign node226 = (inp[0]) ? 9'b000000011 : 9'b000000111;
					assign node230 = (inp[8]) ? node236 : node231;
						assign node231 = (inp[0]) ? node233 : 9'b000000111;
							assign node233 = (inp[2]) ? 9'b000000011 : 9'b000000111;
						assign node236 = (inp[4]) ? node238 : 9'b000000011;
							assign node238 = (inp[1]) ? node244 : node239;
								assign node239 = (inp[0]) ? node241 : 9'b000000011;
									assign node241 = (inp[2]) ? 9'b000000001 : 9'b000000011;
								assign node244 = (inp[2]) ? node246 : 9'b000000001;
									assign node246 = (inp[0]) ? 9'b000000000 : 9'b000000001;

endmodule