module dtc_split66_bm82 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node34;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node63;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node76;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node226;

	assign outp = (inp[0]) ? node112 : node1;
		assign node1 = (inp[3]) ? node59 : node2;
			assign node2 = (inp[6]) ? node28 : node3;
				assign node3 = (inp[4]) ? node15 : node4;
					assign node4 = (inp[7]) ? node10 : node5;
						assign node5 = (inp[11]) ? 3'b001 : node6;
							assign node6 = (inp[2]) ? 3'b001 : 3'b001;
						assign node10 = (inp[1]) ? node12 : 3'b111;
							assign node12 = (inp[9]) ? 3'b001 : 3'b010;
					assign node15 = (inp[1]) ? node21 : node16;
						assign node16 = (inp[7]) ? node18 : 3'b111;
							assign node18 = (inp[9]) ? 3'b111 : 3'b111;
						assign node21 = (inp[9]) ? node25 : node22;
							assign node22 = (inp[7]) ? 3'b001 : 3'b101;
							assign node25 = (inp[7]) ? 3'b111 : 3'b101;
				assign node28 = (inp[1]) ? node44 : node29;
					assign node29 = (inp[9]) ? node37 : node30;
						assign node30 = (inp[7]) ? node34 : node31;
							assign node31 = (inp[2]) ? 3'b011 : 3'b001;
							assign node34 = (inp[4]) ? 3'b010 : 3'b110;
						assign node37 = (inp[7]) ? node41 : node38;
							assign node38 = (inp[4]) ? 3'b111 : 3'b011;
							assign node41 = (inp[2]) ? 3'b110 : 3'b001;
					assign node44 = (inp[9]) ? node52 : node45;
						assign node45 = (inp[4]) ? node49 : node46;
							assign node46 = (inp[7]) ? 3'b000 : 3'b000;
							assign node49 = (inp[7]) ? 3'b000 : 3'b110;
						assign node52 = (inp[7]) ? node56 : node53;
							assign node53 = (inp[8]) ? 3'b110 : 3'b001;
							assign node56 = (inp[2]) ? 3'b110 : 3'b010;
			assign node59 = (inp[6]) ? node81 : node60;
				assign node60 = (inp[1]) ? node68 : node61;
					assign node61 = (inp[2]) ? node63 : 3'b111;
						assign node63 = (inp[8]) ? node65 : 3'b111;
							assign node65 = (inp[7]) ? 3'b111 : 3'b111;
					assign node68 = (inp[9]) ? node76 : node69;
						assign node69 = (inp[4]) ? node73 : node70;
							assign node70 = (inp[7]) ? 3'b011 : 3'b111;
							assign node73 = (inp[5]) ? 3'b111 : 3'b111;
						assign node76 = (inp[2]) ? node78 : 3'b111;
							assign node78 = (inp[11]) ? 3'b111 : 3'b111;
				assign node81 = (inp[9]) ? node97 : node82;
					assign node82 = (inp[1]) ? node90 : node83;
						assign node83 = (inp[7]) ? node87 : node84;
							assign node84 = (inp[4]) ? 3'b111 : 3'b011;
							assign node87 = (inp[4]) ? 3'b011 : 3'b001;
						assign node90 = (inp[7]) ? node94 : node91;
							assign node91 = (inp[8]) ? 3'b011 : 3'b101;
							assign node94 = (inp[4]) ? 3'b001 : 3'b010;
					assign node97 = (inp[1]) ? node105 : node98;
						assign node98 = (inp[4]) ? node102 : node99;
							assign node99 = (inp[2]) ? 3'b111 : 3'b111;
							assign node102 = (inp[10]) ? 3'b111 : 3'b111;
						assign node105 = (inp[7]) ? node109 : node106;
							assign node106 = (inp[4]) ? 3'b111 : 3'b011;
							assign node109 = (inp[4]) ? 3'b101 : 3'b001;
		assign node112 = (inp[6]) ? node176 : node113;
			assign node113 = (inp[3]) ? node145 : node114;
				assign node114 = (inp[1]) ? node130 : node115;
					assign node115 = (inp[4]) ? node123 : node116;
						assign node116 = (inp[7]) ? node120 : node117;
							assign node117 = (inp[9]) ? 3'b001 : 3'b000;
							assign node120 = (inp[9]) ? 3'b110 : 3'b000;
						assign node123 = (inp[7]) ? node127 : node124;
							assign node124 = (inp[8]) ? 3'b011 : 3'b101;
							assign node127 = (inp[9]) ? 3'b001 : 3'b100;
					assign node130 = (inp[7]) ? node138 : node131;
						assign node131 = (inp[4]) ? node135 : node132;
							assign node132 = (inp[9]) ? 3'b010 : 3'b010;
							assign node135 = (inp[9]) ? 3'b110 : 3'b110;
						assign node138 = (inp[9]) ? node142 : node139;
							assign node139 = (inp[4]) ? 3'b000 : 3'b000;
							assign node142 = (inp[4]) ? 3'b010 : 3'b000;
				assign node145 = (inp[1]) ? node161 : node146;
					assign node146 = (inp[9]) ? node154 : node147;
						assign node147 = (inp[7]) ? node151 : node148;
							assign node148 = (inp[4]) ? 3'b111 : 3'b001;
							assign node151 = (inp[4]) ? 3'b001 : 3'b001;
						assign node154 = (inp[7]) ? node158 : node155;
							assign node155 = (inp[10]) ? 3'b111 : 3'b111;
							assign node158 = (inp[4]) ? 3'b111 : 3'b011;
					assign node161 = (inp[9]) ? node169 : node162;
						assign node162 = (inp[7]) ? node166 : node163;
							assign node163 = (inp[4]) ? 3'b001 : 3'b110;
							assign node166 = (inp[4]) ? 3'b110 : 3'b000;
						assign node169 = (inp[7]) ? node173 : node170;
							assign node170 = (inp[4]) ? 3'b111 : 3'b101;
							assign node173 = (inp[10]) ? 3'b001 : 3'b100;
			assign node176 = (inp[3]) ? node198 : node177;
				assign node177 = (inp[9]) ? node185 : node178;
					assign node178 = (inp[4]) ? node180 : 3'b000;
						assign node180 = (inp[1]) ? 3'b000 : node181;
							assign node181 = (inp[7]) ? 3'b000 : 3'b000;
					assign node185 = (inp[1]) ? node193 : node186;
						assign node186 = (inp[7]) ? node190 : node187;
							assign node187 = (inp[4]) ? 3'b010 : 3'b100;
							assign node190 = (inp[4]) ? 3'b000 : 3'b000;
						assign node193 = (inp[7]) ? 3'b000 : node194;
							assign node194 = (inp[4]) ? 3'b000 : 3'b000;
				assign node198 = (inp[1]) ? node214 : node199;
					assign node199 = (inp[9]) ? node207 : node200;
						assign node200 = (inp[7]) ? node204 : node201;
							assign node201 = (inp[4]) ? 3'b010 : 3'b010;
							assign node204 = (inp[4]) ? 3'b010 : 3'b000;
						assign node207 = (inp[7]) ? node211 : node208;
							assign node208 = (inp[4]) ? 3'b101 : 3'b101;
							assign node211 = (inp[4]) ? 3'b011 : 3'b010;
					assign node214 = (inp[9]) ? node222 : node215;
						assign node215 = (inp[7]) ? node219 : node216;
							assign node216 = (inp[10]) ? 3'b000 : 3'b000;
							assign node219 = (inp[4]) ? 3'b000 : 3'b000;
						assign node222 = (inp[7]) ? node226 : node223;
							assign node223 = (inp[4]) ? 3'b110 : 3'b010;
							assign node226 = (inp[4]) ? 3'b000 : 3'b000;

endmodule