module dtc_split05_bm24 (
	input  wire [13-1:0] inp,
	output wire [13-1:0] outp
);

	wire [13-1:0] node1;
	wire [13-1:0] node2;
	wire [13-1:0] node3;
	wire [13-1:0] node4;
	wire [13-1:0] node5;
	wire [13-1:0] node6;
	wire [13-1:0] node7;
	wire [13-1:0] node9;
	wire [13-1:0] node12;
	wire [13-1:0] node13;
	wire [13-1:0] node16;
	wire [13-1:0] node19;
	wire [13-1:0] node22;
	wire [13-1:0] node23;
	wire [13-1:0] node24;
	wire [13-1:0] node27;
	wire [13-1:0] node28;
	wire [13-1:0] node32;
	wire [13-1:0] node33;
	wire [13-1:0] node37;
	wire [13-1:0] node38;
	wire [13-1:0] node39;
	wire [13-1:0] node40;
	wire [13-1:0] node44;
	wire [13-1:0] node45;
	wire [13-1:0] node48;
	wire [13-1:0] node51;
	wire [13-1:0] node52;
	wire [13-1:0] node53;
	wire [13-1:0] node54;
	wire [13-1:0] node59;
	wire [13-1:0] node62;
	wire [13-1:0] node63;
	wire [13-1:0] node64;
	wire [13-1:0] node65;
	wire [13-1:0] node66;
	wire [13-1:0] node68;
	wire [13-1:0] node72;
	wire [13-1:0] node73;
	wire [13-1:0] node74;
	wire [13-1:0] node77;
	wire [13-1:0] node80;
	wire [13-1:0] node83;
	wire [13-1:0] node84;
	wire [13-1:0] node85;
	wire [13-1:0] node86;
	wire [13-1:0] node91;
	wire [13-1:0] node94;
	wire [13-1:0] node95;
	wire [13-1:0] node96;
	wire [13-1:0] node97;
	wire [13-1:0] node99;
	wire [13-1:0] node103;
	wire [13-1:0] node104;
	wire [13-1:0] node106;
	wire [13-1:0] node110;
	wire [13-1:0] node111;
	wire [13-1:0] node113;
	wire [13-1:0] node116;
	wire [13-1:0] node119;
	wire [13-1:0] node120;
	wire [13-1:0] node121;
	wire [13-1:0] node122;
	wire [13-1:0] node123;
	wire [13-1:0] node124;
	wire [13-1:0] node126;
	wire [13-1:0] node129;
	wire [13-1:0] node132;
	wire [13-1:0] node133;
	wire [13-1:0] node137;
	wire [13-1:0] node138;
	wire [13-1:0] node139;
	wire [13-1:0] node141;
	wire [13-1:0] node145;
	wire [13-1:0] node148;
	wire [13-1:0] node149;
	wire [13-1:0] node150;
	wire [13-1:0] node151;
	wire [13-1:0] node152;
	wire [13-1:0] node155;
	wire [13-1:0] node158;
	wire [13-1:0] node159;
	wire [13-1:0] node163;
	wire [13-1:0] node164;
	wire [13-1:0] node165;
	wire [13-1:0] node168;
	wire [13-1:0] node171;
	wire [13-1:0] node173;
	wire [13-1:0] node176;
	wire [13-1:0] node177;
	wire [13-1:0] node178;
	wire [13-1:0] node182;
	wire [13-1:0] node185;
	wire [13-1:0] node186;
	wire [13-1:0] node187;
	wire [13-1:0] node188;
	wire [13-1:0] node191;
	wire [13-1:0] node192;
	wire [13-1:0] node193;
	wire [13-1:0] node197;
	wire [13-1:0] node200;
	wire [13-1:0] node201;
	wire [13-1:0] node202;
	wire [13-1:0] node203;
	wire [13-1:0] node207;
	wire [13-1:0] node210;
	wire [13-1:0] node211;
	wire [13-1:0] node214;
	wire [13-1:0] node217;
	wire [13-1:0] node218;
	wire [13-1:0] node219;
	wire [13-1:0] node220;
	wire [13-1:0] node223;
	wire [13-1:0] node226;
	wire [13-1:0] node228;
	wire [13-1:0] node230;
	wire [13-1:0] node233;
	wire [13-1:0] node234;
	wire [13-1:0] node236;
	wire [13-1:0] node238;
	wire [13-1:0] node241;
	wire [13-1:0] node242;
	wire [13-1:0] node244;
	wire [13-1:0] node247;
	wire [13-1:0] node249;
	wire [13-1:0] node252;
	wire [13-1:0] node253;
	wire [13-1:0] node254;
	wire [13-1:0] node255;
	wire [13-1:0] node256;
	wire [13-1:0] node257;
	wire [13-1:0] node258;
	wire [13-1:0] node259;
	wire [13-1:0] node263;
	wire [13-1:0] node265;
	wire [13-1:0] node268;
	wire [13-1:0] node269;
	wire [13-1:0] node272;
	wire [13-1:0] node275;
	wire [13-1:0] node276;
	wire [13-1:0] node277;
	wire [13-1:0] node279;
	wire [13-1:0] node283;
	wire [13-1:0] node284;
	wire [13-1:0] node287;
	wire [13-1:0] node290;
	wire [13-1:0] node291;
	wire [13-1:0] node292;
	wire [13-1:0] node293;
	wire [13-1:0] node294;
	wire [13-1:0] node297;
	wire [13-1:0] node300;
	wire [13-1:0] node301;
	wire [13-1:0] node304;
	wire [13-1:0] node307;
	wire [13-1:0] node308;
	wire [13-1:0] node310;
	wire [13-1:0] node314;
	wire [13-1:0] node315;
	wire [13-1:0] node318;
	wire [13-1:0] node321;
	wire [13-1:0] node322;
	wire [13-1:0] node323;
	wire [13-1:0] node324;
	wire [13-1:0] node325;
	wire [13-1:0] node326;
	wire [13-1:0] node330;
	wire [13-1:0] node331;
	wire [13-1:0] node335;
	wire [13-1:0] node336;
	wire [13-1:0] node338;
	wire [13-1:0] node341;
	wire [13-1:0] node342;
	wire [13-1:0] node346;
	wire [13-1:0] node347;
	wire [13-1:0] node348;
	wire [13-1:0] node352;
	wire [13-1:0] node353;
	wire [13-1:0] node357;
	wire [13-1:0] node358;
	wire [13-1:0] node360;
	wire [13-1:0] node361;
	wire [13-1:0] node363;
	wire [13-1:0] node366;
	wire [13-1:0] node369;
	wire [13-1:0] node370;
	wire [13-1:0] node371;
	wire [13-1:0] node373;
	wire [13-1:0] node376;
	wire [13-1:0] node378;
	wire [13-1:0] node381;
	wire [13-1:0] node383;
	wire [13-1:0] node386;
	wire [13-1:0] node387;
	wire [13-1:0] node388;
	wire [13-1:0] node389;
	wire [13-1:0] node390;
	wire [13-1:0] node391;
	wire [13-1:0] node394;
	wire [13-1:0] node396;
	wire [13-1:0] node399;
	wire [13-1:0] node402;
	wire [13-1:0] node403;
	wire [13-1:0] node404;
	wire [13-1:0] node407;
	wire [13-1:0] node409;
	wire [13-1:0] node412;
	wire [13-1:0] node414;
	wire [13-1:0] node417;
	wire [13-1:0] node418;
	wire [13-1:0] node419;
	wire [13-1:0] node422;
	wire [13-1:0] node425;
	wire [13-1:0] node426;
	wire [13-1:0] node428;
	wire [13-1:0] node429;
	wire [13-1:0] node432;
	wire [13-1:0] node435;
	wire [13-1:0] node436;
	wire [13-1:0] node438;
	wire [13-1:0] node441;
	wire [13-1:0] node444;
	wire [13-1:0] node445;
	wire [13-1:0] node446;
	wire [13-1:0] node447;
	wire [13-1:0] node448;
	wire [13-1:0] node452;
	wire [13-1:0] node455;
	wire [13-1:0] node456;
	wire [13-1:0] node458;
	wire [13-1:0] node461;
	wire [13-1:0] node462;
	wire [13-1:0] node463;
	wire [13-1:0] node467;
	wire [13-1:0] node468;
	wire [13-1:0] node472;
	wire [13-1:0] node473;
	wire [13-1:0] node474;
	wire [13-1:0] node475;
	wire [13-1:0] node477;
	wire [13-1:0] node480;
	wire [13-1:0] node482;
	wire [13-1:0] node485;
	wire [13-1:0] node486;
	wire [13-1:0] node488;
	wire [13-1:0] node492;
	wire [13-1:0] node493;
	wire [13-1:0] node494;
	wire [13-1:0] node496;
	wire [13-1:0] node499;
	wire [13-1:0] node502;
	wire [13-1:0] node503;
	wire [13-1:0] node504;

	assign outp = (inp[1]) ? node252 : node1;
		assign node1 = (inp[10]) ? node119 : node2;
			assign node2 = (inp[12]) ? node62 : node3;
				assign node3 = (inp[2]) ? node37 : node4;
					assign node4 = (inp[6]) ? node22 : node5;
						assign node5 = (inp[8]) ? node19 : node6;
							assign node6 = (inp[0]) ? node12 : node7;
								assign node7 = (inp[5]) ? node9 : 13'b0011111111111;
									assign node9 = (inp[4]) ? 13'b0000111111111 : 13'b0001111111111;
								assign node12 = (inp[5]) ? node16 : node13;
									assign node13 = (inp[4]) ? 13'b0000111111111 : 13'b0011111111111;
									assign node16 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node19 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
						assign node22 = (inp[8]) ? node32 : node23;
							assign node23 = (inp[9]) ? node27 : node24;
								assign node24 = (inp[5]) ? 13'b0000111111111 : 13'b0001111111111;
								assign node27 = (inp[5]) ? 13'b0000011111111 : node28;
									assign node28 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node32 = (inp[9]) ? 13'b0000000111111 : node33;
								assign node33 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
					assign node37 = (inp[0]) ? node51 : node38;
						assign node38 = (inp[6]) ? node44 : node39;
							assign node39 = (inp[4]) ? 13'b0000011111111 : node40;
								assign node40 = (inp[8]) ? 13'b0001111111111 : 13'b0000111111111;
							assign node44 = (inp[9]) ? node48 : node45;
								assign node45 = (inp[3]) ? 13'b0000111111111 : 13'b0000011111111;
								assign node48 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node51 = (inp[7]) ? node59 : node52;
							assign node52 = (inp[9]) ? 13'b0000000111111 : node53;
								assign node53 = (inp[4]) ? 13'b0000011111111 : node54;
									assign node54 = (inp[11]) ? 13'b0000011111111 : 13'b0000001111111;
							assign node59 = (inp[9]) ? 13'b0000001111111 : 13'b0000000111111;
				assign node62 = (inp[3]) ? node94 : node63;
					assign node63 = (inp[5]) ? node83 : node64;
						assign node64 = (inp[8]) ? node72 : node65;
							assign node65 = (inp[6]) ? 13'b0001111111111 : node66;
								assign node66 = (inp[2]) ? node68 : 13'b0000111111111;
									assign node68 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node72 = (inp[0]) ? node80 : node73;
								assign node73 = (inp[11]) ? node77 : node74;
									assign node74 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node77 = (inp[4]) ? 13'b0000011111111 : 13'b0000001111111;
								assign node80 = (inp[7]) ? 13'b0000000011111 : 13'b0000001111111;
						assign node83 = (inp[7]) ? node91 : node84;
							assign node84 = (inp[8]) ? 13'b0000001111111 : node85;
								assign node85 = (inp[0]) ? 13'b0000001111111 : node86;
									assign node86 = (inp[6]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node91 = (inp[0]) ? 13'b0000000011111 : 13'b0000001111111;
					assign node94 = (inp[11]) ? node110 : node95;
						assign node95 = (inp[9]) ? node103 : node96;
							assign node96 = (inp[8]) ? 13'b0000001111111 : node97;
								assign node97 = (inp[2]) ? node99 : 13'b0000111111111;
									assign node99 = (inp[7]) ? 13'b0000001111111 : 13'b0000001111111;
							assign node103 = (inp[5]) ? 13'b0000000111111 : node104;
								assign node104 = (inp[0]) ? node106 : 13'b0000011111111;
									assign node106 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node110 = (inp[0]) ? node116 : node111;
							assign node111 = (inp[8]) ? node113 : 13'b0000000111111;
								assign node113 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node116 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
			assign node119 = (inp[5]) ? node185 : node120;
				assign node120 = (inp[6]) ? node148 : node121;
					assign node121 = (inp[2]) ? node137 : node122;
						assign node122 = (inp[0]) ? node132 : node123;
							assign node123 = (inp[11]) ? node129 : node124;
								assign node124 = (inp[4]) ? node126 : 13'b0001111111111;
									assign node126 = (inp[12]) ? 13'b0000111111111 : 13'b0011111111111;
								assign node129 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node132 = (inp[4]) ? 13'b0000001111111 : node133;
								assign node133 = (inp[8]) ? 13'b0001111111111 : 13'b0000111111111;
						assign node137 = (inp[11]) ? node145 : node138;
							assign node138 = (inp[3]) ? 13'b0000011111111 : node139;
								assign node139 = (inp[4]) ? node141 : 13'b0000001111111;
									assign node141 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node145 = (inp[7]) ? 13'b0000000111111 : 13'b0000011111111;
					assign node148 = (inp[11]) ? node176 : node149;
						assign node149 = (inp[3]) ? node163 : node150;
							assign node150 = (inp[12]) ? node158 : node151;
								assign node151 = (inp[9]) ? node155 : node152;
									assign node152 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node155 = (inp[2]) ? 13'b0000011111111 : 13'b0000001111111;
								assign node158 = (inp[4]) ? 13'b0000000111111 : node159;
									assign node159 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node163 = (inp[8]) ? node171 : node164;
								assign node164 = (inp[4]) ? node168 : node165;
									assign node165 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node168 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node171 = (inp[2]) ? node173 : 13'b0000000001111;
									assign node173 = (inp[0]) ? 13'b0000001111111 : 13'b0000000111111;
						assign node176 = (inp[7]) ? node182 : node177;
							assign node177 = (inp[0]) ? 13'b0000000111111 : node178;
								assign node178 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node182 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
				assign node185 = (inp[2]) ? node217 : node186;
					assign node186 = (inp[9]) ? node200 : node187;
						assign node187 = (inp[12]) ? node191 : node188;
							assign node188 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node191 = (inp[3]) ? node197 : node192;
								assign node192 = (inp[7]) ? 13'b0000001111111 : node193;
									assign node193 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node197 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node200 = (inp[6]) ? node210 : node201;
							assign node201 = (inp[12]) ? node207 : node202;
								assign node202 = (inp[0]) ? 13'b0000000111111 : node203;
									assign node203 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node207 = (inp[0]) ? 13'b0000000001111 : 13'b0000000111111;
							assign node210 = (inp[11]) ? node214 : node211;
								assign node211 = (inp[4]) ? 13'b0000000111111 : 13'b0000000011111;
								assign node214 = (inp[3]) ? 13'b0000000000011 : 13'b0000000011111;
					assign node217 = (inp[12]) ? node233 : node218;
						assign node218 = (inp[9]) ? node226 : node219;
							assign node219 = (inp[8]) ? node223 : node220;
								assign node220 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node223 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node226 = (inp[3]) ? node228 : 13'b0000000111111;
								assign node228 = (inp[7]) ? node230 : 13'b0000000011111;
									assign node230 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node233 = (inp[11]) ? node241 : node234;
							assign node234 = (inp[6]) ? node236 : 13'b0000000111111;
								assign node236 = (inp[3]) ? node238 : 13'b0000000011111;
									assign node238 = (inp[4]) ? 13'b0000000000111 : 13'b0000000011111;
							assign node241 = (inp[8]) ? node247 : node242;
								assign node242 = (inp[7]) ? node244 : 13'b0000000111111;
									assign node244 = (inp[0]) ? 13'b0000000011111 : 13'b0000000001111;
								assign node247 = (inp[0]) ? node249 : 13'b0000000001111;
									assign node249 = (inp[6]) ? 13'b0000000000011 : 13'b0000000001111;
		assign node252 = (inp[11]) ? node386 : node253;
			assign node253 = (inp[9]) ? node321 : node254;
				assign node254 = (inp[8]) ? node290 : node255;
					assign node255 = (inp[2]) ? node275 : node256;
						assign node256 = (inp[5]) ? node268 : node257;
							assign node257 = (inp[7]) ? node263 : node258;
								assign node258 = (inp[10]) ? 13'b0011111111111 : node259;
									assign node259 = (inp[4]) ? 13'b0000111111111 : 13'b0001111111111;
								assign node263 = (inp[12]) ? node265 : 13'b0000111111111;
									assign node265 = (inp[4]) ? 13'b0000011111111 : 13'b0000011111111;
							assign node268 = (inp[0]) ? node272 : node269;
								assign node269 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node272 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node275 = (inp[10]) ? node283 : node276;
							assign node276 = (inp[0]) ? 13'b0000111111111 : node277;
								assign node277 = (inp[4]) ? node279 : 13'b0000011111111;
									assign node279 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node283 = (inp[7]) ? node287 : node284;
								assign node284 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node287 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node290 = (inp[7]) ? node314 : node291;
						assign node291 = (inp[10]) ? node307 : node292;
							assign node292 = (inp[4]) ? node300 : node293;
								assign node293 = (inp[12]) ? node297 : node294;
									assign node294 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node297 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node300 = (inp[5]) ? node304 : node301;
									assign node301 = (inp[3]) ? 13'b0000001111111 : 13'b0000001111111;
									assign node304 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node307 = (inp[4]) ? 13'b0000000111111 : node308;
								assign node308 = (inp[6]) ? node310 : 13'b0000001111111;
									assign node310 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node314 = (inp[5]) ? node318 : node315;
							assign node315 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node318 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
				assign node321 = (inp[2]) ? node357 : node322;
					assign node322 = (inp[5]) ? node346 : node323;
						assign node323 = (inp[4]) ? node335 : node324;
							assign node324 = (inp[7]) ? node330 : node325;
								assign node325 = (inp[8]) ? 13'b0000011111111 : node326;
									assign node326 = (inp[0]) ? 13'b0000111111111 : 13'b0000011111111;
								assign node330 = (inp[10]) ? 13'b0000001111111 : node331;
									assign node331 = (inp[0]) ? 13'b0000011111111 : 13'b0000001111111;
							assign node335 = (inp[10]) ? node341 : node336;
								assign node336 = (inp[6]) ? node338 : 13'b0000011111111;
									assign node338 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node341 = (inp[7]) ? 13'b0000000111111 : node342;
									assign node342 = (inp[3]) ? 13'b0000000111111 : 13'b0000000011111;
						assign node346 = (inp[3]) ? node352 : node347;
							assign node347 = (inp[4]) ? 13'b0000000111111 : node348;
								assign node348 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node352 = (inp[8]) ? 13'b0000000011111 : node353;
								assign node353 = (inp[0]) ? 13'b0000000001111 : 13'b0000000111111;
					assign node357 = (inp[10]) ? node369 : node358;
						assign node358 = (inp[7]) ? node360 : 13'b0000000111111;
							assign node360 = (inp[6]) ? node366 : node361;
								assign node361 = (inp[5]) ? node363 : 13'b0000000111111;
									assign node363 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node366 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node369 = (inp[0]) ? node381 : node370;
							assign node370 = (inp[12]) ? node376 : node371;
								assign node371 = (inp[3]) ? node373 : 13'b0000001111111;
									assign node373 = (inp[4]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node376 = (inp[4]) ? node378 : 13'b0000000011111;
									assign node378 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node381 = (inp[7]) ? node383 : 13'b0000000011111;
								assign node383 = (inp[6]) ? 13'b0000000000111 : 13'b0000000000011;
			assign node386 = (inp[8]) ? node444 : node387;
				assign node387 = (inp[3]) ? node417 : node388;
					assign node388 = (inp[0]) ? node402 : node389;
						assign node389 = (inp[10]) ? node399 : node390;
							assign node390 = (inp[7]) ? node394 : node391;
								assign node391 = (inp[12]) ? 13'b0000111111111 : 13'b0000011111111;
								assign node394 = (inp[2]) ? node396 : 13'b0000011111111;
									assign node396 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node399 = (inp[5]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node402 = (inp[6]) ? node412 : node403;
							assign node403 = (inp[2]) ? node407 : node404;
								assign node404 = (inp[7]) ? 13'b0000011111111 : 13'b0000001111111;
								assign node407 = (inp[9]) ? node409 : 13'b0000000111111;
									assign node409 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node412 = (inp[12]) ? node414 : 13'b0000000011111;
								assign node414 = (inp[9]) ? 13'b0000000011111 : 13'b0000001111111;
					assign node417 = (inp[2]) ? node425 : node418;
						assign node418 = (inp[0]) ? node422 : node419;
							assign node419 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node422 = (inp[6]) ? 13'b0000000111111 : 13'b0000000001111;
						assign node425 = (inp[0]) ? node435 : node426;
							assign node426 = (inp[7]) ? node428 : 13'b0000000111111;
								assign node428 = (inp[12]) ? node432 : node429;
									assign node429 = (inp[9]) ? 13'b0000000111111 : 13'b0000000011111;
									assign node432 = (inp[4]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node435 = (inp[12]) ? node441 : node436;
								assign node436 = (inp[7]) ? node438 : 13'b0000000011111;
									assign node438 = (inp[4]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node441 = (inp[7]) ? 13'b0000000000011 : 13'b0000000000111;
				assign node444 = (inp[5]) ? node472 : node445;
					assign node445 = (inp[12]) ? node455 : node446;
						assign node446 = (inp[2]) ? node452 : node447;
							assign node447 = (inp[3]) ? 13'b0000001111111 : node448;
								assign node448 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node452 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node455 = (inp[3]) ? node461 : node456;
							assign node456 = (inp[6]) ? node458 : 13'b0000001111111;
								assign node458 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node461 = (inp[0]) ? node467 : node462;
								assign node462 = (inp[6]) ? 13'b0000000011111 : node463;
									assign node463 = (inp[10]) ? 13'b0000000111111 : 13'b0000000011111;
								assign node467 = (inp[7]) ? 13'b0000000001111 : node468;
									assign node468 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node472 = (inp[6]) ? node492 : node473;
						assign node473 = (inp[3]) ? node485 : node474;
							assign node474 = (inp[7]) ? node480 : node475;
								assign node475 = (inp[0]) ? node477 : 13'b0000001111111;
									assign node477 = (inp[10]) ? 13'b0000000111111 : 13'b0000000011111;
								assign node480 = (inp[0]) ? node482 : 13'b0000000011111;
									assign node482 = (inp[4]) ? 13'b0000000001111 : 13'b0000000001111;
							assign node485 = (inp[0]) ? 13'b0000000000111 : node486;
								assign node486 = (inp[4]) ? node488 : 13'b0000000011111;
									assign node488 = (inp[10]) ? 13'b0000000001111 : 13'b0000000001111;
						assign node492 = (inp[10]) ? node502 : node493;
							assign node493 = (inp[4]) ? node499 : node494;
								assign node494 = (inp[0]) ? node496 : 13'b0000000111111;
									assign node496 = (inp[9]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node499 = (inp[3]) ? 13'b0000000001111 : 13'b0000000000111;
							assign node502 = (inp[9]) ? 13'b0000000000011 : node503;
								assign node503 = (inp[2]) ? 13'b0000000000111 : node504;
									assign node504 = (inp[3]) ? 13'b0000000011111 : 13'b0000000001111;

endmodule