module dtc_split125_bm23 (
	input  wire [12-1:0] inp,
	output wire [12-1:0] outp
);

	wire [12-1:0] node1;
	wire [12-1:0] node2;
	wire [12-1:0] node3;
	wire [12-1:0] node4;
	wire [12-1:0] node5;
	wire [12-1:0] node6;
	wire [12-1:0] node7;
	wire [12-1:0] node8;
	wire [12-1:0] node11;
	wire [12-1:0] node14;
	wire [12-1:0] node17;
	wire [12-1:0] node19;
	wire [12-1:0] node22;
	wire [12-1:0] node23;
	wire [12-1:0] node24;
	wire [12-1:0] node27;
	wire [12-1:0] node29;
	wire [12-1:0] node32;
	wire [12-1:0] node33;
	wire [12-1:0] node36;
	wire [12-1:0] node38;
	wire [12-1:0] node41;
	wire [12-1:0] node42;
	wire [12-1:0] node43;
	wire [12-1:0] node45;
	wire [12-1:0] node46;
	wire [12-1:0] node50;
	wire [12-1:0] node51;
	wire [12-1:0] node54;
	wire [12-1:0] node56;
	wire [12-1:0] node59;
	wire [12-1:0] node60;
	wire [12-1:0] node61;
	wire [12-1:0] node65;
	wire [12-1:0] node67;
	wire [12-1:0] node70;
	wire [12-1:0] node71;
	wire [12-1:0] node72;
	wire [12-1:0] node73;
	wire [12-1:0] node74;
	wire [12-1:0] node76;
	wire [12-1:0] node79;
	wire [12-1:0] node82;
	wire [12-1:0] node83;
	wire [12-1:0] node84;
	wire [12-1:0] node88;
	wire [12-1:0] node91;
	wire [12-1:0] node92;
	wire [12-1:0] node93;
	wire [12-1:0] node94;
	wire [12-1:0] node98;
	wire [12-1:0] node101;
	wire [12-1:0] node103;
	wire [12-1:0] node106;
	wire [12-1:0] node107;
	wire [12-1:0] node108;
	wire [12-1:0] node109;
	wire [12-1:0] node110;
	wire [12-1:0] node114;
	wire [12-1:0] node117;
	wire [12-1:0] node118;
	wire [12-1:0] node121;
	wire [12-1:0] node122;
	wire [12-1:0] node125;
	wire [12-1:0] node128;
	wire [12-1:0] node129;
	wire [12-1:0] node131;
	wire [12-1:0] node132;
	wire [12-1:0] node136;
	wire [12-1:0] node138;
	wire [12-1:0] node141;
	wire [12-1:0] node142;
	wire [12-1:0] node143;
	wire [12-1:0] node144;
	wire [12-1:0] node145;
	wire [12-1:0] node146;
	wire [12-1:0] node147;
	wire [12-1:0] node151;
	wire [12-1:0] node153;
	wire [12-1:0] node156;
	wire [12-1:0] node157;
	wire [12-1:0] node159;
	wire [12-1:0] node163;
	wire [12-1:0] node164;
	wire [12-1:0] node165;
	wire [12-1:0] node166;
	wire [12-1:0] node170;
	wire [12-1:0] node171;
	wire [12-1:0] node174;
	wire [12-1:0] node177;
	wire [12-1:0] node178;
	wire [12-1:0] node181;
	wire [12-1:0] node182;
	wire [12-1:0] node186;
	wire [12-1:0] node187;
	wire [12-1:0] node188;
	wire [12-1:0] node189;
	wire [12-1:0] node192;
	wire [12-1:0] node196;
	wire [12-1:0] node197;
	wire [12-1:0] node200;
	wire [12-1:0] node201;
	wire [12-1:0] node203;
	wire [12-1:0] node206;
	wire [12-1:0] node209;
	wire [12-1:0] node210;
	wire [12-1:0] node211;
	wire [12-1:0] node212;
	wire [12-1:0] node213;
	wire [12-1:0] node214;
	wire [12-1:0] node217;
	wire [12-1:0] node220;
	wire [12-1:0] node222;
	wire [12-1:0] node225;
	wire [12-1:0] node226;
	wire [12-1:0] node227;
	wire [12-1:0] node231;
	wire [12-1:0] node233;
	wire [12-1:0] node236;
	wire [12-1:0] node237;
	wire [12-1:0] node238;
	wire [12-1:0] node241;
	wire [12-1:0] node242;
	wire [12-1:0] node246;
	wire [12-1:0] node247;
	wire [12-1:0] node249;
	wire [12-1:0] node252;
	wire [12-1:0] node253;
	wire [12-1:0] node257;
	wire [12-1:0] node258;
	wire [12-1:0] node259;
	wire [12-1:0] node261;
	wire [12-1:0] node263;
	wire [12-1:0] node266;
	wire [12-1:0] node267;
	wire [12-1:0] node268;
	wire [12-1:0] node273;
	wire [12-1:0] node274;
	wire [12-1:0] node275;
	wire [12-1:0] node276;
	wire [12-1:0] node279;
	wire [12-1:0] node282;
	wire [12-1:0] node284;
	wire [12-1:0] node287;
	wire [12-1:0] node288;
	wire [12-1:0] node290;
	wire [12-1:0] node293;
	wire [12-1:0] node295;
	wire [12-1:0] node298;
	wire [12-1:0] node299;
	wire [12-1:0] node300;
	wire [12-1:0] node301;
	wire [12-1:0] node302;
	wire [12-1:0] node303;
	wire [12-1:0] node304;
	wire [12-1:0] node306;
	wire [12-1:0] node309;
	wire [12-1:0] node310;
	wire [12-1:0] node313;
	wire [12-1:0] node316;
	wire [12-1:0] node318;
	wire [12-1:0] node320;
	wire [12-1:0] node323;
	wire [12-1:0] node324;
	wire [12-1:0] node325;
	wire [12-1:0] node326;
	wire [12-1:0] node331;
	wire [12-1:0] node332;
	wire [12-1:0] node333;
	wire [12-1:0] node338;
	wire [12-1:0] node339;
	wire [12-1:0] node340;
	wire [12-1:0] node341;
	wire [12-1:0] node344;
	wire [12-1:0] node346;
	wire [12-1:0] node349;
	wire [12-1:0] node351;
	wire [12-1:0] node353;
	wire [12-1:0] node356;
	wire [12-1:0] node357;
	wire [12-1:0] node358;
	wire [12-1:0] node360;
	wire [12-1:0] node363;
	wire [12-1:0] node364;
	wire [12-1:0] node367;
	wire [12-1:0] node370;
	wire [12-1:0] node372;
	wire [12-1:0] node375;
	wire [12-1:0] node376;
	wire [12-1:0] node377;
	wire [12-1:0] node378;
	wire [12-1:0] node379;
	wire [12-1:0] node381;
	wire [12-1:0] node384;
	wire [12-1:0] node387;
	wire [12-1:0] node388;
	wire [12-1:0] node389;
	wire [12-1:0] node392;
	wire [12-1:0] node395;
	wire [12-1:0] node396;
	wire [12-1:0] node399;
	wire [12-1:0] node402;
	wire [12-1:0] node403;
	wire [12-1:0] node405;
	wire [12-1:0] node407;
	wire [12-1:0] node410;
	wire [12-1:0] node411;
	wire [12-1:0] node415;
	wire [12-1:0] node416;
	wire [12-1:0] node417;
	wire [12-1:0] node419;
	wire [12-1:0] node422;
	wire [12-1:0] node423;
	wire [12-1:0] node427;
	wire [12-1:0] node428;
	wire [12-1:0] node430;
	wire [12-1:0] node431;
	wire [12-1:0] node435;
	wire [12-1:0] node436;
	wire [12-1:0] node437;
	wire [12-1:0] node441;
	wire [12-1:0] node443;
	wire [12-1:0] node446;
	wire [12-1:0] node447;
	wire [12-1:0] node448;
	wire [12-1:0] node449;
	wire [12-1:0] node450;
	wire [12-1:0] node451;
	wire [12-1:0] node453;
	wire [12-1:0] node456;
	wire [12-1:0] node458;
	wire [12-1:0] node461;
	wire [12-1:0] node462;
	wire [12-1:0] node463;
	wire [12-1:0] node467;
	wire [12-1:0] node468;
	wire [12-1:0] node472;
	wire [12-1:0] node473;
	wire [12-1:0] node474;
	wire [12-1:0] node476;
	wire [12-1:0] node479;
	wire [12-1:0] node482;
	wire [12-1:0] node483;
	wire [12-1:0] node484;
	wire [12-1:0] node487;
	wire [12-1:0] node490;
	wire [12-1:0] node493;
	wire [12-1:0] node494;
	wire [12-1:0] node495;
	wire [12-1:0] node496;
	wire [12-1:0] node500;
	wire [12-1:0] node501;
	wire [12-1:0] node502;
	wire [12-1:0] node505;
	wire [12-1:0] node508;
	wire [12-1:0] node510;
	wire [12-1:0] node513;
	wire [12-1:0] node514;
	wire [12-1:0] node516;
	wire [12-1:0] node517;
	wire [12-1:0] node520;
	wire [12-1:0] node523;
	wire [12-1:0] node524;
	wire [12-1:0] node525;
	wire [12-1:0] node528;
	wire [12-1:0] node531;
	wire [12-1:0] node533;
	wire [12-1:0] node536;
	wire [12-1:0] node537;
	wire [12-1:0] node538;
	wire [12-1:0] node539;
	wire [12-1:0] node540;
	wire [12-1:0] node541;
	wire [12-1:0] node546;
	wire [12-1:0] node548;
	wire [12-1:0] node551;
	wire [12-1:0] node552;
	wire [12-1:0] node553;
	wire [12-1:0] node554;
	wire [12-1:0] node558;
	wire [12-1:0] node559;
	wire [12-1:0] node562;
	wire [12-1:0] node565;
	wire [12-1:0] node566;
	wire [12-1:0] node567;
	wire [12-1:0] node571;
	wire [12-1:0] node572;
	wire [12-1:0] node576;
	wire [12-1:0] node577;
	wire [12-1:0] node578;
	wire [12-1:0] node579;
	wire [12-1:0] node582;
	wire [12-1:0] node583;
	wire [12-1:0] node587;
	wire [12-1:0] node588;
	wire [12-1:0] node591;
	wire [12-1:0] node593;
	wire [12-1:0] node596;
	wire [12-1:0] node597;
	wire [12-1:0] node598;
	wire [12-1:0] node599;
	wire [12-1:0] node602;

	assign outp = (inp[4]) ? node298 : node1;
		assign node1 = (inp[11]) ? node141 : node2;
			assign node2 = (inp[5]) ? node70 : node3;
				assign node3 = (inp[6]) ? node41 : node4;
					assign node4 = (inp[8]) ? node22 : node5;
						assign node5 = (inp[0]) ? node17 : node6;
							assign node6 = (inp[9]) ? node14 : node7;
								assign node7 = (inp[3]) ? node11 : node8;
									assign node8 = (inp[2]) ? 12'b001111111111 : 12'b001111111111;
									assign node11 = (inp[1]) ? 12'b000111111111 : 12'b001111111111;
								assign node14 = (inp[10]) ? 12'b000011111111 : 12'b000111111111;
							assign node17 = (inp[10]) ? node19 : 12'b000111111111;
								assign node19 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
						assign node22 = (inp[7]) ? node32 : node23;
							assign node23 = (inp[9]) ? node27 : node24;
								assign node24 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
								assign node27 = (inp[10]) ? node29 : 12'b000011111111;
									assign node29 = (inp[1]) ? 12'b000011111111 : 12'b000001111111;
							assign node32 = (inp[1]) ? node36 : node33;
								assign node33 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
								assign node36 = (inp[9]) ? node38 : 12'b000001111111;
									assign node38 = (inp[0]) ? 12'b000001111111 : 12'b000000111111;
					assign node41 = (inp[0]) ? node59 : node42;
						assign node42 = (inp[10]) ? node50 : node43;
							assign node43 = (inp[2]) ? node45 : 12'b000111111111;
								assign node45 = (inp[9]) ? 12'b000011111111 : node46;
									assign node46 = (inp[7]) ? 12'b000011111111 : 12'b000111111111;
							assign node50 = (inp[7]) ? node54 : node51;
								assign node51 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
								assign node54 = (inp[2]) ? node56 : 12'b000001111111;
									assign node56 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
						assign node59 = (inp[1]) ? node65 : node60;
							assign node60 = (inp[3]) ? 12'b000001111111 : node61;
								assign node61 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
							assign node65 = (inp[2]) ? node67 : 12'b000001111111;
								assign node67 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
				assign node70 = (inp[3]) ? node106 : node71;
					assign node71 = (inp[2]) ? node91 : node72;
						assign node72 = (inp[7]) ? node82 : node73;
							assign node73 = (inp[10]) ? node79 : node74;
								assign node74 = (inp[6]) ? node76 : 12'b000111111111;
									assign node76 = (inp[8]) ? 12'b000011111111 : 12'b000011111111;
								assign node79 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
							assign node82 = (inp[8]) ? node88 : node83;
								assign node83 = (inp[9]) ? 12'b000001111111 : node84;
									assign node84 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
								assign node88 = (inp[10]) ? 12'b000000111111 : 12'b000001111111;
						assign node91 = (inp[0]) ? node101 : node92;
							assign node92 = (inp[9]) ? node98 : node93;
								assign node93 = (inp[6]) ? 12'b000001111111 : node94;
									assign node94 = (inp[8]) ? 12'b000011111111 : 12'b000011111111;
								assign node98 = (inp[10]) ? 12'b000000111111 : 12'b000001111111;
							assign node101 = (inp[1]) ? node103 : 12'b000000111111;
								assign node103 = (inp[6]) ? 12'b000000011111 : 12'b000001111111;
					assign node106 = (inp[2]) ? node128 : node107;
						assign node107 = (inp[7]) ? node117 : node108;
							assign node108 = (inp[6]) ? node114 : node109;
								assign node109 = (inp[10]) ? 12'b000001111111 : node110;
									assign node110 = (inp[1]) ? 12'b000011111111 : 12'b000111111111;
								assign node114 = (inp[1]) ? 12'b000000111111 : 12'b000011111111;
							assign node117 = (inp[8]) ? node121 : node118;
								assign node118 = (inp[10]) ? 12'b000000111111 : 12'b000011111111;
								assign node121 = (inp[6]) ? node125 : node122;
									assign node122 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
									assign node125 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
						assign node128 = (inp[8]) ? node136 : node129;
							assign node129 = (inp[0]) ? node131 : 12'b000000111111;
								assign node131 = (inp[1]) ? 12'b000000011111 : node132;
									assign node132 = (inp[10]) ? 12'b000001111111 : 12'b000000011111;
							assign node136 = (inp[6]) ? node138 : 12'b000000011111;
								assign node138 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
			assign node141 = (inp[2]) ? node209 : node142;
				assign node142 = (inp[3]) ? node186 : node143;
					assign node143 = (inp[5]) ? node163 : node144;
						assign node144 = (inp[7]) ? node156 : node145;
							assign node145 = (inp[8]) ? node151 : node146;
								assign node146 = (inp[10]) ? 12'b000011111111 : node147;
									assign node147 = (inp[1]) ? 12'b000111111111 : 12'b000111111111;
								assign node151 = (inp[6]) ? node153 : 12'b000011111111;
									assign node153 = (inp[9]) ? 12'b000011111111 : 12'b000011111111;
							assign node156 = (inp[8]) ? 12'b000001111111 : node157;
								assign node157 = (inp[1]) ? node159 : 12'b000011111111;
									assign node159 = (inp[6]) ? 12'b000000111111 : 12'b000011111111;
						assign node163 = (inp[0]) ? node177 : node164;
							assign node164 = (inp[8]) ? node170 : node165;
								assign node165 = (inp[9]) ? 12'b000011111111 : node166;
									assign node166 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
								assign node170 = (inp[10]) ? node174 : node171;
									assign node171 = (inp[6]) ? 12'b000001111111 : 12'b000001111111;
									assign node174 = (inp[6]) ? 12'b000000011111 : 12'b000001111111;
							assign node177 = (inp[1]) ? node181 : node178;
								assign node178 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
								assign node181 = (inp[6]) ? 12'b000000011111 : node182;
									assign node182 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
					assign node186 = (inp[7]) ? node196 : node187;
						assign node187 = (inp[1]) ? 12'b000000111111 : node188;
							assign node188 = (inp[9]) ? node192 : node189;
								assign node189 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
								assign node192 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
						assign node196 = (inp[8]) ? node200 : node197;
							assign node197 = (inp[9]) ? 12'b000001111111 : 12'b000000111111;
							assign node200 = (inp[5]) ? node206 : node201;
								assign node201 = (inp[10]) ? node203 : 12'b000000111111;
									assign node203 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
								assign node206 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
				assign node209 = (inp[9]) ? node257 : node210;
					assign node210 = (inp[0]) ? node236 : node211;
						assign node211 = (inp[10]) ? node225 : node212;
							assign node212 = (inp[6]) ? node220 : node213;
								assign node213 = (inp[3]) ? node217 : node214;
									assign node214 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
									assign node217 = (inp[5]) ? 12'b000001111111 : 12'b000001111111;
								assign node220 = (inp[7]) ? node222 : 12'b000001111111;
									assign node222 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
							assign node225 = (inp[5]) ? node231 : node226;
								assign node226 = (inp[7]) ? 12'b000000111111 : node227;
									assign node227 = (inp[1]) ? 12'b000001111111 : 12'b000011111111;
								assign node231 = (inp[6]) ? node233 : 12'b000000111111;
									assign node233 = (inp[1]) ? 12'b000000011111 : 12'b000001111111;
						assign node236 = (inp[1]) ? node246 : node237;
							assign node237 = (inp[5]) ? node241 : node238;
								assign node238 = (inp[10]) ? 12'b000000111111 : 12'b000001111111;
								assign node241 = (inp[8]) ? 12'b000000011111 : node242;
									assign node242 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
							assign node246 = (inp[8]) ? node252 : node247;
								assign node247 = (inp[6]) ? node249 : 12'b000000111111;
									assign node249 = (inp[10]) ? 12'b000000001111 : 12'b000000111111;
								assign node252 = (inp[10]) ? 12'b000000001111 : node253;
									assign node253 = (inp[3]) ? 12'b000000001111 : 12'b000000111111;
					assign node257 = (inp[7]) ? node273 : node258;
						assign node258 = (inp[5]) ? node266 : node259;
							assign node259 = (inp[6]) ? node261 : 12'b000001111111;
								assign node261 = (inp[0]) ? node263 : 12'b000000111111;
									assign node263 = (inp[10]) ? 12'b000000001111 : 12'b000000011111;
							assign node266 = (inp[8]) ? 12'b000000011111 : node267;
								assign node267 = (inp[1]) ? 12'b000000001111 : node268;
									assign node268 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
						assign node273 = (inp[8]) ? node287 : node274;
							assign node274 = (inp[6]) ? node282 : node275;
								assign node275 = (inp[1]) ? node279 : node276;
									assign node276 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
									assign node279 = (inp[10]) ? 12'b000000001111 : 12'b000000011111;
								assign node282 = (inp[5]) ? node284 : 12'b000000011111;
									assign node284 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
							assign node287 = (inp[6]) ? node293 : node288;
								assign node288 = (inp[0]) ? node290 : 12'b000000001111;
									assign node290 = (inp[3]) ? 12'b000000000111 : 12'b000000001111;
								assign node293 = (inp[3]) ? node295 : 12'b000000001111;
									assign node295 = (inp[5]) ? 12'b000000000001 : 12'b000000000011;
		assign node298 = (inp[10]) ? node446 : node299;
			assign node299 = (inp[5]) ? node375 : node300;
				assign node300 = (inp[1]) ? node338 : node301;
					assign node301 = (inp[7]) ? node323 : node302;
						assign node302 = (inp[6]) ? node316 : node303;
							assign node303 = (inp[11]) ? node309 : node304;
								assign node304 = (inp[8]) ? node306 : 12'b000111111111;
									assign node306 = (inp[0]) ? 12'b000011111111 : 12'b000111111111;
								assign node309 = (inp[2]) ? node313 : node310;
									assign node310 = (inp[0]) ? 12'b000011111111 : 12'b000011111111;
									assign node313 = (inp[8]) ? 12'b000000111111 : 12'b000011111111;
							assign node316 = (inp[9]) ? node318 : 12'b000011111111;
								assign node318 = (inp[2]) ? node320 : 12'b000001111111;
									assign node320 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
						assign node323 = (inp[2]) ? node331 : node324;
							assign node324 = (inp[6]) ? 12'b000000111111 : node325;
								assign node325 = (inp[9]) ? 12'b000001111111 : node326;
									assign node326 = (inp[11]) ? 12'b000011111111 : 12'b000011111111;
							assign node331 = (inp[9]) ? 12'b000000011111 : node332;
								assign node332 = (inp[11]) ? 12'b000000011111 : node333;
									assign node333 = (inp[0]) ? 12'b000000111111 : 12'b000001111111;
					assign node338 = (inp[6]) ? node356 : node339;
						assign node339 = (inp[3]) ? node349 : node340;
							assign node340 = (inp[2]) ? node344 : node341;
								assign node341 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
								assign node344 = (inp[8]) ? node346 : 12'b000001111111;
									assign node346 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
							assign node349 = (inp[9]) ? node351 : 12'b000001111111;
								assign node351 = (inp[0]) ? node353 : 12'b000000111111;
									assign node353 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
						assign node356 = (inp[3]) ? node370 : node357;
							assign node357 = (inp[2]) ? node363 : node358;
								assign node358 = (inp[9]) ? node360 : 12'b000001111111;
									assign node360 = (inp[8]) ? 12'b000001111111 : 12'b000000111111;
								assign node363 = (inp[11]) ? node367 : node364;
									assign node364 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
									assign node367 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
							assign node370 = (inp[2]) ? node372 : 12'b000000011111;
								assign node372 = (inp[7]) ? 12'b000000011111 : 12'b000000001111;
				assign node375 = (inp[1]) ? node415 : node376;
					assign node376 = (inp[2]) ? node402 : node377;
						assign node377 = (inp[6]) ? node387 : node378;
							assign node378 = (inp[3]) ? node384 : node379;
								assign node379 = (inp[7]) ? node381 : 12'b000011111111;
									assign node381 = (inp[11]) ? 12'b000000111111 : 12'b000011111111;
								assign node384 = (inp[9]) ? 12'b000001111111 : 12'b000000111111;
							assign node387 = (inp[3]) ? node395 : node388;
								assign node388 = (inp[7]) ? node392 : node389;
									assign node389 = (inp[8]) ? 12'b000001111111 : 12'b000000111111;
									assign node392 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
								assign node395 = (inp[0]) ? node399 : node396;
									assign node396 = (inp[9]) ? 12'b000000011111 : 12'b000001111111;
									assign node399 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
						assign node402 = (inp[8]) ? node410 : node403;
							assign node403 = (inp[3]) ? node405 : 12'b000001111111;
								assign node405 = (inp[9]) ? node407 : 12'b000000111111;
									assign node407 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
							assign node410 = (inp[11]) ? 12'b000000011111 : node411;
								assign node411 = (inp[7]) ? 12'b000000011111 : 12'b000000111111;
					assign node415 = (inp[8]) ? node427 : node416;
						assign node416 = (inp[0]) ? node422 : node417;
							assign node417 = (inp[2]) ? node419 : 12'b000011111111;
								assign node419 = (inp[7]) ? 12'b000000111111 : 12'b000001111111;
							assign node422 = (inp[9]) ? 12'b000000001111 : node423;
								assign node423 = (inp[11]) ? 12'b000000111111 : 12'b000000011111;
						assign node427 = (inp[3]) ? node435 : node428;
							assign node428 = (inp[6]) ? node430 : 12'b000000011111;
								assign node430 = (inp[9]) ? 12'b000000001111 : node431;
									assign node431 = (inp[11]) ? 12'b000000011111 : 12'b000000011111;
							assign node435 = (inp[0]) ? node441 : node436;
								assign node436 = (inp[9]) ? 12'b000000001111 : node437;
									assign node437 = (inp[7]) ? 12'b000000001111 : 12'b000001111111;
								assign node441 = (inp[7]) ? node443 : 12'b000000001111;
									assign node443 = (inp[9]) ? 12'b000000000111 : 12'b000000000011;
			assign node446 = (inp[9]) ? node536 : node447;
				assign node447 = (inp[7]) ? node493 : node448;
					assign node448 = (inp[2]) ? node472 : node449;
						assign node449 = (inp[1]) ? node461 : node450;
							assign node450 = (inp[11]) ? node456 : node451;
								assign node451 = (inp[5]) ? node453 : 12'b000011111111;
									assign node453 = (inp[0]) ? 12'b000001111111 : 12'b000000111111;
								assign node456 = (inp[0]) ? node458 : 12'b000001111111;
									assign node458 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
							assign node461 = (inp[0]) ? node467 : node462;
								assign node462 = (inp[3]) ? 12'b000000111111 : node463;
									assign node463 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
								assign node467 = (inp[6]) ? 12'b000000011111 : node468;
									assign node468 = (inp[5]) ? 12'b000000111111 : 12'b000000011111;
						assign node472 = (inp[6]) ? node482 : node473;
							assign node473 = (inp[11]) ? node479 : node474;
								assign node474 = (inp[3]) ? node476 : 12'b000001111111;
									assign node476 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
								assign node479 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
							assign node482 = (inp[1]) ? node490 : node483;
								assign node483 = (inp[11]) ? node487 : node484;
									assign node484 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
									assign node487 = (inp[5]) ? 12'b000000011111 : 12'b000000011111;
								assign node490 = (inp[8]) ? 12'b000000001111 : 12'b000000111111;
					assign node493 = (inp[8]) ? node513 : node494;
						assign node494 = (inp[0]) ? node500 : node495;
							assign node495 = (inp[5]) ? 12'b000000111111 : node496;
								assign node496 = (inp[6]) ? 12'b000001111111 : 12'b000111111111;
							assign node500 = (inp[6]) ? node508 : node501;
								assign node501 = (inp[5]) ? node505 : node502;
									assign node502 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
									assign node505 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
								assign node508 = (inp[1]) ? node510 : 12'b000000001111;
									assign node510 = (inp[2]) ? 12'b000000000111 : 12'b000000001111;
						assign node513 = (inp[11]) ? node523 : node514;
							assign node514 = (inp[1]) ? node516 : 12'b000000111111;
								assign node516 = (inp[3]) ? node520 : node517;
									assign node517 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
									assign node520 = (inp[5]) ? 12'b000000000111 : 12'b000000011111;
							assign node523 = (inp[0]) ? node531 : node524;
								assign node524 = (inp[3]) ? node528 : node525;
									assign node525 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
									assign node528 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
								assign node531 = (inp[5]) ? node533 : 12'b000000001111;
									assign node533 = (inp[2]) ? 12'b000000000011 : 12'b000000000111;
				assign node536 = (inp[11]) ? node576 : node537;
					assign node537 = (inp[8]) ? node551 : node538;
						assign node538 = (inp[7]) ? node546 : node539;
							assign node539 = (inp[2]) ? 12'b000000011111 : node540;
								assign node540 = (inp[0]) ? 12'b000000011111 : node541;
									assign node541 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
							assign node546 = (inp[3]) ? node548 : 12'b000000011111;
								assign node548 = (inp[2]) ? 12'b000000000111 : 12'b000000011111;
						assign node551 = (inp[6]) ? node565 : node552;
							assign node552 = (inp[3]) ? node558 : node553;
								assign node553 = (inp[0]) ? 12'b000000001111 : node554;
									assign node554 = (inp[7]) ? 12'b000000111111 : 12'b000000011111;
								assign node558 = (inp[5]) ? node562 : node559;
									assign node559 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
									assign node562 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
							assign node565 = (inp[1]) ? node571 : node566;
								assign node566 = (inp[3]) ? 12'b000000001111 : node567;
									assign node567 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
								assign node571 = (inp[7]) ? 12'b000000000111 : node572;
									assign node572 = (inp[0]) ? 12'b000000000111 : 12'b000000001111;
					assign node576 = (inp[2]) ? node596 : node577;
						assign node577 = (inp[3]) ? node587 : node578;
							assign node578 = (inp[7]) ? node582 : node579;
								assign node579 = (inp[6]) ? 12'b000000011111 : 12'b000001111111;
								assign node582 = (inp[6]) ? 12'b000000001111 : node583;
									assign node583 = (inp[0]) ? 12'b000000011111 : 12'b000000001111;
							assign node587 = (inp[5]) ? node591 : node588;
								assign node588 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
								assign node591 = (inp[8]) ? node593 : 12'b000000001111;
									assign node593 = (inp[7]) ? 12'b000000000111 : 12'b000000001111;
						assign node596 = (inp[8]) ? 12'b000000001111 : node597;
							assign node597 = (inp[3]) ? 12'b000000000111 : node598;
								assign node598 = (inp[5]) ? node602 : node599;
									assign node599 = (inp[7]) ? 12'b000000001111 : 12'b000000001111;
									assign node602 = (inp[7]) ? 12'b000000000011 : 12'b000000000111;

endmodule