module dtc_split33_bm96 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node38;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node50;
	wire [3-1:0] node53;
	wire [3-1:0] node55;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node62;
	wire [3-1:0] node64;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node139;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node149;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node183;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node204;

	assign outp = (inp[6]) ? node2 : 3'b000;
		assign node2 = (inp[7]) ? node18 : node3;
			assign node3 = (inp[3]) ? node5 : 3'b000;
				assign node5 = (inp[10]) ? 3'b000 : node6;
					assign node6 = (inp[1]) ? node8 : 3'b000;
						assign node8 = (inp[8]) ? node10 : 3'b000;
							assign node10 = (inp[2]) ? node12 : 3'b000;
								assign node12 = (inp[9]) ? 3'b000 : node13;
									assign node13 = (inp[4]) ? 3'b100 : 3'b000;
			assign node18 = (inp[3]) ? node98 : node19;
				assign node19 = (inp[4]) ? node31 : node20;
					assign node20 = (inp[9]) ? node22 : 3'b011;
						assign node22 = (inp[1]) ? 3'b011 : node23;
							assign node23 = (inp[10]) ? node27 : node24;
								assign node24 = (inp[5]) ? 3'b011 : 3'b111;
								assign node27 = (inp[5]) ? 3'b101 : 3'b011;
					assign node31 = (inp[0]) ? node67 : node32;
						assign node32 = (inp[1]) ? node58 : node33;
							assign node33 = (inp[2]) ? node43 : node34;
								assign node34 = (inp[10]) ? 3'b010 : node35;
									assign node35 = (inp[8]) ? 3'b010 : node36;
										assign node36 = (inp[9]) ? node38 : 3'b001;
											assign node38 = (inp[5]) ? 3'b001 : 3'b010;
								assign node43 = (inp[11]) ? node53 : node44;
									assign node44 = (inp[5]) ? node46 : 3'b010;
										assign node46 = (inp[9]) ? node50 : node47;
											assign node47 = (inp[10]) ? 3'b010 : 3'b001;
											assign node50 = (inp[10]) ? 3'b001 : 3'b010;
									assign node53 = (inp[10]) ? node55 : 3'b001;
										assign node55 = (inp[9]) ? 3'b001 : 3'b010;
							assign node58 = (inp[11]) ? node60 : 3'b010;
								assign node60 = (inp[5]) ? node62 : 3'b010;
									assign node62 = (inp[2]) ? node64 : 3'b010;
										assign node64 = (inp[9]) ? 3'b001 : 3'b010;
						assign node67 = (inp[9]) ? node77 : node68;
							assign node68 = (inp[2]) ? node70 : 3'b001;
								assign node70 = (inp[8]) ? 3'b001 : node71;
									assign node71 = (inp[1]) ? node73 : 3'b001;
										assign node73 = (inp[11]) ? 3'b001 : 3'b010;
							assign node77 = (inp[1]) ? node91 : node78;
								assign node78 = (inp[10]) ? node84 : node79;
									assign node79 = (inp[11]) ? node81 : 3'b110;
										assign node81 = (inp[5]) ? 3'b001 : 3'b101;
									assign node84 = (inp[5]) ? node88 : node85;
										assign node85 = (inp[11]) ? 3'b001 : 3'b101;
										assign node88 = (inp[11]) ? 3'b010 : 3'b001;
								assign node91 = (inp[8]) ? node93 : 3'b010;
									assign node93 = (inp[11]) ? 3'b010 : node94;
										assign node94 = (inp[10]) ? 3'b010 : 3'b001;
				assign node98 = (inp[1]) ? node164 : node99;
					assign node99 = (inp[4]) ? node133 : node100;
						assign node100 = (inp[10]) ? node112 : node101;
							assign node101 = (inp[9]) ? node103 : 3'b111;
								assign node103 = (inp[8]) ? node109 : node104;
									assign node104 = (inp[0]) ? 3'b110 : node105;
										assign node105 = (inp[11]) ? 3'b111 : 3'b110;
									assign node109 = (inp[0]) ? 3'b111 : 3'b110;
							assign node112 = (inp[5]) ? node126 : node113;
								assign node113 = (inp[8]) ? node121 : node114;
									assign node114 = (inp[9]) ? node118 : node115;
										assign node115 = (inp[0]) ? 3'b111 : 3'b110;
										assign node118 = (inp[0]) ? 3'b110 : 3'b111;
									assign node121 = (inp[2]) ? 3'b110 : node122;
										assign node122 = (inp[0]) ? 3'b111 : 3'b110;
								assign node126 = (inp[9]) ? node130 : node127;
									assign node127 = (inp[0]) ? 3'b111 : 3'b110;
									assign node130 = (inp[2]) ? 3'b010 : 3'b011;
						assign node133 = (inp[0]) ? node153 : node134;
							assign node134 = (inp[9]) ? node142 : node135;
								assign node135 = (inp[10]) ? node139 : node136;
									assign node136 = (inp[2]) ? 3'b011 : 3'b111;
									assign node139 = (inp[11]) ? 3'b001 : 3'b101;
								assign node142 = (inp[2]) ? 3'b110 : node143;
									assign node143 = (inp[10]) ? node147 : node144;
										assign node144 = (inp[11]) ? 3'b110 : 3'b001;
										assign node147 = (inp[11]) ? node149 : 3'b110;
											assign node149 = (inp[5]) ? 3'b010 : 3'b110;
							assign node153 = (inp[9]) ? node155 : 3'b110;
								assign node155 = (inp[11]) ? node159 : node156;
									assign node156 = (inp[10]) ? 3'b100 : 3'b010;
									assign node159 = (inp[5]) ? node161 : 3'b100;
										assign node161 = (inp[10]) ? 3'b000 : 3'b100;
					assign node164 = (inp[4]) ? node194 : node165;
						assign node165 = (inp[10]) ? node189 : node166;
							assign node166 = (inp[5]) ? node182 : node167;
								assign node167 = (inp[11]) ? node177 : node168;
									assign node168 = (inp[2]) ? 3'b100 : node169;
										assign node169 = (inp[0]) ? node173 : node170;
											assign node170 = (inp[9]) ? 3'b101 : 3'b100;
											assign node173 = (inp[9]) ? 3'b100 : 3'b101;
									assign node177 = (inp[9]) ? node179 : 3'b100;
										assign node179 = (inp[0]) ? 3'b100 : 3'b101;
								assign node182 = (inp[9]) ? node186 : node183;
									assign node183 = (inp[0]) ? 3'b101 : 3'b100;
									assign node186 = (inp[0]) ? 3'b100 : 3'b101;
							assign node189 = (inp[9]) ? node191 : 3'b100;
								assign node191 = (inp[0]) ? 3'b100 : 3'b101;
						assign node194 = (inp[0]) ? node198 : node195;
							assign node195 = (inp[9]) ? 3'b010 : 3'b001;
							assign node198 = (inp[9]) ? 3'b000 : node199;
								assign node199 = (inp[10]) ? node203 : node200;
									assign node200 = (inp[2]) ? 3'b010 : 3'b100;
									assign node203 = (inp[11]) ? 3'b100 : node204;
										assign node204 = (inp[8]) ? 3'b010 : 3'b100;

endmodule