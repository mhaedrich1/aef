module dtc_split05_bm30 (
	input  wire [14-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node7;
	wire [8-1:0] node8;
	wire [8-1:0] node12;
	wire [8-1:0] node13;
	wire [8-1:0] node16;
	wire [8-1:0] node18;
	wire [8-1:0] node21;
	wire [8-1:0] node22;
	wire [8-1:0] node23;
	wire [8-1:0] node27;
	wire [8-1:0] node28;
	wire [8-1:0] node31;
	wire [8-1:0] node32;
	wire [8-1:0] node35;
	wire [8-1:0] node38;
	wire [8-1:0] node39;
	wire [8-1:0] node40;
	wire [8-1:0] node41;
	wire [8-1:0] node45;
	wire [8-1:0] node46;
	wire [8-1:0] node49;
	wire [8-1:0] node53;
	wire [8-1:0] node54;
	wire [8-1:0] node55;
	wire [8-1:0] node56;
	wire [8-1:0] node58;
	wire [8-1:0] node61;
	wire [8-1:0] node62;
	wire [8-1:0] node65;
	wire [8-1:0] node68;
	wire [8-1:0] node69;
	wire [8-1:0] node72;
	wire [8-1:0] node74;
	wire [8-1:0] node75;
	wire [8-1:0] node78;
	wire [8-1:0] node81;
	wire [8-1:0] node82;
	wire [8-1:0] node83;
	wire [8-1:0] node84;
	wire [8-1:0] node87;
	wire [8-1:0] node90;
	wire [8-1:0] node93;
	wire [8-1:0] node94;
	wire [8-1:0] node96;
	wire [8-1:0] node99;
	wire [8-1:0] node100;
	wire [8-1:0] node103;
	wire [8-1:0] node105;
	wire [8-1:0] node108;
	wire [8-1:0] node109;
	wire [8-1:0] node110;
	wire [8-1:0] node111;
	wire [8-1:0] node112;
	wire [8-1:0] node113;
	wire [8-1:0] node116;
	wire [8-1:0] node119;
	wire [8-1:0] node121;
	wire [8-1:0] node122;
	wire [8-1:0] node125;
	wire [8-1:0] node128;
	wire [8-1:0] node129;
	wire [8-1:0] node131;
	wire [8-1:0] node132;
	wire [8-1:0] node135;
	wire [8-1:0] node138;
	wire [8-1:0] node140;
	wire [8-1:0] node141;
	wire [8-1:0] node144;
	wire [8-1:0] node147;
	wire [8-1:0] node148;
	wire [8-1:0] node149;
	wire [8-1:0] node150;
	wire [8-1:0] node152;
	wire [8-1:0] node155;
	wire [8-1:0] node158;
	wire [8-1:0] node159;
	wire [8-1:0] node161;
	wire [8-1:0] node164;
	wire [8-1:0] node165;
	wire [8-1:0] node167;
	wire [8-1:0] node170;
	wire [8-1:0] node173;
	wire [8-1:0] node174;
	wire [8-1:0] node175;
	wire [8-1:0] node178;
	wire [8-1:0] node181;
	wire [8-1:0] node182;
	wire [8-1:0] node185;
	wire [8-1:0] node188;
	wire [8-1:0] node189;
	wire [8-1:0] node190;
	wire [8-1:0] node191;
	wire [8-1:0] node192;
	wire [8-1:0] node193;
	wire [8-1:0] node197;
	wire [8-1:0] node200;
	wire [8-1:0] node202;
	wire [8-1:0] node204;
	wire [8-1:0] node205;
	wire [8-1:0] node209;
	wire [8-1:0] node210;
	wire [8-1:0] node211;
	wire [8-1:0] node213;
	wire [8-1:0] node216;
	wire [8-1:0] node217;
	wire [8-1:0] node221;
	wire [8-1:0] node222;
	wire [8-1:0] node223;
	wire [8-1:0] node227;
	wire [8-1:0] node230;
	wire [8-1:0] node231;
	wire [8-1:0] node232;
	wire [8-1:0] node233;
	wire [8-1:0] node235;
	wire [8-1:0] node236;
	wire [8-1:0] node241;
	wire [8-1:0] node243;
	wire [8-1:0] node246;
	wire [8-1:0] node247;
	wire [8-1:0] node248;
	wire [8-1:0] node251;
	wire [8-1:0] node253;
	wire [8-1:0] node256;
	wire [8-1:0] node257;
	wire [8-1:0] node260;
	wire [8-1:0] node263;
	wire [8-1:0] node264;
	wire [8-1:0] node265;
	wire [8-1:0] node266;
	wire [8-1:0] node267;
	wire [8-1:0] node268;
	wire [8-1:0] node269;
	wire [8-1:0] node270;
	wire [8-1:0] node271;
	wire [8-1:0] node276;
	wire [8-1:0] node280;
	wire [8-1:0] node281;
	wire [8-1:0] node282;
	wire [8-1:0] node285;
	wire [8-1:0] node288;
	wire [8-1:0] node289;
	wire [8-1:0] node291;
	wire [8-1:0] node295;
	wire [8-1:0] node296;
	wire [8-1:0] node297;
	wire [8-1:0] node298;
	wire [8-1:0] node299;
	wire [8-1:0] node304;
	wire [8-1:0] node306;
	wire [8-1:0] node309;
	wire [8-1:0] node310;
	wire [8-1:0] node311;
	wire [8-1:0] node312;
	wire [8-1:0] node315;
	wire [8-1:0] node316;
	wire [8-1:0] node320;
	wire [8-1:0] node321;
	wire [8-1:0] node324;
	wire [8-1:0] node327;
	wire [8-1:0] node328;
	wire [8-1:0] node329;
	wire [8-1:0] node331;
	wire [8-1:0] node335;
	wire [8-1:0] node336;
	wire [8-1:0] node339;
	wire [8-1:0] node341;
	wire [8-1:0] node344;
	wire [8-1:0] node345;
	wire [8-1:0] node346;
	wire [8-1:0] node347;
	wire [8-1:0] node348;
	wire [8-1:0] node352;
	wire [8-1:0] node353;
	wire [8-1:0] node355;
	wire [8-1:0] node358;
	wire [8-1:0] node360;
	wire [8-1:0] node363;
	wire [8-1:0] node364;
	wire [8-1:0] node365;
	wire [8-1:0] node368;
	wire [8-1:0] node371;
	wire [8-1:0] node372;
	wire [8-1:0] node375;
	wire [8-1:0] node376;
	wire [8-1:0] node377;
	wire [8-1:0] node382;
	wire [8-1:0] node383;
	wire [8-1:0] node384;
	wire [8-1:0] node385;
	wire [8-1:0] node386;
	wire [8-1:0] node390;
	wire [8-1:0] node391;
	wire [8-1:0] node393;
	wire [8-1:0] node397;
	wire [8-1:0] node398;
	wire [8-1:0] node402;
	wire [8-1:0] node403;
	wire [8-1:0] node405;
	wire [8-1:0] node408;
	wire [8-1:0] node409;
	wire [8-1:0] node412;
	wire [8-1:0] node413;
	wire [8-1:0] node416;
	wire [8-1:0] node417;
	wire [8-1:0] node421;
	wire [8-1:0] node422;
	wire [8-1:0] node423;
	wire [8-1:0] node424;
	wire [8-1:0] node426;
	wire [8-1:0] node429;
	wire [8-1:0] node430;
	wire [8-1:0] node432;
	wire [8-1:0] node433;
	wire [8-1:0] node435;
	wire [8-1:0] node438;
	wire [8-1:0] node441;
	wire [8-1:0] node442;
	wire [8-1:0] node443;
	wire [8-1:0] node446;
	wire [8-1:0] node449;
	wire [8-1:0] node452;
	wire [8-1:0] node453;
	wire [8-1:0] node455;
	wire [8-1:0] node457;
	wire [8-1:0] node459;
	wire [8-1:0] node461;
	wire [8-1:0] node464;
	wire [8-1:0] node465;
	wire [8-1:0] node467;
	wire [8-1:0] node468;
	wire [8-1:0] node471;
	wire [8-1:0] node474;
	wire [8-1:0] node475;
	wire [8-1:0] node478;
	wire [8-1:0] node480;
	wire [8-1:0] node483;
	wire [8-1:0] node484;
	wire [8-1:0] node486;
	wire [8-1:0] node487;
	wire [8-1:0] node488;
	wire [8-1:0] node491;
	wire [8-1:0] node492;
	wire [8-1:0] node496;
	wire [8-1:0] node497;
	wire [8-1:0] node499;
	wire [8-1:0] node503;
	wire [8-1:0] node504;
	wire [8-1:0] node506;
	wire [8-1:0] node507;
	wire [8-1:0] node510;
	wire [8-1:0] node511;
	wire [8-1:0] node514;
	wire [8-1:0] node517;
	wire [8-1:0] node518;
	wire [8-1:0] node520;
	wire [8-1:0] node523;
	wire [8-1:0] node524;
	wire [8-1:0] node527;
	wire [8-1:0] node530;
	wire [8-1:0] node531;
	wire [8-1:0] node532;
	wire [8-1:0] node533;
	wire [8-1:0] node534;
	wire [8-1:0] node535;
	wire [8-1:0] node536;
	wire [8-1:0] node537;
	wire [8-1:0] node538;
	wire [8-1:0] node543;
	wire [8-1:0] node545;
	wire [8-1:0] node548;
	wire [8-1:0] node549;
	wire [8-1:0] node550;
	wire [8-1:0] node553;
	wire [8-1:0] node557;
	wire [8-1:0] node558;
	wire [8-1:0] node559;
	wire [8-1:0] node560;
	wire [8-1:0] node561;
	wire [8-1:0] node566;
	wire [8-1:0] node567;
	wire [8-1:0] node571;
	wire [8-1:0] node572;
	wire [8-1:0] node576;
	wire [8-1:0] node577;
	wire [8-1:0] node578;
	wire [8-1:0] node579;
	wire [8-1:0] node581;
	wire [8-1:0] node582;
	wire [8-1:0] node585;
	wire [8-1:0] node589;
	wire [8-1:0] node592;
	wire [8-1:0] node593;
	wire [8-1:0] node594;
	wire [8-1:0] node597;
	wire [8-1:0] node598;
	wire [8-1:0] node603;
	wire [8-1:0] node604;
	wire [8-1:0] node605;
	wire [8-1:0] node606;
	wire [8-1:0] node607;
	wire [8-1:0] node609;
	wire [8-1:0] node612;
	wire [8-1:0] node613;
	wire [8-1:0] node615;
	wire [8-1:0] node618;
	wire [8-1:0] node620;
	wire [8-1:0] node623;
	wire [8-1:0] node624;
	wire [8-1:0] node626;
	wire [8-1:0] node629;
	wire [8-1:0] node630;
	wire [8-1:0] node631;
	wire [8-1:0] node634;
	wire [8-1:0] node638;
	wire [8-1:0] node639;
	wire [8-1:0] node640;
	wire [8-1:0] node641;
	wire [8-1:0] node642;
	wire [8-1:0] node643;
	wire [8-1:0] node647;
	wire [8-1:0] node651;
	wire [8-1:0] node652;
	wire [8-1:0] node653;
	wire [8-1:0] node655;
	wire [8-1:0] node659;
	wire [8-1:0] node662;
	wire [8-1:0] node663;
	wire [8-1:0] node664;
	wire [8-1:0] node665;
	wire [8-1:0] node666;
	wire [8-1:0] node668;
	wire [8-1:0] node671;
	wire [8-1:0] node675;
	wire [8-1:0] node676;
	wire [8-1:0] node680;
	wire [8-1:0] node681;
	wire [8-1:0] node682;
	wire [8-1:0] node687;
	wire [8-1:0] node688;
	wire [8-1:0] node689;
	wire [8-1:0] node690;
	wire [8-1:0] node691;
	wire [8-1:0] node692;
	wire [8-1:0] node694;
	wire [8-1:0] node699;
	wire [8-1:0] node700;
	wire [8-1:0] node703;
	wire [8-1:0] node706;
	wire [8-1:0] node707;
	wire [8-1:0] node708;
	wire [8-1:0] node712;
	wire [8-1:0] node713;
	wire [8-1:0] node716;
	wire [8-1:0] node719;
	wire [8-1:0] node720;
	wire [8-1:0] node721;
	wire [8-1:0] node722;
	wire [8-1:0] node725;
	wire [8-1:0] node728;
	wire [8-1:0] node729;
	wire [8-1:0] node730;
	wire [8-1:0] node735;
	wire [8-1:0] node736;
	wire [8-1:0] node737;
	wire [8-1:0] node739;
	wire [8-1:0] node742;
	wire [8-1:0] node744;
	wire [8-1:0] node745;
	wire [8-1:0] node749;
	wire [8-1:0] node750;
	wire [8-1:0] node751;
	wire [8-1:0] node756;
	wire [8-1:0] node757;
	wire [8-1:0] node758;
	wire [8-1:0] node759;
	wire [8-1:0] node760;
	wire [8-1:0] node761;
	wire [8-1:0] node764;
	wire [8-1:0] node765;
	wire [8-1:0] node768;
	wire [8-1:0] node769;
	wire [8-1:0] node773;
	wire [8-1:0] node774;
	wire [8-1:0] node776;
	wire [8-1:0] node777;
	wire [8-1:0] node781;
	wire [8-1:0] node782;
	wire [8-1:0] node785;
	wire [8-1:0] node788;
	wire [8-1:0] node790;
	wire [8-1:0] node791;
	wire [8-1:0] node792;
	wire [8-1:0] node794;
	wire [8-1:0] node797;
	wire [8-1:0] node800;
	wire [8-1:0] node801;
	wire [8-1:0] node804;
	wire [8-1:0] node807;
	wire [8-1:0] node808;
	wire [8-1:0] node809;
	wire [8-1:0] node810;
	wire [8-1:0] node811;
	wire [8-1:0] node814;
	wire [8-1:0] node816;
	wire [8-1:0] node819;
	wire [8-1:0] node821;
	wire [8-1:0] node822;
	wire [8-1:0] node826;
	wire [8-1:0] node827;
	wire [8-1:0] node828;
	wire [8-1:0] node829;
	wire [8-1:0] node833;
	wire [8-1:0] node836;
	wire [8-1:0] node837;
	wire [8-1:0] node839;
	wire [8-1:0] node840;
	wire [8-1:0] node844;
	wire [8-1:0] node847;
	wire [8-1:0] node848;
	wire [8-1:0] node849;
	wire [8-1:0] node852;
	wire [8-1:0] node853;
	wire [8-1:0] node855;
	wire [8-1:0] node858;
	wire [8-1:0] node861;
	wire [8-1:0] node862;
	wire [8-1:0] node863;
	wire [8-1:0] node867;
	wire [8-1:0] node868;
	wire [8-1:0] node869;
	wire [8-1:0] node871;
	wire [8-1:0] node874;
	wire [8-1:0] node877;
	wire [8-1:0] node878;
	wire [8-1:0] node882;
	wire [8-1:0] node883;
	wire [8-1:0] node884;
	wire [8-1:0] node885;
	wire [8-1:0] node886;
	wire [8-1:0] node887;
	wire [8-1:0] node888;
	wire [8-1:0] node893;
	wire [8-1:0] node894;
	wire [8-1:0] node895;
	wire [8-1:0] node897;
	wire [8-1:0] node900;
	wire [8-1:0] node903;
	wire [8-1:0] node906;
	wire [8-1:0] node907;
	wire [8-1:0] node909;
	wire [8-1:0] node910;
	wire [8-1:0] node913;
	wire [8-1:0] node915;
	wire [8-1:0] node918;
	wire [8-1:0] node919;
	wire [8-1:0] node922;
	wire [8-1:0] node925;
	wire [8-1:0] node926;
	wire [8-1:0] node927;
	wire [8-1:0] node928;
	wire [8-1:0] node929;
	wire [8-1:0] node932;
	wire [8-1:0] node934;
	wire [8-1:0] node937;
	wire [8-1:0] node940;
	wire [8-1:0] node941;
	wire [8-1:0] node944;
	wire [8-1:0] node947;
	wire [8-1:0] node948;
	wire [8-1:0] node950;
	wire [8-1:0] node953;
	wire [8-1:0] node954;
	wire [8-1:0] node957;
	wire [8-1:0] node960;
	wire [8-1:0] node961;
	wire [8-1:0] node962;
	wire [8-1:0] node963;
	wire [8-1:0] node966;
	wire [8-1:0] node967;
	wire [8-1:0] node970;
	wire [8-1:0] node971;
	wire [8-1:0] node975;
	wire [8-1:0] node976;
	wire [8-1:0] node977;
	wire [8-1:0] node980;
	wire [8-1:0] node981;
	wire [8-1:0] node985;
	wire [8-1:0] node986;
	wire [8-1:0] node989;
	wire [8-1:0] node990;
	wire [8-1:0] node994;
	wire [8-1:0] node995;
	wire [8-1:0] node996;
	wire [8-1:0] node999;
	wire [8-1:0] node1002;
	wire [8-1:0] node1003;
	wire [8-1:0] node1004;
	wire [8-1:0] node1005;
	wire [8-1:0] node1008;
	wire [8-1:0] node1010;
	wire [8-1:0] node1013;
	wire [8-1:0] node1016;
	wire [8-1:0] node1018;
	wire [8-1:0] node1020;
	wire [8-1:0] node1021;

	assign outp = (inp[13]) ? node530 : node1;
		assign node1 = (inp[4]) ? node263 : node2;
			assign node2 = (inp[7]) ? node108 : node3;
				assign node3 = (inp[11]) ? node53 : node4;
					assign node4 = (inp[5]) ? node38 : node5;
						assign node5 = (inp[1]) ? node21 : node6;
							assign node6 = (inp[2]) ? node12 : node7;
								assign node7 = (inp[3]) ? 8'b01111111 : node8;
									assign node8 = (inp[12]) ? 8'b01111111 : 8'b00111011;
								assign node12 = (inp[8]) ? node16 : node13;
									assign node13 = (inp[0]) ? 8'b01111111 : 8'b00101111;
									assign node16 = (inp[3]) ? node18 : 8'b00111011;
										assign node18 = (inp[10]) ? 8'b00101011 : 8'b00101111;
							assign node21 = (inp[8]) ? node27 : node22;
								assign node22 = (inp[2]) ? 8'b00101110 : node23;
									assign node23 = (inp[6]) ? 8'b01111111 : 8'b00111110;
								assign node27 = (inp[0]) ? node31 : node28;
									assign node28 = (inp[2]) ? 8'b00101010 : 8'b00111010;
									assign node31 = (inp[12]) ? node35 : node32;
										assign node32 = (inp[3]) ? 8'b00111010 : 8'b00111011;
										assign node35 = (inp[6]) ? 8'b00111110 : 8'b01111111;
						assign node38 = (inp[0]) ? 8'b01111111 : node39;
							assign node39 = (inp[1]) ? node45 : node40;
								assign node40 = (inp[10]) ? 8'b01111111 : node41;
									assign node41 = (inp[3]) ? 8'b01111111 : 8'b00111011;
								assign node45 = (inp[8]) ? node49 : node46;
									assign node46 = (inp[3]) ? 8'b01111111 : 8'b00111110;
									assign node49 = (inp[2]) ? 8'b00101111 : 8'b00111011;
					assign node53 = (inp[8]) ? node81 : node54;
						assign node54 = (inp[12]) ? node68 : node55;
							assign node55 = (inp[2]) ? node61 : node56;
								assign node56 = (inp[1]) ? node58 : 8'b00101111;
									assign node58 = (inp[0]) ? 8'b00101011 : 8'b00101110;
								assign node61 = (inp[10]) ? node65 : node62;
									assign node62 = (inp[0]) ? 8'b00101010 : 8'b00111011;
									assign node65 = (inp[0]) ? 8'b00101110 : 8'b00111110;
							assign node68 = (inp[0]) ? node72 : node69;
								assign node69 = (inp[10]) ? 8'b00101110 : 8'b01111111;
								assign node72 = (inp[1]) ? node74 : 8'b00111110;
									assign node74 = (inp[3]) ? node78 : node75;
										assign node75 = (inp[6]) ? 8'b00101011 : 8'b00111011;
										assign node78 = (inp[6]) ? 8'b00111010 : 8'b00111110;
						assign node81 = (inp[2]) ? node93 : node82;
							assign node82 = (inp[12]) ? node90 : node83;
								assign node83 = (inp[9]) ? node87 : node84;
									assign node84 = (inp[1]) ? 8'b00001011 : 8'b00101011;
									assign node87 = (inp[3]) ? 8'b00001111 : 8'b00001011;
								assign node90 = (inp[5]) ? 8'b00111011 : 8'b00011011;
							assign node93 = (inp[5]) ? node99 : node94;
								assign node94 = (inp[12]) ? node96 : 8'b00011111;
									assign node96 = (inp[10]) ? 8'b00101010 : 8'b00101011;
								assign node99 = (inp[0]) ? node103 : node100;
									assign node100 = (inp[10]) ? 8'b00011110 : 8'b00111010;
									assign node103 = (inp[3]) ? node105 : 8'b00001010;
										assign node105 = (inp[12]) ? 8'b00011110 : 8'b00001110;
				assign node108 = (inp[9]) ? node188 : node109;
					assign node109 = (inp[11]) ? node147 : node110;
						assign node110 = (inp[5]) ? node128 : node111;
							assign node111 = (inp[6]) ? node119 : node112;
								assign node112 = (inp[3]) ? node116 : node113;
									assign node113 = (inp[8]) ? 8'b01111111 : 8'b00101011;
									assign node116 = (inp[0]) ? 8'b00111110 : 8'b00111010;
								assign node119 = (inp[0]) ? node121 : 8'b00101010;
									assign node121 = (inp[10]) ? node125 : node122;
										assign node122 = (inp[12]) ? 8'b00101110 : 8'b00101111;
										assign node125 = (inp[3]) ? 8'b00101010 : 8'b00101011;
							assign node128 = (inp[6]) ? node138 : node129;
								assign node129 = (inp[2]) ? node131 : 8'b01111111;
									assign node131 = (inp[12]) ? node135 : node132;
										assign node132 = (inp[1]) ? 8'b00101111 : 8'b00101011;
										assign node135 = (inp[8]) ? 8'b00101110 : 8'b00101010;
								assign node138 = (inp[2]) ? node140 : 8'b00101110;
									assign node140 = (inp[3]) ? node144 : node141;
										assign node141 = (inp[0]) ? 8'b01111111 : 8'b00111110;
										assign node144 = (inp[1]) ? 8'b01111111 : 8'b00111010;
						assign node147 = (inp[2]) ? node173 : node148;
							assign node148 = (inp[3]) ? node158 : node149;
								assign node149 = (inp[10]) ? node155 : node150;
									assign node150 = (inp[8]) ? node152 : 8'b00111110;
										assign node152 = (inp[1]) ? 8'b00101010 : 8'b00101011;
									assign node155 = (inp[0]) ? 8'b00001111 : 8'b00001110;
								assign node158 = (inp[12]) ? node164 : node159;
									assign node159 = (inp[8]) ? node161 : 8'b00111010;
										assign node161 = (inp[0]) ? 8'b00011011 : 8'b00011010;
									assign node164 = (inp[6]) ? node170 : node165;
										assign node165 = (inp[0]) ? node167 : 8'b00111010;
											assign node167 = (inp[10]) ? 8'b00111010 : 8'b00111110;
										assign node170 = (inp[8]) ? 8'b00101010 : 8'b00101110;
							assign node173 = (inp[10]) ? node181 : node174;
								assign node174 = (inp[8]) ? node178 : node175;
									assign node175 = (inp[1]) ? 8'b00111010 : 8'b00101011;
									assign node178 = (inp[6]) ? 8'b00001111 : 8'b00011011;
								assign node181 = (inp[3]) ? node185 : node182;
									assign node182 = (inp[1]) ? 8'b00011111 : 8'b00111010;
									assign node185 = (inp[12]) ? 8'b00011111 : 8'b00011110;
					assign node188 = (inp[1]) ? node230 : node189;
						assign node189 = (inp[3]) ? node209 : node190;
							assign node190 = (inp[11]) ? node200 : node191;
								assign node191 = (inp[0]) ? node197 : node192;
									assign node192 = (inp[8]) ? 8'b00001011 : node193;
										assign node193 = (inp[10]) ? 8'b00001011 : 8'b00001111;
									assign node197 = (inp[8]) ? 8'b10011101 : 8'b00011111;
								assign node200 = (inp[8]) ? node202 : 8'b00011010;
									assign node202 = (inp[12]) ? node204 : 8'b00001010;
										assign node204 = (inp[0]) ? 8'b00001011 : node205;
											assign node205 = (inp[2]) ? 8'b00001011 : 8'b00011011;
							assign node209 = (inp[8]) ? node221 : node210;
								assign node210 = (inp[11]) ? node216 : node211;
									assign node211 = (inp[10]) ? node213 : 8'b00001110;
										assign node213 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node216 = (inp[6]) ? 8'b00011011 : node217;
										assign node217 = (inp[2]) ? 8'b00001110 : 8'b00011010;
								assign node221 = (inp[11]) ? node227 : node222;
									assign node222 = (inp[2]) ? 8'b10010100 : node223;
										assign node223 = (inp[6]) ? 8'b00000010 : 8'b00011010;
									assign node227 = (inp[12]) ? 8'b10100100 : 8'b11110111;
						assign node230 = (inp[10]) ? node246 : node231;
							assign node231 = (inp[8]) ? node241 : node232;
								assign node232 = (inp[11]) ? 8'b00001010 : node233;
									assign node233 = (inp[6]) ? node235 : 8'b00011111;
										assign node235 = (inp[5]) ? 8'b00001111 : node236;
											assign node236 = (inp[12]) ? 8'b00001111 : 8'b00001110;
								assign node241 = (inp[3]) ? node243 : 8'b10011101;
									assign node243 = (inp[5]) ? 8'b10100000 : 8'b10100100;
							assign node246 = (inp[0]) ? node256 : node247;
								assign node247 = (inp[5]) ? node251 : node248;
									assign node248 = (inp[3]) ? 8'b00000010 : 8'b10000010;
									assign node251 = (inp[8]) ? node253 : 8'b00000010;
										assign node253 = (inp[3]) ? 8'b10010101 : 8'b10000100;
								assign node256 = (inp[11]) ? node260 : node257;
									assign node257 = (inp[3]) ? 8'b00011010 : 8'b10010001;
									assign node260 = (inp[8]) ? 8'b10110100 : 8'b10100101;
			assign node263 = (inp[7]) ? node421 : node264;
				assign node264 = (inp[9]) ? node344 : node265;
					assign node265 = (inp[8]) ? node295 : node266;
						assign node266 = (inp[10]) ? node280 : node267;
							assign node267 = (inp[0]) ? 8'b11110101 : node268;
								assign node268 = (inp[12]) ? node276 : node269;
									assign node269 = (inp[11]) ? 8'b11110111 : node270;
										assign node270 = (inp[5]) ? 8'b10000001 : node271;
											assign node271 = (inp[3]) ? 8'b00001011 : 8'b10000010;
									assign node276 = (inp[1]) ? 8'b00000010 : 8'b00011010;
							assign node280 = (inp[6]) ? node288 : node281;
								assign node281 = (inp[0]) ? node285 : node282;
									assign node282 = (inp[3]) ? 8'b00001111 : 8'b00001110;
									assign node285 = (inp[3]) ? 8'b00011110 : 8'b00001010;
								assign node288 = (inp[11]) ? 8'b00011110 : node289;
									assign node289 = (inp[2]) ? node291 : 8'b00011110;
										assign node291 = (inp[5]) ? 8'b00011111 : 8'b00001111;
						assign node295 = (inp[5]) ? node309 : node296;
							assign node296 = (inp[10]) ? node304 : node297;
								assign node297 = (inp[0]) ? 8'b10011101 : node298;
									assign node298 = (inp[3]) ? 8'b00001011 : node299;
										assign node299 = (inp[11]) ? 8'b00001010 : 8'b10000010;
								assign node304 = (inp[12]) ? node306 : 8'b11110111;
									assign node306 = (inp[3]) ? 8'b00001011 : 8'b10000001;
							assign node309 = (inp[3]) ? node327 : node310;
								assign node310 = (inp[10]) ? node320 : node311;
									assign node311 = (inp[0]) ? node315 : node312;
										assign node312 = (inp[6]) ? 8'b00011010 : 8'b00000010;
										assign node315 = (inp[11]) ? 8'b10100001 : node316;
											assign node316 = (inp[1]) ? 8'b10010101 : 8'b10010100;
									assign node320 = (inp[6]) ? node324 : node321;
										assign node321 = (inp[12]) ? 8'b10100100 : 8'b10000100;
										assign node324 = (inp[11]) ? 8'b10111100 : 8'b10010100;
								assign node327 = (inp[11]) ? node335 : node328;
									assign node328 = (inp[6]) ? 8'b10011101 : node329;
										assign node329 = (inp[1]) ? node331 : 8'b10001101;
											assign node331 = (inp[2]) ? 8'b10010101 : 8'b10000101;
									assign node335 = (inp[12]) ? node339 : node336;
										assign node336 = (inp[0]) ? 8'b10111100 : 8'b10110100;
										assign node339 = (inp[0]) ? node341 : 8'b11111101;
											assign node341 = (inp[6]) ? 8'b10111001 : 8'b10101101;
					assign node344 = (inp[11]) ? node382 : node345;
						assign node345 = (inp[5]) ? node363 : node346;
							assign node346 = (inp[0]) ? node352 : node347;
								assign node347 = (inp[10]) ? 8'b00101110 : node348;
									assign node348 = (inp[6]) ? 8'b00111010 : 8'b00101010;
								assign node352 = (inp[3]) ? node358 : node353;
									assign node353 = (inp[6]) ? node355 : 8'b00111010;
										assign node355 = (inp[10]) ? 8'b00111010 : 8'b00111110;
									assign node358 = (inp[1]) ? node360 : 8'b00101111;
										assign node360 = (inp[12]) ? 8'b00111110 : 8'b00111010;
							assign node363 = (inp[1]) ? node371 : node364;
								assign node364 = (inp[3]) ? node368 : node365;
									assign node365 = (inp[2]) ? 8'b00111110 : 8'b00111010;
									assign node368 = (inp[8]) ? 8'b01111111 : 8'b00111011;
								assign node371 = (inp[0]) ? node375 : node372;
									assign node372 = (inp[6]) ? 8'b00111110 : 8'b00101111;
									assign node375 = (inp[8]) ? 8'b01111111 : node376;
										assign node376 = (inp[6]) ? 8'b01111111 : node377;
											assign node377 = (inp[10]) ? 8'b00101111 : 8'b00111011;
						assign node382 = (inp[8]) ? node402 : node383;
							assign node383 = (inp[1]) ? node397 : node384;
								assign node384 = (inp[0]) ? node390 : node385;
									assign node385 = (inp[6]) ? 8'b00111011 : node386;
										assign node386 = (inp[12]) ? 8'b00101110 : 8'b00111011;
									assign node390 = (inp[6]) ? 8'b00101010 : node391;
										assign node391 = (inp[10]) ? node393 : 8'b00101011;
											assign node393 = (inp[2]) ? 8'b00101011 : 8'b00101111;
								assign node397 = (inp[2]) ? 8'b00011111 : node398;
									assign node398 = (inp[5]) ? 8'b00111010 : 8'b00101010;
							assign node402 = (inp[5]) ? node408 : node403;
								assign node403 = (inp[0]) ? node405 : 8'b00101010;
									assign node405 = (inp[3]) ? 8'b00111010 : 8'b00001011;
								assign node408 = (inp[10]) ? node412 : node409;
									assign node409 = (inp[3]) ? 8'b00011010 : 8'b00101010;
									assign node412 = (inp[3]) ? node416 : node413;
										assign node413 = (inp[6]) ? 8'b00011110 : 8'b00011011;
										assign node416 = (inp[0]) ? 8'b00001110 : node417;
											assign node417 = (inp[6]) ? 8'b00001111 : 8'b00001011;
				assign node421 = (inp[12]) ? node483 : node422;
					assign node422 = (inp[11]) ? node452 : node423;
						assign node423 = (inp[0]) ? node429 : node424;
							assign node424 = (inp[5]) ? node426 : 8'b10000010;
								assign node426 = (inp[1]) ? 8'b10000010 : 8'b10010000;
							assign node429 = (inp[2]) ? node441 : node430;
								assign node430 = (inp[10]) ? node432 : 8'b10000010;
									assign node432 = (inp[6]) ? node438 : node433;
										assign node433 = (inp[8]) ? node435 : 8'b10000001;
											assign node435 = (inp[3]) ? 8'b10000101 : 8'b10000001;
										assign node438 = (inp[3]) ? 8'b10000010 : 8'b10000001;
								assign node441 = (inp[6]) ? node449 : node442;
									assign node442 = (inp[10]) ? node446 : node443;
										assign node443 = (inp[9]) ? 8'b10010101 : 8'b10010100;
										assign node446 = (inp[3]) ? 8'b10010000 : 8'b10010001;
									assign node449 = (inp[5]) ? 8'b10010101 : 8'b10000010;
						assign node452 = (inp[0]) ? node464 : node453;
							assign node453 = (inp[3]) ? node455 : 8'b11110111;
								assign node455 = (inp[1]) ? node457 : 8'b11110111;
									assign node457 = (inp[5]) ? node459 : 8'b11110111;
										assign node459 = (inp[2]) ? node461 : 8'b10110000;
											assign node461 = (inp[6]) ? 8'b10100100 : 8'b10110100;
							assign node464 = (inp[1]) ? node474 : node465;
								assign node465 = (inp[5]) ? node467 : 8'b11110111;
									assign node467 = (inp[8]) ? node471 : node468;
										assign node468 = (inp[3]) ? 8'b10100101 : 8'b11110111;
										assign node471 = (inp[2]) ? 8'b10100001 : 8'b10110001;
								assign node474 = (inp[8]) ? node478 : node475;
									assign node475 = (inp[9]) ? 8'b10110100 : 8'b10100100;
									assign node478 = (inp[10]) ? node480 : 8'b10100000;
										assign node480 = (inp[6]) ? 8'b10100000 : 8'b10100101;
					assign node483 = (inp[5]) ? node503 : node484;
						assign node484 = (inp[0]) ? node486 : 8'b00000010;
							assign node486 = (inp[10]) ? node496 : node487;
								assign node487 = (inp[1]) ? node491 : node488;
									assign node488 = (inp[8]) ? 8'b10100100 : 8'b00000010;
									assign node491 = (inp[11]) ? 8'b10100101 : node492;
										assign node492 = (inp[9]) ? 8'b10000001 : 8'b10000101;
								assign node496 = (inp[2]) ? 8'b10010001 : node497;
									assign node497 = (inp[1]) ? node499 : 8'b00000010;
										assign node499 = (inp[11]) ? 8'b00000010 : 8'b10000001;
						assign node503 = (inp[2]) ? node517 : node504;
							assign node504 = (inp[1]) ? node506 : 8'b00000010;
								assign node506 = (inp[10]) ? node510 : node507;
									assign node507 = (inp[11]) ? 8'b00000010 : 8'b10000101;
									assign node510 = (inp[11]) ? node514 : node511;
										assign node511 = (inp[8]) ? 8'b10000101 : 8'b10000001;
										assign node514 = (inp[8]) ? 8'b10100001 : 8'b10100101;
							assign node517 = (inp[11]) ? node523 : node518;
								assign node518 = (inp[1]) ? node520 : 8'b10010100;
									assign node520 = (inp[9]) ? 8'b10010000 : 8'b10010001;
								assign node523 = (inp[10]) ? node527 : node524;
									assign node524 = (inp[1]) ? 8'b10110000 : 8'b11110101;
									assign node527 = (inp[8]) ? 8'b10100100 : 8'b10110100;
		assign node530 = (inp[5]) ? node756 : node531;
			assign node531 = (inp[0]) ? node603 : node532;
				assign node532 = (inp[12]) ? node576 : node533;
					assign node533 = (inp[11]) ? node557 : node534;
						assign node534 = (inp[8]) ? node548 : node535;
							assign node535 = (inp[2]) ? node543 : node536;
								assign node536 = (inp[4]) ? 8'b00011010 : node537;
									assign node537 = (inp[10]) ? 8'b00011010 : node538;
										assign node538 = (inp[1]) ? 8'b00011110 : 8'b00011111;
								assign node543 = (inp[3]) ? node545 : 8'b10000010;
									assign node545 = (inp[10]) ? 8'b00001111 : 8'b00001110;
							assign node548 = (inp[1]) ? 8'b10000010 : node549;
								assign node549 = (inp[10]) ? node553 : node550;
									assign node550 = (inp[4]) ? 8'b10000010 : 8'b00001011;
									assign node553 = (inp[9]) ? 8'b00001011 : 8'b10000010;
						assign node557 = (inp[4]) ? node571 : node558;
							assign node558 = (inp[8]) ? node566 : node559;
								assign node559 = (inp[1]) ? 8'b00011011 : node560;
									assign node560 = (inp[2]) ? 8'b00011110 : node561;
										assign node561 = (inp[3]) ? 8'b00001111 : 8'b00001011;
								assign node566 = (inp[2]) ? 8'b11110111 : node567;
									assign node567 = (inp[6]) ? 8'b00001011 : 8'b00001010;
							assign node571 = (inp[7]) ? 8'b11110111 : node572;
								assign node572 = (inp[6]) ? 8'b00001010 : 8'b11110111;
					assign node576 = (inp[2]) ? node592 : node577;
						assign node577 = (inp[4]) ? node589 : node578;
							assign node578 = (inp[8]) ? 8'b00011010 : node579;
								assign node579 = (inp[10]) ? node581 : 8'b00011110;
									assign node581 = (inp[9]) ? node585 : node582;
										assign node582 = (inp[3]) ? 8'b00011111 : 8'b00011110;
										assign node585 = (inp[1]) ? 8'b00000010 : 8'b00001011;
							assign node589 = (inp[7]) ? 8'b00000010 : 8'b00011010;
						assign node592 = (inp[8]) ? 8'b00000010 : node593;
							assign node593 = (inp[4]) ? node597 : node594;
								assign node594 = (inp[1]) ? 8'b00001110 : 8'b00001111;
								assign node597 = (inp[7]) ? 8'b00000010 : node598;
									assign node598 = (inp[10]) ? 8'b00001110 : 8'b00000010;
				assign node603 = (inp[9]) ? node687 : node604;
					assign node604 = (inp[4]) ? node638 : node605;
						assign node605 = (inp[10]) ? node623 : node606;
							assign node606 = (inp[11]) ? node612 : node607;
								assign node607 = (inp[2]) ? node609 : 8'b11111101;
									assign node609 = (inp[6]) ? 8'b10101100 : 8'b11111101;
								assign node612 = (inp[12]) ? node618 : node613;
									assign node613 = (inp[7]) ? node615 : 8'b10001001;
										assign node615 = (inp[6]) ? 8'b10111001 : 8'b10101000;
									assign node618 = (inp[6]) ? node620 : 8'b10111100;
										assign node620 = (inp[7]) ? 8'b10101100 : 8'b10101101;
							assign node623 = (inp[8]) ? node629 : node624;
								assign node624 = (inp[7]) ? node626 : 8'b10101100;
									assign node626 = (inp[6]) ? 8'b10100000 : 8'b10110001;
								assign node629 = (inp[7]) ? 8'b10101001 : node630;
									assign node630 = (inp[2]) ? node634 : node631;
										assign node631 = (inp[1]) ? 8'b10111001 : 8'b10101001;
										assign node634 = (inp[12]) ? 8'b10111000 : 8'b10111001;
						assign node638 = (inp[11]) ? node662 : node639;
							assign node639 = (inp[8]) ? node651 : node640;
								assign node640 = (inp[1]) ? 8'b10110001 : node641;
									assign node641 = (inp[10]) ? node647 : node642;
										assign node642 = (inp[6]) ? 8'b10100000 : node643;
											assign node643 = (inp[2]) ? 8'b10110000 : 8'b10100000;
										assign node647 = (inp[7]) ? 8'b10100000 : 8'b10111100;
								assign node651 = (inp[10]) ? node659 : node652;
									assign node652 = (inp[6]) ? 8'b10100100 : node653;
										assign node653 = (inp[2]) ? node655 : 8'b10100100;
											assign node655 = (inp[3]) ? 8'b10110100 : 8'b11110101;
									assign node659 = (inp[1]) ? 8'b10100001 : 8'b10100000;
							assign node662 = (inp[7]) ? node680 : node663;
								assign node663 = (inp[6]) ? node675 : node664;
									assign node664 = (inp[3]) ? 8'b10111000 : node665;
										assign node665 = (inp[1]) ? node671 : node666;
											assign node666 = (inp[10]) ? node668 : 8'b10010101;
												assign node668 = (inp[8]) ? 8'b10000101 : 8'b10101001;
											assign node671 = (inp[12]) ? 8'b10010100 : 8'b10000000;
									assign node675 = (inp[12]) ? 8'b10101001 : node676;
										assign node676 = (inp[1]) ? 8'b10001101 : 8'b10001100;
								assign node680 = (inp[10]) ? 8'b10100000 : node681;
									assign node681 = (inp[12]) ? 8'b10000100 : node682;
										assign node682 = (inp[8]) ? 8'b10010000 : 8'b10010100;
					assign node687 = (inp[4]) ? node719 : node688;
						assign node688 = (inp[8]) ? node706 : node689;
							assign node689 = (inp[7]) ? node699 : node690;
								assign node690 = (inp[3]) ? 8'b00011110 : node691;
									assign node691 = (inp[2]) ? 8'b00001010 : node692;
										assign node692 = (inp[1]) ? node694 : 8'b00001111;
											assign node694 = (inp[11]) ? 8'b00011011 : 8'b00011111;
								assign node699 = (inp[2]) ? node703 : node700;
									assign node700 = (inp[12]) ? 8'b10100101 : 8'b10000010;
									assign node703 = (inp[1]) ? 8'b00011011 : 8'b00001011;
							assign node706 = (inp[2]) ? node712 : node707;
								assign node707 = (inp[1]) ? 8'b10101001 : node708;
									assign node708 = (inp[12]) ? 8'b00011011 : 8'b00001010;
								assign node712 = (inp[10]) ? node716 : node713;
									assign node713 = (inp[11]) ? 8'b10100001 : 8'b10001101;
									assign node716 = (inp[11]) ? 8'b10110100 : 8'b10010000;
						assign node719 = (inp[10]) ? node735 : node720;
							assign node720 = (inp[11]) ? node728 : node721;
								assign node721 = (inp[8]) ? node725 : node722;
									assign node722 = (inp[3]) ? 8'b10010000 : 8'b10000001;
									assign node725 = (inp[6]) ? 8'b10000100 : 8'b10001101;
								assign node728 = (inp[6]) ? 8'b11110111 : node729;
									assign node729 = (inp[7]) ? 8'b10100101 : node730;
										assign node730 = (inp[1]) ? 8'b10110001 : 8'b11110101;
							assign node735 = (inp[1]) ? node749 : node736;
								assign node736 = (inp[11]) ? node742 : node737;
									assign node737 = (inp[2]) ? node739 : 8'b00000010;
										assign node739 = (inp[3]) ? 8'b10000010 : 8'b10010000;
									assign node742 = (inp[3]) ? node744 : 8'b00000010;
										assign node744 = (inp[7]) ? 8'b11110101 : node745;
											assign node745 = (inp[6]) ? 8'b00011111 : 8'b00011110;
								assign node749 = (inp[3]) ? 8'b00000010 : node750;
									assign node750 = (inp[11]) ? 8'b10110100 : node751;
										assign node751 = (inp[6]) ? 8'b10000001 : 8'b10010001;
			assign node756 = (inp[4]) ? node882 : node757;
				assign node757 = (inp[11]) ? node807 : node758;
					assign node758 = (inp[0]) ? node788 : node759;
						assign node759 = (inp[9]) ? node773 : node760;
							assign node760 = (inp[7]) ? node764 : node761;
								assign node761 = (inp[10]) ? 8'b10011101 : 8'b00011110;
								assign node764 = (inp[1]) ? node768 : node765;
									assign node765 = (inp[12]) ? 8'b00000010 : 8'b10010000;
									assign node768 = (inp[6]) ? 8'b00001111 : node769;
										assign node769 = (inp[2]) ? 8'b10000001 : 8'b10011001;
							assign node773 = (inp[7]) ? node781 : node774;
								assign node774 = (inp[8]) ? node776 : 8'b11111101;
									assign node776 = (inp[10]) ? 8'b11111101 : node777;
										assign node777 = (inp[2]) ? 8'b10101001 : 8'b10111001;
								assign node781 = (inp[6]) ? node785 : node782;
									assign node782 = (inp[1]) ? 8'b10100001 : 8'b10100000;
									assign node785 = (inp[12]) ? 8'b10101101 : 8'b10111001;
						assign node788 = (inp[7]) ? node790 : 8'b11111101;
							assign node790 = (inp[1]) ? node800 : node791;
								assign node791 = (inp[3]) ? node797 : node792;
									assign node792 = (inp[6]) ? node794 : 8'b11111101;
										assign node794 = (inp[8]) ? 8'b11111101 : 8'b10101101;
									assign node797 = (inp[8]) ? 8'b10110100 : 8'b10111100;
								assign node800 = (inp[6]) ? node804 : node801;
									assign node801 = (inp[9]) ? 8'b11110101 : 8'b10111001;
									assign node804 = (inp[9]) ? 8'b10100001 : 8'b10100101;
					assign node807 = (inp[1]) ? node847 : node808;
						assign node808 = (inp[12]) ? node826 : node809;
							assign node809 = (inp[2]) ? node819 : node810;
								assign node810 = (inp[10]) ? node814 : node811;
									assign node811 = (inp[0]) ? 8'b10001101 : 8'b00001111;
									assign node814 = (inp[8]) ? node816 : 8'b10101101;
										assign node816 = (inp[9]) ? 8'b10001101 : 8'b10101101;
								assign node819 = (inp[7]) ? node821 : 8'b10101100;
									assign node821 = (inp[0]) ? 8'b10000101 : node822;
										assign node822 = (inp[3]) ? 8'b11110111 : 8'b10111100;
							assign node826 = (inp[8]) ? node836 : node827;
								assign node827 = (inp[7]) ? node833 : node828;
									assign node828 = (inp[2]) ? 8'b10111100 : node829;
										assign node829 = (inp[10]) ? 8'b00011111 : 8'b11111101;
									assign node833 = (inp[10]) ? 8'b10111000 : 8'b10101100;
								assign node836 = (inp[7]) ? node844 : node837;
									assign node837 = (inp[2]) ? node839 : 8'b10011101;
										assign node839 = (inp[3]) ? 8'b10011100 : node840;
											assign node840 = (inp[0]) ? 8'b10011100 : 8'b10111100;
									assign node844 = (inp[2]) ? 8'b10010001 : 8'b10011100;
						assign node847 = (inp[8]) ? node861 : node848;
							assign node848 = (inp[0]) ? node852 : node849;
								assign node849 = (inp[9]) ? 8'b10111001 : 8'b00011010;
								assign node852 = (inp[2]) ? node858 : node853;
									assign node853 = (inp[6]) ? node855 : 8'b10111001;
										assign node855 = (inp[7]) ? 8'b10101001 : 8'b10111001;
									assign node858 = (inp[7]) ? 8'b10010100 : 8'b10101000;
							assign node861 = (inp[9]) ? node867 : node862;
								assign node862 = (inp[7]) ? 8'b00001010 : node863;
									assign node863 = (inp[2]) ? 8'b10100001 : 8'b10101101;
								assign node867 = (inp[7]) ? node877 : node868;
									assign node868 = (inp[2]) ? node874 : node869;
										assign node869 = (inp[0]) ? node871 : 8'b10111000;
											assign node871 = (inp[3]) ? 8'b10001001 : 8'b10011001;
										assign node874 = (inp[12]) ? 8'b10010000 : 8'b10010001;
									assign node877 = (inp[3]) ? 8'b10010000 : node878;
										assign node878 = (inp[0]) ? 8'b10000000 : 8'b10000101;
				assign node882 = (inp[7]) ? node960 : node883;
					assign node883 = (inp[3]) ? node925 : node884;
						assign node884 = (inp[11]) ? node906 : node885;
							assign node885 = (inp[6]) ? node893 : node886;
								assign node886 = (inp[1]) ? 8'b11110101 : node887;
									assign node887 = (inp[2]) ? 8'b10110100 : node888;
										assign node888 = (inp[0]) ? 8'b10100000 : 8'b10100100;
								assign node893 = (inp[10]) ? node903 : node894;
									assign node894 = (inp[2]) ? node900 : node895;
										assign node895 = (inp[9]) ? node897 : 8'b10111000;
											assign node897 = (inp[0]) ? 8'b10111100 : 8'b10111000;
										assign node900 = (inp[0]) ? 8'b10110001 : 8'b10110000;
									assign node903 = (inp[12]) ? 8'b10111100 : 8'b00011110;
							assign node906 = (inp[10]) ? node918 : node907;
								assign node907 = (inp[9]) ? node909 : 8'b10010100;
									assign node909 = (inp[1]) ? node913 : node910;
										assign node910 = (inp[12]) ? 8'b10010101 : 8'b10000101;
										assign node913 = (inp[0]) ? node915 : 8'b10100000;
											assign node915 = (inp[8]) ? 8'b10000001 : 8'b10000101;
								assign node918 = (inp[8]) ? node922 : node919;
									assign node919 = (inp[6]) ? 8'b10111000 : 8'b10101001;
									assign node922 = (inp[0]) ? 8'b10010000 : 8'b10000001;
						assign node925 = (inp[8]) ? node947 : node926;
							assign node926 = (inp[9]) ? node940 : node927;
								assign node927 = (inp[0]) ? node937 : node928;
									assign node928 = (inp[6]) ? node932 : node929;
										assign node929 = (inp[2]) ? 8'b00011110 : 8'b00011010;
										assign node932 = (inp[2]) ? node934 : 8'b00001111;
											assign node934 = (inp[12]) ? 8'b00011011 : 8'b00011111;
									assign node937 = (inp[11]) ? 8'b10101001 : 8'b10111001;
								assign node940 = (inp[6]) ? node944 : node941;
									assign node941 = (inp[10]) ? 8'b10101101 : 8'b10110001;
									assign node944 = (inp[10]) ? 8'b11111101 : 8'b10011101;
							assign node947 = (inp[1]) ? node953 : node948;
								assign node948 = (inp[9]) ? node950 : 8'b00001011;
									assign node950 = (inp[11]) ? 8'b10001100 : 8'b10101001;
								assign node953 = (inp[10]) ? node957 : node954;
									assign node954 = (inp[0]) ? 8'b10100101 : 8'b10101101;
									assign node957 = (inp[12]) ? 8'b10100001 : 8'b10001001;
					assign node960 = (inp[11]) ? node994 : node961;
						assign node961 = (inp[8]) ? node975 : node962;
							assign node962 = (inp[1]) ? node966 : node963;
								assign node963 = (inp[2]) ? 8'b10110000 : 8'b10100000;
								assign node966 = (inp[9]) ? node970 : node967;
									assign node967 = (inp[2]) ? 8'b10110001 : 8'b10100001;
									assign node970 = (inp[0]) ? 8'b10100001 : node971;
										assign node971 = (inp[3]) ? 8'b10100001 : 8'b10100000;
							assign node975 = (inp[1]) ? node985 : node976;
								assign node976 = (inp[2]) ? node980 : node977;
									assign node977 = (inp[12]) ? 8'b10100000 : 8'b10100100;
									assign node980 = (inp[0]) ? 8'b10110100 : node981;
										assign node981 = (inp[6]) ? 8'b10010100 : 8'b10000100;
								assign node985 = (inp[2]) ? node989 : node986;
									assign node986 = (inp[0]) ? 8'b10100101 : 8'b10000101;
									assign node989 = (inp[0]) ? 8'b11110101 : node990;
										assign node990 = (inp[6]) ? 8'b10010000 : 8'b10100101;
						assign node994 = (inp[9]) ? node1002 : node995;
							assign node995 = (inp[0]) ? node999 : node996;
								assign node996 = (inp[6]) ? 8'b10100101 : 8'b10110100;
								assign node999 = (inp[1]) ? 8'b10010100 : 8'b10000101;
							assign node1002 = (inp[6]) ? node1016 : node1003;
								assign node1003 = (inp[3]) ? node1013 : node1004;
									assign node1004 = (inp[0]) ? node1008 : node1005;
										assign node1005 = (inp[10]) ? 8'b10010001 : 8'b10010101;
										assign node1008 = (inp[10]) ? node1010 : 8'b10000101;
											assign node1010 = (inp[1]) ? 8'b10010100 : 8'b10010101;
									assign node1013 = (inp[0]) ? 8'b10010000 : 8'b10010100;
								assign node1016 = (inp[0]) ? node1018 : 8'b10100000;
									assign node1018 = (inp[8]) ? node1020 : 8'b10010100;
										assign node1020 = (inp[2]) ? 8'b10000000 : node1021;
											assign node1021 = (inp[1]) ? 8'b10000001 : 8'b10010001;

endmodule