module dtc_split5_bm30 (
	input  wire [14-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node7;
	wire [8-1:0] node9;
	wire [8-1:0] node11;
	wire [8-1:0] node14;
	wire [8-1:0] node15;
	wire [8-1:0] node17;
	wire [8-1:0] node20;
	wire [8-1:0] node22;
	wire [8-1:0] node23;
	wire [8-1:0] node26;
	wire [8-1:0] node29;
	wire [8-1:0] node30;
	wire [8-1:0] node31;
	wire [8-1:0] node33;
	wire [8-1:0] node36;
	wire [8-1:0] node38;
	wire [8-1:0] node39;
	wire [8-1:0] node42;
	wire [8-1:0] node45;
	wire [8-1:0] node46;
	wire [8-1:0] node49;
	wire [8-1:0] node50;
	wire [8-1:0] node51;
	wire [8-1:0] node52;
	wire [8-1:0] node56;
	wire [8-1:0] node57;
	wire [8-1:0] node61;
	wire [8-1:0] node62;
	wire [8-1:0] node64;
	wire [8-1:0] node67;
	wire [8-1:0] node68;
	wire [8-1:0] node72;
	wire [8-1:0] node73;
	wire [8-1:0] node74;
	wire [8-1:0] node75;
	wire [8-1:0] node77;
	wire [8-1:0] node80;
	wire [8-1:0] node81;
	wire [8-1:0] node83;
	wire [8-1:0] node86;
	wire [8-1:0] node88;
	wire [8-1:0] node91;
	wire [8-1:0] node92;
	wire [8-1:0] node93;
	wire [8-1:0] node95;
	wire [8-1:0] node98;
	wire [8-1:0] node100;
	wire [8-1:0] node102;
	wire [8-1:0] node105;
	wire [8-1:0] node106;
	wire [8-1:0] node108;
	wire [8-1:0] node111;
	wire [8-1:0] node112;
	wire [8-1:0] node114;
	wire [8-1:0] node117;
	wire [8-1:0] node119;
	wire [8-1:0] node121;
	wire [8-1:0] node125;
	wire [8-1:0] node126;
	wire [8-1:0] node127;
	wire [8-1:0] node128;
	wire [8-1:0] node131;
	wire [8-1:0] node132;
	wire [8-1:0] node133;
	wire [8-1:0] node134;
	wire [8-1:0] node138;
	wire [8-1:0] node139;
	wire [8-1:0] node143;
	wire [8-1:0] node144;
	wire [8-1:0] node146;
	wire [8-1:0] node149;
	wire [8-1:0] node150;
	wire [8-1:0] node154;
	wire [8-1:0] node155;
	wire [8-1:0] node156;
	wire [8-1:0] node157;
	wire [8-1:0] node158;
	wire [8-1:0] node162;
	wire [8-1:0] node163;
	wire [8-1:0] node167;
	wire [8-1:0] node168;
	wire [8-1:0] node170;
	wire [8-1:0] node171;
	wire [8-1:0] node174;
	wire [8-1:0] node177;
	wire [8-1:0] node178;
	wire [8-1:0] node179;
	wire [8-1:0] node182;
	wire [8-1:0] node186;
	wire [8-1:0] node187;
	wire [8-1:0] node188;
	wire [8-1:0] node190;
	wire [8-1:0] node192;
	wire [8-1:0] node195;
	wire [8-1:0] node197;
	wire [8-1:0] node198;
	wire [8-1:0] node201;
	wire [8-1:0] node204;
	wire [8-1:0] node205;
	wire [8-1:0] node206;
	wire [8-1:0] node210;
	wire [8-1:0] node211;
	wire [8-1:0] node215;
	wire [8-1:0] node216;
	wire [8-1:0] node217;
	wire [8-1:0] node218;
	wire [8-1:0] node219;
	wire [8-1:0] node222;
	wire [8-1:0] node225;
	wire [8-1:0] node226;
	wire [8-1:0] node229;
	wire [8-1:0] node232;
	wire [8-1:0] node233;
	wire [8-1:0] node234;
	wire [8-1:0] node235;
	wire [8-1:0] node238;
	wire [8-1:0] node239;
	wire [8-1:0] node242;
	wire [8-1:0] node245;
	wire [8-1:0] node246;
	wire [8-1:0] node247;
	wire [8-1:0] node250;
	wire [8-1:0] node251;
	wire [8-1:0] node254;
	wire [8-1:0] node257;
	wire [8-1:0] node258;
	wire [8-1:0] node261;
	wire [8-1:0] node262;
	wire [8-1:0] node266;
	wire [8-1:0] node267;
	wire [8-1:0] node268;
	wire [8-1:0] node271;
	wire [8-1:0] node273;
	wire [8-1:0] node275;
	wire [8-1:0] node278;
	wire [8-1:0] node279;
	wire [8-1:0] node280;
	wire [8-1:0] node283;
	wire [8-1:0] node284;
	wire [8-1:0] node288;
	wire [8-1:0] node289;
	wire [8-1:0] node293;
	wire [8-1:0] node294;
	wire [8-1:0] node295;
	wire [8-1:0] node296;
	wire [8-1:0] node297;
	wire [8-1:0] node301;
	wire [8-1:0] node302;
	wire [8-1:0] node303;
	wire [8-1:0] node306;
	wire [8-1:0] node310;
	wire [8-1:0] node311;
	wire [8-1:0] node312;
	wire [8-1:0] node313;
	wire [8-1:0] node317;
	wire [8-1:0] node318;
	wire [8-1:0] node322;
	wire [8-1:0] node323;
	wire [8-1:0] node324;
	wire [8-1:0] node327;
	wire [8-1:0] node330;
	wire [8-1:0] node331;
	wire [8-1:0] node333;
	wire [8-1:0] node337;
	wire [8-1:0] node338;
	wire [8-1:0] node339;
	wire [8-1:0] node340;
	wire [8-1:0] node344;
	wire [8-1:0] node345;
	wire [8-1:0] node346;
	wire [8-1:0] node349;
	wire [8-1:0] node353;
	wire [8-1:0] node354;
	wire [8-1:0] node355;
	wire [8-1:0] node356;
	wire [8-1:0] node359;
	wire [8-1:0] node362;
	wire [8-1:0] node363;
	wire [8-1:0] node366;
	wire [8-1:0] node369;
	wire [8-1:0] node372;
	wire [8-1:0] node373;
	wire [8-1:0] node374;
	wire [8-1:0] node375;
	wire [8-1:0] node376;
	wire [8-1:0] node377;
	wire [8-1:0] node378;
	wire [8-1:0] node379;
	wire [8-1:0] node382;
	wire [8-1:0] node383;
	wire [8-1:0] node387;
	wire [8-1:0] node388;
	wire [8-1:0] node389;
	wire [8-1:0] node390;
	wire [8-1:0] node394;
	wire [8-1:0] node397;
	wire [8-1:0] node398;
	wire [8-1:0] node400;
	wire [8-1:0] node404;
	wire [8-1:0] node405;
	wire [8-1:0] node406;
	wire [8-1:0] node407;
	wire [8-1:0] node410;
	wire [8-1:0] node412;
	wire [8-1:0] node415;
	wire [8-1:0] node416;
	wire [8-1:0] node420;
	wire [8-1:0] node421;
	wire [8-1:0] node422;
	wire [8-1:0] node425;
	wire [8-1:0] node427;
	wire [8-1:0] node430;
	wire [8-1:0] node431;
	wire [8-1:0] node434;
	wire [8-1:0] node436;
	wire [8-1:0] node439;
	wire [8-1:0] node440;
	wire [8-1:0] node442;
	wire [8-1:0] node444;
	wire [8-1:0] node447;
	wire [8-1:0] node448;
	wire [8-1:0] node451;
	wire [8-1:0] node452;
	wire [8-1:0] node454;
	wire [8-1:0] node457;
	wire [8-1:0] node458;
	wire [8-1:0] node462;
	wire [8-1:0] node463;
	wire [8-1:0] node464;
	wire [8-1:0] node465;
	wire [8-1:0] node466;
	wire [8-1:0] node468;
	wire [8-1:0] node472;
	wire [8-1:0] node473;
	wire [8-1:0] node474;
	wire [8-1:0] node478;
	wire [8-1:0] node481;
	wire [8-1:0] node482;
	wire [8-1:0] node484;
	wire [8-1:0] node488;
	wire [8-1:0] node489;
	wire [8-1:0] node490;
	wire [8-1:0] node491;
	wire [8-1:0] node492;
	wire [8-1:0] node493;
	wire [8-1:0] node496;
	wire [8-1:0] node499;
	wire [8-1:0] node500;
	wire [8-1:0] node504;
	wire [8-1:0] node505;
	wire [8-1:0] node506;
	wire [8-1:0] node510;
	wire [8-1:0] node513;
	wire [8-1:0] node514;
	wire [8-1:0] node516;
	wire [8-1:0] node519;
	wire [8-1:0] node522;
	wire [8-1:0] node523;
	wire [8-1:0] node524;
	wire [8-1:0] node527;
	wire [8-1:0] node528;
	wire [8-1:0] node531;
	wire [8-1:0] node532;
	wire [8-1:0] node535;
	wire [8-1:0] node538;
	wire [8-1:0] node539;
	wire [8-1:0] node540;
	wire [8-1:0] node544;
	wire [8-1:0] node546;
	wire [8-1:0] node548;
	wire [8-1:0] node551;
	wire [8-1:0] node552;
	wire [8-1:0] node553;
	wire [8-1:0] node554;
	wire [8-1:0] node555;
	wire [8-1:0] node556;
	wire [8-1:0] node557;
	wire [8-1:0] node560;
	wire [8-1:0] node563;
	wire [8-1:0] node564;
	wire [8-1:0] node566;
	wire [8-1:0] node570;
	wire [8-1:0] node571;
	wire [8-1:0] node572;
	wire [8-1:0] node575;
	wire [8-1:0] node578;
	wire [8-1:0] node580;
	wire [8-1:0] node581;
	wire [8-1:0] node585;
	wire [8-1:0] node586;
	wire [8-1:0] node587;
	wire [8-1:0] node589;
	wire [8-1:0] node590;
	wire [8-1:0] node592;
	wire [8-1:0] node595;
	wire [8-1:0] node598;
	wire [8-1:0] node599;
	wire [8-1:0] node602;
	wire [8-1:0] node603;
	wire [8-1:0] node607;
	wire [8-1:0] node608;
	wire [8-1:0] node609;
	wire [8-1:0] node613;
	wire [8-1:0] node614;
	wire [8-1:0] node615;
	wire [8-1:0] node619;
	wire [8-1:0] node621;
	wire [8-1:0] node624;
	wire [8-1:0] node625;
	wire [8-1:0] node626;
	wire [8-1:0] node627;
	wire [8-1:0] node628;
	wire [8-1:0] node630;
	wire [8-1:0] node633;
	wire [8-1:0] node635;
	wire [8-1:0] node638;
	wire [8-1:0] node639;
	wire [8-1:0] node642;
	wire [8-1:0] node644;
	wire [8-1:0] node647;
	wire [8-1:0] node648;
	wire [8-1:0] node649;
	wire [8-1:0] node651;
	wire [8-1:0] node654;
	wire [8-1:0] node656;
	wire [8-1:0] node659;
	wire [8-1:0] node660;
	wire [8-1:0] node663;
	wire [8-1:0] node666;
	wire [8-1:0] node667;
	wire [8-1:0] node668;
	wire [8-1:0] node670;
	wire [8-1:0] node671;
	wire [8-1:0] node675;
	wire [8-1:0] node676;
	wire [8-1:0] node679;
	wire [8-1:0] node680;
	wire [8-1:0] node684;
	wire [8-1:0] node685;
	wire [8-1:0] node686;
	wire [8-1:0] node688;
	wire [8-1:0] node689;
	wire [8-1:0] node693;
	wire [8-1:0] node696;
	wire [8-1:0] node697;
	wire [8-1:0] node699;
	wire [8-1:0] node701;
	wire [8-1:0] node704;
	wire [8-1:0] node706;
	wire [8-1:0] node707;
	wire [8-1:0] node711;
	wire [8-1:0] node712;
	wire [8-1:0] node713;
	wire [8-1:0] node714;
	wire [8-1:0] node716;
	wire [8-1:0] node717;
	wire [8-1:0] node719;
	wire [8-1:0] node723;
	wire [8-1:0] node725;
	wire [8-1:0] node726;
	wire [8-1:0] node729;
	wire [8-1:0] node730;
	wire [8-1:0] node731;
	wire [8-1:0] node736;
	wire [8-1:0] node737;
	wire [8-1:0] node738;
	wire [8-1:0] node739;
	wire [8-1:0] node740;
	wire [8-1:0] node745;
	wire [8-1:0] node746;
	wire [8-1:0] node750;
	wire [8-1:0] node751;
	wire [8-1:0] node752;
	wire [8-1:0] node753;
	wire [8-1:0] node754;
	wire [8-1:0] node757;
	wire [8-1:0] node761;
	wire [8-1:0] node762;
	wire [8-1:0] node765;
	wire [8-1:0] node766;
	wire [8-1:0] node770;
	wire [8-1:0] node771;
	wire [8-1:0] node772;
	wire [8-1:0] node775;
	wire [8-1:0] node776;
	wire [8-1:0] node780;
	wire [8-1:0] node781;
	wire [8-1:0] node783;
	wire [8-1:0] node786;
	wire [8-1:0] node789;
	wire [8-1:0] node790;
	wire [8-1:0] node791;
	wire [8-1:0] node792;
	wire [8-1:0] node793;
	wire [8-1:0] node796;
	wire [8-1:0] node797;
	wire [8-1:0] node799;
	wire [8-1:0] node803;
	wire [8-1:0] node804;
	wire [8-1:0] node805;
	wire [8-1:0] node808;
	wire [8-1:0] node811;
	wire [8-1:0] node812;
	wire [8-1:0] node816;
	wire [8-1:0] node817;
	wire [8-1:0] node818;
	wire [8-1:0] node819;
	wire [8-1:0] node823;
	wire [8-1:0] node824;
	wire [8-1:0] node826;
	wire [8-1:0] node829;
	wire [8-1:0] node830;
	wire [8-1:0] node834;
	wire [8-1:0] node835;
	wire [8-1:0] node836;
	wire [8-1:0] node839;
	wire [8-1:0] node840;
	wire [8-1:0] node844;
	wire [8-1:0] node847;
	wire [8-1:0] node848;
	wire [8-1:0] node849;
	wire [8-1:0] node850;
	wire [8-1:0] node851;
	wire [8-1:0] node852;
	wire [8-1:0] node855;
	wire [8-1:0] node859;
	wire [8-1:0] node860;
	wire [8-1:0] node864;
	wire [8-1:0] node865;
	wire [8-1:0] node866;
	wire [8-1:0] node867;
	wire [8-1:0] node871;
	wire [8-1:0] node874;
	wire [8-1:0] node875;
	wire [8-1:0] node879;
	wire [8-1:0] node880;
	wire [8-1:0] node881;
	wire [8-1:0] node882;
	wire [8-1:0] node886;
	wire [8-1:0] node887;
	wire [8-1:0] node891;
	wire [8-1:0] node894;
	wire [8-1:0] node895;
	wire [8-1:0] node896;
	wire [8-1:0] node897;
	wire [8-1:0] node898;
	wire [8-1:0] node899;
	wire [8-1:0] node900;
	wire [8-1:0] node901;
	wire [8-1:0] node904;
	wire [8-1:0] node908;
	wire [8-1:0] node909;
	wire [8-1:0] node911;
	wire [8-1:0] node914;
	wire [8-1:0] node915;
	wire [8-1:0] node916;
	wire [8-1:0] node920;
	wire [8-1:0] node921;
	wire [8-1:0] node925;
	wire [8-1:0] node926;
	wire [8-1:0] node927;
	wire [8-1:0] node929;
	wire [8-1:0] node933;
	wire [8-1:0] node934;
	wire [8-1:0] node935;
	wire [8-1:0] node937;
	wire [8-1:0] node940;
	wire [8-1:0] node942;
	wire [8-1:0] node945;
	wire [8-1:0] node946;
	wire [8-1:0] node947;
	wire [8-1:0] node950;
	wire [8-1:0] node954;
	wire [8-1:0] node955;
	wire [8-1:0] node956;
	wire [8-1:0] node957;
	wire [8-1:0] node958;
	wire [8-1:0] node960;
	wire [8-1:0] node964;
	wire [8-1:0] node965;
	wire [8-1:0] node968;
	wire [8-1:0] node971;
	wire [8-1:0] node972;
	wire [8-1:0] node973;
	wire [8-1:0] node976;
	wire [8-1:0] node979;
	wire [8-1:0] node980;
	wire [8-1:0] node983;
	wire [8-1:0] node985;
	wire [8-1:0] node988;
	wire [8-1:0] node989;
	wire [8-1:0] node990;
	wire [8-1:0] node992;
	wire [8-1:0] node994;
	wire [8-1:0] node997;
	wire [8-1:0] node998;
	wire [8-1:0] node1000;
	wire [8-1:0] node1003;
	wire [8-1:0] node1006;
	wire [8-1:0] node1007;
	wire [8-1:0] node1008;
	wire [8-1:0] node1009;
	wire [8-1:0] node1013;
	wire [8-1:0] node1014;
	wire [8-1:0] node1017;
	wire [8-1:0] node1020;
	wire [8-1:0] node1021;
	wire [8-1:0] node1022;
	wire [8-1:0] node1026;
	wire [8-1:0] node1028;
	wire [8-1:0] node1029;
	wire [8-1:0] node1033;
	wire [8-1:0] node1034;
	wire [8-1:0] node1035;
	wire [8-1:0] node1036;
	wire [8-1:0] node1037;
	wire [8-1:0] node1038;
	wire [8-1:0] node1041;
	wire [8-1:0] node1043;
	wire [8-1:0] node1046;
	wire [8-1:0] node1048;
	wire [8-1:0] node1049;
	wire [8-1:0] node1053;
	wire [8-1:0] node1054;
	wire [8-1:0] node1056;
	wire [8-1:0] node1058;
	wire [8-1:0] node1061;
	wire [8-1:0] node1063;
	wire [8-1:0] node1066;
	wire [8-1:0] node1067;
	wire [8-1:0] node1068;
	wire [8-1:0] node1070;
	wire [8-1:0] node1073;
	wire [8-1:0] node1074;
	wire [8-1:0] node1078;
	wire [8-1:0] node1079;
	wire [8-1:0] node1080;
	wire [8-1:0] node1081;
	wire [8-1:0] node1084;
	wire [8-1:0] node1088;
	wire [8-1:0] node1089;
	wire [8-1:0] node1091;
	wire [8-1:0] node1094;
	wire [8-1:0] node1097;
	wire [8-1:0] node1098;
	wire [8-1:0] node1099;
	wire [8-1:0] node1100;
	wire [8-1:0] node1101;
	wire [8-1:0] node1104;
	wire [8-1:0] node1107;
	wire [8-1:0] node1108;
	wire [8-1:0] node1110;
	wire [8-1:0] node1113;
	wire [8-1:0] node1115;
	wire [8-1:0] node1118;
	wire [8-1:0] node1119;
	wire [8-1:0] node1120;
	wire [8-1:0] node1122;
	wire [8-1:0] node1126;
	wire [8-1:0] node1128;
	wire [8-1:0] node1131;
	wire [8-1:0] node1132;
	wire [8-1:0] node1133;
	wire [8-1:0] node1134;
	wire [8-1:0] node1136;
	wire [8-1:0] node1137;
	wire [8-1:0] node1141;
	wire [8-1:0] node1144;
	wire [8-1:0] node1145;
	wire [8-1:0] node1146;
	wire [8-1:0] node1151;
	wire [8-1:0] node1152;
	wire [8-1:0] node1153;
	wire [8-1:0] node1154;
	wire [8-1:0] node1155;
	wire [8-1:0] node1158;
	wire [8-1:0] node1161;
	wire [8-1:0] node1162;
	wire [8-1:0] node1166;
	wire [8-1:0] node1167;
	wire [8-1:0] node1170;
	wire [8-1:0] node1173;
	wire [8-1:0] node1174;
	wire [8-1:0] node1175;
	wire [8-1:0] node1178;
	wire [8-1:0] node1181;
	wire [8-1:0] node1184;
	wire [8-1:0] node1185;
	wire [8-1:0] node1186;
	wire [8-1:0] node1187;
	wire [8-1:0] node1188;
	wire [8-1:0] node1189;
	wire [8-1:0] node1192;
	wire [8-1:0] node1193;
	wire [8-1:0] node1197;
	wire [8-1:0] node1198;
	wire [8-1:0] node1200;
	wire [8-1:0] node1201;
	wire [8-1:0] node1206;
	wire [8-1:0] node1207;
	wire [8-1:0] node1208;
	wire [8-1:0] node1209;
	wire [8-1:0] node1213;
	wire [8-1:0] node1214;
	wire [8-1:0] node1218;
	wire [8-1:0] node1219;
	wire [8-1:0] node1223;
	wire [8-1:0] node1224;
	wire [8-1:0] node1225;
	wire [8-1:0] node1226;
	wire [8-1:0] node1227;
	wire [8-1:0] node1229;
	wire [8-1:0] node1233;
	wire [8-1:0] node1234;
	wire [8-1:0] node1235;
	wire [8-1:0] node1236;
	wire [8-1:0] node1240;
	wire [8-1:0] node1241;
	wire [8-1:0] node1245;
	wire [8-1:0] node1246;
	wire [8-1:0] node1249;
	wire [8-1:0] node1252;
	wire [8-1:0] node1253;
	wire [8-1:0] node1255;
	wire [8-1:0] node1257;
	wire [8-1:0] node1260;
	wire [8-1:0] node1261;
	wire [8-1:0] node1263;
	wire [8-1:0] node1266;
	wire [8-1:0] node1267;
	wire [8-1:0] node1271;
	wire [8-1:0] node1272;
	wire [8-1:0] node1273;
	wire [8-1:0] node1274;
	wire [8-1:0] node1277;
	wire [8-1:0] node1280;
	wire [8-1:0] node1282;
	wire [8-1:0] node1284;
	wire [8-1:0] node1287;
	wire [8-1:0] node1288;
	wire [8-1:0] node1289;
	wire [8-1:0] node1290;
	wire [8-1:0] node1291;
	wire [8-1:0] node1295;
	wire [8-1:0] node1298;
	wire [8-1:0] node1301;
	wire [8-1:0] node1302;
	wire [8-1:0] node1304;
	wire [8-1:0] node1307;
	wire [8-1:0] node1308;
	wire [8-1:0] node1309;
	wire [8-1:0] node1312;
	wire [8-1:0] node1316;
	wire [8-1:0] node1317;
	wire [8-1:0] node1318;
	wire [8-1:0] node1319;
	wire [8-1:0] node1320;
	wire [8-1:0] node1322;
	wire [8-1:0] node1324;
	wire [8-1:0] node1327;
	wire [8-1:0] node1329;
	wire [8-1:0] node1332;
	wire [8-1:0] node1333;
	wire [8-1:0] node1334;
	wire [8-1:0] node1337;
	wire [8-1:0] node1340;
	wire [8-1:0] node1341;
	wire [8-1:0] node1344;
	wire [8-1:0] node1347;
	wire [8-1:0] node1348;
	wire [8-1:0] node1349;
	wire [8-1:0] node1352;
	wire [8-1:0] node1353;
	wire [8-1:0] node1356;
	wire [8-1:0] node1359;
	wire [8-1:0] node1360;
	wire [8-1:0] node1362;
	wire [8-1:0] node1365;
	wire [8-1:0] node1366;
	wire [8-1:0] node1369;
	wire [8-1:0] node1372;
	wire [8-1:0] node1373;
	wire [8-1:0] node1374;
	wire [8-1:0] node1375;
	wire [8-1:0] node1376;
	wire [8-1:0] node1377;
	wire [8-1:0] node1381;
	wire [8-1:0] node1382;
	wire [8-1:0] node1383;
	wire [8-1:0] node1388;
	wire [8-1:0] node1389;
	wire [8-1:0] node1391;
	wire [8-1:0] node1394;
	wire [8-1:0] node1396;
	wire [8-1:0] node1398;
	wire [8-1:0] node1401;
	wire [8-1:0] node1402;
	wire [8-1:0] node1403;
	wire [8-1:0] node1405;
	wire [8-1:0] node1408;
	wire [8-1:0] node1409;
	wire [8-1:0] node1412;
	wire [8-1:0] node1413;
	wire [8-1:0] node1417;
	wire [8-1:0] node1418;
	wire [8-1:0] node1419;
	wire [8-1:0] node1420;
	wire [8-1:0] node1424;
	wire [8-1:0] node1427;
	wire [8-1:0] node1429;
	wire [8-1:0] node1432;
	wire [8-1:0] node1433;
	wire [8-1:0] node1434;
	wire [8-1:0] node1435;
	wire [8-1:0] node1438;
	wire [8-1:0] node1441;
	wire [8-1:0] node1442;
	wire [8-1:0] node1444;
	wire [8-1:0] node1447;
	wire [8-1:0] node1450;
	wire [8-1:0] node1451;
	wire [8-1:0] node1452;
	wire [8-1:0] node1455;
	wire [8-1:0] node1458;
	wire [8-1:0] node1461;
	wire [8-1:0] node1462;
	wire [8-1:0] node1463;
	wire [8-1:0] node1464;
	wire [8-1:0] node1465;
	wire [8-1:0] node1466;
	wire [8-1:0] node1467;
	wire [8-1:0] node1469;
	wire [8-1:0] node1472;
	wire [8-1:0] node1473;
	wire [8-1:0] node1477;
	wire [8-1:0] node1478;
	wire [8-1:0] node1479;
	wire [8-1:0] node1480;
	wire [8-1:0] node1481;
	wire [8-1:0] node1483;
	wire [8-1:0] node1486;
	wire [8-1:0] node1489;
	wire [8-1:0] node1491;
	wire [8-1:0] node1494;
	wire [8-1:0] node1495;
	wire [8-1:0] node1496;
	wire [8-1:0] node1499;
	wire [8-1:0] node1500;
	wire [8-1:0] node1505;
	wire [8-1:0] node1506;
	wire [8-1:0] node1507;
	wire [8-1:0] node1508;
	wire [8-1:0] node1509;
	wire [8-1:0] node1510;
	wire [8-1:0] node1515;
	wire [8-1:0] node1516;
	wire [8-1:0] node1520;
	wire [8-1:0] node1522;
	wire [8-1:0] node1525;
	wire [8-1:0] node1526;
	wire [8-1:0] node1528;
	wire [8-1:0] node1531;
	wire [8-1:0] node1533;
	wire [8-1:0] node1536;
	wire [8-1:0] node1537;
	wire [8-1:0] node1538;
	wire [8-1:0] node1540;
	wire [8-1:0] node1543;
	wire [8-1:0] node1544;
	wire [8-1:0] node1548;
	wire [8-1:0] node1549;
	wire [8-1:0] node1550;
	wire [8-1:0] node1551;
	wire [8-1:0] node1552;
	wire [8-1:0] node1556;
	wire [8-1:0] node1557;
	wire [8-1:0] node1561;
	wire [8-1:0] node1562;
	wire [8-1:0] node1566;
	wire [8-1:0] node1567;
	wire [8-1:0] node1568;
	wire [8-1:0] node1569;
	wire [8-1:0] node1572;
	wire [8-1:0] node1575;
	wire [8-1:0] node1578;
	wire [8-1:0] node1579;
	wire [8-1:0] node1583;
	wire [8-1:0] node1584;
	wire [8-1:0] node1585;
	wire [8-1:0] node1586;
	wire [8-1:0] node1587;
	wire [8-1:0] node1588;
	wire [8-1:0] node1590;
	wire [8-1:0] node1593;
	wire [8-1:0] node1595;
	wire [8-1:0] node1598;
	wire [8-1:0] node1600;
	wire [8-1:0] node1603;
	wire [8-1:0] node1604;
	wire [8-1:0] node1608;
	wire [8-1:0] node1609;
	wire [8-1:0] node1610;
	wire [8-1:0] node1611;
	wire [8-1:0] node1615;
	wire [8-1:0] node1616;
	wire [8-1:0] node1617;
	wire [8-1:0] node1622;
	wire [8-1:0] node1623;
	wire [8-1:0] node1624;
	wire [8-1:0] node1625;
	wire [8-1:0] node1630;
	wire [8-1:0] node1631;
	wire [8-1:0] node1635;
	wire [8-1:0] node1636;
	wire [8-1:0] node1637;
	wire [8-1:0] node1638;
	wire [8-1:0] node1642;
	wire [8-1:0] node1643;
	wire [8-1:0] node1645;
	wire [8-1:0] node1648;
	wire [8-1:0] node1649;
	wire [8-1:0] node1653;
	wire [8-1:0] node1654;
	wire [8-1:0] node1658;
	wire [8-1:0] node1659;
	wire [8-1:0] node1660;
	wire [8-1:0] node1661;
	wire [8-1:0] node1662;
	wire [8-1:0] node1663;
	wire [8-1:0] node1665;
	wire [8-1:0] node1668;
	wire [8-1:0] node1669;
	wire [8-1:0] node1672;
	wire [8-1:0] node1673;
	wire [8-1:0] node1676;
	wire [8-1:0] node1679;
	wire [8-1:0] node1680;
	wire [8-1:0] node1681;
	wire [8-1:0] node1683;
	wire [8-1:0] node1686;
	wire [8-1:0] node1687;
	wire [8-1:0] node1690;
	wire [8-1:0] node1692;
	wire [8-1:0] node1695;
	wire [8-1:0] node1696;
	wire [8-1:0] node1698;
	wire [8-1:0] node1701;
	wire [8-1:0] node1702;
	wire [8-1:0] node1705;
	wire [8-1:0] node1706;
	wire [8-1:0] node1709;
	wire [8-1:0] node1712;
	wire [8-1:0] node1713;
	wire [8-1:0] node1714;
	wire [8-1:0] node1715;
	wire [8-1:0] node1717;
	wire [8-1:0] node1718;
	wire [8-1:0] node1722;
	wire [8-1:0] node1723;
	wire [8-1:0] node1724;
	wire [8-1:0] node1726;
	wire [8-1:0] node1729;
	wire [8-1:0] node1730;
	wire [8-1:0] node1734;
	wire [8-1:0] node1737;
	wire [8-1:0] node1738;
	wire [8-1:0] node1739;
	wire [8-1:0] node1740;
	wire [8-1:0] node1742;
	wire [8-1:0] node1745;
	wire [8-1:0] node1746;
	wire [8-1:0] node1749;
	wire [8-1:0] node1752;
	wire [8-1:0] node1754;
	wire [8-1:0] node1756;
	wire [8-1:0] node1759;
	wire [8-1:0] node1760;
	wire [8-1:0] node1762;
	wire [8-1:0] node1765;
	wire [8-1:0] node1768;
	wire [8-1:0] node1769;
	wire [8-1:0] node1770;
	wire [8-1:0] node1771;
	wire [8-1:0] node1772;
	wire [8-1:0] node1773;
	wire [8-1:0] node1776;
	wire [8-1:0] node1779;
	wire [8-1:0] node1781;
	wire [8-1:0] node1784;
	wire [8-1:0] node1785;
	wire [8-1:0] node1787;
	wire [8-1:0] node1791;
	wire [8-1:0] node1792;
	wire [8-1:0] node1793;
	wire [8-1:0] node1796;
	wire [8-1:0] node1799;
	wire [8-1:0] node1801;
	wire [8-1:0] node1804;
	wire [8-1:0] node1805;
	wire [8-1:0] node1806;
	wire [8-1:0] node1808;
	wire [8-1:0] node1811;
	wire [8-1:0] node1812;
	wire [8-1:0] node1815;
	wire [8-1:0] node1818;
	wire [8-1:0] node1819;
	wire [8-1:0] node1821;
	wire [8-1:0] node1824;
	wire [8-1:0] node1825;
	wire [8-1:0] node1828;
	wire [8-1:0] node1829;
	wire [8-1:0] node1833;
	wire [8-1:0] node1834;
	wire [8-1:0] node1835;
	wire [8-1:0] node1836;
	wire [8-1:0] node1837;
	wire [8-1:0] node1838;
	wire [8-1:0] node1842;
	wire [8-1:0] node1843;
	wire [8-1:0] node1846;
	wire [8-1:0] node1847;
	wire [8-1:0] node1850;
	wire [8-1:0] node1853;
	wire [8-1:0] node1854;
	wire [8-1:0] node1855;
	wire [8-1:0] node1857;
	wire [8-1:0] node1858;
	wire [8-1:0] node1862;
	wire [8-1:0] node1864;
	wire [8-1:0] node1866;
	wire [8-1:0] node1869;
	wire [8-1:0] node1870;
	wire [8-1:0] node1871;
	wire [8-1:0] node1875;
	wire [8-1:0] node1876;
	wire [8-1:0] node1877;
	wire [8-1:0] node1882;
	wire [8-1:0] node1883;
	wire [8-1:0] node1884;
	wire [8-1:0] node1885;
	wire [8-1:0] node1888;
	wire [8-1:0] node1890;
	wire [8-1:0] node1893;
	wire [8-1:0] node1895;
	wire [8-1:0] node1897;
	wire [8-1:0] node1900;
	wire [8-1:0] node1901;
	wire [8-1:0] node1902;
	wire [8-1:0] node1905;
	wire [8-1:0] node1908;
	wire [8-1:0] node1909;
	wire [8-1:0] node1910;
	wire [8-1:0] node1913;
	wire [8-1:0] node1916;
	wire [8-1:0] node1918;
	wire [8-1:0] node1921;
	wire [8-1:0] node1922;
	wire [8-1:0] node1923;
	wire [8-1:0] node1924;
	wire [8-1:0] node1925;
	wire [8-1:0] node1926;
	wire [8-1:0] node1930;
	wire [8-1:0] node1932;
	wire [8-1:0] node1934;
	wire [8-1:0] node1937;
	wire [8-1:0] node1938;
	wire [8-1:0] node1939;
	wire [8-1:0] node1943;
	wire [8-1:0] node1944;
	wire [8-1:0] node1947;
	wire [8-1:0] node1950;
	wire [8-1:0] node1951;
	wire [8-1:0] node1952;
	wire [8-1:0] node1955;
	wire [8-1:0] node1957;
	wire [8-1:0] node1960;
	wire [8-1:0] node1961;
	wire [8-1:0] node1963;
	wire [8-1:0] node1966;
	wire [8-1:0] node1969;
	wire [8-1:0] node1970;
	wire [8-1:0] node1971;
	wire [8-1:0] node1972;
	wire [8-1:0] node1976;
	wire [8-1:0] node1977;
	wire [8-1:0] node1978;
	wire [8-1:0] node1980;
	wire [8-1:0] node1983;
	wire [8-1:0] node1984;
	wire [8-1:0] node1988;
	wire [8-1:0] node1990;
	wire [8-1:0] node1993;
	wire [8-1:0] node1994;
	wire [8-1:0] node1995;
	wire [8-1:0] node1997;
	wire [8-1:0] node1999;
	wire [8-1:0] node2003;
	wire [8-1:0] node2004;
	wire [8-1:0] node2005;
	wire [8-1:0] node2006;
	wire [8-1:0] node2009;
	wire [8-1:0] node2012;
	wire [8-1:0] node2016;
	wire [8-1:0] node2017;
	wire [8-1:0] node2018;
	wire [8-1:0] node2019;
	wire [8-1:0] node2020;
	wire [8-1:0] node2021;
	wire [8-1:0] node2023;
	wire [8-1:0] node2026;
	wire [8-1:0] node2029;
	wire [8-1:0] node2031;
	wire [8-1:0] node2032;
	wire [8-1:0] node2036;
	wire [8-1:0] node2037;
	wire [8-1:0] node2038;
	wire [8-1:0] node2040;
	wire [8-1:0] node2043;
	wire [8-1:0] node2044;
	wire [8-1:0] node2047;
	wire [8-1:0] node2048;
	wire [8-1:0] node2051;
	wire [8-1:0] node2054;
	wire [8-1:0] node2055;
	wire [8-1:0] node2057;
	wire [8-1:0] node2060;
	wire [8-1:0] node2061;
	wire [8-1:0] node2065;
	wire [8-1:0] node2066;
	wire [8-1:0] node2067;
	wire [8-1:0] node2068;
	wire [8-1:0] node2071;
	wire [8-1:0] node2072;
	wire [8-1:0] node2074;
	wire [8-1:0] node2077;
	wire [8-1:0] node2079;
	wire [8-1:0] node2082;
	wire [8-1:0] node2083;
	wire [8-1:0] node2084;
	wire [8-1:0] node2085;
	wire [8-1:0] node2088;
	wire [8-1:0] node2089;
	wire [8-1:0] node2092;
	wire [8-1:0] node2095;
	wire [8-1:0] node2096;
	wire [8-1:0] node2099;
	wire [8-1:0] node2100;
	wire [8-1:0] node2104;
	wire [8-1:0] node2105;
	wire [8-1:0] node2106;
	wire [8-1:0] node2110;
	wire [8-1:0] node2113;
	wire [8-1:0] node2114;
	wire [8-1:0] node2115;
	wire [8-1:0] node2116;
	wire [8-1:0] node2118;
	wire [8-1:0] node2121;
	wire [8-1:0] node2122;
	wire [8-1:0] node2123;
	wire [8-1:0] node2126;
	wire [8-1:0] node2130;
	wire [8-1:0] node2131;
	wire [8-1:0] node2132;
	wire [8-1:0] node2133;
	wire [8-1:0] node2138;
	wire [8-1:0] node2140;
	wire [8-1:0] node2143;
	wire [8-1:0] node2144;
	wire [8-1:0] node2145;
	wire [8-1:0] node2148;
	wire [8-1:0] node2149;
	wire [8-1:0] node2153;
	wire [8-1:0] node2154;
	wire [8-1:0] node2156;
	wire [8-1:0] node2158;
	wire [8-1:0] node2161;
	wire [8-1:0] node2163;
	wire [8-1:0] node2164;
	wire [8-1:0] node2168;
	wire [8-1:0] node2169;
	wire [8-1:0] node2170;
	wire [8-1:0] node2171;
	wire [8-1:0] node2172;
	wire [8-1:0] node2173;
	wire [8-1:0] node2177;
	wire [8-1:0] node2178;
	wire [8-1:0] node2181;
	wire [8-1:0] node2183;
	wire [8-1:0] node2186;
	wire [8-1:0] node2187;
	wire [8-1:0] node2188;
	wire [8-1:0] node2191;
	wire [8-1:0] node2194;
	wire [8-1:0] node2196;
	wire [8-1:0] node2199;
	wire [8-1:0] node2200;
	wire [8-1:0] node2201;
	wire [8-1:0] node2203;
	wire [8-1:0] node2206;
	wire [8-1:0] node2207;
	wire [8-1:0] node2209;
	wire [8-1:0] node2212;
	wire [8-1:0] node2215;
	wire [8-1:0] node2216;
	wire [8-1:0] node2217;
	wire [8-1:0] node2218;
	wire [8-1:0] node2222;
	wire [8-1:0] node2223;
	wire [8-1:0] node2226;
	wire [8-1:0] node2229;
	wire [8-1:0] node2230;
	wire [8-1:0] node2231;
	wire [8-1:0] node2234;
	wire [8-1:0] node2238;
	wire [8-1:0] node2239;
	wire [8-1:0] node2240;
	wire [8-1:0] node2241;
	wire [8-1:0] node2242;
	wire [8-1:0] node2244;
	wire [8-1:0] node2245;
	wire [8-1:0] node2249;
	wire [8-1:0] node2252;
	wire [8-1:0] node2253;
	wire [8-1:0] node2254;
	wire [8-1:0] node2256;
	wire [8-1:0] node2259;
	wire [8-1:0] node2261;
	wire [8-1:0] node2264;
	wire [8-1:0] node2267;
	wire [8-1:0] node2268;
	wire [8-1:0] node2270;
	wire [8-1:0] node2272;
	wire [8-1:0] node2275;
	wire [8-1:0] node2276;
	wire [8-1:0] node2278;
	wire [8-1:0] node2281;
	wire [8-1:0] node2283;
	wire [8-1:0] node2284;
	wire [8-1:0] node2288;
	wire [8-1:0] node2289;
	wire [8-1:0] node2290;
	wire [8-1:0] node2292;
	wire [8-1:0] node2293;
	wire [8-1:0] node2296;
	wire [8-1:0] node2299;
	wire [8-1:0] node2300;
	wire [8-1:0] node2303;
	wire [8-1:0] node2304;
	wire [8-1:0] node2305;
	wire [8-1:0] node2309;
	wire [8-1:0] node2312;
	wire [8-1:0] node2313;
	wire [8-1:0] node2314;
	wire [8-1:0] node2315;
	wire [8-1:0] node2316;
	wire [8-1:0] node2320;
	wire [8-1:0] node2322;
	wire [8-1:0] node2326;
	wire [8-1:0] node2327;
	wire [8-1:0] node2330;
	wire [8-1:0] node2331;
	wire [8-1:0] node2334;
	wire [8-1:0] node2337;
	wire [8-1:0] node2338;
	wire [8-1:0] node2339;
	wire [8-1:0] node2340;
	wire [8-1:0] node2341;
	wire [8-1:0] node2342;
	wire [8-1:0] node2343;
	wire [8-1:0] node2345;
	wire [8-1:0] node2347;
	wire [8-1:0] node2350;
	wire [8-1:0] node2351;
	wire [8-1:0] node2353;
	wire [8-1:0] node2356;
	wire [8-1:0] node2357;
	wire [8-1:0] node2361;
	wire [8-1:0] node2362;
	wire [8-1:0] node2363;
	wire [8-1:0] node2365;
	wire [8-1:0] node2368;
	wire [8-1:0] node2370;
	wire [8-1:0] node2373;
	wire [8-1:0] node2374;
	wire [8-1:0] node2375;
	wire [8-1:0] node2378;
	wire [8-1:0] node2381;
	wire [8-1:0] node2384;
	wire [8-1:0] node2385;
	wire [8-1:0] node2386;
	wire [8-1:0] node2387;
	wire [8-1:0] node2389;
	wire [8-1:0] node2392;
	wire [8-1:0] node2393;
	wire [8-1:0] node2394;
	wire [8-1:0] node2399;
	wire [8-1:0] node2400;
	wire [8-1:0] node2402;
	wire [8-1:0] node2405;
	wire [8-1:0] node2406;
	wire [8-1:0] node2409;
	wire [8-1:0] node2411;
	wire [8-1:0] node2414;
	wire [8-1:0] node2415;
	wire [8-1:0] node2416;
	wire [8-1:0] node2419;
	wire [8-1:0] node2422;
	wire [8-1:0] node2423;
	wire [8-1:0] node2427;
	wire [8-1:0] node2428;
	wire [8-1:0] node2429;
	wire [8-1:0] node2430;
	wire [8-1:0] node2432;
	wire [8-1:0] node2434;
	wire [8-1:0] node2437;
	wire [8-1:0] node2438;
	wire [8-1:0] node2440;
	wire [8-1:0] node2443;
	wire [8-1:0] node2445;
	wire [8-1:0] node2448;
	wire [8-1:0] node2449;
	wire [8-1:0] node2450;
	wire [8-1:0] node2452;
	wire [8-1:0] node2455;
	wire [8-1:0] node2458;
	wire [8-1:0] node2459;
	wire [8-1:0] node2462;
	wire [8-1:0] node2463;
	wire [8-1:0] node2466;
	wire [8-1:0] node2469;
	wire [8-1:0] node2470;
	wire [8-1:0] node2471;
	wire [8-1:0] node2472;
	wire [8-1:0] node2474;
	wire [8-1:0] node2477;
	wire [8-1:0] node2479;
	wire [8-1:0] node2482;
	wire [8-1:0] node2483;
	wire [8-1:0] node2485;
	wire [8-1:0] node2486;
	wire [8-1:0] node2490;
	wire [8-1:0] node2491;
	wire [8-1:0] node2492;
	wire [8-1:0] node2495;
	wire [8-1:0] node2499;
	wire [8-1:0] node2500;
	wire [8-1:0] node2501;
	wire [8-1:0] node2503;
	wire [8-1:0] node2504;
	wire [8-1:0] node2508;
	wire [8-1:0] node2509;
	wire [8-1:0] node2511;
	wire [8-1:0] node2514;
	wire [8-1:0] node2517;
	wire [8-1:0] node2518;
	wire [8-1:0] node2521;
	wire [8-1:0] node2523;
	wire [8-1:0] node2524;
	wire [8-1:0] node2528;
	wire [8-1:0] node2529;
	wire [8-1:0] node2531;
	wire [8-1:0] node2533;
	wire [8-1:0] node2536;
	wire [8-1:0] node2537;
	wire [8-1:0] node2538;
	wire [8-1:0] node2539;
	wire [8-1:0] node2540;
	wire [8-1:0] node2542;
	wire [8-1:0] node2545;
	wire [8-1:0] node2546;
	wire [8-1:0] node2550;
	wire [8-1:0] node2551;
	wire [8-1:0] node2555;
	wire [8-1:0] node2556;
	wire [8-1:0] node2557;
	wire [8-1:0] node2558;
	wire [8-1:0] node2562;
	wire [8-1:0] node2565;
	wire [8-1:0] node2566;
	wire [8-1:0] node2567;
	wire [8-1:0] node2570;
	wire [8-1:0] node2573;
	wire [8-1:0] node2574;
	wire [8-1:0] node2578;
	wire [8-1:0] node2579;
	wire [8-1:0] node2580;
	wire [8-1:0] node2581;
	wire [8-1:0] node2585;
	wire [8-1:0] node2586;
	wire [8-1:0] node2590;
	wire [8-1:0] node2591;
	wire [8-1:0] node2594;
	wire [8-1:0] node2597;
	wire [8-1:0] node2598;
	wire [8-1:0] node2599;
	wire [8-1:0] node2600;
	wire [8-1:0] node2601;
	wire [8-1:0] node2602;
	wire [8-1:0] node2604;
	wire [8-1:0] node2605;
	wire [8-1:0] node2606;
	wire [8-1:0] node2609;
	wire [8-1:0] node2612;
	wire [8-1:0] node2613;
	wire [8-1:0] node2616;
	wire [8-1:0] node2619;
	wire [8-1:0] node2621;
	wire [8-1:0] node2622;
	wire [8-1:0] node2625;
	wire [8-1:0] node2626;
	wire [8-1:0] node2630;
	wire [8-1:0] node2631;
	wire [8-1:0] node2632;
	wire [8-1:0] node2633;
	wire [8-1:0] node2637;
	wire [8-1:0] node2639;
	wire [8-1:0] node2642;
	wire [8-1:0] node2643;
	wire [8-1:0] node2644;
	wire [8-1:0] node2645;
	wire [8-1:0] node2649;
	wire [8-1:0] node2651;
	wire [8-1:0] node2654;
	wire [8-1:0] node2655;
	wire [8-1:0] node2656;
	wire [8-1:0] node2657;
	wire [8-1:0] node2662;
	wire [8-1:0] node2664;
	wire [8-1:0] node2667;
	wire [8-1:0] node2668;
	wire [8-1:0] node2669;
	wire [8-1:0] node2670;
	wire [8-1:0] node2671;
	wire [8-1:0] node2674;
	wire [8-1:0] node2677;
	wire [8-1:0] node2678;
	wire [8-1:0] node2679;
	wire [8-1:0] node2682;
	wire [8-1:0] node2685;
	wire [8-1:0] node2686;
	wire [8-1:0] node2690;
	wire [8-1:0] node2691;
	wire [8-1:0] node2692;
	wire [8-1:0] node2693;
	wire [8-1:0] node2696;
	wire [8-1:0] node2698;
	wire [8-1:0] node2701;
	wire [8-1:0] node2702;
	wire [8-1:0] node2705;
	wire [8-1:0] node2708;
	wire [8-1:0] node2709;
	wire [8-1:0] node2712;
	wire [8-1:0] node2714;
	wire [8-1:0] node2717;
	wire [8-1:0] node2718;
	wire [8-1:0] node2719;
	wire [8-1:0] node2720;
	wire [8-1:0] node2722;
	wire [8-1:0] node2726;
	wire [8-1:0] node2727;
	wire [8-1:0] node2730;
	wire [8-1:0] node2732;
	wire [8-1:0] node2735;
	wire [8-1:0] node2736;
	wire [8-1:0] node2737;
	wire [8-1:0] node2738;
	wire [8-1:0] node2742;
	wire [8-1:0] node2745;
	wire [8-1:0] node2747;
	wire [8-1:0] node2750;
	wire [8-1:0] node2751;
	wire [8-1:0] node2752;
	wire [8-1:0] node2753;
	wire [8-1:0] node2754;
	wire [8-1:0] node2757;
	wire [8-1:0] node2758;
	wire [8-1:0] node2761;
	wire [8-1:0] node2764;
	wire [8-1:0] node2765;
	wire [8-1:0] node2766;
	wire [8-1:0] node2767;
	wire [8-1:0] node2770;
	wire [8-1:0] node2771;
	wire [8-1:0] node2775;
	wire [8-1:0] node2776;
	wire [8-1:0] node2779;
	wire [8-1:0] node2780;
	wire [8-1:0] node2784;
	wire [8-1:0] node2785;
	wire [8-1:0] node2786;
	wire [8-1:0] node2789;
	wire [8-1:0] node2793;
	wire [8-1:0] node2794;
	wire [8-1:0] node2795;
	wire [8-1:0] node2796;
	wire [8-1:0] node2799;
	wire [8-1:0] node2801;
	wire [8-1:0] node2804;
	wire [8-1:0] node2805;
	wire [8-1:0] node2806;
	wire [8-1:0] node2809;
	wire [8-1:0] node2812;
	wire [8-1:0] node2813;
	wire [8-1:0] node2816;
	wire [8-1:0] node2817;
	wire [8-1:0] node2820;
	wire [8-1:0] node2823;
	wire [8-1:0] node2824;
	wire [8-1:0] node2825;
	wire [8-1:0] node2827;
	wire [8-1:0] node2830;
	wire [8-1:0] node2832;
	wire [8-1:0] node2835;
	wire [8-1:0] node2836;
	wire [8-1:0] node2838;
	wire [8-1:0] node2841;
	wire [8-1:0] node2843;
	wire [8-1:0] node2846;
	wire [8-1:0] node2847;
	wire [8-1:0] node2848;
	wire [8-1:0] node2849;
	wire [8-1:0] node2852;
	wire [8-1:0] node2854;
	wire [8-1:0] node2857;
	wire [8-1:0] node2858;
	wire [8-1:0] node2861;
	wire [8-1:0] node2862;
	wire [8-1:0] node2863;
	wire [8-1:0] node2867;
	wire [8-1:0] node2868;
	wire [8-1:0] node2872;
	wire [8-1:0] node2873;
	wire [8-1:0] node2874;
	wire [8-1:0] node2876;
	wire [8-1:0] node2877;
	wire [8-1:0] node2881;
	wire [8-1:0] node2883;
	wire [8-1:0] node2886;
	wire [8-1:0] node2887;
	wire [8-1:0] node2889;
	wire [8-1:0] node2892;
	wire [8-1:0] node2894;
	wire [8-1:0] node2897;
	wire [8-1:0] node2898;
	wire [8-1:0] node2899;
	wire [8-1:0] node2900;
	wire [8-1:0] node2901;
	wire [8-1:0] node2902;
	wire [8-1:0] node2903;
	wire [8-1:0] node2906;
	wire [8-1:0] node2907;
	wire [8-1:0] node2911;
	wire [8-1:0] node2912;
	wire [8-1:0] node2915;
	wire [8-1:0] node2916;
	wire [8-1:0] node2920;
	wire [8-1:0] node2921;
	wire [8-1:0] node2923;
	wire [8-1:0] node2926;
	wire [8-1:0] node2927;
	wire [8-1:0] node2929;
	wire [8-1:0] node2932;
	wire [8-1:0] node2933;
	wire [8-1:0] node2936;
	wire [8-1:0] node2939;
	wire [8-1:0] node2940;
	wire [8-1:0] node2941;
	wire [8-1:0] node2942;
	wire [8-1:0] node2945;
	wire [8-1:0] node2946;
	wire [8-1:0] node2950;
	wire [8-1:0] node2951;
	wire [8-1:0] node2954;
	wire [8-1:0] node2955;
	wire [8-1:0] node2958;
	wire [8-1:0] node2961;
	wire [8-1:0] node2962;
	wire [8-1:0] node2964;
	wire [8-1:0] node2967;
	wire [8-1:0] node2968;
	wire [8-1:0] node2971;
	wire [8-1:0] node2972;
	wire [8-1:0] node2975;
	wire [8-1:0] node2978;
	wire [8-1:0] node2979;
	wire [8-1:0] node2980;
	wire [8-1:0] node2983;
	wire [8-1:0] node2984;
	wire [8-1:0] node2985;
	wire [8-1:0] node2988;
	wire [8-1:0] node2991;
	wire [8-1:0] node2993;
	wire [8-1:0] node2996;
	wire [8-1:0] node2997;
	wire [8-1:0] node2999;
	wire [8-1:0] node3002;
	wire [8-1:0] node3004;
	wire [8-1:0] node3007;
	wire [8-1:0] node3008;
	wire [8-1:0] node3009;
	wire [8-1:0] node3010;
	wire [8-1:0] node3011;
	wire [8-1:0] node3013;
	wire [8-1:0] node3014;
	wire [8-1:0] node3017;
	wire [8-1:0] node3020;
	wire [8-1:0] node3021;
	wire [8-1:0] node3024;
	wire [8-1:0] node3027;
	wire [8-1:0] node3028;
	wire [8-1:0] node3029;
	wire [8-1:0] node3032;
	wire [8-1:0] node3033;
	wire [8-1:0] node3036;
	wire [8-1:0] node3039;
	wire [8-1:0] node3040;
	wire [8-1:0] node3041;
	wire [8-1:0] node3045;
	wire [8-1:0] node3047;
	wire [8-1:0] node3048;
	wire [8-1:0] node3052;
	wire [8-1:0] node3053;
	wire [8-1:0] node3056;
	wire [8-1:0] node3057;
	wire [8-1:0] node3060;
	wire [8-1:0] node3063;
	wire [8-1:0] node3064;
	wire [8-1:0] node3065;
	wire [8-1:0] node3066;
	wire [8-1:0] node3067;
	wire [8-1:0] node3068;
	wire [8-1:0] node3071;
	wire [8-1:0] node3074;
	wire [8-1:0] node3075;
	wire [8-1:0] node3078;
	wire [8-1:0] node3081;
	wire [8-1:0] node3082;
	wire [8-1:0] node3083;
	wire [8-1:0] node3084;
	wire [8-1:0] node3089;
	wire [8-1:0] node3090;
	wire [8-1:0] node3093;
	wire [8-1:0] node3096;
	wire [8-1:0] node3097;
	wire [8-1:0] node3098;
	wire [8-1:0] node3099;
	wire [8-1:0] node3102;
	wire [8-1:0] node3105;
	wire [8-1:0] node3106;
	wire [8-1:0] node3110;
	wire [8-1:0] node3111;
	wire [8-1:0] node3113;
	wire [8-1:0] node3114;
	wire [8-1:0] node3118;
	wire [8-1:0] node3121;
	wire [8-1:0] node3124;
	wire [8-1:0] node3125;
	wire [8-1:0] node3126;
	wire [8-1:0] node3127;
	wire [8-1:0] node3128;
	wire [8-1:0] node3129;
	wire [8-1:0] node3130;
	wire [8-1:0] node3131;
	wire [8-1:0] node3132;
	wire [8-1:0] node3133;
	wire [8-1:0] node3135;
	wire [8-1:0] node3138;
	wire [8-1:0] node3140;
	wire [8-1:0] node3141;
	wire [8-1:0] node3145;
	wire [8-1:0] node3146;
	wire [8-1:0] node3147;
	wire [8-1:0] node3150;
	wire [8-1:0] node3151;
	wire [8-1:0] node3155;
	wire [8-1:0] node3156;
	wire [8-1:0] node3158;
	wire [8-1:0] node3160;
	wire [8-1:0] node3164;
	wire [8-1:0] node3165;
	wire [8-1:0] node3166;
	wire [8-1:0] node3168;
	wire [8-1:0] node3171;
	wire [8-1:0] node3172;
	wire [8-1:0] node3176;
	wire [8-1:0] node3177;
	wire [8-1:0] node3178;
	wire [8-1:0] node3180;
	wire [8-1:0] node3183;
	wire [8-1:0] node3185;
	wire [8-1:0] node3188;
	wire [8-1:0] node3189;
	wire [8-1:0] node3192;
	wire [8-1:0] node3195;
	wire [8-1:0] node3196;
	wire [8-1:0] node3197;
	wire [8-1:0] node3198;
	wire [8-1:0] node3199;
	wire [8-1:0] node3201;
	wire [8-1:0] node3205;
	wire [8-1:0] node3206;
	wire [8-1:0] node3208;
	wire [8-1:0] node3211;
	wire [8-1:0] node3212;
	wire [8-1:0] node3216;
	wire [8-1:0] node3217;
	wire [8-1:0] node3218;
	wire [8-1:0] node3221;
	wire [8-1:0] node3224;
	wire [8-1:0] node3225;
	wire [8-1:0] node3226;
	wire [8-1:0] node3229;
	wire [8-1:0] node3232;
	wire [8-1:0] node3235;
	wire [8-1:0] node3236;
	wire [8-1:0] node3237;
	wire [8-1:0] node3238;
	wire [8-1:0] node3240;
	wire [8-1:0] node3243;
	wire [8-1:0] node3244;
	wire [8-1:0] node3247;
	wire [8-1:0] node3250;
	wire [8-1:0] node3251;
	wire [8-1:0] node3254;
	wire [8-1:0] node3255;
	wire [8-1:0] node3256;
	wire [8-1:0] node3259;
	wire [8-1:0] node3262;
	wire [8-1:0] node3265;
	wire [8-1:0] node3266;
	wire [8-1:0] node3267;
	wire [8-1:0] node3268;
	wire [8-1:0] node3272;
	wire [8-1:0] node3274;
	wire [8-1:0] node3277;
	wire [8-1:0] node3278;
	wire [8-1:0] node3280;
	wire [8-1:0] node3283;
	wire [8-1:0] node3286;
	wire [8-1:0] node3287;
	wire [8-1:0] node3288;
	wire [8-1:0] node3289;
	wire [8-1:0] node3290;
	wire [8-1:0] node3292;
	wire [8-1:0] node3293;
	wire [8-1:0] node3296;
	wire [8-1:0] node3299;
	wire [8-1:0] node3300;
	wire [8-1:0] node3302;
	wire [8-1:0] node3306;
	wire [8-1:0] node3307;
	wire [8-1:0] node3309;
	wire [8-1:0] node3310;
	wire [8-1:0] node3314;
	wire [8-1:0] node3315;
	wire [8-1:0] node3318;
	wire [8-1:0] node3320;
	wire [8-1:0] node3323;
	wire [8-1:0] node3324;
	wire [8-1:0] node3325;
	wire [8-1:0] node3326;
	wire [8-1:0] node3328;
	wire [8-1:0] node3331;
	wire [8-1:0] node3332;
	wire [8-1:0] node3336;
	wire [8-1:0] node3337;
	wire [8-1:0] node3339;
	wire [8-1:0] node3342;
	wire [8-1:0] node3343;
	wire [8-1:0] node3346;
	wire [8-1:0] node3349;
	wire [8-1:0] node3350;
	wire [8-1:0] node3352;
	wire [8-1:0] node3356;
	wire [8-1:0] node3357;
	wire [8-1:0] node3358;
	wire [8-1:0] node3359;
	wire [8-1:0] node3360;
	wire [8-1:0] node3362;
	wire [8-1:0] node3366;
	wire [8-1:0] node3367;
	wire [8-1:0] node3368;
	wire [8-1:0] node3372;
	wire [8-1:0] node3375;
	wire [8-1:0] node3376;
	wire [8-1:0] node3378;
	wire [8-1:0] node3380;
	wire [8-1:0] node3383;
	wire [8-1:0] node3384;
	wire [8-1:0] node3386;
	wire [8-1:0] node3389;
	wire [8-1:0] node3390;
	wire [8-1:0] node3393;
	wire [8-1:0] node3396;
	wire [8-1:0] node3397;
	wire [8-1:0] node3398;
	wire [8-1:0] node3400;
	wire [8-1:0] node3401;
	wire [8-1:0] node3404;
	wire [8-1:0] node3405;
	wire [8-1:0] node3408;
	wire [8-1:0] node3411;
	wire [8-1:0] node3412;
	wire [8-1:0] node3414;
	wire [8-1:0] node3417;
	wire [8-1:0] node3420;
	wire [8-1:0] node3421;
	wire [8-1:0] node3422;
	wire [8-1:0] node3423;
	wire [8-1:0] node3427;
	wire [8-1:0] node3428;
	wire [8-1:0] node3431;
	wire [8-1:0] node3433;
	wire [8-1:0] node3436;
	wire [8-1:0] node3437;
	wire [8-1:0] node3440;
	wire [8-1:0] node3443;
	wire [8-1:0] node3444;
	wire [8-1:0] node3445;
	wire [8-1:0] node3446;
	wire [8-1:0] node3447;
	wire [8-1:0] node3448;
	wire [8-1:0] node3451;
	wire [8-1:0] node3452;
	wire [8-1:0] node3456;
	wire [8-1:0] node3457;
	wire [8-1:0] node3458;
	wire [8-1:0] node3459;
	wire [8-1:0] node3463;
	wire [8-1:0] node3464;
	wire [8-1:0] node3468;
	wire [8-1:0] node3469;
	wire [8-1:0] node3473;
	wire [8-1:0] node3474;
	wire [8-1:0] node3475;
	wire [8-1:0] node3478;
	wire [8-1:0] node3480;
	wire [8-1:0] node3483;
	wire [8-1:0] node3484;
	wire [8-1:0] node3488;
	wire [8-1:0] node3489;
	wire [8-1:0] node3490;
	wire [8-1:0] node3491;
	wire [8-1:0] node3492;
	wire [8-1:0] node3495;
	wire [8-1:0] node3498;
	wire [8-1:0] node3500;
	wire [8-1:0] node3503;
	wire [8-1:0] node3504;
	wire [8-1:0] node3505;
	wire [8-1:0] node3506;
	wire [8-1:0] node3510;
	wire [8-1:0] node3513;
	wire [8-1:0] node3514;
	wire [8-1:0] node3516;
	wire [8-1:0] node3519;
	wire [8-1:0] node3520;
	wire [8-1:0] node3522;
	wire [8-1:0] node3526;
	wire [8-1:0] node3527;
	wire [8-1:0] node3528;
	wire [8-1:0] node3530;
	wire [8-1:0] node3533;
	wire [8-1:0] node3534;
	wire [8-1:0] node3537;
	wire [8-1:0] node3540;
	wire [8-1:0] node3541;
	wire [8-1:0] node3542;
	wire [8-1:0] node3544;
	wire [8-1:0] node3545;
	wire [8-1:0] node3549;
	wire [8-1:0] node3551;
	wire [8-1:0] node3553;
	wire [8-1:0] node3556;
	wire [8-1:0] node3557;
	wire [8-1:0] node3558;
	wire [8-1:0] node3561;
	wire [8-1:0] node3564;
	wire [8-1:0] node3566;
	wire [8-1:0] node3569;
	wire [8-1:0] node3570;
	wire [8-1:0] node3571;
	wire [8-1:0] node3572;
	wire [8-1:0] node3573;
	wire [8-1:0] node3574;
	wire [8-1:0] node3575;
	wire [8-1:0] node3579;
	wire [8-1:0] node3581;
	wire [8-1:0] node3584;
	wire [8-1:0] node3585;
	wire [8-1:0] node3589;
	wire [8-1:0] node3590;
	wire [8-1:0] node3591;
	wire [8-1:0] node3595;
	wire [8-1:0] node3596;
	wire [8-1:0] node3597;
	wire [8-1:0] node3600;
	wire [8-1:0] node3603;
	wire [8-1:0] node3606;
	wire [8-1:0] node3607;
	wire [8-1:0] node3608;
	wire [8-1:0] node3609;
	wire [8-1:0] node3613;
	wire [8-1:0] node3614;
	wire [8-1:0] node3618;
	wire [8-1:0] node3619;
	wire [8-1:0] node3620;
	wire [8-1:0] node3624;
	wire [8-1:0] node3627;
	wire [8-1:0] node3628;
	wire [8-1:0] node3629;
	wire [8-1:0] node3630;
	wire [8-1:0] node3631;
	wire [8-1:0] node3634;
	wire [8-1:0] node3636;
	wire [8-1:0] node3639;
	wire [8-1:0] node3640;
	wire [8-1:0] node3641;
	wire [8-1:0] node3643;
	wire [8-1:0] node3646;
	wire [8-1:0] node3647;
	wire [8-1:0] node3651;
	wire [8-1:0] node3654;
	wire [8-1:0] node3655;
	wire [8-1:0] node3656;
	wire [8-1:0] node3658;
	wire [8-1:0] node3659;
	wire [8-1:0] node3663;
	wire [8-1:0] node3665;
	wire [8-1:0] node3666;
	wire [8-1:0] node3670;
	wire [8-1:0] node3671;
	wire [8-1:0] node3672;
	wire [8-1:0] node3676;
	wire [8-1:0] node3679;
	wire [8-1:0] node3680;
	wire [8-1:0] node3681;
	wire [8-1:0] node3682;
	wire [8-1:0] node3684;
	wire [8-1:0] node3686;
	wire [8-1:0] node3689;
	wire [8-1:0] node3692;
	wire [8-1:0] node3693;
	wire [8-1:0] node3694;
	wire [8-1:0] node3696;
	wire [8-1:0] node3700;
	wire [8-1:0] node3703;
	wire [8-1:0] node3704;
	wire [8-1:0] node3705;
	wire [8-1:0] node3706;
	wire [8-1:0] node3708;
	wire [8-1:0] node3711;
	wire [8-1:0] node3712;
	wire [8-1:0] node3716;
	wire [8-1:0] node3717;
	wire [8-1:0] node3720;
	wire [8-1:0] node3723;
	wire [8-1:0] node3724;
	wire [8-1:0] node3727;
	wire [8-1:0] node3730;
	wire [8-1:0] node3731;
	wire [8-1:0] node3732;
	wire [8-1:0] node3733;
	wire [8-1:0] node3734;
	wire [8-1:0] node3736;
	wire [8-1:0] node3737;
	wire [8-1:0] node3741;
	wire [8-1:0] node3742;
	wire [8-1:0] node3744;
	wire [8-1:0] node3747;
	wire [8-1:0] node3748;
	wire [8-1:0] node3749;
	wire [8-1:0] node3752;
	wire [8-1:0] node3756;
	wire [8-1:0] node3757;
	wire [8-1:0] node3758;
	wire [8-1:0] node3759;
	wire [8-1:0] node3760;
	wire [8-1:0] node3761;
	wire [8-1:0] node3764;
	wire [8-1:0] node3766;
	wire [8-1:0] node3769;
	wire [8-1:0] node3770;
	wire [8-1:0] node3771;
	wire [8-1:0] node3774;
	wire [8-1:0] node3777;
	wire [8-1:0] node3779;
	wire [8-1:0] node3782;
	wire [8-1:0] node3783;
	wire [8-1:0] node3786;
	wire [8-1:0] node3788;
	wire [8-1:0] node3790;
	wire [8-1:0] node3793;
	wire [8-1:0] node3794;
	wire [8-1:0] node3795;
	wire [8-1:0] node3796;
	wire [8-1:0] node3800;
	wire [8-1:0] node3803;
	wire [8-1:0] node3804;
	wire [8-1:0] node3808;
	wire [8-1:0] node3809;
	wire [8-1:0] node3810;
	wire [8-1:0] node3811;
	wire [8-1:0] node3812;
	wire [8-1:0] node3817;
	wire [8-1:0] node3818;
	wire [8-1:0] node3819;
	wire [8-1:0] node3822;
	wire [8-1:0] node3825;
	wire [8-1:0] node3826;
	wire [8-1:0] node3830;
	wire [8-1:0] node3831;
	wire [8-1:0] node3833;
	wire [8-1:0] node3837;
	wire [8-1:0] node3838;
	wire [8-1:0] node3839;
	wire [8-1:0] node3840;
	wire [8-1:0] node3841;
	wire [8-1:0] node3845;
	wire [8-1:0] node3846;
	wire [8-1:0] node3847;
	wire [8-1:0] node3850;
	wire [8-1:0] node3854;
	wire [8-1:0] node3855;
	wire [8-1:0] node3856;
	wire [8-1:0] node3857;
	wire [8-1:0] node3861;
	wire [8-1:0] node3862;
	wire [8-1:0] node3866;
	wire [8-1:0] node3867;
	wire [8-1:0] node3868;
	wire [8-1:0] node3870;
	wire [8-1:0] node3874;
	wire [8-1:0] node3876;
	wire [8-1:0] node3877;
	wire [8-1:0] node3881;
	wire [8-1:0] node3882;
	wire [8-1:0] node3883;
	wire [8-1:0] node3884;
	wire [8-1:0] node3886;
	wire [8-1:0] node3887;
	wire [8-1:0] node3890;
	wire [8-1:0] node3892;
	wire [8-1:0] node3895;
	wire [8-1:0] node3897;
	wire [8-1:0] node3898;
	wire [8-1:0] node3902;
	wire [8-1:0] node3903;
	wire [8-1:0] node3905;
	wire [8-1:0] node3906;
	wire [8-1:0] node3907;
	wire [8-1:0] node3910;
	wire [8-1:0] node3913;
	wire [8-1:0] node3914;
	wire [8-1:0] node3918;
	wire [8-1:0] node3920;
	wire [8-1:0] node3921;
	wire [8-1:0] node3924;
	wire [8-1:0] node3927;
	wire [8-1:0] node3928;
	wire [8-1:0] node3930;
	wire [8-1:0] node3934;
	wire [8-1:0] node3935;
	wire [8-1:0] node3936;
	wire [8-1:0] node3937;
	wire [8-1:0] node3938;
	wire [8-1:0] node3939;
	wire [8-1:0] node3940;
	wire [8-1:0] node3944;
	wire [8-1:0] node3945;
	wire [8-1:0] node3946;
	wire [8-1:0] node3950;
	wire [8-1:0] node3951;
	wire [8-1:0] node3955;
	wire [8-1:0] node3956;
	wire [8-1:0] node3957;
	wire [8-1:0] node3959;
	wire [8-1:0] node3962;
	wire [8-1:0] node3964;
	wire [8-1:0] node3967;
	wire [8-1:0] node3969;
	wire [8-1:0] node3970;
	wire [8-1:0] node3973;
	wire [8-1:0] node3976;
	wire [8-1:0] node3977;
	wire [8-1:0] node3978;
	wire [8-1:0] node3979;
	wire [8-1:0] node3981;
	wire [8-1:0] node3984;
	wire [8-1:0] node3985;
	wire [8-1:0] node3989;
	wire [8-1:0] node3990;
	wire [8-1:0] node3991;
	wire [8-1:0] node3995;
	wire [8-1:0] node3996;
	wire [8-1:0] node3998;
	wire [8-1:0] node4001;
	wire [8-1:0] node4003;
	wire [8-1:0] node4006;
	wire [8-1:0] node4007;
	wire [8-1:0] node4008;
	wire [8-1:0] node4011;
	wire [8-1:0] node4014;
	wire [8-1:0] node4015;
	wire [8-1:0] node4017;
	wire [8-1:0] node4020;
	wire [8-1:0] node4022;
	wire [8-1:0] node4025;
	wire [8-1:0] node4026;
	wire [8-1:0] node4027;
	wire [8-1:0] node4028;
	wire [8-1:0] node4029;
	wire [8-1:0] node4032;
	wire [8-1:0] node4035;
	wire [8-1:0] node4036;
	wire [8-1:0] node4039;
	wire [8-1:0] node4042;
	wire [8-1:0] node4043;
	wire [8-1:0] node4044;
	wire [8-1:0] node4046;
	wire [8-1:0] node4049;
	wire [8-1:0] node4051;
	wire [8-1:0] node4054;
	wire [8-1:0] node4055;
	wire [8-1:0] node4057;
	wire [8-1:0] node4060;
	wire [8-1:0] node4063;
	wire [8-1:0] node4064;
	wire [8-1:0] node4065;
	wire [8-1:0] node4066;
	wire [8-1:0] node4068;
	wire [8-1:0] node4071;
	wire [8-1:0] node4072;
	wire [8-1:0] node4075;
	wire [8-1:0] node4076;
	wire [8-1:0] node4079;
	wire [8-1:0] node4082;
	wire [8-1:0] node4083;
	wire [8-1:0] node4084;
	wire [8-1:0] node4087;
	wire [8-1:0] node4090;
	wire [8-1:0] node4093;
	wire [8-1:0] node4094;
	wire [8-1:0] node4096;
	wire [8-1:0] node4097;
	wire [8-1:0] node4100;
	wire [8-1:0] node4103;
	wire [8-1:0] node4104;
	wire [8-1:0] node4105;
	wire [8-1:0] node4106;
	wire [8-1:0] node4109;
	wire [8-1:0] node4112;
	wire [8-1:0] node4115;
	wire [8-1:0] node4118;
	wire [8-1:0] node4119;
	wire [8-1:0] node4120;
	wire [8-1:0] node4121;
	wire [8-1:0] node4122;
	wire [8-1:0] node4123;
	wire [8-1:0] node4125;
	wire [8-1:0] node4128;
	wire [8-1:0] node4130;
	wire [8-1:0] node4132;
	wire [8-1:0] node4135;
	wire [8-1:0] node4137;
	wire [8-1:0] node4139;
	wire [8-1:0] node4140;
	wire [8-1:0] node4144;
	wire [8-1:0] node4145;
	wire [8-1:0] node4146;
	wire [8-1:0] node4150;
	wire [8-1:0] node4151;
	wire [8-1:0] node4155;
	wire [8-1:0] node4156;
	wire [8-1:0] node4157;
	wire [8-1:0] node4158;
	wire [8-1:0] node4161;
	wire [8-1:0] node4162;
	wire [8-1:0] node4166;
	wire [8-1:0] node4167;
	wire [8-1:0] node4171;
	wire [8-1:0] node4172;
	wire [8-1:0] node4173;
	wire [8-1:0] node4175;
	wire [8-1:0] node4176;
	wire [8-1:0] node4180;
	wire [8-1:0] node4181;
	wire [8-1:0] node4183;
	wire [8-1:0] node4187;
	wire [8-1:0] node4188;
	wire [8-1:0] node4189;
	wire [8-1:0] node4193;
	wire [8-1:0] node4196;
	wire [8-1:0] node4197;
	wire [8-1:0] node4198;
	wire [8-1:0] node4199;
	wire [8-1:0] node4201;
	wire [8-1:0] node4204;
	wire [8-1:0] node4205;
	wire [8-1:0] node4206;
	wire [8-1:0] node4208;
	wire [8-1:0] node4212;
	wire [8-1:0] node4214;
	wire [8-1:0] node4217;
	wire [8-1:0] node4218;
	wire [8-1:0] node4219;
	wire [8-1:0] node4220;
	wire [8-1:0] node4224;
	wire [8-1:0] node4225;
	wire [8-1:0] node4228;
	wire [8-1:0] node4231;
	wire [8-1:0] node4232;
	wire [8-1:0] node4233;
	wire [8-1:0] node4237;
	wire [8-1:0] node4238;
	wire [8-1:0] node4242;
	wire [8-1:0] node4243;
	wire [8-1:0] node4244;
	wire [8-1:0] node4246;
	wire [8-1:0] node4247;
	wire [8-1:0] node4250;
	wire [8-1:0] node4253;
	wire [8-1:0] node4254;
	wire [8-1:0] node4256;
	wire [8-1:0] node4259;
	wire [8-1:0] node4260;
	wire [8-1:0] node4263;
	wire [8-1:0] node4265;
	wire [8-1:0] node4268;
	wire [8-1:0] node4269;
	wire [8-1:0] node4270;
	wire [8-1:0] node4274;
	wire [8-1:0] node4277;
	wire [8-1:0] node4278;
	wire [8-1:0] node4279;
	wire [8-1:0] node4280;
	wire [8-1:0] node4281;
	wire [8-1:0] node4282;
	wire [8-1:0] node4283;
	wire [8-1:0] node4285;
	wire [8-1:0] node4288;
	wire [8-1:0] node4289;
	wire [8-1:0] node4291;
	wire [8-1:0] node4294;
	wire [8-1:0] node4296;
	wire [8-1:0] node4299;
	wire [8-1:0] node4300;
	wire [8-1:0] node4301;
	wire [8-1:0] node4302;
	wire [8-1:0] node4305;
	wire [8-1:0] node4307;
	wire [8-1:0] node4310;
	wire [8-1:0] node4311;
	wire [8-1:0] node4315;
	wire [8-1:0] node4316;
	wire [8-1:0] node4317;
	wire [8-1:0] node4319;
	wire [8-1:0] node4323;
	wire [8-1:0] node4325;
	wire [8-1:0] node4328;
	wire [8-1:0] node4329;
	wire [8-1:0] node4330;
	wire [8-1:0] node4332;
	wire [8-1:0] node4335;
	wire [8-1:0] node4336;
	wire [8-1:0] node4337;
	wire [8-1:0] node4341;
	wire [8-1:0] node4342;
	wire [8-1:0] node4346;
	wire [8-1:0] node4347;
	wire [8-1:0] node4348;
	wire [8-1:0] node4349;
	wire [8-1:0] node4350;
	wire [8-1:0] node4355;
	wire [8-1:0] node4356;
	wire [8-1:0] node4360;
	wire [8-1:0] node4361;
	wire [8-1:0] node4363;
	wire [8-1:0] node4366;
	wire [8-1:0] node4368;
	wire [8-1:0] node4371;
	wire [8-1:0] node4372;
	wire [8-1:0] node4373;
	wire [8-1:0] node4374;
	wire [8-1:0] node4375;
	wire [8-1:0] node4376;
	wire [8-1:0] node4381;
	wire [8-1:0] node4382;
	wire [8-1:0] node4386;
	wire [8-1:0] node4387;
	wire [8-1:0] node4389;
	wire [8-1:0] node4392;
	wire [8-1:0] node4394;
	wire [8-1:0] node4397;
	wire [8-1:0] node4398;
	wire [8-1:0] node4399;
	wire [8-1:0] node4401;
	wire [8-1:0] node4404;
	wire [8-1:0] node4405;
	wire [8-1:0] node4409;
	wire [8-1:0] node4410;
	wire [8-1:0] node4414;
	wire [8-1:0] node4415;
	wire [8-1:0] node4416;
	wire [8-1:0] node4417;
	wire [8-1:0] node4418;
	wire [8-1:0] node4419;
	wire [8-1:0] node4420;
	wire [8-1:0] node4422;
	wire [8-1:0] node4425;
	wire [8-1:0] node4426;
	wire [8-1:0] node4430;
	wire [8-1:0] node4432;
	wire [8-1:0] node4434;
	wire [8-1:0] node4435;
	wire [8-1:0] node4438;
	wire [8-1:0] node4441;
	wire [8-1:0] node4442;
	wire [8-1:0] node4443;
	wire [8-1:0] node4444;
	wire [8-1:0] node4449;
	wire [8-1:0] node4450;
	wire [8-1:0] node4451;
	wire [8-1:0] node4454;
	wire [8-1:0] node4457;
	wire [8-1:0] node4458;
	wire [8-1:0] node4462;
	wire [8-1:0] node4463;
	wire [8-1:0] node4464;
	wire [8-1:0] node4465;
	wire [8-1:0] node4467;
	wire [8-1:0] node4468;
	wire [8-1:0] node4472;
	wire [8-1:0] node4474;
	wire [8-1:0] node4477;
	wire [8-1:0] node4478;
	wire [8-1:0] node4479;
	wire [8-1:0] node4481;
	wire [8-1:0] node4484;
	wire [8-1:0] node4485;
	wire [8-1:0] node4488;
	wire [8-1:0] node4491;
	wire [8-1:0] node4493;
	wire [8-1:0] node4496;
	wire [8-1:0] node4497;
	wire [8-1:0] node4498;
	wire [8-1:0] node4500;
	wire [8-1:0] node4501;
	wire [8-1:0] node4504;
	wire [8-1:0] node4508;
	wire [8-1:0] node4509;
	wire [8-1:0] node4511;
	wire [8-1:0] node4514;
	wire [8-1:0] node4515;
	wire [8-1:0] node4518;
	wire [8-1:0] node4521;
	wire [8-1:0] node4522;
	wire [8-1:0] node4523;
	wire [8-1:0] node4524;
	wire [8-1:0] node4525;
	wire [8-1:0] node4526;
	wire [8-1:0] node4529;
	wire [8-1:0] node4532;
	wire [8-1:0] node4533;
	wire [8-1:0] node4537;
	wire [8-1:0] node4538;
	wire [8-1:0] node4541;
	wire [8-1:0] node4542;
	wire [8-1:0] node4543;
	wire [8-1:0] node4546;
	wire [8-1:0] node4549;
	wire [8-1:0] node4550;
	wire [8-1:0] node4554;
	wire [8-1:0] node4555;
	wire [8-1:0] node4556;
	wire [8-1:0] node4558;
	wire [8-1:0] node4560;
	wire [8-1:0] node4563;
	wire [8-1:0] node4565;
	wire [8-1:0] node4568;
	wire [8-1:0] node4570;
	wire [8-1:0] node4571;
	wire [8-1:0] node4573;
	wire [8-1:0] node4576;
	wire [8-1:0] node4578;
	wire [8-1:0] node4581;
	wire [8-1:0] node4582;
	wire [8-1:0] node4583;
	wire [8-1:0] node4584;
	wire [8-1:0] node4585;
	wire [8-1:0] node4586;
	wire [8-1:0] node4589;
	wire [8-1:0] node4592;
	wire [8-1:0] node4595;
	wire [8-1:0] node4596;
	wire [8-1:0] node4599;
	wire [8-1:0] node4602;
	wire [8-1:0] node4603;
	wire [8-1:0] node4605;
	wire [8-1:0] node4608;
	wire [8-1:0] node4609;
	wire [8-1:0] node4610;
	wire [8-1:0] node4615;
	wire [8-1:0] node4616;
	wire [8-1:0] node4617;
	wire [8-1:0] node4618;
	wire [8-1:0] node4619;
	wire [8-1:0] node4623;
	wire [8-1:0] node4626;
	wire [8-1:0] node4628;
	wire [8-1:0] node4629;
	wire [8-1:0] node4633;
	wire [8-1:0] node4634;
	wire [8-1:0] node4636;
	wire [8-1:0] node4638;
	wire [8-1:0] node4641;
	wire [8-1:0] node4643;
	wire [8-1:0] node4646;
	wire [8-1:0] node4647;
	wire [8-1:0] node4648;
	wire [8-1:0] node4649;
	wire [8-1:0] node4650;
	wire [8-1:0] node4651;
	wire [8-1:0] node4654;
	wire [8-1:0] node4657;
	wire [8-1:0] node4658;
	wire [8-1:0] node4660;
	wire [8-1:0] node4663;
	wire [8-1:0] node4666;
	wire [8-1:0] node4667;
	wire [8-1:0] node4668;
	wire [8-1:0] node4669;
	wire [8-1:0] node4673;
	wire [8-1:0] node4676;
	wire [8-1:0] node4678;
	wire [8-1:0] node4679;
	wire [8-1:0] node4681;
	wire [8-1:0] node4684;
	wire [8-1:0] node4687;
	wire [8-1:0] node4688;
	wire [8-1:0] node4689;
	wire [8-1:0] node4690;
	wire [8-1:0] node4691;
	wire [8-1:0] node4692;
	wire [8-1:0] node4696;
	wire [8-1:0] node4697;
	wire [8-1:0] node4701;
	wire [8-1:0] node4702;
	wire [8-1:0] node4705;
	wire [8-1:0] node4708;
	wire [8-1:0] node4709;
	wire [8-1:0] node4710;
	wire [8-1:0] node4712;
	wire [8-1:0] node4715;
	wire [8-1:0] node4716;
	wire [8-1:0] node4720;
	wire [8-1:0] node4721;
	wire [8-1:0] node4722;
	wire [8-1:0] node4727;
	wire [8-1:0] node4728;
	wire [8-1:0] node4729;
	wire [8-1:0] node4730;
	wire [8-1:0] node4732;
	wire [8-1:0] node4736;
	wire [8-1:0] node4737;
	wire [8-1:0] node4738;
	wire [8-1:0] node4741;
	wire [8-1:0] node4744;
	wire [8-1:0] node4746;
	wire [8-1:0] node4749;
	wire [8-1:0] node4750;
	wire [8-1:0] node4752;
	wire [8-1:0] node4755;
	wire [8-1:0] node4756;
	wire [8-1:0] node4758;
	wire [8-1:0] node4761;
	wire [8-1:0] node4764;
	wire [8-1:0] node4765;
	wire [8-1:0] node4766;
	wire [8-1:0] node4767;
	wire [8-1:0] node4768;
	wire [8-1:0] node4771;
	wire [8-1:0] node4772;
	wire [8-1:0] node4774;
	wire [8-1:0] node4777;
	wire [8-1:0] node4778;
	wire [8-1:0] node4782;
	wire [8-1:0] node4784;
	wire [8-1:0] node4785;
	wire [8-1:0] node4788;
	wire [8-1:0] node4791;
	wire [8-1:0] node4792;
	wire [8-1:0] node4794;
	wire [8-1:0] node4797;
	wire [8-1:0] node4799;
	wire [8-1:0] node4802;
	wire [8-1:0] node4803;
	wire [8-1:0] node4804;
	wire [8-1:0] node4805;
	wire [8-1:0] node4806;
	wire [8-1:0] node4809;
	wire [8-1:0] node4812;
	wire [8-1:0] node4813;
	wire [8-1:0] node4815;
	wire [8-1:0] node4818;
	wire [8-1:0] node4821;
	wire [8-1:0] node4822;
	wire [8-1:0] node4823;
	wire [8-1:0] node4826;
	wire [8-1:0] node4829;
	wire [8-1:0] node4832;
	wire [8-1:0] node4833;
	wire [8-1:0] node4834;
	wire [8-1:0] node4836;
	wire [8-1:0] node4839;
	wire [8-1:0] node4841;
	wire [8-1:0] node4844;
	wire [8-1:0] node4845;
	wire [8-1:0] node4847;
	wire [8-1:0] node4848;
	wire [8-1:0] node4852;
	wire [8-1:0] node4855;
	wire [8-1:0] node4856;
	wire [8-1:0] node4857;
	wire [8-1:0] node4858;
	wire [8-1:0] node4859;
	wire [8-1:0] node4860;
	wire [8-1:0] node4861;
	wire [8-1:0] node4864;
	wire [8-1:0] node4867;
	wire [8-1:0] node4869;
	wire [8-1:0] node4872;
	wire [8-1:0] node4873;
	wire [8-1:0] node4874;
	wire [8-1:0] node4875;
	wire [8-1:0] node4879;
	wire [8-1:0] node4880;
	wire [8-1:0] node4884;
	wire [8-1:0] node4885;
	wire [8-1:0] node4886;
	wire [8-1:0] node4890;
	wire [8-1:0] node4893;
	wire [8-1:0] node4894;
	wire [8-1:0] node4895;
	wire [8-1:0] node4896;
	wire [8-1:0] node4899;
	wire [8-1:0] node4901;
	wire [8-1:0] node4904;
	wire [8-1:0] node4905;
	wire [8-1:0] node4908;
	wire [8-1:0] node4910;
	wire [8-1:0] node4913;
	wire [8-1:0] node4914;
	wire [8-1:0] node4915;
	wire [8-1:0] node4916;
	wire [8-1:0] node4920;
	wire [8-1:0] node4921;
	wire [8-1:0] node4924;
	wire [8-1:0] node4927;
	wire [8-1:0] node4928;
	wire [8-1:0] node4929;
	wire [8-1:0] node4932;
	wire [8-1:0] node4936;
	wire [8-1:0] node4937;
	wire [8-1:0] node4938;
	wire [8-1:0] node4939;
	wire [8-1:0] node4940;
	wire [8-1:0] node4943;
	wire [8-1:0] node4945;
	wire [8-1:0] node4948;
	wire [8-1:0] node4949;
	wire [8-1:0] node4952;
	wire [8-1:0] node4954;
	wire [8-1:0] node4957;
	wire [8-1:0] node4958;
	wire [8-1:0] node4959;
	wire [8-1:0] node4960;
	wire [8-1:0] node4964;
	wire [8-1:0] node4965;
	wire [8-1:0] node4969;
	wire [8-1:0] node4970;
	wire [8-1:0] node4971;
	wire [8-1:0] node4975;
	wire [8-1:0] node4978;
	wire [8-1:0] node4979;
	wire [8-1:0] node4980;
	wire [8-1:0] node4981;
	wire [8-1:0] node4983;
	wire [8-1:0] node4986;
	wire [8-1:0] node4988;
	wire [8-1:0] node4991;
	wire [8-1:0] node4993;
	wire [8-1:0] node4995;
	wire [8-1:0] node4998;
	wire [8-1:0] node4999;
	wire [8-1:0] node5000;
	wire [8-1:0] node5002;
	wire [8-1:0] node5005;
	wire [8-1:0] node5007;
	wire [8-1:0] node5010;
	wire [8-1:0] node5012;
	wire [8-1:0] node5014;
	wire [8-1:0] node5017;
	wire [8-1:0] node5018;
	wire [8-1:0] node5019;
	wire [8-1:0] node5020;
	wire [8-1:0] node5021;
	wire [8-1:0] node5022;
	wire [8-1:0] node5023;
	wire [8-1:0] node5024;
	wire [8-1:0] node5028;
	wire [8-1:0] node5030;
	wire [8-1:0] node5033;
	wire [8-1:0] node5034;
	wire [8-1:0] node5036;
	wire [8-1:0] node5039;
	wire [8-1:0] node5041;
	wire [8-1:0] node5044;
	wire [8-1:0] node5045;
	wire [8-1:0] node5046;
	wire [8-1:0] node5049;
	wire [8-1:0] node5050;
	wire [8-1:0] node5051;
	wire [8-1:0] node5054;
	wire [8-1:0] node5058;
	wire [8-1:0] node5059;
	wire [8-1:0] node5060;
	wire [8-1:0] node5064;
	wire [8-1:0] node5067;
	wire [8-1:0] node5068;
	wire [8-1:0] node5069;
	wire [8-1:0] node5070;
	wire [8-1:0] node5071;
	wire [8-1:0] node5072;
	wire [8-1:0] node5076;
	wire [8-1:0] node5077;
	wire [8-1:0] node5080;
	wire [8-1:0] node5083;
	wire [8-1:0] node5084;
	wire [8-1:0] node5087;
	wire [8-1:0] node5090;
	wire [8-1:0] node5092;
	wire [8-1:0] node5093;
	wire [8-1:0] node5095;
	wire [8-1:0] node5099;
	wire [8-1:0] node5100;
	wire [8-1:0] node5101;
	wire [8-1:0] node5104;
	wire [8-1:0] node5107;
	wire [8-1:0] node5110;
	wire [8-1:0] node5111;
	wire [8-1:0] node5112;
	wire [8-1:0] node5113;
	wire [8-1:0] node5114;
	wire [8-1:0] node5115;
	wire [8-1:0] node5118;
	wire [8-1:0] node5121;
	wire [8-1:0] node5123;
	wire [8-1:0] node5124;
	wire [8-1:0] node5128;
	wire [8-1:0] node5130;
	wire [8-1:0] node5131;
	wire [8-1:0] node5134;
	wire [8-1:0] node5137;
	wire [8-1:0] node5138;
	wire [8-1:0] node5139;
	wire [8-1:0] node5141;
	wire [8-1:0] node5142;
	wire [8-1:0] node5146;
	wire [8-1:0] node5147;
	wire [8-1:0] node5148;
	wire [8-1:0] node5153;
	wire [8-1:0] node5154;
	wire [8-1:0] node5155;
	wire [8-1:0] node5157;
	wire [8-1:0] node5160;
	wire [8-1:0] node5161;
	wire [8-1:0] node5165;
	wire [8-1:0] node5166;
	wire [8-1:0] node5167;
	wire [8-1:0] node5172;
	wire [8-1:0] node5173;
	wire [8-1:0] node5174;
	wire [8-1:0] node5175;
	wire [8-1:0] node5176;
	wire [8-1:0] node5177;
	wire [8-1:0] node5182;
	wire [8-1:0] node5185;
	wire [8-1:0] node5186;
	wire [8-1:0] node5189;
	wire [8-1:0] node5192;
	wire [8-1:0] node5193;
	wire [8-1:0] node5194;
	wire [8-1:0] node5197;
	wire [8-1:0] node5200;
	wire [8-1:0] node5203;
	wire [8-1:0] node5204;
	wire [8-1:0] node5205;
	wire [8-1:0] node5206;
	wire [8-1:0] node5207;
	wire [8-1:0] node5208;
	wire [8-1:0] node5212;
	wire [8-1:0] node5213;
	wire [8-1:0] node5216;
	wire [8-1:0] node5219;
	wire [8-1:0] node5220;
	wire [8-1:0] node5221;
	wire [8-1:0] node5223;
	wire [8-1:0] node5226;
	wire [8-1:0] node5227;
	wire [8-1:0] node5231;
	wire [8-1:0] node5232;
	wire [8-1:0] node5233;
	wire [8-1:0] node5234;
	wire [8-1:0] node5238;
	wire [8-1:0] node5242;
	wire [8-1:0] node5243;
	wire [8-1:0] node5244;
	wire [8-1:0] node5245;
	wire [8-1:0] node5246;
	wire [8-1:0] node5249;
	wire [8-1:0] node5252;
	wire [8-1:0] node5255;
	wire [8-1:0] node5256;
	wire [8-1:0] node5257;
	wire [8-1:0] node5259;
	wire [8-1:0] node5262;
	wire [8-1:0] node5265;
	wire [8-1:0] node5268;
	wire [8-1:0] node5269;
	wire [8-1:0] node5270;
	wire [8-1:0] node5271;
	wire [8-1:0] node5274;
	wire [8-1:0] node5277;
	wire [8-1:0] node5280;
	wire [8-1:0] node5281;
	wire [8-1:0] node5282;
	wire [8-1:0] node5285;
	wire [8-1:0] node5286;
	wire [8-1:0] node5290;
	wire [8-1:0] node5291;
	wire [8-1:0] node5294;
	wire [8-1:0] node5297;
	wire [8-1:0] node5298;
	wire [8-1:0] node5299;
	wire [8-1:0] node5300;
	wire [8-1:0] node5301;
	wire [8-1:0] node5302;
	wire [8-1:0] node5305;
	wire [8-1:0] node5308;
	wire [8-1:0] node5309;
	wire [8-1:0] node5313;
	wire [8-1:0] node5314;
	wire [8-1:0] node5315;
	wire [8-1:0] node5318;
	wire [8-1:0] node5321;
	wire [8-1:0] node5322;
	wire [8-1:0] node5325;
	wire [8-1:0] node5328;
	wire [8-1:0] node5329;
	wire [8-1:0] node5332;
	wire [8-1:0] node5335;
	wire [8-1:0] node5336;
	wire [8-1:0] node5337;
	wire [8-1:0] node5339;
	wire [8-1:0] node5342;
	wire [8-1:0] node5345;
	wire [8-1:0] node5346;
	wire [8-1:0] node5347;
	wire [8-1:0] node5348;
	wire [8-1:0] node5350;
	wire [8-1:0] node5353;
	wire [8-1:0] node5357;
	wire [8-1:0] node5358;
	wire [8-1:0] node5362;
	wire [8-1:0] node5363;
	wire [8-1:0] node5364;
	wire [8-1:0] node5365;
	wire [8-1:0] node5367;
	wire [8-1:0] node5368;
	wire [8-1:0] node5369;
	wire [8-1:0] node5370;
	wire [8-1:0] node5371;
	wire [8-1:0] node5372;
	wire [8-1:0] node5377;
	wire [8-1:0] node5379;
	wire [8-1:0] node5382;
	wire [8-1:0] node5383;
	wire [8-1:0] node5384;
	wire [8-1:0] node5386;
	wire [8-1:0] node5389;
	wire [8-1:0] node5391;
	wire [8-1:0] node5394;
	wire [8-1:0] node5395;
	wire [8-1:0] node5397;
	wire [8-1:0] node5400;
	wire [8-1:0] node5401;
	wire [8-1:0] node5403;
	wire [8-1:0] node5407;
	wire [8-1:0] node5408;
	wire [8-1:0] node5409;
	wire [8-1:0] node5410;
	wire [8-1:0] node5411;
	wire [8-1:0] node5414;
	wire [8-1:0] node5417;
	wire [8-1:0] node5419;
	wire [8-1:0] node5422;
	wire [8-1:0] node5424;
	wire [8-1:0] node5425;
	wire [8-1:0] node5427;
	wire [8-1:0] node5430;
	wire [8-1:0] node5433;
	wire [8-1:0] node5434;
	wire [8-1:0] node5435;
	wire [8-1:0] node5436;
	wire [8-1:0] node5441;
	wire [8-1:0] node5442;
	wire [8-1:0] node5446;
	wire [8-1:0] node5447;
	wire [8-1:0] node5448;
	wire [8-1:0] node5449;
	wire [8-1:0] node5451;
	wire [8-1:0] node5452;
	wire [8-1:0] node5456;
	wire [8-1:0] node5457;
	wire [8-1:0] node5458;
	wire [8-1:0] node5462;
	wire [8-1:0] node5463;
	wire [8-1:0] node5464;
	wire [8-1:0] node5469;
	wire [8-1:0] node5470;
	wire [8-1:0] node5471;
	wire [8-1:0] node5472;
	wire [8-1:0] node5476;
	wire [8-1:0] node5477;
	wire [8-1:0] node5478;
	wire [8-1:0] node5481;
	wire [8-1:0] node5485;
	wire [8-1:0] node5486;
	wire [8-1:0] node5487;
	wire [8-1:0] node5488;
	wire [8-1:0] node5491;
	wire [8-1:0] node5495;
	wire [8-1:0] node5496;
	wire [8-1:0] node5498;
	wire [8-1:0] node5502;
	wire [8-1:0] node5503;
	wire [8-1:0] node5504;
	wire [8-1:0] node5505;
	wire [8-1:0] node5506;
	wire [8-1:0] node5510;
	wire [8-1:0] node5511;
	wire [8-1:0] node5513;
	wire [8-1:0] node5517;
	wire [8-1:0] node5518;
	wire [8-1:0] node5519;
	wire [8-1:0] node5520;
	wire [8-1:0] node5523;
	wire [8-1:0] node5526;
	wire [8-1:0] node5527;
	wire [8-1:0] node5529;
	wire [8-1:0] node5532;
	wire [8-1:0] node5535;
	wire [8-1:0] node5538;
	wire [8-1:0] node5539;
	wire [8-1:0] node5540;
	wire [8-1:0] node5541;
	wire [8-1:0] node5544;
	wire [8-1:0] node5545;
	wire [8-1:0] node5549;
	wire [8-1:0] node5550;
	wire [8-1:0] node5551;
	wire [8-1:0] node5554;
	wire [8-1:0] node5555;
	wire [8-1:0] node5558;
	wire [8-1:0] node5562;
	wire [8-1:0] node5563;
	wire [8-1:0] node5564;
	wire [8-1:0] node5565;
	wire [8-1:0] node5568;
	wire [8-1:0] node5569;
	wire [8-1:0] node5574;
	wire [8-1:0] node5575;
	wire [8-1:0] node5576;
	wire [8-1:0] node5578;
	wire [8-1:0] node5581;
	wire [8-1:0] node5582;
	wire [8-1:0] node5585;
	wire [8-1:0] node5589;
	wire [8-1:0] node5590;
	wire [8-1:0] node5592;
	wire [8-1:0] node5593;
	wire [8-1:0] node5594;
	wire [8-1:0] node5595;
	wire [8-1:0] node5597;
	wire [8-1:0] node5600;
	wire [8-1:0] node5601;
	wire [8-1:0] node5603;
	wire [8-1:0] node5606;
	wire [8-1:0] node5608;
	wire [8-1:0] node5611;
	wire [8-1:0] node5612;
	wire [8-1:0] node5614;
	wire [8-1:0] node5615;
	wire [8-1:0] node5617;
	wire [8-1:0] node5620;
	wire [8-1:0] node5622;
	wire [8-1:0] node5625;
	wire [8-1:0] node5626;
	wire [8-1:0] node5628;
	wire [8-1:0] node5631;
	wire [8-1:0] node5634;
	wire [8-1:0] node5635;
	wire [8-1:0] node5636;
	wire [8-1:0] node5637;
	wire [8-1:0] node5639;
	wire [8-1:0] node5642;
	wire [8-1:0] node5643;
	wire [8-1:0] node5645;
	wire [8-1:0] node5648;
	wire [8-1:0] node5650;
	wire [8-1:0] node5653;
	wire [8-1:0] node5654;
	wire [8-1:0] node5657;
	wire [8-1:0] node5658;
	wire [8-1:0] node5660;
	wire [8-1:0] node5663;
	wire [8-1:0] node5666;
	wire [8-1:0] node5667;
	wire [8-1:0] node5668;
	wire [8-1:0] node5670;
	wire [8-1:0] node5673;
	wire [8-1:0] node5676;
	wire [8-1:0] node5677;
	wire [8-1:0] node5678;
	wire [8-1:0] node5680;
	wire [8-1:0] node5684;
	wire [8-1:0] node5685;
	wire [8-1:0] node5687;
	wire [8-1:0] node5690;
	wire [8-1:0] node5693;
	wire [8-1:0] node5694;
	wire [8-1:0] node5695;
	wire [8-1:0] node5696;
	wire [8-1:0] node5698;
	wire [8-1:0] node5700;
	wire [8-1:0] node5703;
	wire [8-1:0] node5704;
	wire [8-1:0] node5706;
	wire [8-1:0] node5707;
	wire [8-1:0] node5711;
	wire [8-1:0] node5712;
	wire [8-1:0] node5714;
	wire [8-1:0] node5717;
	wire [8-1:0] node5720;
	wire [8-1:0] node5721;
	wire [8-1:0] node5722;
	wire [8-1:0] node5723;
	wire [8-1:0] node5724;
	wire [8-1:0] node5728;
	wire [8-1:0] node5729;
	wire [8-1:0] node5733;
	wire [8-1:0] node5736;
	wire [8-1:0] node5737;
	wire [8-1:0] node5738;
	wire [8-1:0] node5739;
	wire [8-1:0] node5742;
	wire [8-1:0] node5745;
	wire [8-1:0] node5746;
	wire [8-1:0] node5747;
	wire [8-1:0] node5751;
	wire [8-1:0] node5754;
	wire [8-1:0] node5757;
	wire [8-1:0] node5758;
	wire [8-1:0] node5759;
	wire [8-1:0] node5760;
	wire [8-1:0] node5761;
	wire [8-1:0] node5762;
	wire [8-1:0] node5767;
	wire [8-1:0] node5768;
	wire [8-1:0] node5769;
	wire [8-1:0] node5772;
	wire [8-1:0] node5776;
	wire [8-1:0] node5777;
	wire [8-1:0] node5778;
	wire [8-1:0] node5780;
	wire [8-1:0] node5782;
	wire [8-1:0] node5785;
	wire [8-1:0] node5786;
	wire [8-1:0] node5790;
	wire [8-1:0] node5793;
	wire [8-1:0] node5794;
	wire [8-1:0] node5795;
	wire [8-1:0] node5796;
	wire [8-1:0] node5797;
	wire [8-1:0] node5798;
	wire [8-1:0] node5801;
	wire [8-1:0] node5805;
	wire [8-1:0] node5806;
	wire [8-1:0] node5809;
	wire [8-1:0] node5811;
	wire [8-1:0] node5814;
	wire [8-1:0] node5815;
	wire [8-1:0] node5816;
	wire [8-1:0] node5819;
	wire [8-1:0] node5820;
	wire [8-1:0] node5824;
	wire [8-1:0] node5826;
	wire [8-1:0] node5827;
	wire [8-1:0] node5831;
	wire [8-1:0] node5832;
	wire [8-1:0] node5835;
	wire [8-1:0] node5838;
	wire [8-1:0] node5839;
	wire [8-1:0] node5841;
	wire [8-1:0] node5842;
	wire [8-1:0] node5843;
	wire [8-1:0] node5844;
	wire [8-1:0] node5846;
	wire [8-1:0] node5849;
	wire [8-1:0] node5850;
	wire [8-1:0] node5852;
	wire [8-1:0] node5855;
	wire [8-1:0] node5856;
	wire [8-1:0] node5858;
	wire [8-1:0] node5862;
	wire [8-1:0] node5863;
	wire [8-1:0] node5864;
	wire [8-1:0] node5866;
	wire [8-1:0] node5868;
	wire [8-1:0] node5871;
	wire [8-1:0] node5872;
	wire [8-1:0] node5875;
	wire [8-1:0] node5877;
	wire [8-1:0] node5879;
	wire [8-1:0] node5882;
	wire [8-1:0] node5883;
	wire [8-1:0] node5885;
	wire [8-1:0] node5886;
	wire [8-1:0] node5890;
	wire [8-1:0] node5891;
	wire [8-1:0] node5893;
	wire [8-1:0] node5896;
	wire [8-1:0] node5897;
	wire [8-1:0] node5898;
	wire [8-1:0] node5903;
	wire [8-1:0] node5904;
	wire [8-1:0] node5905;
	wire [8-1:0] node5906;
	wire [8-1:0] node5908;
	wire [8-1:0] node5911;
	wire [8-1:0] node5912;
	wire [8-1:0] node5915;
	wire [8-1:0] node5917;
	wire [8-1:0] node5920;
	wire [8-1:0] node5921;
	wire [8-1:0] node5922;
	wire [8-1:0] node5924;
	wire [8-1:0] node5927;
	wire [8-1:0] node5928;
	wire [8-1:0] node5931;
	wire [8-1:0] node5932;
	wire [8-1:0] node5935;
	wire [8-1:0] node5938;
	wire [8-1:0] node5939;
	wire [8-1:0] node5940;
	wire [8-1:0] node5942;
	wire [8-1:0] node5945;
	wire [8-1:0] node5947;
	wire [8-1:0] node5950;
	wire [8-1:0] node5951;
	wire [8-1:0] node5954;
	wire [8-1:0] node5955;
	wire [8-1:0] node5959;
	wire [8-1:0] node5960;
	wire [8-1:0] node5961;
	wire [8-1:0] node5962;
	wire [8-1:0] node5964;
	wire [8-1:0] node5967;
	wire [8-1:0] node5968;
	wire [8-1:0] node5971;
	wire [8-1:0] node5973;
	wire [8-1:0] node5976;
	wire [8-1:0] node5977;
	wire [8-1:0] node5979;
	wire [8-1:0] node5981;
	wire [8-1:0] node5984;
	wire [8-1:0] node5986;
	wire [8-1:0] node5989;
	wire [8-1:0] node5990;
	wire [8-1:0] node5991;
	wire [8-1:0] node5993;
	wire [8-1:0] node5996;
	wire [8-1:0] node5998;
	wire [8-1:0] node6000;
	wire [8-1:0] node6003;
	wire [8-1:0] node6004;
	wire [8-1:0] node6006;
	wire [8-1:0] node6009;
	wire [8-1:0] node6010;
	wire [8-1:0] node6012;
	wire [8-1:0] node6015;
	wire [8-1:0] node6017;
	wire [8-1:0] node6019;
	wire [8-1:0] node6022;
	wire [8-1:0] node6023;
	wire [8-1:0] node6024;
	wire [8-1:0] node6025;
	wire [8-1:0] node6027;
	wire [8-1:0] node6028;
	wire [8-1:0] node6029;
	wire [8-1:0] node6033;
	wire [8-1:0] node6036;
	wire [8-1:0] node6037;
	wire [8-1:0] node6039;
	wire [8-1:0] node6042;
	wire [8-1:0] node6043;
	wire [8-1:0] node6044;
	wire [8-1:0] node6045;
	wire [8-1:0] node6046;
	wire [8-1:0] node6047;
	wire [8-1:0] node6050;
	wire [8-1:0] node6055;
	wire [8-1:0] node6058;
	wire [8-1:0] node6061;
	wire [8-1:0] node6062;
	wire [8-1:0] node6063;
	wire [8-1:0] node6064;
	wire [8-1:0] node6066;
	wire [8-1:0] node6068;
	wire [8-1:0] node6071;
	wire [8-1:0] node6072;
	wire [8-1:0] node6073;
	wire [8-1:0] node6077;
	wire [8-1:0] node6078;
	wire [8-1:0] node6082;
	wire [8-1:0] node6083;
	wire [8-1:0] node6085;
	wire [8-1:0] node6087;
	wire [8-1:0] node6090;
	wire [8-1:0] node6091;
	wire [8-1:0] node6092;
	wire [8-1:0] node6096;
	wire [8-1:0] node6097;
	wire [8-1:0] node6099;
	wire [8-1:0] node6103;
	wire [8-1:0] node6104;
	wire [8-1:0] node6105;
	wire [8-1:0] node6106;
	wire [8-1:0] node6110;
	wire [8-1:0] node6111;
	wire [8-1:0] node6113;
	wire [8-1:0] node6115;
	wire [8-1:0] node6118;
	wire [8-1:0] node6121;
	wire [8-1:0] node6122;
	wire [8-1:0] node6123;
	wire [8-1:0] node6124;
	wire [8-1:0] node6127;
	wire [8-1:0] node6130;
	wire [8-1:0] node6133;
	wire [8-1:0] node6134;
	wire [8-1:0] node6135;
	wire [8-1:0] node6138;
	wire [8-1:0] node6139;
	wire [8-1:0] node6142;
	wire [8-1:0] node6145;
	wire [8-1:0] node6146;
	wire [8-1:0] node6149;
	wire [8-1:0] node6152;
	wire [8-1:0] node6153;
	wire [8-1:0] node6154;
	wire [8-1:0] node6155;
	wire [8-1:0] node6156;
	wire [8-1:0] node6158;
	wire [8-1:0] node6159;
	wire [8-1:0] node6162;
	wire [8-1:0] node6164;
	wire [8-1:0] node6167;
	wire [8-1:0] node6168;
	wire [8-1:0] node6170;
	wire [8-1:0] node6173;
	wire [8-1:0] node6175;
	wire [8-1:0] node6178;
	wire [8-1:0] node6179;
	wire [8-1:0] node6180;
	wire [8-1:0] node6181;
	wire [8-1:0] node6184;
	wire [8-1:0] node6185;
	wire [8-1:0] node6189;
	wire [8-1:0] node6191;
	wire [8-1:0] node6194;
	wire [8-1:0] node6195;
	wire [8-1:0] node6196;
	wire [8-1:0] node6197;
	wire [8-1:0] node6201;
	wire [8-1:0] node6204;
	wire [8-1:0] node6205;
	wire [8-1:0] node6209;
	wire [8-1:0] node6210;
	wire [8-1:0] node6211;
	wire [8-1:0] node6212;
	wire [8-1:0] node6213;
	wire [8-1:0] node6217;
	wire [8-1:0] node6218;
	wire [8-1:0] node6221;
	wire [8-1:0] node6224;
	wire [8-1:0] node6225;
	wire [8-1:0] node6226;
	wire [8-1:0] node6227;
	wire [8-1:0] node6230;
	wire [8-1:0] node6233;
	wire [8-1:0] node6235;
	wire [8-1:0] node6238;
	wire [8-1:0] node6239;
	wire [8-1:0] node6240;
	wire [8-1:0] node6244;
	wire [8-1:0] node6247;
	wire [8-1:0] node6248;
	wire [8-1:0] node6249;
	wire [8-1:0] node6250;
	wire [8-1:0] node6254;
	wire [8-1:0] node6257;
	wire [8-1:0] node6258;
	wire [8-1:0] node6262;
	wire [8-1:0] node6263;
	wire [8-1:0] node6264;
	wire [8-1:0] node6265;
	wire [8-1:0] node6266;
	wire [8-1:0] node6267;
	wire [8-1:0] node6270;
	wire [8-1:0] node6273;
	wire [8-1:0] node6274;
	wire [8-1:0] node6277;
	wire [8-1:0] node6280;
	wire [8-1:0] node6281;
	wire [8-1:0] node6284;
	wire [8-1:0] node6285;
	wire [8-1:0] node6289;
	wire [8-1:0] node6290;
	wire [8-1:0] node6291;
	wire [8-1:0] node6292;
	wire [8-1:0] node6295;
	wire [8-1:0] node6298;
	wire [8-1:0] node6301;
	wire [8-1:0] node6302;
	wire [8-1:0] node6303;
	wire [8-1:0] node6306;
	wire [8-1:0] node6309;
	wire [8-1:0] node6311;
	wire [8-1:0] node6314;
	wire [8-1:0] node6315;
	wire [8-1:0] node6316;
	wire [8-1:0] node6317;
	wire [8-1:0] node6320;
	wire [8-1:0] node6323;
	wire [8-1:0] node6324;
	wire [8-1:0] node6327;
	wire [8-1:0] node6330;
	wire [8-1:0] node6331;
	wire [8-1:0] node6332;
	wire [8-1:0] node6335;
	wire [8-1:0] node6338;
	wire [8-1:0] node6339;
	wire [8-1:0] node6342;

	assign outp = (inp[4]) ? node3124 : node1;
		assign node1 = (inp[13]) ? node1461 : node2;
			assign node2 = (inp[7]) ? node372 : node3;
				assign node3 = (inp[11]) ? node125 : node4;
					assign node4 = (inp[0]) ? node72 : node5;
						assign node5 = (inp[2]) ? node29 : node6;
							assign node6 = (inp[1]) ? node14 : node7;
								assign node7 = (inp[8]) ? node9 : 8'b01111111;
									assign node9 = (inp[5]) ? node11 : 8'b00111011;
										assign node11 = (inp[10]) ? 8'b01111111 : 8'b00111011;
								assign node14 = (inp[8]) ? node20 : node15;
									assign node15 = (inp[3]) ? node17 : 8'b00111110;
										assign node17 = (inp[5]) ? 8'b01111111 : 8'b00111110;
									assign node20 = (inp[5]) ? node22 : 8'b00111010;
										assign node22 = (inp[3]) ? node26 : node23;
											assign node23 = (inp[10]) ? 8'b00111110 : 8'b00111010;
											assign node26 = (inp[10]) ? 8'b01111111 : 8'b00111011;
							assign node29 = (inp[8]) ? node45 : node30;
								assign node30 = (inp[1]) ? node36 : node31;
									assign node31 = (inp[5]) ? node33 : 8'b00101111;
										assign node33 = (inp[6]) ? 8'b01111111 : 8'b00101111;
									assign node36 = (inp[5]) ? node38 : 8'b00101110;
										assign node38 = (inp[6]) ? node42 : node39;
											assign node39 = (inp[3]) ? 8'b00101111 : 8'b00101110;
											assign node42 = (inp[3]) ? 8'b01111111 : 8'b00111110;
								assign node45 = (inp[5]) ? node49 : node46;
									assign node46 = (inp[1]) ? 8'b00101010 : 8'b00101011;
									assign node49 = (inp[10]) ? node61 : node50;
										assign node50 = (inp[6]) ? node56 : node51;
											assign node51 = (inp[3]) ? 8'b00101011 : node52;
												assign node52 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node56 = (inp[3]) ? 8'b00111011 : node57;
												assign node57 = (inp[1]) ? 8'b00111010 : 8'b00111011;
										assign node61 = (inp[6]) ? node67 : node62;
											assign node62 = (inp[1]) ? node64 : 8'b00101111;
												assign node64 = (inp[3]) ? 8'b00101111 : 8'b00101110;
											assign node67 = (inp[3]) ? 8'b01111111 : node68;
												assign node68 = (inp[1]) ? 8'b00111110 : 8'b01111111;
						assign node72 = (inp[5]) ? 8'b01111111 : node73;
							assign node73 = (inp[6]) ? node91 : node74;
								assign node74 = (inp[3]) ? node80 : node75;
									assign node75 = (inp[8]) ? node77 : 8'b01111111;
										assign node77 = (inp[10]) ? 8'b00111011 : 8'b01111111;
									assign node80 = (inp[1]) ? node86 : node81;
										assign node81 = (inp[10]) ? node83 : 8'b01111111;
											assign node83 = (inp[8]) ? 8'b00111011 : 8'b01111111;
										assign node86 = (inp[8]) ? node88 : 8'b00111110;
											assign node88 = (inp[10]) ? 8'b00111010 : 8'b00111110;
								assign node91 = (inp[2]) ? node105 : node92;
									assign node92 = (inp[10]) ? node98 : node93;
										assign node93 = (inp[1]) ? node95 : 8'b01111111;
											assign node95 = (inp[3]) ? 8'b00111110 : 8'b01111111;
										assign node98 = (inp[8]) ? node100 : 8'b01111111;
											assign node100 = (inp[1]) ? node102 : 8'b00111011;
												assign node102 = (inp[3]) ? 8'b00111010 : 8'b00111011;
									assign node105 = (inp[8]) ? node111 : node106;
										assign node106 = (inp[1]) ? node108 : 8'b00101111;
											assign node108 = (inp[3]) ? 8'b00101110 : 8'b00101111;
										assign node111 = (inp[10]) ? node117 : node112;
											assign node112 = (inp[3]) ? node114 : 8'b00101111;
												assign node114 = (inp[1]) ? 8'b00101110 : 8'b00101111;
											assign node117 = (inp[12]) ? node119 : 8'b00101011;
												assign node119 = (inp[3]) ? node121 : 8'b00101011;
													assign node121 = (inp[1]) ? 8'b00101010 : 8'b00101011;
					assign node125 = (inp[8]) ? node215 : node126;
						assign node126 = (inp[1]) ? node154 : node127;
							assign node127 = (inp[2]) ? node131 : node128;
								assign node128 = (inp[12]) ? 8'b01111111 : 8'b00101111;
								assign node131 = (inp[12]) ? node143 : node132;
									assign node132 = (inp[5]) ? node138 : node133;
										assign node133 = (inp[6]) ? 8'b00111110 : node134;
											assign node134 = (inp[0]) ? 8'b00101110 : 8'b00111110;
										assign node138 = (inp[6]) ? 8'b00101110 : node139;
											assign node139 = (inp[0]) ? 8'b00101110 : 8'b00111110;
									assign node143 = (inp[5]) ? node149 : node144;
										assign node144 = (inp[0]) ? node146 : 8'b00101111;
											assign node146 = (inp[6]) ? 8'b00101111 : 8'b00111110;
										assign node149 = (inp[0]) ? 8'b00111110 : node150;
											assign node150 = (inp[6]) ? 8'b00111110 : 8'b00101111;
							assign node154 = (inp[12]) ? node186 : node155;
								assign node155 = (inp[2]) ? node167 : node156;
									assign node156 = (inp[5]) ? node162 : node157;
										assign node157 = (inp[3]) ? 8'b00101110 : node158;
											assign node158 = (inp[0]) ? 8'b00101011 : 8'b00101110;
										assign node162 = (inp[3]) ? 8'b00101011 : node163;
											assign node163 = (inp[0]) ? 8'b00101011 : 8'b00101110;
									assign node167 = (inp[0]) ? node177 : node168;
										assign node168 = (inp[5]) ? node170 : 8'b00111011;
											assign node170 = (inp[3]) ? node174 : node171;
												assign node171 = (inp[6]) ? 8'b00101011 : 8'b00111011;
												assign node174 = (inp[6]) ? 8'b00101010 : 8'b00111010;
										assign node177 = (inp[5]) ? 8'b00101010 : node178;
											assign node178 = (inp[6]) ? node182 : node179;
												assign node179 = (inp[3]) ? 8'b00101011 : 8'b00101010;
												assign node182 = (inp[3]) ? 8'b00111011 : 8'b00111010;
								assign node186 = (inp[5]) ? node204 : node187;
									assign node187 = (inp[2]) ? node195 : node188;
										assign node188 = (inp[6]) ? node190 : 8'b00111110;
											assign node190 = (inp[0]) ? node192 : 8'b00111110;
												assign node192 = (inp[3]) ? 8'b00111110 : 8'b00111011;
										assign node195 = (inp[0]) ? node197 : 8'b00101110;
											assign node197 = (inp[6]) ? node201 : node198;
												assign node198 = (inp[3]) ? 8'b00111011 : 8'b00111010;
												assign node201 = (inp[3]) ? 8'b00101110 : 8'b00101011;
									assign node204 = (inp[2]) ? node210 : node205;
										assign node205 = (inp[3]) ? 8'b00111011 : node206;
											assign node206 = (inp[0]) ? 8'b00111011 : 8'b00111110;
										assign node210 = (inp[0]) ? 8'b00111010 : node211;
											assign node211 = (inp[6]) ? 8'b00111010 : 8'b00101011;
						assign node215 = (inp[5]) ? node293 : node216;
							assign node216 = (inp[0]) ? node232 : node217;
								assign node217 = (inp[1]) ? node225 : node218;
									assign node218 = (inp[12]) ? node222 : node219;
										assign node219 = (inp[2]) ? 8'b00111010 : 8'b00101011;
										assign node222 = (inp[2]) ? 8'b00101011 : 8'b00111011;
									assign node225 = (inp[2]) ? node229 : node226;
										assign node226 = (inp[12]) ? 8'b00111010 : 8'b00101010;
										assign node229 = (inp[12]) ? 8'b00101010 : 8'b00011111;
								assign node232 = (inp[10]) ? node266 : node233;
									assign node233 = (inp[1]) ? node245 : node234;
										assign node234 = (inp[2]) ? node238 : node235;
											assign node235 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node238 = (inp[12]) ? node242 : node239;
												assign node239 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node242 = (inp[6]) ? 8'b00001111 : 8'b00011110;
										assign node245 = (inp[3]) ? node257 : node246;
											assign node246 = (inp[2]) ? node250 : node247;
												assign node247 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node250 = (inp[12]) ? node254 : node251;
													assign node251 = (inp[9]) ? 8'b00001010 : 8'b00011010;
													assign node254 = (inp[9]) ? 8'b00011010 : 8'b00001011;
											assign node257 = (inp[2]) ? node261 : node258;
												assign node258 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node261 = (inp[9]) ? 8'b00011011 : node262;
													assign node262 = (inp[12]) ? 8'b00001110 : 8'b00011011;
									assign node266 = (inp[1]) ? node278 : node267;
										assign node267 = (inp[2]) ? node271 : node268;
											assign node268 = (inp[12]) ? 8'b00111011 : 8'b00101011;
											assign node271 = (inp[9]) ? node273 : 8'b00111010;
												assign node273 = (inp[6]) ? node275 : 8'b00111010;
													assign node275 = (inp[12]) ? 8'b00101011 : 8'b00111010;
										assign node278 = (inp[3]) ? node288 : node279;
											assign node279 = (inp[2]) ? node283 : node280;
												assign node280 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node283 = (inp[12]) ? 8'b00011110 : node284;
													assign node284 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node288 = (inp[12]) ? 8'b00101010 : node289;
												assign node289 = (inp[2]) ? 8'b00011111 : 8'b00101010;
							assign node293 = (inp[12]) ? node337 : node294;
								assign node294 = (inp[2]) ? node310 : node295;
									assign node295 = (inp[1]) ? node301 : node296;
										assign node296 = (inp[10]) ? 8'b00001111 : node297;
											assign node297 = (inp[0]) ? 8'b00001111 : 8'b00101011;
										assign node301 = (inp[0]) ? 8'b00001011 : node302;
											assign node302 = (inp[3]) ? node306 : node303;
												assign node303 = (inp[10]) ? 8'b00001110 : 8'b00101010;
												assign node306 = (inp[10]) ? 8'b00001011 : 8'b00001111;
									assign node310 = (inp[1]) ? node322 : node311;
										assign node311 = (inp[10]) ? node317 : node312;
											assign node312 = (inp[0]) ? 8'b00001110 : node313;
												assign node313 = (inp[6]) ? 8'b00101010 : 8'b00111010;
											assign node317 = (inp[0]) ? 8'b00001110 : node318;
												assign node318 = (inp[6]) ? 8'b00001110 : 8'b00011110;
										assign node322 = (inp[3]) ? node330 : node323;
											assign node323 = (inp[6]) ? node327 : node324;
												assign node324 = (inp[10]) ? 8'b00011011 : 8'b00011111;
												assign node327 = (inp[0]) ? 8'b00001010 : 8'b00001111;
											assign node330 = (inp[0]) ? 8'b00001010 : node331;
												assign node331 = (inp[6]) ? node333 : 8'b00011010;
													assign node333 = (inp[10]) ? 8'b00001010 : 8'b00001110;
								assign node337 = (inp[2]) ? node353 : node338;
									assign node338 = (inp[1]) ? node344 : node339;
										assign node339 = (inp[10]) ? 8'b00011111 : node340;
											assign node340 = (inp[0]) ? 8'b00011111 : 8'b00111011;
										assign node344 = (inp[0]) ? 8'b00011011 : node345;
											assign node345 = (inp[3]) ? node349 : node346;
												assign node346 = (inp[6]) ? 8'b00111010 : 8'b00011110;
												assign node349 = (inp[10]) ? 8'b00011011 : 8'b00011111;
									assign node353 = (inp[0]) ? node369 : node354;
										assign node354 = (inp[6]) ? node362 : node355;
											assign node355 = (inp[10]) ? node359 : node356;
												assign node356 = (inp[1]) ? 8'b00001111 : 8'b00101011;
												assign node359 = (inp[1]) ? 8'b00001110 : 8'b00001111;
											assign node362 = (inp[10]) ? node366 : node363;
												assign node363 = (inp[1]) ? 8'b00011110 : 8'b00111010;
												assign node366 = (inp[1]) ? 8'b00011011 : 8'b00011110;
										assign node369 = (inp[1]) ? 8'b00011010 : 8'b00011110;
				assign node372 = (inp[9]) ? node894 : node373;
					assign node373 = (inp[11]) ? node551 : node374;
						assign node374 = (inp[6]) ? node462 : node375;
							assign node375 = (inp[0]) ? node439 : node376;
								assign node376 = (inp[2]) ? node404 : node377;
									assign node377 = (inp[5]) ? node387 : node378;
										assign node378 = (inp[8]) ? node382 : node379;
											assign node379 = (inp[10]) ? 8'b00111010 : 8'b00111110;
											assign node382 = (inp[3]) ? 8'b00111010 : node383;
												assign node383 = (inp[1]) ? 8'b00111010 : 8'b00111011;
										assign node387 = (inp[3]) ? node397 : node388;
											assign node388 = (inp[1]) ? node394 : node389;
												assign node389 = (inp[10]) ? 8'b01111111 : node390;
													assign node390 = (inp[8]) ? 8'b00111011 : 8'b01111111;
												assign node394 = (inp[8]) ? 8'b00111110 : 8'b00111010;
											assign node397 = (inp[1]) ? 8'b01111111 : node398;
												assign node398 = (inp[8]) ? node400 : 8'b00111010;
													assign node400 = (inp[10]) ? 8'b00111110 : 8'b00111010;
									assign node404 = (inp[10]) ? node420 : node405;
										assign node405 = (inp[8]) ? node415 : node406;
											assign node406 = (inp[3]) ? node410 : node407;
												assign node407 = (inp[1]) ? 8'b00101110 : 8'b00101111;
												assign node410 = (inp[1]) ? node412 : 8'b00101110;
													assign node412 = (inp[5]) ? 8'b00101111 : 8'b00101110;
											assign node415 = (inp[12]) ? 8'b00101010 : node416;
												assign node416 = (inp[3]) ? 8'b00101010 : 8'b00101011;
										assign node420 = (inp[8]) ? node430 : node421;
											assign node421 = (inp[3]) ? node425 : node422;
												assign node422 = (inp[1]) ? 8'b00101010 : 8'b00101011;
												assign node425 = (inp[1]) ? node427 : 8'b00101010;
													assign node427 = (inp[5]) ? 8'b00101011 : 8'b00101010;
											assign node430 = (inp[5]) ? node434 : node431;
												assign node431 = (inp[3]) ? 8'b00101010 : 8'b00101011;
												assign node434 = (inp[1]) ? node436 : 8'b00101110;
													assign node436 = (inp[3]) ? 8'b00101111 : 8'b00101110;
								assign node439 = (inp[3]) ? node447 : node440;
									assign node440 = (inp[10]) ? node442 : 8'b01111111;
										assign node442 = (inp[5]) ? node444 : 8'b00111011;
											assign node444 = (inp[8]) ? 8'b01111111 : 8'b00111011;
									assign node447 = (inp[5]) ? node451 : node448;
										assign node448 = (inp[10]) ? 8'b00111010 : 8'b00111110;
										assign node451 = (inp[1]) ? node457 : node452;
											assign node452 = (inp[10]) ? node454 : 8'b00111110;
												assign node454 = (inp[8]) ? 8'b00111110 : 8'b00111010;
											assign node457 = (inp[8]) ? 8'b01111111 : node458;
												assign node458 = (inp[10]) ? 8'b00111011 : 8'b01111111;
							assign node462 = (inp[5]) ? node488 : node463;
								assign node463 = (inp[10]) ? node481 : node464;
									assign node464 = (inp[8]) ? node472 : node465;
										assign node465 = (inp[3]) ? 8'b00101110 : node466;
											assign node466 = (inp[1]) ? node468 : 8'b00101111;
												assign node468 = (inp[0]) ? 8'b00101111 : 8'b00101110;
										assign node472 = (inp[0]) ? node478 : node473;
											assign node473 = (inp[3]) ? 8'b00101010 : node474;
												assign node474 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node478 = (inp[3]) ? 8'b00101110 : 8'b00101111;
									assign node481 = (inp[3]) ? 8'b00101010 : node482;
										assign node482 = (inp[1]) ? node484 : 8'b00101011;
											assign node484 = (inp[0]) ? 8'b00101011 : 8'b00101010;
								assign node488 = (inp[2]) ? node522 : node489;
									assign node489 = (inp[0]) ? node513 : node490;
										assign node490 = (inp[10]) ? node504 : node491;
											assign node491 = (inp[8]) ? node499 : node492;
												assign node492 = (inp[3]) ? node496 : node493;
													assign node493 = (inp[1]) ? 8'b00101110 : 8'b00101111;
													assign node496 = (inp[1]) ? 8'b00101111 : 8'b00101110;
												assign node499 = (inp[3]) ? 8'b00101011 : node500;
													assign node500 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node504 = (inp[8]) ? node510 : node505;
												assign node505 = (inp[3]) ? 8'b00101010 : node506;
													assign node506 = (inp[1]) ? 8'b00101010 : 8'b00101011;
												assign node510 = (inp[1]) ? 8'b00101110 : 8'b00101111;
										assign node513 = (inp[3]) ? node519 : node514;
											assign node514 = (inp[10]) ? node516 : 8'b00101111;
												assign node516 = (inp[8]) ? 8'b00101111 : 8'b00101011;
											assign node519 = (inp[1]) ? 8'b00101111 : 8'b00101110;
									assign node522 = (inp[0]) ? node538 : node523;
										assign node523 = (inp[3]) ? node527 : node524;
											assign node524 = (inp[1]) ? 8'b00111010 : 8'b00111011;
											assign node527 = (inp[1]) ? node531 : node528;
												assign node528 = (inp[10]) ? 8'b00111110 : 8'b00111010;
												assign node531 = (inp[12]) ? node535 : node532;
													assign node532 = (inp[8]) ? 8'b01111111 : 8'b00111011;
													assign node535 = (inp[8]) ? 8'b00111011 : 8'b01111111;
										assign node538 = (inp[10]) ? node544 : node539;
											assign node539 = (inp[1]) ? 8'b01111111 : node540;
												assign node540 = (inp[3]) ? 8'b00111110 : 8'b01111111;
											assign node544 = (inp[8]) ? node546 : 8'b00111011;
												assign node546 = (inp[12]) ? node548 : 8'b01111111;
													assign node548 = (inp[3]) ? 8'b00111110 : 8'b01111111;
						assign node551 = (inp[8]) ? node711 : node552;
							assign node552 = (inp[10]) ? node624 : node553;
								assign node553 = (inp[1]) ? node585 : node554;
									assign node554 = (inp[3]) ? node570 : node555;
										assign node555 = (inp[12]) ? node563 : node556;
											assign node556 = (inp[6]) ? node560 : node557;
												assign node557 = (inp[0]) ? 8'b00101110 : 8'b00101111;
												assign node560 = (inp[5]) ? 8'b00101110 : 8'b00111110;
											assign node563 = (inp[6]) ? 8'b00101111 : node564;
												assign node564 = (inp[2]) ? node566 : 8'b01111111;
													assign node566 = (inp[0]) ? 8'b00111110 : 8'b00101111;
										assign node570 = (inp[2]) ? node578 : node571;
											assign node571 = (inp[6]) ? node575 : node572;
												assign node572 = (inp[12]) ? 8'b00111110 : 8'b00101110;
												assign node575 = (inp[12]) ? 8'b00101110 : 8'b00111011;
											assign node578 = (inp[12]) ? node580 : 8'b00101011;
												assign node580 = (inp[0]) ? 8'b00111011 : node581;
													assign node581 = (inp[5]) ? 8'b00111011 : 8'b00101110;
									assign node585 = (inp[0]) ? node607 : node586;
										assign node586 = (inp[12]) ? node598 : node587;
											assign node587 = (inp[5]) ? node589 : 8'b00111011;
												assign node589 = (inp[3]) ? node595 : node590;
													assign node590 = (inp[6]) ? node592 : 8'b00111011;
														assign node592 = (inp[2]) ? 8'b00101011 : 8'b00111011;
													assign node595 = (inp[2]) ? 8'b00111010 : 8'b00101011;
											assign node598 = (inp[5]) ? node602 : node599;
												assign node599 = (inp[2]) ? 8'b00101110 : 8'b00111110;
												assign node602 = (inp[2]) ? 8'b00111011 : node603;
													assign node603 = (inp[3]) ? 8'b00111011 : 8'b00101110;
										assign node607 = (inp[3]) ? node613 : node608;
											assign node608 = (inp[12]) ? 8'b00111010 : node609;
												assign node609 = (inp[5]) ? 8'b00101010 : 8'b00111010;
											assign node613 = (inp[5]) ? node619 : node614;
												assign node614 = (inp[6]) ? 8'b00111011 : node615;
													assign node615 = (inp[2]) ? 8'b00111011 : 8'b00101110;
												assign node619 = (inp[2]) ? node621 : 8'b00101011;
													assign node621 = (inp[12]) ? 8'b00111010 : 8'b00101010;
								assign node624 = (inp[1]) ? node666 : node625;
									assign node625 = (inp[3]) ? node647 : node626;
										assign node626 = (inp[12]) ? node638 : node627;
											assign node627 = (inp[6]) ? node633 : node628;
												assign node628 = (inp[2]) ? node630 : 8'b00101011;
													assign node630 = (inp[0]) ? 8'b00101010 : 8'b00111010;
												assign node633 = (inp[2]) ? node635 : 8'b00111010;
													assign node635 = (inp[5]) ? 8'b00101010 : 8'b00111010;
											assign node638 = (inp[2]) ? node642 : node639;
												assign node639 = (inp[6]) ? 8'b00101011 : 8'b00111011;
												assign node642 = (inp[0]) ? node644 : 8'b00101011;
													assign node644 = (inp[5]) ? 8'b00111010 : 8'b00101011;
										assign node647 = (inp[12]) ? node659 : node648;
											assign node648 = (inp[6]) ? node654 : node649;
												assign node649 = (inp[2]) ? node651 : 8'b00101010;
													assign node651 = (inp[0]) ? 8'b00001111 : 8'b00011111;
												assign node654 = (inp[2]) ? node656 : 8'b00011111;
													assign node656 = (inp[5]) ? 8'b00001111 : 8'b00011111;
											assign node659 = (inp[5]) ? node663 : node660;
												assign node660 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node663 = (inp[6]) ? 8'b00011111 : 8'b00101010;
									assign node666 = (inp[2]) ? node684 : node667;
										assign node667 = (inp[6]) ? node675 : node668;
											assign node668 = (inp[12]) ? node670 : 8'b00101010;
												assign node670 = (inp[5]) ? 8'b00011111 : node671;
													assign node671 = (inp[3]) ? 8'b00111010 : 8'b00011111;
											assign node675 = (inp[12]) ? node679 : node676;
												assign node676 = (inp[5]) ? 8'b00011110 : 8'b00011111;
												assign node679 = (inp[5]) ? 8'b00001111 : node680;
													assign node680 = (inp[3]) ? 8'b00101010 : 8'b00001111;
										assign node684 = (inp[12]) ? node696 : node685;
											assign node685 = (inp[5]) ? node693 : node686;
												assign node686 = (inp[0]) ? node688 : 8'b00011111;
													assign node688 = (inp[3]) ? 8'b00001111 : node689;
														assign node689 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node693 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node696 = (inp[0]) ? node704 : node697;
												assign node697 = (inp[5]) ? node699 : 8'b00101010;
													assign node699 = (inp[3]) ? node701 : 8'b00101010;
														assign node701 = (inp[6]) ? 8'b00011110 : 8'b00001111;
												assign node704 = (inp[6]) ? node706 : 8'b00011110;
													assign node706 = (inp[3]) ? 8'b00101010 : node707;
														assign node707 = (inp[5]) ? 8'b00011110 : 8'b00001111;
							assign node711 = (inp[0]) ? node789 : node712;
								assign node712 = (inp[12]) ? node736 : node713;
									assign node713 = (inp[2]) ? node723 : node714;
										assign node714 = (inp[6]) ? node716 : 8'b00101010;
											assign node716 = (inp[3]) ? 8'b00011111 : node717;
												assign node717 = (inp[1]) ? node719 : 8'b00111010;
													assign node719 = (inp[5]) ? 8'b00011011 : 8'b00011111;
										assign node723 = (inp[5]) ? node725 : 8'b00011111;
											assign node725 = (inp[6]) ? node729 : node726;
												assign node726 = (inp[3]) ? 8'b00011110 : 8'b00111010;
												assign node729 = (inp[3]) ? 8'b00001010 : node730;
													assign node730 = (inp[1]) ? 8'b00001111 : node731;
														assign node731 = (inp[10]) ? 8'b00001110 : 8'b00101010;
									assign node736 = (inp[5]) ? node750 : node737;
										assign node737 = (inp[6]) ? node745 : node738;
											assign node738 = (inp[2]) ? 8'b00101010 : node739;
												assign node739 = (inp[1]) ? 8'b00111010 : node740;
													assign node740 = (inp[3]) ? 8'b00111010 : 8'b00111011;
											assign node745 = (inp[1]) ? 8'b00101010 : node746;
												assign node746 = (inp[3]) ? 8'b00101010 : 8'b00101011;
										assign node750 = (inp[10]) ? node770 : node751;
											assign node751 = (inp[3]) ? node761 : node752;
												assign node752 = (inp[1]) ? 8'b00101010 : node753;
													assign node753 = (inp[2]) ? node757 : node754;
														assign node754 = (inp[6]) ? 8'b00101011 : 8'b00111011;
														assign node757 = (inp[6]) ? 8'b00111010 : 8'b00101011;
												assign node761 = (inp[2]) ? node765 : node762;
													assign node762 = (inp[6]) ? 8'b00101010 : 8'b00111010;
													assign node765 = (inp[6]) ? 8'b00011111 : node766;
														assign node766 = (inp[1]) ? 8'b00001111 : 8'b00101010;
											assign node770 = (inp[1]) ? node780 : node771;
												assign node771 = (inp[3]) ? node775 : node772;
													assign node772 = (inp[6]) ? 8'b00011110 : 8'b00011111;
													assign node775 = (inp[2]) ? 8'b00001110 : node776;
														assign node776 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node780 = (inp[3]) ? node786 : node781;
													assign node781 = (inp[6]) ? node783 : 8'b00001110;
														assign node783 = (inp[2]) ? 8'b00011011 : 8'b00001110;
													assign node786 = (inp[6]) ? 8'b00011010 : 8'b00011011;
								assign node789 = (inp[1]) ? node847 : node790;
									assign node790 = (inp[10]) ? node816 : node791;
										assign node791 = (inp[3]) ? node803 : node792;
											assign node792 = (inp[2]) ? node796 : node793;
												assign node793 = (inp[6]) ? 8'b00001111 : 8'b00011111;
												assign node796 = (inp[12]) ? 8'b00011110 : node797;
													assign node797 = (inp[6]) ? node799 : 8'b00001110;
														assign node799 = (inp[5]) ? 8'b00001110 : 8'b00011110;
											assign node803 = (inp[2]) ? node811 : node804;
												assign node804 = (inp[12]) ? node808 : node805;
													assign node805 = (inp[6]) ? 8'b00011011 : 8'b00001110;
													assign node808 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node811 = (inp[6]) ? 8'b00001110 : node812;
													assign node812 = (inp[12]) ? 8'b00011011 : 8'b00001011;
										assign node816 = (inp[5]) ? node834 : node817;
											assign node817 = (inp[3]) ? node823 : node818;
												assign node818 = (inp[6]) ? 8'b00111010 : node819;
													assign node819 = (inp[12]) ? 8'b00111011 : 8'b00101011;
												assign node823 = (inp[2]) ? node829 : node824;
													assign node824 = (inp[6]) ? node826 : 8'b00101010;
														assign node826 = (inp[12]) ? 8'b00101010 : 8'b00011111;
													assign node829 = (inp[12]) ? 8'b00011111 : node830;
														assign node830 = (inp[6]) ? 8'b00011111 : 8'b00001111;
											assign node834 = (inp[2]) ? node844 : node835;
												assign node835 = (inp[3]) ? node839 : node836;
													assign node836 = (inp[12]) ? 8'b00011111 : 8'b00011110;
													assign node839 = (inp[6]) ? 8'b00001110 : node840;
														assign node840 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node844 = (inp[3]) ? 8'b00001011 : 8'b00001110;
									assign node847 = (inp[5]) ? node879 : node848;
										assign node848 = (inp[10]) ? node864 : node849;
											assign node849 = (inp[12]) ? node859 : node850;
												assign node850 = (inp[6]) ? 8'b00011011 : node851;
													assign node851 = (inp[2]) ? node855 : node852;
														assign node852 = (inp[3]) ? 8'b00001110 : 8'b00001011;
														assign node855 = (inp[3]) ? 8'b00001011 : 8'b00001010;
												assign node859 = (inp[6]) ? 8'b00001110 : node860;
													assign node860 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node864 = (inp[3]) ? node874 : node865;
												assign node865 = (inp[12]) ? node871 : node866;
													assign node866 = (inp[6]) ? 8'b00011110 : node867;
														assign node867 = (inp[2]) ? 8'b00001110 : 8'b00001111;
													assign node871 = (inp[6]) ? 8'b00001111 : 8'b00011111;
												assign node874 = (inp[6]) ? 8'b00011111 : node875;
													assign node875 = (inp[12]) ? 8'b00111010 : 8'b00101010;
										assign node879 = (inp[2]) ? node891 : node880;
											assign node880 = (inp[10]) ? node886 : node881;
												assign node881 = (inp[12]) ? 8'b00001011 : node882;
													assign node882 = (inp[6]) ? 8'b00011010 : 8'b00001011;
												assign node886 = (inp[3]) ? 8'b00001011 : node887;
													assign node887 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node891 = (inp[12]) ? 8'b00011010 : 8'b00001010;
					assign node894 = (inp[8]) ? node1184 : node895;
						assign node895 = (inp[10]) ? node1033 : node896;
							assign node896 = (inp[11]) ? node954 : node897;
								assign node897 = (inp[6]) ? node925 : node898;
									assign node898 = (inp[3]) ? node908 : node899;
										assign node899 = (inp[0]) ? 8'b00011111 : node900;
											assign node900 = (inp[2]) ? node904 : node901;
												assign node901 = (inp[1]) ? 8'b00011110 : 8'b00011111;
												assign node904 = (inp[1]) ? 8'b00001110 : 8'b00001111;
										assign node908 = (inp[1]) ? node914 : node909;
											assign node909 = (inp[2]) ? node911 : 8'b00011110;
												assign node911 = (inp[12]) ? 8'b00001110 : 8'b00011110;
											assign node914 = (inp[5]) ? node920 : node915;
												assign node915 = (inp[0]) ? 8'b00011110 : node916;
													assign node916 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node920 = (inp[0]) ? 8'b00011111 : node921;
													assign node921 = (inp[12]) ? 8'b00011111 : 8'b00001111;
									assign node925 = (inp[5]) ? node933 : node926;
										assign node926 = (inp[3]) ? 8'b00001110 : node927;
											assign node927 = (inp[1]) ? node929 : 8'b00001111;
												assign node929 = (inp[12]) ? 8'b00001110 : 8'b00001111;
										assign node933 = (inp[2]) ? node945 : node934;
											assign node934 = (inp[0]) ? node940 : node935;
												assign node935 = (inp[1]) ? node937 : 8'b00001111;
													assign node937 = (inp[3]) ? 8'b00001111 : 8'b00001110;
												assign node940 = (inp[3]) ? node942 : 8'b00001111;
													assign node942 = (inp[1]) ? 8'b00001111 : 8'b00001110;
											assign node945 = (inp[0]) ? 8'b00011111 : node946;
												assign node946 = (inp[1]) ? node950 : node947;
													assign node947 = (inp[3]) ? 8'b00011110 : 8'b00011111;
													assign node950 = (inp[3]) ? 8'b00011111 : 8'b00011110;
								assign node954 = (inp[1]) ? node988 : node955;
									assign node955 = (inp[6]) ? node971 : node956;
										assign node956 = (inp[12]) ? node964 : node957;
											assign node957 = (inp[5]) ? 8'b00001011 : node958;
												assign node958 = (inp[2]) ? node960 : 8'b00001110;
													assign node960 = (inp[0]) ? 8'b00001110 : 8'b00011110;
											assign node964 = (inp[3]) ? node968 : node965;
												assign node965 = (inp[2]) ? 8'b00011110 : 8'b00011111;
												assign node968 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node971 = (inp[3]) ? node979 : node972;
											assign node972 = (inp[12]) ? node976 : node973;
												assign node973 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node976 = (inp[2]) ? 8'b00011110 : 8'b00001111;
											assign node979 = (inp[12]) ? node983 : node980;
												assign node980 = (inp[0]) ? 8'b00001011 : 8'b00011011;
												assign node983 = (inp[2]) ? node985 : 8'b00001110;
													assign node985 = (inp[5]) ? 8'b00011011 : 8'b00001110;
									assign node988 = (inp[12]) ? node1006 : node989;
										assign node989 = (inp[6]) ? node997 : node990;
											assign node990 = (inp[2]) ? node992 : 8'b00001110;
												assign node992 = (inp[3]) ? node994 : 8'b00011011;
													assign node994 = (inp[5]) ? 8'b00001010 : 8'b00001011;
											assign node997 = (inp[5]) ? node1003 : node998;
												assign node998 = (inp[0]) ? node1000 : 8'b00011011;
													assign node1000 = (inp[3]) ? 8'b00011011 : 8'b00011010;
												assign node1003 = (inp[2]) ? 8'b00001011 : 8'b00011011;
										assign node1006 = (inp[5]) ? node1020 : node1007;
											assign node1007 = (inp[0]) ? node1013 : node1008;
												assign node1008 = (inp[2]) ? 8'b00001110 : node1009;
													assign node1009 = (inp[3]) ? 8'b00011110 : 8'b00001110;
												assign node1013 = (inp[3]) ? node1017 : node1014;
													assign node1014 = (inp[6]) ? 8'b00001011 : 8'b00011010;
													assign node1017 = (inp[2]) ? 8'b00001110 : 8'b00011110;
											assign node1020 = (inp[2]) ? node1026 : node1021;
												assign node1021 = (inp[6]) ? 8'b00001011 : node1022;
													assign node1022 = (inp[0]) ? 8'b00011011 : 8'b00011110;
												assign node1026 = (inp[3]) ? node1028 : 8'b00001110;
													assign node1028 = (inp[0]) ? 8'b00011010 : node1029;
														assign node1029 = (inp[6]) ? 8'b00011010 : 8'b00001011;
							assign node1033 = (inp[1]) ? node1097 : node1034;
								assign node1034 = (inp[3]) ? node1066 : node1035;
									assign node1035 = (inp[6]) ? node1053 : node1036;
										assign node1036 = (inp[0]) ? node1046 : node1037;
											assign node1037 = (inp[2]) ? node1041 : node1038;
												assign node1038 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node1041 = (inp[11]) ? node1043 : 8'b00001011;
													assign node1043 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node1046 = (inp[11]) ? node1048 : 8'b00011011;
												assign node1048 = (inp[2]) ? 8'b00011010 : node1049;
													assign node1049 = (inp[12]) ? 8'b00011011 : 8'b00001011;
										assign node1053 = (inp[12]) ? node1061 : node1054;
											assign node1054 = (inp[11]) ? node1056 : 8'b00001011;
												assign node1056 = (inp[2]) ? node1058 : 8'b00011010;
													assign node1058 = (inp[5]) ? 8'b00001010 : 8'b00011010;
											assign node1061 = (inp[5]) ? node1063 : 8'b00001011;
												assign node1063 = (inp[2]) ? 8'b00011011 : 8'b00001011;
									assign node1066 = (inp[2]) ? node1078 : node1067;
										assign node1067 = (inp[6]) ? node1073 : node1068;
											assign node1068 = (inp[11]) ? node1070 : 8'b00011010;
												assign node1070 = (inp[12]) ? 8'b00011010 : 8'b00001010;
											assign node1073 = (inp[12]) ? 8'b00000010 : node1074;
												assign node1074 = (inp[11]) ? 8'b11110111 : 8'b10000010;
										assign node1078 = (inp[11]) ? node1088 : node1079;
											assign node1079 = (inp[0]) ? 8'b10010000 : node1080;
												assign node1080 = (inp[6]) ? node1084 : node1081;
													assign node1081 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node1084 = (inp[12]) ? 8'b10010000 : 8'b10000010;
											assign node1088 = (inp[12]) ? node1094 : node1089;
												assign node1089 = (inp[5]) ? node1091 : 8'b11110111;
													assign node1091 = (inp[0]) ? 8'b10100101 : 8'b11110111;
												assign node1094 = (inp[0]) ? 8'b11110101 : 8'b00000010;
								assign node1097 = (inp[11]) ? node1131 : node1098;
									assign node1098 = (inp[0]) ? node1118 : node1099;
										assign node1099 = (inp[5]) ? node1107 : node1100;
											assign node1100 = (inp[2]) ? node1104 : node1101;
												assign node1101 = (inp[6]) ? 8'b00000010 : 8'b00011010;
												assign node1104 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node1107 = (inp[3]) ? node1113 : node1108;
												assign node1108 = (inp[6]) ? node1110 : 8'b00011010;
													assign node1110 = (inp[2]) ? 8'b10010000 : 8'b10000010;
												assign node1113 = (inp[2]) ? node1115 : 8'b10011001;
													assign node1115 = (inp[6]) ? 8'b10010001 : 8'b10000001;
										assign node1118 = (inp[6]) ? node1126 : node1119;
											assign node1119 = (inp[2]) ? 8'b10010001 : node1120;
												assign node1120 = (inp[3]) ? node1122 : 8'b10011001;
													assign node1122 = (inp[5]) ? 8'b10011001 : 8'b00011010;
											assign node1126 = (inp[3]) ? node1128 : 8'b10000001;
												assign node1128 = (inp[5]) ? 8'b10000001 : 8'b10000010;
									assign node1131 = (inp[5]) ? node1151 : node1132;
										assign node1132 = (inp[2]) ? node1144 : node1133;
											assign node1133 = (inp[6]) ? node1141 : node1134;
												assign node1134 = (inp[12]) ? node1136 : 8'b00001010;
													assign node1136 = (inp[3]) ? 8'b00011010 : node1137;
														assign node1137 = (inp[0]) ? 8'b11111101 : 8'b00011010;
												assign node1141 = (inp[12]) ? 8'b00000010 : 8'b11110111;
											assign node1144 = (inp[12]) ? 8'b00000010 : node1145;
												assign node1145 = (inp[3]) ? 8'b11110111 : node1146;
													assign node1146 = (inp[6]) ? 8'b10110100 : 8'b10100100;
										assign node1151 = (inp[0]) ? node1173 : node1152;
											assign node1152 = (inp[3]) ? node1166 : node1153;
												assign node1153 = (inp[6]) ? node1161 : node1154;
													assign node1154 = (inp[2]) ? node1158 : node1155;
														assign node1155 = (inp[12]) ? 8'b00011010 : 8'b00001010;
														assign node1158 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node1161 = (inp[2]) ? 8'b11110101 : node1162;
														assign node1162 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node1166 = (inp[12]) ? node1170 : node1167;
													assign node1167 = (inp[2]) ? 8'b10100100 : 8'b10110100;
													assign node1170 = (inp[2]) ? 8'b10110100 : 8'b10100101;
											assign node1173 = (inp[2]) ? node1181 : node1174;
												assign node1174 = (inp[6]) ? node1178 : node1175;
													assign node1175 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node1178 = (inp[12]) ? 8'b10100101 : 8'b10110100;
												assign node1181 = (inp[12]) ? 8'b10110100 : 8'b10100100;
						assign node1184 = (inp[0]) ? node1316 : node1185;
							assign node1185 = (inp[5]) ? node1223 : node1186;
								assign node1186 = (inp[12]) ? node1206 : node1187;
									assign node1187 = (inp[11]) ? node1197 : node1188;
										assign node1188 = (inp[2]) ? node1192 : node1189;
											assign node1189 = (inp[6]) ? 8'b10000010 : 8'b00011010;
											assign node1192 = (inp[3]) ? 8'b10000010 : node1193;
												assign node1193 = (inp[1]) ? 8'b10000010 : 8'b00001011;
										assign node1197 = (inp[3]) ? 8'b11110111 : node1198;
											assign node1198 = (inp[1]) ? node1200 : 8'b00011010;
												assign node1200 = (inp[2]) ? 8'b11110111 : node1201;
													assign node1201 = (inp[6]) ? 8'b11110111 : 8'b00001010;
									assign node1206 = (inp[3]) ? node1218 : node1207;
										assign node1207 = (inp[1]) ? node1213 : node1208;
											assign node1208 = (inp[6]) ? 8'b00001011 : node1209;
												assign node1209 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node1213 = (inp[6]) ? 8'b00000010 : node1214;
												assign node1214 = (inp[2]) ? 8'b00000010 : 8'b00011010;
										assign node1218 = (inp[6]) ? 8'b00000010 : node1219;
											assign node1219 = (inp[2]) ? 8'b00000010 : 8'b00011010;
								assign node1223 = (inp[10]) ? node1271 : node1224;
									assign node1224 = (inp[3]) ? node1252 : node1225;
										assign node1225 = (inp[1]) ? node1233 : node1226;
											assign node1226 = (inp[11]) ? 8'b00001010 : node1227;
												assign node1227 = (inp[6]) ? node1229 : 8'b00011011;
													assign node1229 = (inp[2]) ? 8'b00011011 : 8'b00001011;
											assign node1233 = (inp[12]) ? node1245 : node1234;
												assign node1234 = (inp[11]) ? node1240 : node1235;
													assign node1235 = (inp[6]) ? 8'b10000010 : node1236;
														assign node1236 = (inp[2]) ? 8'b10000010 : 8'b00011010;
													assign node1240 = (inp[2]) ? 8'b11110111 : node1241;
														assign node1241 = (inp[6]) ? 8'b11110111 : 8'b00001010;
												assign node1245 = (inp[2]) ? node1249 : node1246;
													assign node1246 = (inp[6]) ? 8'b00000010 : 8'b00011010;
													assign node1249 = (inp[6]) ? 8'b10010000 : 8'b00000010;
										assign node1252 = (inp[1]) ? node1260 : node1253;
											assign node1253 = (inp[12]) ? node1255 : 8'b11110111;
												assign node1255 = (inp[11]) ? node1257 : 8'b00000010;
													assign node1257 = (inp[6]) ? 8'b00000010 : 8'b00011010;
											assign node1260 = (inp[11]) ? node1266 : node1261;
												assign node1261 = (inp[6]) ? node1263 : 8'b10011001;
													assign node1263 = (inp[2]) ? 8'b10010001 : 8'b10000001;
												assign node1266 = (inp[12]) ? 8'b10100101 : node1267;
													assign node1267 = (inp[6]) ? 8'b10110100 : 8'b10101101;
									assign node1271 = (inp[11]) ? node1287 : node1272;
										assign node1272 = (inp[6]) ? node1280 : node1273;
											assign node1273 = (inp[2]) ? node1277 : node1274;
												assign node1274 = (inp[3]) ? 8'b10011101 : 8'b10011100;
												assign node1277 = (inp[12]) ? 8'b10001101 : 8'b10000100;
											assign node1280 = (inp[3]) ? node1282 : 8'b10011101;
												assign node1282 = (inp[12]) ? node1284 : 8'b10000101;
													assign node1284 = (inp[2]) ? 8'b10010100 : 8'b10000100;
										assign node1287 = (inp[2]) ? node1301 : node1288;
											assign node1288 = (inp[3]) ? node1298 : node1289;
												assign node1289 = (inp[1]) ? node1295 : node1290;
													assign node1290 = (inp[12]) ? 8'b10101101 : node1291;
														assign node1291 = (inp[6]) ? 8'b10111100 : 8'b10101101;
													assign node1295 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node1298 = (inp[6]) ? 8'b10110000 : 8'b10101001;
											assign node1301 = (inp[1]) ? node1307 : node1302;
												assign node1302 = (inp[3]) ? node1304 : 8'b10101101;
													assign node1304 = (inp[6]) ? 8'b10100001 : 8'b10100100;
												assign node1307 = (inp[3]) ? 8'b10110000 : node1308;
													assign node1308 = (inp[12]) ? node1312 : node1309;
														assign node1309 = (inp[6]) ? 8'b10100001 : 8'b10110001;
														assign node1312 = (inp[6]) ? 8'b10110001 : 8'b10100100;
							assign node1316 = (inp[11]) ? node1372 : node1317;
								assign node1317 = (inp[3]) ? node1347 : node1318;
									assign node1318 = (inp[6]) ? node1332 : node1319;
										assign node1319 = (inp[5]) ? node1327 : node1320;
											assign node1320 = (inp[10]) ? node1322 : 8'b10011101;
												assign node1322 = (inp[1]) ? node1324 : 8'b00011011;
													assign node1324 = (inp[12]) ? 8'b10011001 : 8'b10010001;
											assign node1327 = (inp[1]) ? node1329 : 8'b10011101;
												assign node1329 = (inp[2]) ? 8'b10010101 : 8'b10011101;
										assign node1332 = (inp[1]) ? node1340 : node1333;
											assign node1333 = (inp[5]) ? node1337 : node1334;
												assign node1334 = (inp[10]) ? 8'b00001011 : 8'b10001101;
												assign node1337 = (inp[2]) ? 8'b10011101 : 8'b10001101;
											assign node1340 = (inp[5]) ? node1344 : node1341;
												assign node1341 = (inp[10]) ? 8'b10000001 : 8'b10000101;
												assign node1344 = (inp[2]) ? 8'b10010101 : 8'b10000101;
									assign node1347 = (inp[6]) ? node1359 : node1348;
										assign node1348 = (inp[2]) ? node1352 : node1349;
											assign node1349 = (inp[1]) ? 8'b10011101 : 8'b10011100;
											assign node1352 = (inp[10]) ? node1356 : node1353;
												assign node1353 = (inp[5]) ? 8'b10010101 : 8'b10010100;
												assign node1356 = (inp[12]) ? 8'b10010000 : 8'b10010100;
										assign node1359 = (inp[5]) ? node1365 : node1360;
											assign node1360 = (inp[10]) ? node1362 : 8'b10000100;
												assign node1362 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node1365 = (inp[2]) ? node1369 : node1366;
												assign node1366 = (inp[1]) ? 8'b10000101 : 8'b10000100;
												assign node1369 = (inp[1]) ? 8'b10010101 : 8'b10010100;
								assign node1372 = (inp[5]) ? node1432 : node1373;
									assign node1373 = (inp[10]) ? node1401 : node1374;
										assign node1374 = (inp[1]) ? node1388 : node1375;
											assign node1375 = (inp[3]) ? node1381 : node1376;
												assign node1376 = (inp[6]) ? 8'b10101101 : node1377;
													assign node1377 = (inp[2]) ? 8'b10101100 : 8'b10101101;
												assign node1381 = (inp[2]) ? 8'b10100001 : node1382;
													assign node1382 = (inp[6]) ? 8'b10100100 : node1383;
														assign node1383 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node1388 = (inp[2]) ? node1394 : node1389;
												assign node1389 = (inp[3]) ? node1391 : 8'b10111001;
													assign node1391 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node1394 = (inp[3]) ? node1396 : 8'b10110000;
													assign node1396 = (inp[6]) ? node1398 : 8'b10110001;
														assign node1398 = (inp[12]) ? 8'b10100100 : 8'b10110001;
										assign node1401 = (inp[1]) ? node1417 : node1402;
											assign node1402 = (inp[3]) ? node1408 : node1403;
												assign node1403 = (inp[12]) ? node1405 : 8'b00001010;
													assign node1405 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node1408 = (inp[12]) ? node1412 : node1409;
													assign node1409 = (inp[6]) ? 8'b11110111 : 8'b10100101;
													assign node1412 = (inp[6]) ? 8'b00000010 : node1413;
														assign node1413 = (inp[2]) ? 8'b11110101 : 8'b00011010;
											assign node1417 = (inp[3]) ? node1427 : node1418;
												assign node1418 = (inp[12]) ? node1424 : node1419;
													assign node1419 = (inp[6]) ? 8'b10110100 : node1420;
														assign node1420 = (inp[2]) ? 8'b10100100 : 8'b10101101;
													assign node1424 = (inp[6]) ? 8'b10100101 : 8'b11111101;
												assign node1427 = (inp[2]) ? node1429 : 8'b00000010;
													assign node1429 = (inp[6]) ? 8'b11110111 : 8'b10100101;
									assign node1432 = (inp[1]) ? node1450 : node1433;
										assign node1433 = (inp[3]) ? node1441 : node1434;
											assign node1434 = (inp[2]) ? node1438 : node1435;
												assign node1435 = (inp[10]) ? 8'b10111100 : 8'b10101101;
												assign node1438 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node1441 = (inp[2]) ? node1447 : node1442;
												assign node1442 = (inp[12]) ? node1444 : 8'b10110001;
													assign node1444 = (inp[6]) ? 8'b10100100 : 8'b10111100;
												assign node1447 = (inp[12]) ? 8'b10110001 : 8'b10100001;
										assign node1450 = (inp[2]) ? node1458 : node1451;
											assign node1451 = (inp[6]) ? node1455 : node1452;
												assign node1452 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node1455 = (inp[12]) ? 8'b10100001 : 8'b10110000;
											assign node1458 = (inp[12]) ? 8'b10110000 : 8'b10100000;
			assign node1461 = (inp[0]) ? node2337 : node1462;
				assign node1462 = (inp[5]) ? node1658 : node1463;
					assign node1463 = (inp[8]) ? node1583 : node1464;
						assign node1464 = (inp[1]) ? node1536 : node1465;
							assign node1465 = (inp[7]) ? node1477 : node1466;
								assign node1466 = (inp[2]) ? node1472 : node1467;
									assign node1467 = (inp[11]) ? node1469 : 8'b00011111;
										assign node1469 = (inp[12]) ? 8'b00011111 : 8'b00001111;
									assign node1472 = (inp[12]) ? 8'b00001111 : node1473;
										assign node1473 = (inp[11]) ? 8'b00011110 : 8'b00001111;
								assign node1477 = (inp[10]) ? node1505 : node1478;
									assign node1478 = (inp[3]) ? node1494 : node1479;
										assign node1479 = (inp[2]) ? node1489 : node1480;
											assign node1480 = (inp[6]) ? node1486 : node1481;
												assign node1481 = (inp[11]) ? node1483 : 8'b00011111;
													assign node1483 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node1486 = (inp[11]) ? 8'b00011110 : 8'b00001111;
											assign node1489 = (inp[11]) ? node1491 : 8'b00001111;
												assign node1491 = (inp[12]) ? 8'b00001111 : 8'b00011110;
										assign node1494 = (inp[6]) ? 8'b00001110 : node1495;
											assign node1495 = (inp[2]) ? node1499 : node1496;
												assign node1496 = (inp[11]) ? 8'b00001110 : 8'b00011110;
												assign node1499 = (inp[12]) ? 8'b00001110 : node1500;
													assign node1500 = (inp[11]) ? 8'b00011011 : 8'b00001110;
									assign node1505 = (inp[3]) ? node1525 : node1506;
										assign node1506 = (inp[6]) ? node1520 : node1507;
											assign node1507 = (inp[9]) ? node1515 : node1508;
												assign node1508 = (inp[2]) ? 8'b00011010 : node1509;
													assign node1509 = (inp[12]) ? 8'b00011011 : node1510;
														assign node1510 = (inp[11]) ? 8'b00001011 : 8'b00011011;
												assign node1515 = (inp[11]) ? 8'b00001011 : node1516;
													assign node1516 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node1520 = (inp[11]) ? node1522 : 8'b00001011;
												assign node1522 = (inp[12]) ? 8'b00001011 : 8'b00011010;
										assign node1525 = (inp[11]) ? node1531 : node1526;
											assign node1526 = (inp[6]) ? node1528 : 8'b00011010;
												assign node1528 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node1531 = (inp[9]) ? node1533 : 8'b11110111;
												assign node1533 = (inp[2]) ? 8'b11110111 : 8'b00001010;
							assign node1536 = (inp[7]) ? node1548 : node1537;
								assign node1537 = (inp[2]) ? node1543 : node1538;
									assign node1538 = (inp[11]) ? node1540 : 8'b00011110;
										assign node1540 = (inp[12]) ? 8'b00011110 : 8'b00001110;
									assign node1543 = (inp[12]) ? 8'b00001110 : node1544;
										assign node1544 = (inp[11]) ? 8'b00011011 : 8'b00001110;
								assign node1548 = (inp[10]) ? node1566 : node1549;
									assign node1549 = (inp[12]) ? node1561 : node1550;
										assign node1550 = (inp[11]) ? node1556 : node1551;
											assign node1551 = (inp[6]) ? 8'b00001110 : node1552;
												assign node1552 = (inp[2]) ? 8'b00001110 : 8'b00011110;
											assign node1556 = (inp[2]) ? 8'b00011011 : node1557;
												assign node1557 = (inp[6]) ? 8'b00011011 : 8'b00001110;
										assign node1561 = (inp[2]) ? 8'b00001110 : node1562;
											assign node1562 = (inp[6]) ? 8'b00001110 : 8'b00011110;
									assign node1566 = (inp[12]) ? node1578 : node1567;
										assign node1567 = (inp[2]) ? node1575 : node1568;
											assign node1568 = (inp[6]) ? node1572 : node1569;
												assign node1569 = (inp[11]) ? 8'b00001010 : 8'b00011010;
												assign node1572 = (inp[11]) ? 8'b11110111 : 8'b10000010;
											assign node1575 = (inp[11]) ? 8'b11110111 : 8'b10000010;
										assign node1578 = (inp[2]) ? 8'b00000010 : node1579;
											assign node1579 = (inp[6]) ? 8'b00000010 : 8'b00011010;
						assign node1583 = (inp[1]) ? node1635 : node1584;
							assign node1584 = (inp[3]) ? node1608 : node1585;
								assign node1585 = (inp[2]) ? node1603 : node1586;
									assign node1586 = (inp[12]) ? node1598 : node1587;
										assign node1587 = (inp[11]) ? node1593 : node1588;
											assign node1588 = (inp[6]) ? node1590 : 8'b00011011;
												assign node1590 = (inp[10]) ? 8'b00011011 : 8'b00001011;
											assign node1593 = (inp[6]) ? node1595 : 8'b00001011;
												assign node1595 = (inp[7]) ? 8'b00011010 : 8'b00001011;
										assign node1598 = (inp[6]) ? node1600 : 8'b00011011;
											assign node1600 = (inp[7]) ? 8'b00001011 : 8'b00011011;
									assign node1603 = (inp[12]) ? 8'b00001011 : node1604;
										assign node1604 = (inp[11]) ? 8'b00011010 : 8'b00001011;
								assign node1608 = (inp[7]) ? node1622 : node1609;
									assign node1609 = (inp[2]) ? node1615 : node1610;
										assign node1610 = (inp[12]) ? 8'b00011011 : node1611;
											assign node1611 = (inp[11]) ? 8'b00001011 : 8'b00011011;
										assign node1615 = (inp[9]) ? 8'b00001011 : node1616;
											assign node1616 = (inp[12]) ? 8'b00001011 : node1617;
												assign node1617 = (inp[11]) ? 8'b00011010 : 8'b00001011;
									assign node1622 = (inp[12]) ? node1630 : node1623;
										assign node1623 = (inp[11]) ? 8'b11110111 : node1624;
											assign node1624 = (inp[6]) ? 8'b10000010 : node1625;
												assign node1625 = (inp[2]) ? 8'b10000010 : 8'b00011010;
										assign node1630 = (inp[6]) ? 8'b00000010 : node1631;
											assign node1631 = (inp[2]) ? 8'b00000010 : 8'b00011010;
							assign node1635 = (inp[2]) ? node1653 : node1636;
								assign node1636 = (inp[7]) ? node1642 : node1637;
									assign node1637 = (inp[12]) ? 8'b00011010 : node1638;
										assign node1638 = (inp[11]) ? 8'b00001010 : 8'b00011010;
									assign node1642 = (inp[6]) ? node1648 : node1643;
										assign node1643 = (inp[11]) ? node1645 : 8'b00011010;
											assign node1645 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node1648 = (inp[12]) ? 8'b00000010 : node1649;
											assign node1649 = (inp[11]) ? 8'b11110111 : 8'b10000010;
								assign node1653 = (inp[12]) ? 8'b00000010 : node1654;
									assign node1654 = (inp[11]) ? 8'b11110111 : 8'b10000010;
					assign node1658 = (inp[9]) ? node2016 : node1659;
						assign node1659 = (inp[8]) ? node1833 : node1660;
							assign node1660 = (inp[7]) ? node1712 : node1661;
								assign node1661 = (inp[1]) ? node1679 : node1662;
									assign node1662 = (inp[11]) ? node1668 : node1663;
										assign node1663 = (inp[2]) ? node1665 : 8'b00011111;
											assign node1665 = (inp[6]) ? 8'b00011111 : 8'b00001111;
										assign node1668 = (inp[2]) ? node1672 : node1669;
											assign node1669 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node1672 = (inp[6]) ? node1676 : node1673;
												assign node1673 = (inp[12]) ? 8'b00001111 : 8'b00011110;
												assign node1676 = (inp[12]) ? 8'b00011110 : 8'b00001110;
									assign node1679 = (inp[3]) ? node1695 : node1680;
										assign node1680 = (inp[11]) ? node1686 : node1681;
											assign node1681 = (inp[2]) ? node1683 : 8'b00011110;
												assign node1683 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node1686 = (inp[2]) ? node1690 : node1687;
												assign node1687 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node1690 = (inp[6]) ? node1692 : 8'b00001110;
													assign node1692 = (inp[12]) ? 8'b00011011 : 8'b00001011;
										assign node1695 = (inp[11]) ? node1701 : node1696;
											assign node1696 = (inp[2]) ? node1698 : 8'b00011111;
												assign node1698 = (inp[6]) ? 8'b00011111 : 8'b00001111;
											assign node1701 = (inp[2]) ? node1705 : node1702;
												assign node1702 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node1705 = (inp[6]) ? node1709 : node1706;
													assign node1706 = (inp[12]) ? 8'b00001011 : 8'b00011010;
													assign node1709 = (inp[12]) ? 8'b00011010 : 8'b00001010;
								assign node1712 = (inp[10]) ? node1768 : node1713;
									assign node1713 = (inp[11]) ? node1737 : node1714;
										assign node1714 = (inp[1]) ? node1722 : node1715;
											assign node1715 = (inp[3]) ? node1717 : 8'b00011111;
												assign node1717 = (inp[2]) ? 8'b00011110 : node1718;
													assign node1718 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node1722 = (inp[3]) ? node1734 : node1723;
												assign node1723 = (inp[12]) ? node1729 : node1724;
													assign node1724 = (inp[2]) ? node1726 : 8'b00001110;
														assign node1726 = (inp[6]) ? 8'b00011110 : 8'b00001110;
													assign node1729 = (inp[2]) ? 8'b00001110 : node1730;
														assign node1730 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node1734 = (inp[12]) ? 8'b00001111 : 8'b00011111;
										assign node1737 = (inp[3]) ? node1759 : node1738;
											assign node1738 = (inp[1]) ? node1752 : node1739;
												assign node1739 = (inp[12]) ? node1745 : node1740;
													assign node1740 = (inp[2]) ? node1742 : 8'b00011110;
														assign node1742 = (inp[6]) ? 8'b00001110 : 8'b00011110;
													assign node1745 = (inp[2]) ? node1749 : node1746;
														assign node1746 = (inp[6]) ? 8'b00001111 : 8'b00011111;
														assign node1749 = (inp[6]) ? 8'b00011110 : 8'b00001111;
												assign node1752 = (inp[2]) ? node1754 : 8'b00001110;
													assign node1754 = (inp[12]) ? node1756 : 8'b00011011;
														assign node1756 = (inp[6]) ? 8'b00011011 : 8'b00001110;
											assign node1759 = (inp[2]) ? node1765 : node1760;
												assign node1760 = (inp[1]) ? node1762 : 8'b00001110;
													assign node1762 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node1765 = (inp[1]) ? 8'b00011010 : 8'b00011011;
									assign node1768 = (inp[3]) ? node1804 : node1769;
										assign node1769 = (inp[1]) ? node1791 : node1770;
											assign node1770 = (inp[11]) ? node1784 : node1771;
												assign node1771 = (inp[12]) ? node1779 : node1772;
													assign node1772 = (inp[2]) ? node1776 : node1773;
														assign node1773 = (inp[6]) ? 8'b00001011 : 8'b00011011;
														assign node1776 = (inp[6]) ? 8'b00011011 : 8'b00001011;
													assign node1779 = (inp[2]) ? node1781 : 8'b00011011;
														assign node1781 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node1784 = (inp[12]) ? 8'b00011011 : node1785;
													assign node1785 = (inp[6]) ? node1787 : 8'b00011010;
														assign node1787 = (inp[2]) ? 8'b00001010 : 8'b00011010;
											assign node1791 = (inp[2]) ? node1799 : node1792;
												assign node1792 = (inp[6]) ? node1796 : node1793;
													assign node1793 = (inp[11]) ? 8'b00001010 : 8'b00011010;
													assign node1796 = (inp[11]) ? 8'b00000010 : 8'b10000010;
												assign node1799 = (inp[11]) ? node1801 : 8'b10010000;
													assign node1801 = (inp[6]) ? 8'b10100101 : 8'b11110111;
										assign node1804 = (inp[1]) ? node1818 : node1805;
											assign node1805 = (inp[2]) ? node1811 : node1806;
												assign node1806 = (inp[6]) ? node1808 : 8'b00011010;
													assign node1808 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node1811 = (inp[6]) ? node1815 : node1812;
													assign node1812 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node1815 = (inp[12]) ? 8'b11110101 : 8'b10010000;
											assign node1818 = (inp[11]) ? node1824 : node1819;
												assign node1819 = (inp[2]) ? node1821 : 8'b10000001;
													assign node1821 = (inp[6]) ? 8'b10010001 : 8'b10000001;
												assign node1824 = (inp[2]) ? node1828 : node1825;
													assign node1825 = (inp[6]) ? 8'b10100101 : 8'b11111101;
													assign node1828 = (inp[6]) ? 8'b10110100 : node1829;
														assign node1829 = (inp[12]) ? 8'b10100101 : 8'b10110100;
							assign node1833 = (inp[10]) ? node1921 : node1834;
								assign node1834 = (inp[1]) ? node1882 : node1835;
									assign node1835 = (inp[7]) ? node1853 : node1836;
										assign node1836 = (inp[11]) ? node1842 : node1837;
											assign node1837 = (inp[6]) ? 8'b00011011 : node1838;
												assign node1838 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node1842 = (inp[2]) ? node1846 : node1843;
												assign node1843 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node1846 = (inp[12]) ? node1850 : node1847;
													assign node1847 = (inp[6]) ? 8'b00001010 : 8'b00011010;
													assign node1850 = (inp[6]) ? 8'b00011010 : 8'b00001011;
										assign node1853 = (inp[3]) ? node1869 : node1854;
											assign node1854 = (inp[2]) ? node1862 : node1855;
												assign node1855 = (inp[11]) ? node1857 : 8'b00011011;
													assign node1857 = (inp[6]) ? 8'b00001011 : node1858;
														assign node1858 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node1862 = (inp[11]) ? node1864 : 8'b00011011;
													assign node1864 = (inp[6]) ? node1866 : 8'b00011010;
														assign node1866 = (inp[12]) ? 8'b00011010 : 8'b00001010;
											assign node1869 = (inp[6]) ? node1875 : node1870;
												assign node1870 = (inp[2]) ? 8'b00000010 : node1871;
													assign node1871 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node1875 = (inp[11]) ? 8'b10100101 : node1876;
													assign node1876 = (inp[2]) ? 8'b10010000 : node1877;
														assign node1877 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node1882 = (inp[3]) ? node1900 : node1883;
										assign node1883 = (inp[2]) ? node1893 : node1884;
											assign node1884 = (inp[12]) ? node1888 : node1885;
												assign node1885 = (inp[11]) ? 8'b00001010 : 8'b00011010;
												assign node1888 = (inp[7]) ? node1890 : 8'b00011010;
													assign node1890 = (inp[6]) ? 8'b00000010 : 8'b00011010;
											assign node1893 = (inp[6]) ? node1895 : 8'b00000010;
												assign node1895 = (inp[11]) ? node1897 : 8'b10010000;
													assign node1897 = (inp[12]) ? 8'b11110101 : 8'b10100101;
										assign node1900 = (inp[11]) ? node1908 : node1901;
											assign node1901 = (inp[2]) ? node1905 : node1902;
												assign node1902 = (inp[6]) ? 8'b10000001 : 8'b10011001;
												assign node1905 = (inp[6]) ? 8'b10010001 : 8'b10000001;
											assign node1908 = (inp[7]) ? node1916 : node1909;
												assign node1909 = (inp[2]) ? node1913 : node1910;
													assign node1910 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node1913 = (inp[12]) ? 8'b10100101 : 8'b10110100;
												assign node1916 = (inp[2]) ? node1918 : 8'b10110100;
													assign node1918 = (inp[12]) ? 8'b10110100 : 8'b10100100;
								assign node1921 = (inp[11]) ? node1969 : node1922;
									assign node1922 = (inp[1]) ? node1950 : node1923;
										assign node1923 = (inp[3]) ? node1937 : node1924;
											assign node1924 = (inp[12]) ? node1930 : node1925;
												assign node1925 = (inp[2]) ? 8'b10001101 : node1926;
													assign node1926 = (inp[6]) ? 8'b10001101 : 8'b10011101;
												assign node1930 = (inp[7]) ? node1932 : 8'b10011101;
													assign node1932 = (inp[2]) ? node1934 : 8'b10011101;
														assign node1934 = (inp[6]) ? 8'b10011101 : 8'b10001101;
											assign node1937 = (inp[7]) ? node1943 : node1938;
												assign node1938 = (inp[6]) ? 8'b10011101 : node1939;
													assign node1939 = (inp[2]) ? 8'b10001101 : 8'b10011101;
												assign node1943 = (inp[6]) ? node1947 : node1944;
													assign node1944 = (inp[2]) ? 8'b10000100 : 8'b10011100;
													assign node1947 = (inp[2]) ? 8'b10010100 : 8'b10000100;
										assign node1950 = (inp[3]) ? node1960 : node1951;
											assign node1951 = (inp[7]) ? node1955 : node1952;
												assign node1952 = (inp[2]) ? 8'b10010100 : 8'b10011100;
												assign node1955 = (inp[2]) ? node1957 : 8'b10000100;
													assign node1957 = (inp[6]) ? 8'b10010100 : 8'b10000100;
											assign node1960 = (inp[2]) ? node1966 : node1961;
												assign node1961 = (inp[6]) ? node1963 : 8'b10011101;
													assign node1963 = (inp[7]) ? 8'b10000101 : 8'b10011101;
												assign node1966 = (inp[7]) ? 8'b10010101 : 8'b10000101;
									assign node1969 = (inp[1]) ? node1993 : node1970;
										assign node1970 = (inp[2]) ? node1976 : node1971;
											assign node1971 = (inp[12]) ? 8'b11111101 : node1972;
												assign node1972 = (inp[7]) ? 8'b10101100 : 8'b10101101;
											assign node1976 = (inp[7]) ? node1988 : node1977;
												assign node1977 = (inp[3]) ? node1983 : node1978;
													assign node1978 = (inp[12]) ? node1980 : 8'b10111100;
														assign node1980 = (inp[6]) ? 8'b10111100 : 8'b10101101;
													assign node1983 = (inp[12]) ? 8'b10111100 : node1984;
														assign node1984 = (inp[6]) ? 8'b10101100 : 8'b10111100;
												assign node1988 = (inp[3]) ? node1990 : 8'b10111100;
													assign node1990 = (inp[6]) ? 8'b10100001 : 8'b10110001;
										assign node1993 = (inp[2]) ? node2003 : node1994;
											assign node1994 = (inp[3]) ? 8'b10111001 : node1995;
												assign node1995 = (inp[12]) ? node1997 : 8'b10110001;
													assign node1997 = (inp[6]) ? node1999 : 8'b10111100;
														assign node1999 = (inp[7]) ? 8'b10100100 : 8'b10111100;
											assign node2003 = (inp[7]) ? 8'b10110001 : node2004;
												assign node2004 = (inp[3]) ? node2012 : node2005;
													assign node2005 = (inp[6]) ? node2009 : node2006;
														assign node2006 = (inp[12]) ? 8'b10100100 : 8'b10110001;
														assign node2009 = (inp[12]) ? 8'b10110001 : 8'b10100001;
													assign node2012 = (inp[6]) ? 8'b10100000 : 8'b10100001;
						assign node2016 = (inp[8]) ? node2168 : node2017;
							assign node2017 = (inp[7]) ? node2065 : node2018;
								assign node2018 = (inp[1]) ? node2036 : node2019;
									assign node2019 = (inp[12]) ? node2029 : node2020;
										assign node2020 = (inp[11]) ? node2026 : node2021;
											assign node2021 = (inp[2]) ? node2023 : 8'b11111101;
												assign node2023 = (inp[6]) ? 8'b11111101 : 8'b10101101;
											assign node2026 = (inp[2]) ? 8'b10101100 : 8'b10101101;
										assign node2029 = (inp[2]) ? node2031 : 8'b11111101;
											assign node2031 = (inp[11]) ? 8'b10111100 : node2032;
												assign node2032 = (inp[3]) ? 8'b11111101 : 8'b10101101;
									assign node2036 = (inp[3]) ? node2054 : node2037;
										assign node2037 = (inp[11]) ? node2043 : node2038;
											assign node2038 = (inp[2]) ? node2040 : 8'b10111100;
												assign node2040 = (inp[6]) ? 8'b10111100 : 8'b10101100;
											assign node2043 = (inp[2]) ? node2047 : node2044;
												assign node2044 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node2047 = (inp[6]) ? node2051 : node2048;
													assign node2048 = (inp[12]) ? 8'b10101100 : 8'b10111001;
													assign node2051 = (inp[12]) ? 8'b10111001 : 8'b10101001;
										assign node2054 = (inp[11]) ? node2060 : node2055;
											assign node2055 = (inp[2]) ? node2057 : 8'b11111101;
												assign node2057 = (inp[6]) ? 8'b11111101 : 8'b10101101;
											assign node2060 = (inp[2]) ? 8'b10111000 : node2061;
												assign node2061 = (inp[12]) ? 8'b10111001 : 8'b10101001;
								assign node2065 = (inp[10]) ? node2113 : node2066;
									assign node2066 = (inp[11]) ? node2082 : node2067;
										assign node2067 = (inp[6]) ? node2071 : node2068;
											assign node2068 = (inp[2]) ? 8'b10101101 : 8'b11111101;
											assign node2071 = (inp[2]) ? node2077 : node2072;
												assign node2072 = (inp[1]) ? node2074 : 8'b10101101;
													assign node2074 = (inp[3]) ? 8'b10101101 : 8'b10101100;
												assign node2077 = (inp[1]) ? node2079 : 8'b10111100;
													assign node2079 = (inp[3]) ? 8'b11111101 : 8'b10111100;
										assign node2082 = (inp[1]) ? node2104 : node2083;
											assign node2083 = (inp[3]) ? node2095 : node2084;
												assign node2084 = (inp[6]) ? node2088 : node2085;
													assign node2085 = (inp[2]) ? 8'b10101101 : 8'b11111101;
													assign node2088 = (inp[2]) ? node2092 : node2089;
														assign node2089 = (inp[12]) ? 8'b10101101 : 8'b10111100;
														assign node2092 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node2095 = (inp[2]) ? node2099 : node2096;
													assign node2096 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node2099 = (inp[6]) ? 8'b10111001 : node2100;
														assign node2100 = (inp[12]) ? 8'b10101100 : 8'b10111001;
											assign node2104 = (inp[6]) ? node2110 : node2105;
												assign node2105 = (inp[3]) ? 8'b10111000 : node2106;
													assign node2106 = (inp[2]) ? 8'b10101100 : 8'b10111100;
												assign node2110 = (inp[3]) ? 8'b10101001 : 8'b10111001;
									assign node2113 = (inp[1]) ? node2143 : node2114;
										assign node2114 = (inp[3]) ? node2130 : node2115;
											assign node2115 = (inp[11]) ? node2121 : node2116;
												assign node2116 = (inp[6]) ? node2118 : 8'b10101001;
													assign node2118 = (inp[2]) ? 8'b10111001 : 8'b10101001;
												assign node2121 = (inp[2]) ? 8'b10111000 : node2122;
													assign node2122 = (inp[6]) ? node2126 : node2123;
														assign node2123 = (inp[12]) ? 8'b10111001 : 8'b10101001;
														assign node2126 = (inp[12]) ? 8'b10101001 : 8'b10111000;
											assign node2130 = (inp[6]) ? node2138 : node2131;
												assign node2131 = (inp[2]) ? 8'b10100000 : node2132;
													assign node2132 = (inp[12]) ? 8'b10111000 : node2133;
														assign node2133 = (inp[11]) ? 8'b10101000 : 8'b10111000;
												assign node2138 = (inp[2]) ? node2140 : 8'b10100000;
													assign node2140 = (inp[11]) ? 8'b10000101 : 8'b10110000;
										assign node2143 = (inp[11]) ? node2153 : node2144;
											assign node2144 = (inp[6]) ? node2148 : node2145;
												assign node2145 = (inp[12]) ? 8'b10111000 : 8'b10111001;
												assign node2148 = (inp[3]) ? 8'b10100001 : node2149;
													assign node2149 = (inp[2]) ? 8'b10110000 : 8'b10100000;
											assign node2153 = (inp[6]) ? node2161 : node2154;
												assign node2154 = (inp[3]) ? node2156 : 8'b10100000;
													assign node2156 = (inp[2]) ? node2158 : 8'b10001101;
														assign node2158 = (inp[12]) ? 8'b10000101 : 8'b10010100;
												assign node2161 = (inp[3]) ? node2163 : 8'b10010101;
													assign node2163 = (inp[12]) ? 8'b10010100 : node2164;
														assign node2164 = (inp[2]) ? 8'b10000100 : 8'b10010100;
							assign node2168 = (inp[11]) ? node2238 : node2169;
								assign node2169 = (inp[10]) ? node2199 : node2170;
									assign node2170 = (inp[1]) ? node2186 : node2171;
										assign node2171 = (inp[7]) ? node2177 : node2172;
											assign node2172 = (inp[6]) ? 8'b10111001 : node2173;
												assign node2173 = (inp[2]) ? 8'b10101001 : 8'b10111001;
											assign node2177 = (inp[3]) ? node2181 : node2178;
												assign node2178 = (inp[2]) ? 8'b10111001 : 8'b10101001;
												assign node2181 = (inp[6]) ? node2183 : 8'b10111000;
													assign node2183 = (inp[2]) ? 8'b10110000 : 8'b10100000;
										assign node2186 = (inp[3]) ? node2194 : node2187;
											assign node2187 = (inp[2]) ? node2191 : node2188;
												assign node2188 = (inp[7]) ? 8'b10100000 : 8'b10111000;
												assign node2191 = (inp[6]) ? 8'b10110000 : 8'b10100000;
											assign node2194 = (inp[2]) ? node2196 : 8'b10111001;
												assign node2196 = (inp[6]) ? 8'b10110001 : 8'b10100001;
									assign node2199 = (inp[7]) ? node2215 : node2200;
										assign node2200 = (inp[2]) ? node2206 : node2201;
											assign node2201 = (inp[1]) ? node2203 : 8'b11111101;
												assign node2203 = (inp[3]) ? 8'b11111101 : 8'b10111100;
											assign node2206 = (inp[6]) ? node2212 : node2207;
												assign node2207 = (inp[1]) ? node2209 : 8'b10101101;
													assign node2209 = (inp[3]) ? 8'b10100101 : 8'b10100100;
												assign node2212 = (inp[12]) ? 8'b11110101 : 8'b11111101;
										assign node2215 = (inp[3]) ? node2229 : node2216;
											assign node2216 = (inp[1]) ? node2222 : node2217;
												assign node2217 = (inp[6]) ? 8'b11111101 : node2218;
													assign node2218 = (inp[2]) ? 8'b10101101 : 8'b11111101;
												assign node2222 = (inp[6]) ? node2226 : node2223;
													assign node2223 = (inp[2]) ? 8'b10100100 : 8'b10111100;
													assign node2226 = (inp[2]) ? 8'b10110100 : 8'b10100100;
											assign node2229 = (inp[1]) ? 8'b10100101 : node2230;
												assign node2230 = (inp[6]) ? node2234 : node2231;
													assign node2231 = (inp[2]) ? 8'b10100100 : 8'b10111100;
													assign node2234 = (inp[2]) ? 8'b10110100 : 8'b10100100;
								assign node2238 = (inp[1]) ? node2288 : node2239;
									assign node2239 = (inp[10]) ? node2267 : node2240;
										assign node2240 = (inp[12]) ? node2252 : node2241;
											assign node2241 = (inp[2]) ? node2249 : node2242;
												assign node2242 = (inp[7]) ? node2244 : 8'b10101001;
													assign node2244 = (inp[6]) ? 8'b10111000 : node2245;
														assign node2245 = (inp[3]) ? 8'b10101000 : 8'b10101001;
												assign node2249 = (inp[6]) ? 8'b10101000 : 8'b10111000;
											assign node2252 = (inp[6]) ? node2264 : node2253;
												assign node2253 = (inp[2]) ? node2259 : node2254;
													assign node2254 = (inp[7]) ? node2256 : 8'b10111001;
														assign node2256 = (inp[3]) ? 8'b10111000 : 8'b10111001;
													assign node2259 = (inp[3]) ? node2261 : 8'b10101001;
														assign node2261 = (inp[7]) ? 8'b10100000 : 8'b10101001;
												assign node2264 = (inp[3]) ? 8'b10010101 : 8'b10111000;
										assign node2267 = (inp[7]) ? node2275 : node2268;
											assign node2268 = (inp[2]) ? node2270 : 8'b10001101;
												assign node2270 = (inp[3]) ? node2272 : 8'b10011100;
													assign node2272 = (inp[6]) ? 8'b10001100 : 8'b10011100;
											assign node2275 = (inp[6]) ? node2281 : node2276;
												assign node2276 = (inp[12]) ? node2278 : 8'b10001100;
													assign node2278 = (inp[2]) ? 8'b10001101 : 8'b10011101;
												assign node2281 = (inp[3]) ? node2283 : 8'b10011100;
													assign node2283 = (inp[2]) ? 8'b10010001 : node2284;
														assign node2284 = (inp[12]) ? 8'b10000100 : 8'b10010001;
									assign node2288 = (inp[2]) ? node2312 : node2289;
										assign node2289 = (inp[7]) ? node2299 : node2290;
											assign node2290 = (inp[3]) ? node2292 : 8'b10111000;
												assign node2292 = (inp[10]) ? node2296 : node2293;
													assign node2293 = (inp[6]) ? 8'b10011101 : 8'b10001101;
													assign node2296 = (inp[12]) ? 8'b10011001 : 8'b10001001;
											assign node2299 = (inp[6]) ? node2303 : node2300;
												assign node2300 = (inp[3]) ? 8'b10001001 : 8'b10001100;
												assign node2303 = (inp[12]) ? node2309 : node2304;
													assign node2304 = (inp[3]) ? 8'b10010000 : node2305;
														assign node2305 = (inp[10]) ? 8'b10010001 : 8'b10010101;
													assign node2309 = (inp[3]) ? 8'b10000001 : 8'b10000100;
										assign node2312 = (inp[10]) ? node2326 : node2313;
											assign node2313 = (inp[7]) ? 8'b10000101 : node2314;
												assign node2314 = (inp[3]) ? node2320 : node2315;
													assign node2315 = (inp[12]) ? 8'b10100000 : node2316;
														assign node2316 = (inp[6]) ? 8'b10000101 : 8'b10010101;
													assign node2320 = (inp[6]) ? node2322 : 8'b10000101;
														assign node2322 = (inp[12]) ? 8'b10010100 : 8'b10000100;
											assign node2326 = (inp[12]) ? node2330 : node2327;
												assign node2327 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node2330 = (inp[6]) ? node2334 : node2331;
													assign node2331 = (inp[3]) ? 8'b10000001 : 8'b10000100;
													assign node2334 = (inp[3]) ? 8'b10010000 : 8'b10010001;
				assign node2337 = (inp[11]) ? node2597 : node2338;
					assign node2338 = (inp[5]) ? node2528 : node2339;
						assign node2339 = (inp[9]) ? node2427 : node2340;
							assign node2340 = (inp[3]) ? node2384 : node2341;
								assign node2341 = (inp[6]) ? node2361 : node2342;
									assign node2342 = (inp[10]) ? node2350 : node2343;
										assign node2343 = (inp[2]) ? node2345 : 8'b11111101;
											assign node2345 = (inp[8]) ? node2347 : 8'b11111101;
												assign node2347 = (inp[1]) ? 8'b11110101 : 8'b11111101;
										assign node2350 = (inp[8]) ? node2356 : node2351;
											assign node2351 = (inp[7]) ? node2353 : 8'b11111101;
												assign node2353 = (inp[2]) ? 8'b10110001 : 8'b10111001;
											assign node2356 = (inp[12]) ? 8'b10111001 : node2357;
												assign node2357 = (inp[2]) ? 8'b10110001 : 8'b10111001;
									assign node2361 = (inp[10]) ? node2373 : node2362;
										assign node2362 = (inp[2]) ? node2368 : node2363;
											assign node2363 = (inp[7]) ? node2365 : 8'b11111101;
												assign node2365 = (inp[1]) ? 8'b10100101 : 8'b10101101;
											assign node2368 = (inp[1]) ? node2370 : 8'b10101101;
												assign node2370 = (inp[7]) ? 8'b10101101 : 8'b10100101;
										assign node2373 = (inp[7]) ? node2381 : node2374;
											assign node2374 = (inp[2]) ? node2378 : node2375;
												assign node2375 = (inp[8]) ? 8'b10111001 : 8'b11111101;
												assign node2378 = (inp[8]) ? 8'b10101001 : 8'b10101101;
											assign node2381 = (inp[1]) ? 8'b10100001 : 8'b10101001;
								assign node2384 = (inp[7]) ? node2414 : node2385;
									assign node2385 = (inp[1]) ? node2399 : node2386;
										assign node2386 = (inp[2]) ? node2392 : node2387;
											assign node2387 = (inp[8]) ? node2389 : 8'b11111101;
												assign node2389 = (inp[10]) ? 8'b10111001 : 8'b11111101;
											assign node2392 = (inp[6]) ? 8'b10101101 : node2393;
												assign node2393 = (inp[12]) ? 8'b11111101 : node2394;
													assign node2394 = (inp[8]) ? 8'b10111001 : 8'b11111101;
										assign node2399 = (inp[2]) ? node2405 : node2400;
											assign node2400 = (inp[8]) ? node2402 : 8'b10111100;
												assign node2402 = (inp[10]) ? 8'b10111000 : 8'b10111100;
											assign node2405 = (inp[8]) ? node2409 : node2406;
												assign node2406 = (inp[6]) ? 8'b10101100 : 8'b10111100;
												assign node2409 = (inp[6]) ? node2411 : 8'b10110100;
													assign node2411 = (inp[10]) ? 8'b10100000 : 8'b10100100;
									assign node2414 = (inp[10]) ? node2422 : node2415;
										assign node2415 = (inp[6]) ? node2419 : node2416;
											assign node2416 = (inp[2]) ? 8'b10110100 : 8'b10111100;
											assign node2419 = (inp[8]) ? 8'b10100100 : 8'b10101100;
										assign node2422 = (inp[6]) ? 8'b10100000 : node2423;
											assign node2423 = (inp[2]) ? 8'b10110000 : 8'b10111000;
							assign node2427 = (inp[8]) ? node2469 : node2428;
								assign node2428 = (inp[6]) ? node2448 : node2429;
									assign node2429 = (inp[3]) ? node2437 : node2430;
										assign node2430 = (inp[10]) ? node2432 : 8'b00011111;
											assign node2432 = (inp[7]) ? node2434 : 8'b00011111;
												assign node2434 = (inp[1]) ? 8'b10011001 : 8'b00011011;
										assign node2437 = (inp[1]) ? node2443 : node2438;
											assign node2438 = (inp[7]) ? node2440 : 8'b00011111;
												assign node2440 = (inp[10]) ? 8'b00011010 : 8'b00011110;
											assign node2443 = (inp[7]) ? node2445 : 8'b00011110;
												assign node2445 = (inp[2]) ? 8'b00011110 : 8'b00011010;
									assign node2448 = (inp[7]) ? node2458 : node2449;
										assign node2449 = (inp[2]) ? node2455 : node2450;
											assign node2450 = (inp[1]) ? node2452 : 8'b00011111;
												assign node2452 = (inp[3]) ? 8'b00011110 : 8'b00011111;
											assign node2455 = (inp[3]) ? 8'b00001110 : 8'b00001111;
										assign node2458 = (inp[10]) ? node2462 : node2459;
											assign node2459 = (inp[3]) ? 8'b00001110 : 8'b00001111;
											assign node2462 = (inp[3]) ? node2466 : node2463;
												assign node2463 = (inp[1]) ? 8'b10000001 : 8'b00001011;
												assign node2466 = (inp[12]) ? 8'b00000010 : 8'b10000010;
								assign node2469 = (inp[10]) ? node2499 : node2470;
									assign node2470 = (inp[3]) ? node2482 : node2471;
										assign node2471 = (inp[6]) ? node2477 : node2472;
											assign node2472 = (inp[2]) ? node2474 : 8'b10011101;
												assign node2474 = (inp[1]) ? 8'b10010101 : 8'b10011101;
											assign node2477 = (inp[1]) ? node2479 : 8'b10001101;
												assign node2479 = (inp[7]) ? 8'b10000101 : 8'b10011101;
										assign node2482 = (inp[6]) ? node2490 : node2483;
											assign node2483 = (inp[2]) ? node2485 : 8'b10011100;
												assign node2485 = (inp[7]) ? 8'b10010100 : node2486;
													assign node2486 = (inp[1]) ? 8'b10010100 : 8'b10011101;
											assign node2490 = (inp[7]) ? 8'b10000100 : node2491;
												assign node2491 = (inp[2]) ? node2495 : node2492;
													assign node2492 = (inp[1]) ? 8'b10011100 : 8'b10011101;
													assign node2495 = (inp[1]) ? 8'b10000100 : 8'b10001101;
									assign node2499 = (inp[3]) ? node2517 : node2500;
										assign node2500 = (inp[1]) ? node2508 : node2501;
											assign node2501 = (inp[6]) ? node2503 : 8'b00011011;
												assign node2503 = (inp[7]) ? 8'b00001011 : node2504;
													assign node2504 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node2508 = (inp[2]) ? node2514 : node2509;
												assign node2509 = (inp[6]) ? node2511 : 8'b10011001;
													assign node2511 = (inp[7]) ? 8'b10000001 : 8'b10011001;
												assign node2514 = (inp[6]) ? 8'b10000001 : 8'b10010001;
										assign node2517 = (inp[6]) ? node2521 : node2518;
											assign node2518 = (inp[2]) ? 8'b10010000 : 8'b00011010;
											assign node2521 = (inp[12]) ? node2523 : 8'b10000010;
												assign node2523 = (inp[7]) ? 8'b00000010 : node2524;
													assign node2524 = (inp[1]) ? 8'b00000010 : 8'b00001011;
						assign node2528 = (inp[7]) ? node2536 : node2529;
							assign node2529 = (inp[2]) ? node2531 : 8'b11111101;
								assign node2531 = (inp[1]) ? node2533 : 8'b11111101;
									assign node2533 = (inp[8]) ? 8'b11110101 : 8'b11111101;
							assign node2536 = (inp[8]) ? node2578 : node2537;
								assign node2537 = (inp[10]) ? node2555 : node2538;
									assign node2538 = (inp[1]) ? node2550 : node2539;
										assign node2539 = (inp[3]) ? node2545 : node2540;
											assign node2540 = (inp[6]) ? node2542 : 8'b11111101;
												assign node2542 = (inp[2]) ? 8'b11111101 : 8'b10101101;
											assign node2545 = (inp[2]) ? 8'b10111100 : node2546;
												assign node2546 = (inp[6]) ? 8'b10101100 : 8'b10111100;
										assign node2550 = (inp[2]) ? 8'b11111101 : node2551;
											assign node2551 = (inp[6]) ? 8'b10101101 : 8'b11111101;
									assign node2555 = (inp[6]) ? node2565 : node2556;
										assign node2556 = (inp[2]) ? node2562 : node2557;
											assign node2557 = (inp[1]) ? 8'b10111001 : node2558;
												assign node2558 = (inp[3]) ? 8'b10111000 : 8'b10111001;
											assign node2562 = (inp[1]) ? 8'b10110001 : 8'b10110000;
										assign node2565 = (inp[2]) ? node2573 : node2566;
											assign node2566 = (inp[3]) ? node2570 : node2567;
												assign node2567 = (inp[1]) ? 8'b10100001 : 8'b10101001;
												assign node2570 = (inp[1]) ? 8'b10100001 : 8'b10100000;
											assign node2573 = (inp[1]) ? 8'b10110001 : node2574;
												assign node2574 = (inp[3]) ? 8'b10110000 : 8'b10111001;
								assign node2578 = (inp[1]) ? node2590 : node2579;
									assign node2579 = (inp[3]) ? node2585 : node2580;
										assign node2580 = (inp[2]) ? 8'b11111101 : node2581;
											assign node2581 = (inp[6]) ? 8'b10101101 : 8'b11111101;
										assign node2585 = (inp[2]) ? 8'b10110100 : node2586;
											assign node2586 = (inp[6]) ? 8'b10100100 : 8'b10111100;
									assign node2590 = (inp[6]) ? node2594 : node2591;
										assign node2591 = (inp[2]) ? 8'b11110101 : 8'b11111101;
										assign node2594 = (inp[2]) ? 8'b11110101 : 8'b10100101;
					assign node2597 = (inp[1]) ? node2897 : node2598;
						assign node2598 = (inp[9]) ? node2750 : node2599;
							assign node2599 = (inp[8]) ? node2667 : node2600;
								assign node2600 = (inp[2]) ? node2630 : node2601;
									assign node2601 = (inp[12]) ? node2619 : node2602;
										assign node2602 = (inp[7]) ? node2604 : 8'b10101101;
											assign node2604 = (inp[6]) ? node2612 : node2605;
												assign node2605 = (inp[3]) ? node2609 : node2606;
													assign node2606 = (inp[10]) ? 8'b10101001 : 8'b10101101;
													assign node2609 = (inp[10]) ? 8'b10101000 : 8'b10101100;
												assign node2612 = (inp[3]) ? node2616 : node2613;
													assign node2613 = (inp[10]) ? 8'b10111000 : 8'b10111100;
													assign node2616 = (inp[10]) ? 8'b10010101 : 8'b10111001;
										assign node2619 = (inp[7]) ? node2621 : 8'b11111101;
											assign node2621 = (inp[10]) ? node2625 : node2622;
												assign node2622 = (inp[3]) ? 8'b10111100 : 8'b11111101;
												assign node2625 = (inp[3]) ? 8'b10111000 : node2626;
													assign node2626 = (inp[6]) ? 8'b10101001 : 8'b10111001;
									assign node2630 = (inp[7]) ? node2642 : node2631;
										assign node2631 = (inp[12]) ? node2637 : node2632;
											assign node2632 = (inp[5]) ? 8'b10101100 : node2633;
												assign node2633 = (inp[6]) ? 8'b10111100 : 8'b10101100;
											assign node2637 = (inp[6]) ? node2639 : 8'b10111100;
												assign node2639 = (inp[5]) ? 8'b10111100 : 8'b10101101;
										assign node2642 = (inp[3]) ? node2654 : node2643;
											assign node2643 = (inp[10]) ? node2649 : node2644;
												assign node2644 = (inp[12]) ? 8'b10111100 : node2645;
													assign node2645 = (inp[5]) ? 8'b10101100 : 8'b10111100;
												assign node2649 = (inp[6]) ? node2651 : 8'b10111000;
													assign node2651 = (inp[12]) ? 8'b10101001 : 8'b10101000;
											assign node2654 = (inp[10]) ? node2662 : node2655;
												assign node2655 = (inp[12]) ? 8'b10101100 : node2656;
													assign node2656 = (inp[5]) ? 8'b10101001 : node2657;
														assign node2657 = (inp[6]) ? 8'b10111001 : 8'b10101001;
												assign node2662 = (inp[12]) ? node2664 : 8'b10010101;
													assign node2664 = (inp[6]) ? 8'b10100000 : 8'b10010101;
								assign node2667 = (inp[5]) ? node2717 : node2668;
									assign node2668 = (inp[10]) ? node2690 : node2669;
										assign node2669 = (inp[7]) ? node2677 : node2670;
											assign node2670 = (inp[12]) ? node2674 : node2671;
												assign node2671 = (inp[2]) ? 8'b10001100 : 8'b10001101;
												assign node2674 = (inp[2]) ? 8'b10001101 : 8'b10011101;
											assign node2677 = (inp[3]) ? node2685 : node2678;
												assign node2678 = (inp[6]) ? node2682 : node2679;
													assign node2679 = (inp[12]) ? 8'b10011101 : 8'b10001101;
													assign node2682 = (inp[12]) ? 8'b10001101 : 8'b10011100;
												assign node2685 = (inp[6]) ? 8'b10010001 : node2686;
													assign node2686 = (inp[12]) ? 8'b10011100 : 8'b10001100;
										assign node2690 = (inp[12]) ? node2708 : node2691;
											assign node2691 = (inp[6]) ? node2701 : node2692;
												assign node2692 = (inp[2]) ? node2696 : node2693;
													assign node2693 = (inp[7]) ? 8'b10101000 : 8'b10101001;
													assign node2696 = (inp[7]) ? node2698 : 8'b10101000;
														assign node2698 = (inp[3]) ? 8'b10000101 : 8'b10101000;
												assign node2701 = (inp[3]) ? node2705 : node2702;
													assign node2702 = (inp[7]) ? 8'b10111000 : 8'b10101001;
													assign node2705 = (inp[7]) ? 8'b10010101 : 8'b10111000;
											assign node2708 = (inp[6]) ? node2712 : node2709;
												assign node2709 = (inp[3]) ? 8'b10111000 : 8'b10111001;
												assign node2712 = (inp[3]) ? node2714 : 8'b10101001;
													assign node2714 = (inp[2]) ? 8'b10101001 : 8'b10111001;
									assign node2717 = (inp[12]) ? node2735 : node2718;
										assign node2718 = (inp[6]) ? node2726 : node2719;
											assign node2719 = (inp[2]) ? 8'b10001100 : node2720;
												assign node2720 = (inp[7]) ? node2722 : 8'b10001101;
													assign node2722 = (inp[3]) ? 8'b10001100 : 8'b10001101;
											assign node2726 = (inp[7]) ? node2730 : node2727;
												assign node2727 = (inp[2]) ? 8'b10001100 : 8'b10001101;
												assign node2730 = (inp[3]) ? node2732 : 8'b10011100;
													assign node2732 = (inp[10]) ? 8'b10000001 : 8'b10010001;
										assign node2735 = (inp[2]) ? node2745 : node2736;
											assign node2736 = (inp[6]) ? node2742 : node2737;
												assign node2737 = (inp[10]) ? 8'b10011101 : node2738;
													assign node2738 = (inp[3]) ? 8'b10011100 : 8'b10011101;
												assign node2742 = (inp[7]) ? 8'b10001101 : 8'b10011101;
											assign node2745 = (inp[3]) ? node2747 : 8'b10011100;
												assign node2747 = (inp[7]) ? 8'b10010001 : 8'b10011100;
							assign node2750 = (inp[5]) ? node2846 : node2751;
								assign node2751 = (inp[8]) ? node2793 : node2752;
									assign node2752 = (inp[7]) ? node2764 : node2753;
										assign node2753 = (inp[2]) ? node2757 : node2754;
											assign node2754 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node2757 = (inp[6]) ? node2761 : node2758;
												assign node2758 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node2761 = (inp[12]) ? 8'b00001111 : 8'b00011110;
										assign node2764 = (inp[10]) ? node2784 : node2765;
											assign node2765 = (inp[3]) ? node2775 : node2766;
												assign node2766 = (inp[2]) ? node2770 : node2767;
													assign node2767 = (inp[6]) ? 8'b00011110 : 8'b00011111;
													assign node2770 = (inp[12]) ? 8'b00011110 : node2771;
														assign node2771 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node2775 = (inp[12]) ? node2779 : node2776;
													assign node2776 = (inp[6]) ? 8'b00011011 : 8'b00001110;
													assign node2779 = (inp[6]) ? 8'b00001110 : node2780;
														assign node2780 = (inp[2]) ? 8'b00011011 : 8'b00011110;
											assign node2784 = (inp[2]) ? 8'b11110111 : node2785;
												assign node2785 = (inp[6]) ? node2789 : node2786;
													assign node2786 = (inp[3]) ? 8'b00011010 : 8'b00001011;
													assign node2789 = (inp[12]) ? 8'b00000010 : 8'b00011010;
									assign node2793 = (inp[10]) ? node2823 : node2794;
										assign node2794 = (inp[7]) ? node2804 : node2795;
											assign node2795 = (inp[2]) ? node2799 : node2796;
												assign node2796 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node2799 = (inp[12]) ? node2801 : 8'b10111100;
													assign node2801 = (inp[6]) ? 8'b10101101 : 8'b10111100;
											assign node2804 = (inp[3]) ? node2812 : node2805;
												assign node2805 = (inp[2]) ? node2809 : node2806;
													assign node2806 = (inp[6]) ? 8'b10111100 : 8'b10101101;
													assign node2809 = (inp[6]) ? 8'b10101101 : 8'b10111100;
												assign node2812 = (inp[2]) ? node2816 : node2813;
													assign node2813 = (inp[6]) ? 8'b10100100 : 8'b10111100;
													assign node2816 = (inp[12]) ? node2820 : node2817;
														assign node2817 = (inp[6]) ? 8'b10110001 : 8'b10100001;
														assign node2820 = (inp[6]) ? 8'b10100100 : 8'b10110001;
										assign node2823 = (inp[2]) ? node2835 : node2824;
											assign node2824 = (inp[12]) ? node2830 : node2825;
												assign node2825 = (inp[7]) ? node2827 : 8'b00001011;
													assign node2827 = (inp[6]) ? 8'b11110111 : 8'b00001011;
												assign node2830 = (inp[6]) ? node2832 : 8'b00011011;
													assign node2832 = (inp[7]) ? 8'b00001011 : 8'b00011011;
											assign node2835 = (inp[7]) ? node2841 : node2836;
												assign node2836 = (inp[6]) ? node2838 : 8'b00011010;
													assign node2838 = (inp[3]) ? 8'b00011010 : 8'b00001011;
												assign node2841 = (inp[3]) ? node2843 : 8'b00001010;
													assign node2843 = (inp[12]) ? 8'b00000010 : 8'b10100101;
								assign node2846 = (inp[8]) ? node2872 : node2847;
									assign node2847 = (inp[12]) ? node2857 : node2848;
										assign node2848 = (inp[7]) ? node2852 : node2849;
											assign node2849 = (inp[2]) ? 8'b10101100 : 8'b10101101;
											assign node2852 = (inp[3]) ? node2854 : 8'b10101000;
												assign node2854 = (inp[10]) ? 8'b10000101 : 8'b10101001;
										assign node2857 = (inp[7]) ? node2861 : node2858;
											assign node2858 = (inp[2]) ? 8'b10111100 : 8'b11111101;
											assign node2861 = (inp[6]) ? node2867 : node2862;
												assign node2862 = (inp[2]) ? 8'b10111100 : node2863;
													assign node2863 = (inp[3]) ? 8'b10111000 : 8'b10111001;
												assign node2867 = (inp[2]) ? 8'b10111001 : node2868;
													assign node2868 = (inp[3]) ? 8'b10100000 : 8'b10101001;
									assign node2872 = (inp[12]) ? node2886 : node2873;
										assign node2873 = (inp[2]) ? node2881 : node2874;
											assign node2874 = (inp[7]) ? node2876 : 8'b10001101;
												assign node2876 = (inp[6]) ? 8'b10011100 : node2877;
													assign node2877 = (inp[3]) ? 8'b10001100 : 8'b10001101;
											assign node2881 = (inp[7]) ? node2883 : 8'b10001100;
												assign node2883 = (inp[6]) ? 8'b10000001 : 8'b10001100;
										assign node2886 = (inp[2]) ? node2892 : node2887;
											assign node2887 = (inp[7]) ? node2889 : 8'b10011101;
												assign node2889 = (inp[6]) ? 8'b10001101 : 8'b10011100;
											assign node2892 = (inp[7]) ? node2894 : 8'b10011100;
												assign node2894 = (inp[3]) ? 8'b10010001 : 8'b10011100;
						assign node2897 = (inp[8]) ? node3007 : node2898;
							assign node2898 = (inp[5]) ? node2978 : node2899;
								assign node2899 = (inp[9]) ? node2939 : node2900;
									assign node2900 = (inp[7]) ? node2920 : node2901;
										assign node2901 = (inp[12]) ? node2911 : node2902;
											assign node2902 = (inp[2]) ? node2906 : node2903;
												assign node2903 = (inp[3]) ? 8'b10101100 : 8'b10101001;
												assign node2906 = (inp[6]) ? 8'b10111001 : node2907;
													assign node2907 = (inp[3]) ? 8'b10101001 : 8'b10101000;
											assign node2911 = (inp[3]) ? node2915 : node2912;
												assign node2912 = (inp[2]) ? 8'b10111000 : 8'b10111001;
												assign node2915 = (inp[6]) ? 8'b10101100 : node2916;
													assign node2916 = (inp[2]) ? 8'b10111001 : 8'b10111100;
										assign node2920 = (inp[10]) ? node2926 : node2921;
											assign node2921 = (inp[12]) ? node2923 : 8'b10111000;
												assign node2923 = (inp[3]) ? 8'b10101100 : 8'b10101001;
											assign node2926 = (inp[6]) ? node2932 : node2927;
												assign node2927 = (inp[3]) ? node2929 : 8'b10001101;
													assign node2929 = (inp[12]) ? 8'b10010101 : 8'b10000101;
												assign node2932 = (inp[12]) ? node2936 : node2933;
													assign node2933 = (inp[2]) ? 8'b10010101 : 8'b10010100;
													assign node2936 = (inp[3]) ? 8'b10100000 : 8'b10000101;
									assign node2939 = (inp[7]) ? node2961 : node2940;
										assign node2940 = (inp[3]) ? node2950 : node2941;
											assign node2941 = (inp[2]) ? node2945 : node2942;
												assign node2942 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node2945 = (inp[12]) ? 8'b00011010 : node2946;
													assign node2946 = (inp[6]) ? 8'b00011010 : 8'b00001010;
											assign node2950 = (inp[2]) ? node2954 : node2951;
												assign node2951 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node2954 = (inp[6]) ? node2958 : node2955;
													assign node2955 = (inp[12]) ? 8'b00011011 : 8'b00001011;
													assign node2958 = (inp[12]) ? 8'b00001110 : 8'b00011011;
										assign node2961 = (inp[10]) ? node2967 : node2962;
											assign node2962 = (inp[6]) ? node2964 : 8'b00001011;
												assign node2964 = (inp[2]) ? 8'b00011010 : 8'b00011011;
											assign node2967 = (inp[2]) ? node2971 : node2968;
												assign node2968 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node2971 = (inp[6]) ? node2975 : node2972;
													assign node2972 = (inp[12]) ? 8'b10110100 : 8'b10100101;
													assign node2975 = (inp[12]) ? 8'b00000010 : 8'b11110111;
								assign node2978 = (inp[2]) ? node2996 : node2979;
									assign node2979 = (inp[7]) ? node2983 : node2980;
										assign node2980 = (inp[12]) ? 8'b10111001 : 8'b10101001;
										assign node2983 = (inp[10]) ? node2991 : node2984;
											assign node2984 = (inp[12]) ? node2988 : node2985;
												assign node2985 = (inp[6]) ? 8'b10111000 : 8'b10101001;
												assign node2988 = (inp[6]) ? 8'b10101001 : 8'b10111001;
											assign node2991 = (inp[6]) ? node2993 : 8'b10001101;
												assign node2993 = (inp[12]) ? 8'b10000101 : 8'b10010100;
									assign node2996 = (inp[12]) ? node3002 : node2997;
										assign node2997 = (inp[7]) ? node2999 : 8'b10101000;
											assign node2999 = (inp[10]) ? 8'b10000100 : 8'b10101000;
										assign node3002 = (inp[10]) ? node3004 : 8'b10111000;
											assign node3004 = (inp[7]) ? 8'b10010100 : 8'b10111000;
							assign node3007 = (inp[2]) ? node3063 : node3008;
								assign node3008 = (inp[5]) ? node3052 : node3009;
									assign node3009 = (inp[3]) ? node3027 : node3010;
										assign node3010 = (inp[9]) ? node3020 : node3011;
											assign node3011 = (inp[10]) ? node3013 : 8'b10011001;
												assign node3013 = (inp[6]) ? node3017 : node3014;
													assign node3014 = (inp[7]) ? 8'b10011101 : 8'b10001101;
													assign node3017 = (inp[12]) ? 8'b10011101 : 8'b10010100;
											assign node3020 = (inp[10]) ? node3024 : node3021;
												assign node3021 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node3024 = (inp[12]) ? 8'b11111101 : 8'b10101101;
										assign node3027 = (inp[10]) ? node3039 : node3028;
											assign node3028 = (inp[9]) ? node3032 : node3029;
												assign node3029 = (inp[12]) ? 8'b10011100 : 8'b10001100;
												assign node3032 = (inp[6]) ? node3036 : node3033;
													assign node3033 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node3036 = (inp[7]) ? 8'b10110001 : 8'b10101100;
											assign node3039 = (inp[9]) ? node3045 : node3040;
												assign node3040 = (inp[6]) ? 8'b10100000 : node3041;
													assign node3041 = (inp[12]) ? 8'b10111000 : 8'b10101000;
												assign node3045 = (inp[7]) ? node3047 : 8'b00011010;
													assign node3047 = (inp[6]) ? 8'b00000010 : node3048;
														assign node3048 = (inp[12]) ? 8'b00011010 : 8'b00001010;
									assign node3052 = (inp[7]) ? node3056 : node3053;
										assign node3053 = (inp[12]) ? 8'b10011001 : 8'b10001001;
										assign node3056 = (inp[6]) ? node3060 : node3057;
											assign node3057 = (inp[12]) ? 8'b10011001 : 8'b10001001;
											assign node3060 = (inp[12]) ? 8'b10000001 : 8'b10010000;
								assign node3063 = (inp[5]) ? node3121 : node3064;
									assign node3064 = (inp[9]) ? node3096 : node3065;
										assign node3065 = (inp[10]) ? node3081 : node3066;
											assign node3066 = (inp[3]) ? node3074 : node3067;
												assign node3067 = (inp[6]) ? node3071 : node3068;
													assign node3068 = (inp[12]) ? 8'b10010000 : 8'b10000000;
													assign node3071 = (inp[12]) ? 8'b10000001 : 8'b10010000;
												assign node3074 = (inp[6]) ? node3078 : node3075;
													assign node3075 = (inp[7]) ? 8'b10000001 : 8'b10010001;
													assign node3078 = (inp[12]) ? 8'b10000100 : 8'b10010001;
											assign node3081 = (inp[3]) ? node3089 : node3082;
												assign node3082 = (inp[7]) ? 8'b10010100 : node3083;
													assign node3083 = (inp[12]) ? 8'b10010100 : node3084;
														assign node3084 = (inp[6]) ? 8'b10010100 : 8'b10000100;
												assign node3089 = (inp[6]) ? node3093 : node3090;
													assign node3090 = (inp[7]) ? 8'b10000101 : 8'b10010101;
													assign node3093 = (inp[12]) ? 8'b10100000 : 8'b10010101;
										assign node3096 = (inp[10]) ? node3110 : node3097;
											assign node3097 = (inp[3]) ? node3105 : node3098;
												assign node3098 = (inp[12]) ? node3102 : node3099;
													assign node3099 = (inp[6]) ? 8'b10110000 : 8'b10100000;
													assign node3102 = (inp[6]) ? 8'b10100001 : 8'b10110000;
												assign node3105 = (inp[6]) ? 8'b10110001 : node3106;
													assign node3106 = (inp[12]) ? 8'b10110001 : 8'b10100001;
											assign node3110 = (inp[3]) ? node3118 : node3111;
												assign node3111 = (inp[7]) ? node3113 : 8'b10100100;
													assign node3113 = (inp[6]) ? 8'b10110100 : node3114;
														assign node3114 = (inp[12]) ? 8'b10110100 : 8'b10100100;
												assign node3118 = (inp[6]) ? 8'b11110111 : 8'b10100101;
									assign node3121 = (inp[12]) ? 8'b10010000 : 8'b10000000;
		assign node3124 = (inp[7]) ? node5362 : node3125;
			assign node3125 = (inp[13]) ? node4277 : node3126;
				assign node3126 = (inp[9]) ? node3730 : node3127;
					assign node3127 = (inp[8]) ? node3443 : node3128;
						assign node3128 = (inp[10]) ? node3286 : node3129;
							assign node3129 = (inp[1]) ? node3195 : node3130;
								assign node3130 = (inp[3]) ? node3164 : node3131;
									assign node3131 = (inp[11]) ? node3145 : node3132;
										assign node3132 = (inp[6]) ? node3138 : node3133;
											assign node3133 = (inp[12]) ? node3135 : 8'b10000010;
												assign node3135 = (inp[0]) ? 8'b10010000 : 8'b00000010;
											assign node3138 = (inp[2]) ? node3140 : 8'b00011010;
												assign node3140 = (inp[5]) ? 8'b10010000 : node3141;
													assign node3141 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node3145 = (inp[5]) ? node3155 : node3146;
											assign node3146 = (inp[12]) ? node3150 : node3147;
												assign node3147 = (inp[6]) ? 8'b00001010 : 8'b11110111;
												assign node3150 = (inp[2]) ? 8'b00000010 : node3151;
													assign node3151 = (inp[6]) ? 8'b00011010 : 8'b00000010;
											assign node3155 = (inp[6]) ? 8'b11110101 : node3156;
												assign node3156 = (inp[12]) ? node3158 : 8'b11110111;
													assign node3158 = (inp[2]) ? node3160 : 8'b00000010;
														assign node3160 = (inp[0]) ? 8'b11110101 : 8'b00000010;
									assign node3164 = (inp[11]) ? node3176 : node3165;
										assign node3165 = (inp[6]) ? node3171 : node3166;
											assign node3166 = (inp[2]) ? node3168 : 8'b00001011;
												assign node3168 = (inp[0]) ? 8'b00011011 : 8'b00001011;
											assign node3171 = (inp[5]) ? 8'b00011011 : node3172;
												assign node3172 = (inp[2]) ? 8'b00001011 : 8'b00011011;
										assign node3176 = (inp[2]) ? node3188 : node3177;
											assign node3177 = (inp[0]) ? node3183 : node3178;
												assign node3178 = (inp[6]) ? node3180 : 8'b00001011;
													assign node3180 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node3183 = (inp[12]) ? node3185 : 8'b00011010;
													assign node3185 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node3188 = (inp[12]) ? node3192 : node3189;
												assign node3189 = (inp[0]) ? 8'b00001010 : 8'b00011010;
												assign node3192 = (inp[0]) ? 8'b00011010 : 8'b00001011;
								assign node3195 = (inp[11]) ? node3235 : node3196;
									assign node3196 = (inp[0]) ? node3216 : node3197;
										assign node3197 = (inp[6]) ? node3205 : node3198;
											assign node3198 = (inp[12]) ? 8'b00000010 : node3199;
												assign node3199 = (inp[3]) ? node3201 : 8'b10000010;
													assign node3201 = (inp[5]) ? 8'b10000001 : 8'b10000010;
											assign node3205 = (inp[2]) ? node3211 : node3206;
												assign node3206 = (inp[3]) ? node3208 : 8'b00011010;
													assign node3208 = (inp[5]) ? 8'b10011001 : 8'b00011010;
												assign node3211 = (inp[5]) ? 8'b10010001 : node3212;
													assign node3212 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node3216 = (inp[3]) ? node3224 : node3217;
											assign node3217 = (inp[6]) ? node3221 : node3218;
												assign node3218 = (inp[2]) ? 8'b10010001 : 8'b10000001;
												assign node3221 = (inp[2]) ? 8'b10000001 : 8'b10011001;
											assign node3224 = (inp[5]) ? node3232 : node3225;
												assign node3225 = (inp[6]) ? node3229 : node3226;
													assign node3226 = (inp[2]) ? 8'b10010000 : 8'b10000010;
													assign node3229 = (inp[2]) ? 8'b00000010 : 8'b00011010;
												assign node3232 = (inp[6]) ? 8'b10011001 : 8'b10010001;
									assign node3235 = (inp[5]) ? node3265 : node3236;
										assign node3236 = (inp[2]) ? node3250 : node3237;
											assign node3237 = (inp[3]) ? node3243 : node3238;
												assign node3238 = (inp[0]) ? node3240 : 8'b00011010;
													assign node3240 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node3243 = (inp[6]) ? node3247 : node3244;
													assign node3244 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node3247 = (inp[12]) ? 8'b00011010 : 8'b00001010;
											assign node3250 = (inp[0]) ? node3254 : node3251;
												assign node3251 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node3254 = (inp[3]) ? node3262 : node3255;
													assign node3255 = (inp[6]) ? node3259 : node3256;
														assign node3256 = (inp[12]) ? 8'b10110100 : 8'b10100100;
														assign node3259 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node3262 = (inp[6]) ? 8'b11110111 : 8'b11110101;
										assign node3265 = (inp[2]) ? node3277 : node3266;
											assign node3266 = (inp[6]) ? node3272 : node3267;
												assign node3267 = (inp[12]) ? 8'b10100101 : node3268;
													assign node3268 = (inp[3]) ? 8'b10110100 : 8'b11110111;
												assign node3272 = (inp[3]) ? node3274 : 8'b00001010;
													assign node3274 = (inp[12]) ? 8'b11111101 : 8'b10101101;
											assign node3277 = (inp[0]) ? node3283 : node3278;
												assign node3278 = (inp[3]) ? node3280 : 8'b11110111;
													assign node3280 = (inp[6]) ? 8'b10110100 : 8'b10100101;
												assign node3283 = (inp[12]) ? 8'b10110100 : 8'b10100100;
							assign node3286 = (inp[11]) ? node3356 : node3287;
								assign node3287 = (inp[6]) ? node3323 : node3288;
									assign node3288 = (inp[2]) ? node3306 : node3289;
										assign node3289 = (inp[5]) ? node3299 : node3290;
											assign node3290 = (inp[0]) ? node3292 : 8'b00001110;
												assign node3292 = (inp[1]) ? node3296 : node3293;
													assign node3293 = (inp[3]) ? 8'b00001111 : 8'b00001110;
													assign node3296 = (inp[3]) ? 8'b00001110 : 8'b00001111;
											assign node3299 = (inp[3]) ? 8'b00001111 : node3300;
												assign node3300 = (inp[0]) ? node3302 : 8'b00001110;
													assign node3302 = (inp[1]) ? 8'b00001111 : 8'b00001110;
										assign node3306 = (inp[0]) ? node3314 : node3307;
											assign node3307 = (inp[3]) ? node3309 : 8'b00001110;
												assign node3309 = (inp[5]) ? 8'b00001111 : node3310;
													assign node3310 = (inp[1]) ? 8'b00001110 : 8'b00001111;
											assign node3314 = (inp[1]) ? node3318 : node3315;
												assign node3315 = (inp[3]) ? 8'b00011111 : 8'b00011110;
												assign node3318 = (inp[3]) ? node3320 : 8'b00011111;
													assign node3320 = (inp[5]) ? 8'b00011111 : 8'b00011110;
									assign node3323 = (inp[5]) ? node3349 : node3324;
										assign node3324 = (inp[2]) ? node3336 : node3325;
											assign node3325 = (inp[12]) ? node3331 : node3326;
												assign node3326 = (inp[3]) ? node3328 : 8'b00011111;
													assign node3328 = (inp[1]) ? 8'b00011110 : 8'b00011111;
												assign node3331 = (inp[1]) ? 8'b00011110 : node3332;
													assign node3332 = (inp[3]) ? 8'b00011111 : 8'b00011110;
											assign node3336 = (inp[12]) ? node3342 : node3337;
												assign node3337 = (inp[3]) ? node3339 : 8'b00001110;
													assign node3339 = (inp[1]) ? 8'b00001110 : 8'b00001111;
												assign node3342 = (inp[1]) ? node3346 : node3343;
													assign node3343 = (inp[3]) ? 8'b00001111 : 8'b00001110;
													assign node3346 = (inp[3]) ? 8'b00001110 : 8'b00001111;
										assign node3349 = (inp[3]) ? 8'b00011111 : node3350;
											assign node3350 = (inp[0]) ? node3352 : 8'b00011110;
												assign node3352 = (inp[1]) ? 8'b00011111 : 8'b00011110;
								assign node3356 = (inp[1]) ? node3396 : node3357;
									assign node3357 = (inp[3]) ? node3375 : node3358;
										assign node3358 = (inp[2]) ? node3366 : node3359;
											assign node3359 = (inp[5]) ? 8'b00001110 : node3360;
												assign node3360 = (inp[12]) ? node3362 : 8'b00011011;
													assign node3362 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node3366 = (inp[12]) ? node3372 : node3367;
												assign node3367 = (inp[5]) ? 8'b00001011 : node3368;
													assign node3368 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node3372 = (inp[0]) ? 8'b00011011 : 8'b00001110;
										assign node3375 = (inp[12]) ? node3383 : node3376;
											assign node3376 = (inp[6]) ? node3378 : 8'b00011110;
												assign node3378 = (inp[5]) ? node3380 : 8'b00011110;
													assign node3380 = (inp[2]) ? 8'b00001110 : 8'b00001111;
											assign node3383 = (inp[6]) ? node3389 : node3384;
												assign node3384 = (inp[2]) ? node3386 : 8'b00001111;
													assign node3386 = (inp[0]) ? 8'b00011110 : 8'b00001111;
												assign node3389 = (inp[5]) ? node3393 : node3390;
													assign node3390 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node3393 = (inp[2]) ? 8'b00011110 : 8'b00011111;
									assign node3396 = (inp[0]) ? node3420 : node3397;
										assign node3397 = (inp[12]) ? node3411 : node3398;
											assign node3398 = (inp[5]) ? node3400 : 8'b00011011;
												assign node3400 = (inp[6]) ? node3404 : node3401;
													assign node3401 = (inp[3]) ? 8'b00011010 : 8'b00011011;
													assign node3404 = (inp[3]) ? node3408 : node3405;
														assign node3405 = (inp[2]) ? 8'b00001011 : 8'b00001110;
														assign node3408 = (inp[2]) ? 8'b00001010 : 8'b00001011;
											assign node3411 = (inp[5]) ? node3417 : node3412;
												assign node3412 = (inp[6]) ? node3414 : 8'b00001110;
													assign node3414 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node3417 = (inp[6]) ? 8'b00011011 : 8'b00001011;
										assign node3420 = (inp[5]) ? node3436 : node3421;
											assign node3421 = (inp[2]) ? node3427 : node3422;
												assign node3422 = (inp[3]) ? 8'b00011011 : node3423;
													assign node3423 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node3427 = (inp[3]) ? node3431 : node3428;
													assign node3428 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node3431 = (inp[6]) ? node3433 : 8'b00011011;
														assign node3433 = (inp[12]) ? 8'b00001110 : 8'b00011011;
											assign node3436 = (inp[12]) ? node3440 : node3437;
												assign node3437 = (inp[2]) ? 8'b00001010 : 8'b00011010;
												assign node3440 = (inp[2]) ? 8'b00011010 : 8'b00011011;
						assign node3443 = (inp[0]) ? node3569 : node3444;
							assign node3444 = (inp[5]) ? node3488 : node3445;
								assign node3445 = (inp[1]) ? node3473 : node3446;
									assign node3446 = (inp[3]) ? node3456 : node3447;
										assign node3447 = (inp[6]) ? node3451 : node3448;
											assign node3448 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node3451 = (inp[2]) ? 8'b10000010 : node3452;
												assign node3452 = (inp[11]) ? 8'b00001010 : 8'b00011010;
										assign node3456 = (inp[12]) ? node3468 : node3457;
											assign node3457 = (inp[11]) ? node3463 : node3458;
												assign node3458 = (inp[2]) ? 8'b00001011 : node3459;
													assign node3459 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node3463 = (inp[2]) ? 8'b00011010 : node3464;
													assign node3464 = (inp[6]) ? 8'b00001011 : 8'b00011010;
											assign node3468 = (inp[2]) ? 8'b00001011 : node3469;
												assign node3469 = (inp[6]) ? 8'b00011011 : 8'b00001011;
									assign node3473 = (inp[12]) ? node3483 : node3474;
										assign node3474 = (inp[11]) ? node3478 : node3475;
											assign node3475 = (inp[10]) ? 8'b10000010 : 8'b00011010;
											assign node3478 = (inp[6]) ? node3480 : 8'b11110111;
												assign node3480 = (inp[2]) ? 8'b11110111 : 8'b00001010;
										assign node3483 = (inp[2]) ? 8'b00000010 : node3484;
											assign node3484 = (inp[6]) ? 8'b00011010 : 8'b00000010;
								assign node3488 = (inp[10]) ? node3526 : node3489;
									assign node3489 = (inp[6]) ? node3503 : node3490;
										assign node3490 = (inp[12]) ? node3498 : node3491;
											assign node3491 = (inp[11]) ? node3495 : node3492;
												assign node3492 = (inp[3]) ? 8'b10000001 : 8'b10000010;
												assign node3495 = (inp[3]) ? 8'b00011010 : 8'b11110111;
											assign node3498 = (inp[3]) ? node3500 : 8'b00000010;
												assign node3500 = (inp[1]) ? 8'b10100101 : 8'b00001011;
										assign node3503 = (inp[2]) ? node3513 : node3504;
											assign node3504 = (inp[3]) ? node3510 : node3505;
												assign node3505 = (inp[12]) ? 8'b00011010 : node3506;
													assign node3506 = (inp[11]) ? 8'b00001010 : 8'b00011010;
												assign node3510 = (inp[1]) ? 8'b10011001 : 8'b00011011;
											assign node3513 = (inp[12]) ? node3519 : node3514;
												assign node3514 = (inp[11]) ? node3516 : 8'b10010001;
													assign node3516 = (inp[3]) ? 8'b10100100 : 8'b10100101;
												assign node3519 = (inp[1]) ? 8'b10110100 : node3520;
													assign node3520 = (inp[3]) ? node3522 : 8'b10010000;
														assign node3522 = (inp[11]) ? 8'b00011010 : 8'b00011011;
									assign node3526 = (inp[11]) ? node3540 : node3527;
										assign node3527 = (inp[3]) ? node3533 : node3528;
											assign node3528 = (inp[6]) ? node3530 : 8'b10000100;
												assign node3530 = (inp[1]) ? 8'b10010100 : 8'b10011100;
											assign node3533 = (inp[6]) ? node3537 : node3534;
												assign node3534 = (inp[1]) ? 8'b10000101 : 8'b10001101;
												assign node3537 = (inp[2]) ? 8'b10010101 : 8'b10011101;
										assign node3540 = (inp[1]) ? node3556 : node3541;
											assign node3541 = (inp[3]) ? node3549 : node3542;
												assign node3542 = (inp[6]) ? node3544 : 8'b10110001;
													assign node3544 = (inp[2]) ? 8'b10110001 : node3545;
														assign node3545 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node3549 = (inp[2]) ? node3551 : 8'b10101101;
													assign node3551 = (inp[6]) ? node3553 : 8'b10111100;
														assign node3553 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node3556 = (inp[12]) ? node3564 : node3557;
												assign node3557 = (inp[6]) ? node3561 : node3558;
													assign node3558 = (inp[3]) ? 8'b10110000 : 8'b10110001;
													assign node3561 = (inp[2]) ? 8'b10100000 : 8'b10101001;
												assign node3564 = (inp[6]) ? node3566 : 8'b10100100;
													assign node3566 = (inp[3]) ? 8'b10110000 : 8'b10111100;
							assign node3569 = (inp[11]) ? node3627 : node3570;
								assign node3570 = (inp[5]) ? node3606 : node3571;
									assign node3571 = (inp[10]) ? node3589 : node3572;
										assign node3572 = (inp[1]) ? node3584 : node3573;
											assign node3573 = (inp[3]) ? node3579 : node3574;
												assign node3574 = (inp[2]) ? 8'b10000100 : node3575;
													assign node3575 = (inp[6]) ? 8'b10011100 : 8'b10000100;
												assign node3579 = (inp[2]) ? node3581 : 8'b10011101;
													assign node3581 = (inp[6]) ? 8'b10001101 : 8'b10011101;
											assign node3584 = (inp[3]) ? 8'b10000100 : node3585;
												assign node3585 = (inp[2]) ? 8'b10010101 : 8'b10000101;
										assign node3589 = (inp[1]) ? node3595 : node3590;
											assign node3590 = (inp[12]) ? 8'b00000010 : node3591;
												assign node3591 = (inp[6]) ? 8'b00011010 : 8'b00011011;
											assign node3595 = (inp[3]) ? node3603 : node3596;
												assign node3596 = (inp[6]) ? node3600 : node3597;
													assign node3597 = (inp[2]) ? 8'b10010001 : 8'b10000001;
													assign node3600 = (inp[2]) ? 8'b10000001 : 8'b10011001;
												assign node3603 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node3606 = (inp[6]) ? node3618 : node3607;
										assign node3607 = (inp[2]) ? node3613 : node3608;
											assign node3608 = (inp[1]) ? 8'b10000101 : node3609;
												assign node3609 = (inp[3]) ? 8'b10001101 : 8'b10000100;
											assign node3613 = (inp[1]) ? 8'b10010101 : node3614;
												assign node3614 = (inp[3]) ? 8'b10011101 : 8'b10010100;
										assign node3618 = (inp[2]) ? node3624 : node3619;
											assign node3619 = (inp[3]) ? 8'b10011101 : node3620;
												assign node3620 = (inp[1]) ? 8'b10011101 : 8'b10011100;
											assign node3624 = (inp[1]) ? 8'b10010101 : 8'b10011101;
								assign node3627 = (inp[1]) ? node3679 : node3628;
									assign node3628 = (inp[3]) ? node3654 : node3629;
										assign node3629 = (inp[2]) ? node3639 : node3630;
											assign node3630 = (inp[10]) ? node3634 : node3631;
												assign node3631 = (inp[6]) ? 8'b10111100 : 8'b10100100;
												assign node3634 = (inp[12]) ? node3636 : 8'b11110111;
													assign node3636 = (inp[6]) ? 8'b00011010 : 8'b00000010;
											assign node3639 = (inp[5]) ? node3651 : node3640;
												assign node3640 = (inp[12]) ? node3646 : node3641;
													assign node3641 = (inp[10]) ? node3643 : 8'b10110001;
														assign node3643 = (inp[6]) ? 8'b11110111 : 8'b10100101;
													assign node3646 = (inp[10]) ? 8'b00000010 : node3647;
														assign node3647 = (inp[6]) ? 8'b10100100 : 8'b10110001;
												assign node3651 = (inp[12]) ? 8'b10110001 : 8'b10100001;
										assign node3654 = (inp[5]) ? node3670 : node3655;
											assign node3655 = (inp[10]) ? node3663 : node3656;
												assign node3656 = (inp[2]) ? node3658 : 8'b10101101;
													assign node3658 = (inp[12]) ? 8'b10111100 : node3659;
														assign node3659 = (inp[6]) ? 8'b10111100 : 8'b10101100;
												assign node3663 = (inp[12]) ? node3665 : 8'b00011010;
													assign node3665 = (inp[2]) ? 8'b00001011 : node3666;
														assign node3666 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node3670 = (inp[12]) ? node3676 : node3671;
												assign node3671 = (inp[2]) ? 8'b10101100 : node3672;
													assign node3672 = (inp[6]) ? 8'b10101101 : 8'b10111100;
												assign node3676 = (inp[2]) ? 8'b10111100 : 8'b11111101;
									assign node3679 = (inp[10]) ? node3703 : node3680;
										assign node3680 = (inp[2]) ? node3692 : node3681;
											assign node3681 = (inp[6]) ? node3689 : node3682;
												assign node3682 = (inp[12]) ? node3684 : 8'b10110000;
													assign node3684 = (inp[3]) ? node3686 : 8'b10100001;
														assign node3686 = (inp[5]) ? 8'b10100001 : 8'b10100100;
												assign node3689 = (inp[12]) ? 8'b10111001 : 8'b10101001;
											assign node3692 = (inp[5]) ? node3700 : node3693;
												assign node3693 = (inp[12]) ? 8'b10100001 : node3694;
													assign node3694 = (inp[3]) ? node3696 : 8'b10110000;
														assign node3696 = (inp[6]) ? 8'b10110001 : 8'b10100001;
												assign node3700 = (inp[12]) ? 8'b10110000 : 8'b10100000;
										assign node3703 = (inp[5]) ? node3723 : node3704;
											assign node3704 = (inp[3]) ? node3716 : node3705;
												assign node3705 = (inp[12]) ? node3711 : node3706;
													assign node3706 = (inp[2]) ? node3708 : 8'b10110100;
														assign node3708 = (inp[6]) ? 8'b10110100 : 8'b10100100;
													assign node3711 = (inp[6]) ? 8'b10100101 : node3712;
														assign node3712 = (inp[2]) ? 8'b10110100 : 8'b10100101;
												assign node3716 = (inp[6]) ? node3720 : node3717;
													assign node3717 = (inp[12]) ? 8'b11110101 : 8'b11110111;
													assign node3720 = (inp[2]) ? 8'b00000010 : 8'b00001010;
											assign node3723 = (inp[12]) ? node3727 : node3724;
												assign node3724 = (inp[2]) ? 8'b10100000 : 8'b10110000;
												assign node3727 = (inp[2]) ? 8'b10110000 : 8'b10100001;
					assign node3730 = (inp[11]) ? node3934 : node3731;
						assign node3731 = (inp[10]) ? node3837 : node3732;
							assign node3732 = (inp[0]) ? node3756 : node3733;
								assign node3733 = (inp[3]) ? node3741 : node3734;
									assign node3734 = (inp[6]) ? node3736 : 8'b00101010;
										assign node3736 = (inp[5]) ? 8'b00111010 : node3737;
											assign node3737 = (inp[2]) ? 8'b00101010 : 8'b00111010;
									assign node3741 = (inp[6]) ? node3747 : node3742;
										assign node3742 = (inp[1]) ? node3744 : 8'b00101011;
											assign node3744 = (inp[5]) ? 8'b00101011 : 8'b00101010;
										assign node3747 = (inp[5]) ? 8'b00111011 : node3748;
											assign node3748 = (inp[1]) ? node3752 : node3749;
												assign node3749 = (inp[2]) ? 8'b00101011 : 8'b00111011;
												assign node3752 = (inp[2]) ? 8'b00101010 : 8'b00111010;
								assign node3756 = (inp[8]) ? node3808 : node3757;
									assign node3757 = (inp[5]) ? node3793 : node3758;
										assign node3758 = (inp[12]) ? node3782 : node3759;
											assign node3759 = (inp[6]) ? node3769 : node3760;
												assign node3760 = (inp[2]) ? node3764 : node3761;
													assign node3761 = (inp[1]) ? 8'b00101011 : 8'b00101010;
													assign node3764 = (inp[3]) ? node3766 : 8'b00111010;
														assign node3766 = (inp[1]) ? 8'b00111010 : 8'b00111011;
												assign node3769 = (inp[2]) ? node3777 : node3770;
													assign node3770 = (inp[3]) ? node3774 : node3771;
														assign node3771 = (inp[1]) ? 8'b00111011 : 8'b00111010;
														assign node3774 = (inp[1]) ? 8'b00111010 : 8'b00111011;
													assign node3777 = (inp[3]) ? node3779 : 8'b00101011;
														assign node3779 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node3782 = (inp[1]) ? node3786 : node3783;
												assign node3783 = (inp[3]) ? 8'b00101011 : 8'b00101010;
												assign node3786 = (inp[3]) ? node3788 : 8'b00101011;
													assign node3788 = (inp[6]) ? node3790 : 8'b00101010;
														assign node3790 = (inp[2]) ? 8'b00101010 : 8'b00111010;
										assign node3793 = (inp[3]) ? node3803 : node3794;
											assign node3794 = (inp[1]) ? node3800 : node3795;
												assign node3795 = (inp[6]) ? 8'b00111010 : node3796;
													assign node3796 = (inp[2]) ? 8'b00111010 : 8'b00101010;
												assign node3800 = (inp[2]) ? 8'b00111011 : 8'b00101011;
											assign node3803 = (inp[6]) ? 8'b00111011 : node3804;
												assign node3804 = (inp[2]) ? 8'b00111011 : 8'b00101011;
									assign node3808 = (inp[5]) ? node3830 : node3809;
										assign node3809 = (inp[2]) ? node3817 : node3810;
											assign node3810 = (inp[6]) ? 8'b01111111 : node3811;
												assign node3811 = (inp[3]) ? 8'b00101111 : node3812;
													assign node3812 = (inp[1]) ? 8'b00101111 : 8'b00101110;
											assign node3817 = (inp[6]) ? node3825 : node3818;
												assign node3818 = (inp[1]) ? node3822 : node3819;
													assign node3819 = (inp[3]) ? 8'b01111111 : 8'b00111110;
													assign node3822 = (inp[3]) ? 8'b00111110 : 8'b01111111;
												assign node3825 = (inp[3]) ? 8'b00101110 : node3826;
													assign node3826 = (inp[1]) ? 8'b00101111 : 8'b00101110;
										assign node3830 = (inp[1]) ? 8'b01111111 : node3831;
											assign node3831 = (inp[3]) ? node3833 : 8'b00111110;
												assign node3833 = (inp[2]) ? 8'b01111111 : 8'b00101111;
							assign node3837 = (inp[3]) ? node3881 : node3838;
								assign node3838 = (inp[0]) ? node3854 : node3839;
									assign node3839 = (inp[6]) ? node3845 : node3840;
										assign node3840 = (inp[5]) ? 8'b00101110 : node3841;
											assign node3841 = (inp[8]) ? 8'b00101010 : 8'b00101110;
										assign node3845 = (inp[5]) ? 8'b00111110 : node3846;
											assign node3846 = (inp[2]) ? node3850 : node3847;
												assign node3847 = (inp[8]) ? 8'b00111010 : 8'b00111110;
												assign node3850 = (inp[8]) ? 8'b00101010 : 8'b00101110;
									assign node3854 = (inp[1]) ? node3866 : node3855;
										assign node3855 = (inp[5]) ? node3861 : node3856;
											assign node3856 = (inp[2]) ? 8'b00101010 : node3857;
												assign node3857 = (inp[8]) ? 8'b00111010 : 8'b00111110;
											assign node3861 = (inp[6]) ? 8'b00111110 : node3862;
												assign node3862 = (inp[2]) ? 8'b00111110 : 8'b00101110;
										assign node3866 = (inp[6]) ? node3874 : node3867;
											assign node3867 = (inp[2]) ? 8'b01111111 : node3868;
												assign node3868 = (inp[8]) ? node3870 : 8'b00101111;
													assign node3870 = (inp[5]) ? 8'b00101111 : 8'b00101011;
											assign node3874 = (inp[2]) ? node3876 : 8'b01111111;
												assign node3876 = (inp[5]) ? 8'b01111111 : node3877;
													assign node3877 = (inp[8]) ? 8'b00101011 : 8'b00101111;
								assign node3881 = (inp[5]) ? node3927 : node3882;
									assign node3882 = (inp[8]) ? node3902 : node3883;
										assign node3883 = (inp[1]) ? node3895 : node3884;
											assign node3884 = (inp[12]) ? node3886 : 8'b00101111;
												assign node3886 = (inp[0]) ? node3890 : node3887;
													assign node3887 = (inp[2]) ? 8'b00101111 : 8'b01111111;
													assign node3890 = (inp[2]) ? node3892 : 8'b00101111;
														assign node3892 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node3895 = (inp[0]) ? node3897 : 8'b00101110;
												assign node3897 = (inp[6]) ? 8'b00101110 : node3898;
													assign node3898 = (inp[2]) ? 8'b00111110 : 8'b00101110;
										assign node3902 = (inp[1]) ? node3918 : node3903;
											assign node3903 = (inp[0]) ? node3905 : 8'b00101011;
												assign node3905 = (inp[12]) ? node3913 : node3906;
													assign node3906 = (inp[2]) ? node3910 : node3907;
														assign node3907 = (inp[6]) ? 8'b00111011 : 8'b00101011;
														assign node3910 = (inp[6]) ? 8'b00101011 : 8'b00111011;
													assign node3913 = (inp[6]) ? 8'b00101011 : node3914;
														assign node3914 = (inp[2]) ? 8'b00111011 : 8'b00101011;
											assign node3918 = (inp[12]) ? node3920 : 8'b00101010;
												assign node3920 = (inp[6]) ? node3924 : node3921;
													assign node3921 = (inp[2]) ? 8'b00111010 : 8'b00101010;
													assign node3924 = (inp[0]) ? 8'b00101010 : 8'b00111010;
									assign node3927 = (inp[6]) ? 8'b01111111 : node3928;
										assign node3928 = (inp[2]) ? node3930 : 8'b00101111;
											assign node3930 = (inp[0]) ? 8'b01111111 : 8'b00101111;
						assign node3934 = (inp[8]) ? node4118 : node3935;
							assign node3935 = (inp[10]) ? node4025 : node3936;
								assign node3936 = (inp[1]) ? node3976 : node3937;
									assign node3937 = (inp[3]) ? node3955 : node3938;
										assign node3938 = (inp[2]) ? node3944 : node3939;
											assign node3939 = (inp[6]) ? 8'b00101010 : node3940;
												assign node3940 = (inp[12]) ? 8'b00101010 : 8'b00011111;
											assign node3944 = (inp[12]) ? node3950 : node3945;
												assign node3945 = (inp[0]) ? 8'b00001111 : node3946;
													assign node3946 = (inp[5]) ? 8'b00001111 : 8'b00011111;
												assign node3950 = (inp[5]) ? 8'b00011111 : node3951;
													assign node3951 = (inp[0]) ? 8'b00011111 : 8'b00101010;
										assign node3955 = (inp[12]) ? node3967 : node3956;
											assign node3956 = (inp[6]) ? node3962 : node3957;
												assign node3957 = (inp[2]) ? node3959 : 8'b00111010;
													assign node3959 = (inp[0]) ? 8'b00101010 : 8'b00111010;
												assign node3962 = (inp[2]) ? node3964 : 8'b00101011;
													assign node3964 = (inp[5]) ? 8'b00101010 : 8'b00111010;
											assign node3967 = (inp[6]) ? node3969 : 8'b00101011;
												assign node3969 = (inp[5]) ? node3973 : node3970;
													assign node3970 = (inp[2]) ? 8'b00101011 : 8'b00111011;
													assign node3973 = (inp[2]) ? 8'b00111010 : 8'b00111011;
									assign node3976 = (inp[5]) ? node4006 : node3977;
										assign node3977 = (inp[12]) ? node3989 : node3978;
											assign node3978 = (inp[6]) ? node3984 : node3979;
												assign node3979 = (inp[0]) ? node3981 : 8'b00011111;
													assign node3981 = (inp[2]) ? 8'b00001111 : 8'b00011111;
												assign node3984 = (inp[3]) ? 8'b00101010 : node3985;
													assign node3985 = (inp[0]) ? 8'b00011110 : 8'b00011111;
											assign node3989 = (inp[0]) ? node3995 : node3990;
												assign node3990 = (inp[2]) ? 8'b00101010 : node3991;
													assign node3991 = (inp[6]) ? 8'b00111010 : 8'b00101010;
												assign node3995 = (inp[3]) ? node4001 : node3996;
													assign node3996 = (inp[6]) ? node3998 : 8'b00011110;
														assign node3998 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node4001 = (inp[6]) ? node4003 : 8'b00011111;
														assign node4003 = (inp[2]) ? 8'b00101010 : 8'b00111010;
										assign node4006 = (inp[6]) ? node4014 : node4007;
											assign node4007 = (inp[3]) ? node4011 : node4008;
												assign node4008 = (inp[0]) ? 8'b00001111 : 8'b00101010;
												assign node4011 = (inp[12]) ? 8'b00001111 : 8'b00001110;
											assign node4014 = (inp[12]) ? node4020 : node4015;
												assign node4015 = (inp[2]) ? node4017 : 8'b00001111;
													assign node4017 = (inp[3]) ? 8'b00001110 : 8'b00001111;
												assign node4020 = (inp[2]) ? node4022 : 8'b00011111;
													assign node4022 = (inp[0]) ? 8'b00011110 : 8'b00011111;
								assign node4025 = (inp[1]) ? node4063 : node4026;
									assign node4026 = (inp[3]) ? node4042 : node4027;
										assign node4027 = (inp[2]) ? node4035 : node4028;
											assign node4028 = (inp[6]) ? node4032 : node4029;
												assign node4029 = (inp[12]) ? 8'b00101110 : 8'b00111011;
												assign node4032 = (inp[12]) ? 8'b00111110 : 8'b00101110;
											assign node4035 = (inp[0]) ? node4039 : node4036;
												assign node4036 = (inp[12]) ? 8'b00101110 : 8'b00111011;
												assign node4039 = (inp[12]) ? 8'b00111011 : 8'b00101011;
										assign node4042 = (inp[12]) ? node4054 : node4043;
											assign node4043 = (inp[6]) ? node4049 : node4044;
												assign node4044 = (inp[0]) ? node4046 : 8'b00111110;
													assign node4046 = (inp[2]) ? 8'b00101110 : 8'b00111110;
												assign node4049 = (inp[2]) ? node4051 : 8'b00101111;
													assign node4051 = (inp[0]) ? 8'b00101110 : 8'b00111110;
											assign node4054 = (inp[6]) ? node4060 : node4055;
												assign node4055 = (inp[0]) ? node4057 : 8'b00101111;
													assign node4057 = (inp[5]) ? 8'b00111110 : 8'b00101111;
												assign node4060 = (inp[2]) ? 8'b00111110 : 8'b01111111;
									assign node4063 = (inp[5]) ? node4093 : node4064;
										assign node4064 = (inp[2]) ? node4082 : node4065;
											assign node4065 = (inp[0]) ? node4071 : node4066;
												assign node4066 = (inp[6]) ? node4068 : 8'b00101110;
													assign node4068 = (inp[12]) ? 8'b00111110 : 8'b00101110;
												assign node4071 = (inp[3]) ? node4075 : node4072;
													assign node4072 = (inp[12]) ? 8'b00111011 : 8'b00101011;
													assign node4075 = (inp[6]) ? node4079 : node4076;
														assign node4076 = (inp[12]) ? 8'b00101110 : 8'b00111011;
														assign node4079 = (inp[12]) ? 8'b00111110 : 8'b00101110;
											assign node4082 = (inp[6]) ? node4090 : node4083;
												assign node4083 = (inp[12]) ? node4087 : node4084;
													assign node4084 = (inp[0]) ? 8'b00101010 : 8'b00111011;
													assign node4087 = (inp[0]) ? 8'b00111010 : 8'b00101110;
												assign node4090 = (inp[3]) ? 8'b00111011 : 8'b00101011;
										assign node4093 = (inp[2]) ? node4103 : node4094;
											assign node4094 = (inp[0]) ? node4096 : 8'b00111110;
												assign node4096 = (inp[12]) ? node4100 : node4097;
													assign node4097 = (inp[6]) ? 8'b00101011 : 8'b00111010;
													assign node4100 = (inp[6]) ? 8'b00111011 : 8'b00101011;
											assign node4103 = (inp[0]) ? node4115 : node4104;
												assign node4104 = (inp[6]) ? node4112 : node4105;
													assign node4105 = (inp[12]) ? node4109 : node4106;
														assign node4106 = (inp[3]) ? 8'b00111010 : 8'b00111011;
														assign node4109 = (inp[3]) ? 8'b00101011 : 8'b00101110;
													assign node4112 = (inp[12]) ? 8'b00111010 : 8'b00101010;
												assign node4115 = (inp[12]) ? 8'b00111010 : 8'b00101010;
							assign node4118 = (inp[5]) ? node4196 : node4119;
								assign node4119 = (inp[12]) ? node4155 : node4120;
									assign node4120 = (inp[6]) ? node4144 : node4121;
										assign node4121 = (inp[10]) ? node4135 : node4122;
											assign node4122 = (inp[1]) ? node4128 : node4123;
												assign node4123 = (inp[3]) ? node4125 : 8'b00011111;
													assign node4125 = (inp[0]) ? 8'b00001110 : 8'b00111010;
												assign node4128 = (inp[0]) ? node4130 : 8'b00011111;
													assign node4130 = (inp[3]) ? node4132 : 8'b00011010;
														assign node4132 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node4135 = (inp[2]) ? node4137 : 8'b00011111;
												assign node4137 = (inp[0]) ? node4139 : 8'b00011111;
													assign node4139 = (inp[3]) ? 8'b00001111 : node4140;
														assign node4140 = (inp[1]) ? 8'b00001110 : 8'b00001111;
										assign node4144 = (inp[2]) ? node4150 : node4145;
											assign node4145 = (inp[10]) ? 8'b00101010 : node4146;
												assign node4146 = (inp[3]) ? 8'b00101011 : 8'b00001011;
											assign node4150 = (inp[3]) ? 8'b00111010 : node4151;
												assign node4151 = (inp[10]) ? 8'b00011111 : 8'b00011011;
									assign node4155 = (inp[0]) ? node4171 : node4156;
										assign node4156 = (inp[2]) ? node4166 : node4157;
											assign node4157 = (inp[6]) ? node4161 : node4158;
												assign node4158 = (inp[10]) ? 8'b00101010 : 8'b00101011;
												assign node4161 = (inp[1]) ? 8'b00111010 : node4162;
													assign node4162 = (inp[10]) ? 8'b00111010 : 8'b00111011;
											assign node4166 = (inp[1]) ? 8'b00101010 : node4167;
												assign node4167 = (inp[10]) ? 8'b00101010 : 8'b00101011;
										assign node4171 = (inp[10]) ? node4187 : node4172;
											assign node4172 = (inp[1]) ? node4180 : node4173;
												assign node4173 = (inp[3]) ? node4175 : 8'b00001110;
													assign node4175 = (inp[2]) ? 8'b00011110 : node4176;
														assign node4176 = (inp[6]) ? 8'b00011111 : 8'b00001111;
												assign node4180 = (inp[6]) ? 8'b00001110 : node4181;
													assign node4181 = (inp[2]) ? node4183 : 8'b00001011;
														assign node4183 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node4187 = (inp[2]) ? node4193 : node4188;
												assign node4188 = (inp[6]) ? 8'b00111010 : node4189;
													assign node4189 = (inp[1]) ? 8'b00101010 : 8'b00101011;
												assign node4193 = (inp[3]) ? 8'b00111010 : 8'b00011111;
								assign node4196 = (inp[1]) ? node4242 : node4197;
									assign node4197 = (inp[12]) ? node4217 : node4198;
										assign node4198 = (inp[10]) ? node4204 : node4199;
											assign node4199 = (inp[6]) ? node4201 : 8'b00111010;
												assign node4201 = (inp[3]) ? 8'b00101011 : 8'b00101010;
											assign node4204 = (inp[3]) ? node4212 : node4205;
												assign node4205 = (inp[6]) ? 8'b00001011 : node4206;
													assign node4206 = (inp[0]) ? node4208 : 8'b00011011;
														assign node4208 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node4212 = (inp[6]) ? node4214 : 8'b00011110;
													assign node4214 = (inp[0]) ? 8'b00001111 : 8'b00001110;
										assign node4217 = (inp[10]) ? node4231 : node4218;
											assign node4218 = (inp[0]) ? node4224 : node4219;
												assign node4219 = (inp[3]) ? 8'b00111010 : node4220;
													assign node4220 = (inp[2]) ? 8'b00011111 : 8'b00111010;
												assign node4224 = (inp[3]) ? node4228 : node4225;
													assign node4225 = (inp[6]) ? 8'b00011110 : 8'b00011011;
													assign node4228 = (inp[2]) ? 8'b00011110 : 8'b00011111;
											assign node4231 = (inp[6]) ? node4237 : node4232;
												assign node4232 = (inp[0]) ? 8'b00011110 : node4233;
													assign node4233 = (inp[3]) ? 8'b00001111 : 8'b00001110;
												assign node4237 = (inp[2]) ? 8'b00011110 : node4238;
													assign node4238 = (inp[3]) ? 8'b00011111 : 8'b00011110;
									assign node4242 = (inp[0]) ? node4268 : node4243;
										assign node4243 = (inp[10]) ? node4253 : node4244;
											assign node4244 = (inp[2]) ? node4246 : 8'b00011111;
												assign node4246 = (inp[12]) ? node4250 : node4247;
													assign node4247 = (inp[3]) ? 8'b00011110 : 8'b00011111;
													assign node4250 = (inp[6]) ? 8'b00011111 : 8'b00101010;
											assign node4253 = (inp[3]) ? node4259 : node4254;
												assign node4254 = (inp[6]) ? node4256 : 8'b00001110;
													assign node4256 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node4259 = (inp[12]) ? node4263 : node4260;
													assign node4260 = (inp[6]) ? 8'b00001010 : 8'b00011010;
													assign node4263 = (inp[6]) ? node4265 : 8'b00001011;
														assign node4265 = (inp[2]) ? 8'b00011010 : 8'b00011011;
										assign node4268 = (inp[2]) ? node4274 : node4269;
											assign node4269 = (inp[6]) ? 8'b00001011 : node4270;
												assign node4270 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node4274 = (inp[12]) ? 8'b00011010 : 8'b00001010;
				assign node4277 = (inp[5]) ? node4855 : node4278;
					assign node4278 = (inp[0]) ? node4414 : node4279;
						assign node4279 = (inp[12]) ? node4371 : node4280;
							assign node4280 = (inp[11]) ? node4328 : node4281;
								assign node4281 = (inp[10]) ? node4299 : node4282;
									assign node4282 = (inp[6]) ? node4288 : node4283;
										assign node4283 = (inp[3]) ? node4285 : 8'b10000010;
											assign node4285 = (inp[1]) ? 8'b10000010 : 8'b00001011;
										assign node4288 = (inp[2]) ? node4294 : node4289;
											assign node4289 = (inp[3]) ? node4291 : 8'b00011010;
												assign node4291 = (inp[1]) ? 8'b00011010 : 8'b00011011;
											assign node4294 = (inp[3]) ? node4296 : 8'b10000010;
												assign node4296 = (inp[1]) ? 8'b10000010 : 8'b00001011;
									assign node4299 = (inp[8]) ? node4315 : node4300;
										assign node4300 = (inp[2]) ? node4310 : node4301;
											assign node4301 = (inp[6]) ? node4305 : node4302;
												assign node4302 = (inp[3]) ? 8'b00001111 : 8'b00001110;
												assign node4305 = (inp[3]) ? node4307 : 8'b00011110;
													assign node4307 = (inp[1]) ? 8'b00011110 : 8'b00011111;
											assign node4310 = (inp[1]) ? 8'b00001110 : node4311;
												assign node4311 = (inp[3]) ? 8'b00001111 : 8'b00001110;
										assign node4315 = (inp[2]) ? node4323 : node4316;
											assign node4316 = (inp[6]) ? 8'b00011010 : node4317;
												assign node4317 = (inp[3]) ? node4319 : 8'b10000010;
													assign node4319 = (inp[1]) ? 8'b10000010 : 8'b00001011;
											assign node4323 = (inp[3]) ? node4325 : 8'b10000010;
												assign node4325 = (inp[1]) ? 8'b10000010 : 8'b00001011;
								assign node4328 = (inp[6]) ? node4346 : node4329;
									assign node4329 = (inp[3]) ? node4335 : node4330;
										assign node4330 = (inp[10]) ? node4332 : 8'b11110111;
											assign node4332 = (inp[8]) ? 8'b11110111 : 8'b00011011;
										assign node4335 = (inp[1]) ? node4341 : node4336;
											assign node4336 = (inp[8]) ? 8'b00011010 : node4337;
												assign node4337 = (inp[10]) ? 8'b00011110 : 8'b00011010;
											assign node4341 = (inp[2]) ? 8'b11110111 : node4342;
												assign node4342 = (inp[8]) ? 8'b11110111 : 8'b00011011;
									assign node4346 = (inp[2]) ? node4360 : node4347;
										assign node4347 = (inp[1]) ? node4355 : node4348;
											assign node4348 = (inp[3]) ? 8'b00001011 : node4349;
												assign node4349 = (inp[8]) ? 8'b00001010 : node4350;
													assign node4350 = (inp[10]) ? 8'b00001110 : 8'b00001010;
											assign node4355 = (inp[8]) ? 8'b00001010 : node4356;
												assign node4356 = (inp[10]) ? 8'b00001110 : 8'b00001010;
										assign node4360 = (inp[1]) ? node4366 : node4361;
											assign node4361 = (inp[3]) ? node4363 : 8'b11110111;
												assign node4363 = (inp[8]) ? 8'b00011010 : 8'b00011110;
											assign node4366 = (inp[10]) ? node4368 : 8'b11110111;
												assign node4368 = (inp[8]) ? 8'b11110111 : 8'b00011011;
							assign node4371 = (inp[1]) ? node4397 : node4372;
								assign node4372 = (inp[3]) ? node4386 : node4373;
									assign node4373 = (inp[8]) ? node4381 : node4374;
										assign node4374 = (inp[10]) ? 8'b00001110 : node4375;
											assign node4375 = (inp[2]) ? 8'b00000010 : node4376;
												assign node4376 = (inp[6]) ? 8'b00011010 : 8'b00000010;
										assign node4381 = (inp[2]) ? 8'b00000010 : node4382;
											assign node4382 = (inp[6]) ? 8'b00011010 : 8'b00000010;
									assign node4386 = (inp[2]) ? node4392 : node4387;
										assign node4387 = (inp[6]) ? node4389 : 8'b00001011;
											assign node4389 = (inp[8]) ? 8'b00011011 : 8'b00011111;
										assign node4392 = (inp[10]) ? node4394 : 8'b00001011;
											assign node4394 = (inp[8]) ? 8'b00001011 : 8'b00001111;
								assign node4397 = (inp[2]) ? node4409 : node4398;
									assign node4398 = (inp[6]) ? node4404 : node4399;
										assign node4399 = (inp[10]) ? node4401 : 8'b00000010;
											assign node4401 = (inp[8]) ? 8'b00000010 : 8'b00001110;
										assign node4404 = (inp[8]) ? 8'b00011010 : node4405;
											assign node4405 = (inp[10]) ? 8'b00011110 : 8'b00011010;
									assign node4409 = (inp[8]) ? 8'b00000010 : node4410;
										assign node4410 = (inp[10]) ? 8'b00001110 : 8'b00000010;
						assign node4414 = (inp[9]) ? node4646 : node4415;
							assign node4415 = (inp[11]) ? node4521 : node4416;
								assign node4416 = (inp[8]) ? node4462 : node4417;
									assign node4417 = (inp[10]) ? node4441 : node4418;
										assign node4418 = (inp[1]) ? node4430 : node4419;
											assign node4419 = (inp[3]) ? node4425 : node4420;
												assign node4420 = (inp[2]) ? node4422 : 8'b10100000;
													assign node4422 = (inp[6]) ? 8'b10100000 : 8'b10110000;
												assign node4425 = (inp[6]) ? 8'b10101001 : node4426;
													assign node4426 = (inp[2]) ? 8'b10111001 : 8'b10101001;
											assign node4430 = (inp[3]) ? node4432 : 8'b10100001;
												assign node4432 = (inp[12]) ? node4434 : 8'b10100000;
													assign node4434 = (inp[6]) ? node4438 : node4435;
														assign node4435 = (inp[2]) ? 8'b10110000 : 8'b10100000;
														assign node4438 = (inp[2]) ? 8'b10100000 : 8'b10111000;
										assign node4441 = (inp[2]) ? node4449 : node4442;
											assign node4442 = (inp[6]) ? 8'b10111100 : node4443;
												assign node4443 = (inp[3]) ? 8'b10101100 : node4444;
													assign node4444 = (inp[1]) ? 8'b10101101 : 8'b10101100;
											assign node4449 = (inp[6]) ? node4457 : node4450;
												assign node4450 = (inp[3]) ? node4454 : node4451;
													assign node4451 = (inp[1]) ? 8'b11111101 : 8'b10111100;
													assign node4454 = (inp[12]) ? 8'b10111100 : 8'b11111101;
												assign node4457 = (inp[1]) ? 8'b10101101 : node4458;
													assign node4458 = (inp[3]) ? 8'b10101101 : 8'b10101100;
									assign node4462 = (inp[10]) ? node4496 : node4463;
										assign node4463 = (inp[6]) ? node4477 : node4464;
											assign node4464 = (inp[2]) ? node4472 : node4465;
												assign node4465 = (inp[12]) ? node4467 : 8'b10101101;
													assign node4467 = (inp[3]) ? 8'b10100100 : node4468;
														assign node4468 = (inp[1]) ? 8'b10100101 : 8'b10100100;
												assign node4472 = (inp[1]) ? node4474 : 8'b10110100;
													assign node4474 = (inp[3]) ? 8'b10110100 : 8'b11110101;
											assign node4477 = (inp[2]) ? node4491 : node4478;
												assign node4478 = (inp[12]) ? node4484 : node4479;
													assign node4479 = (inp[1]) ? node4481 : 8'b10111100;
														assign node4481 = (inp[3]) ? 8'b10111100 : 8'b11111101;
													assign node4484 = (inp[1]) ? node4488 : node4485;
														assign node4485 = (inp[3]) ? 8'b11111101 : 8'b10111100;
														assign node4488 = (inp[3]) ? 8'b10111100 : 8'b11111101;
												assign node4491 = (inp[12]) ? node4493 : 8'b10100100;
													assign node4493 = (inp[1]) ? 8'b10100101 : 8'b10101101;
										assign node4496 = (inp[1]) ? node4508 : node4497;
											assign node4497 = (inp[3]) ? 8'b10101001 : node4498;
												assign node4498 = (inp[12]) ? node4500 : 8'b10111000;
													assign node4500 = (inp[6]) ? node4504 : node4501;
														assign node4501 = (inp[2]) ? 8'b10110000 : 8'b10100000;
														assign node4504 = (inp[2]) ? 8'b10100000 : 8'b10111000;
											assign node4508 = (inp[3]) ? node4514 : node4509;
												assign node4509 = (inp[2]) ? node4511 : 8'b10100001;
													assign node4511 = (inp[6]) ? 8'b10100001 : 8'b10110001;
												assign node4514 = (inp[6]) ? node4518 : node4515;
													assign node4515 = (inp[2]) ? 8'b10110000 : 8'b10100000;
													assign node4518 = (inp[2]) ? 8'b10100000 : 8'b10111000;
								assign node4521 = (inp[10]) ? node4581 : node4522;
									assign node4522 = (inp[6]) ? node4554 : node4523;
										assign node4523 = (inp[3]) ? node4537 : node4524;
											assign node4524 = (inp[8]) ? node4532 : node4525;
												assign node4525 = (inp[12]) ? node4529 : node4526;
													assign node4526 = (inp[2]) ? 8'b10000100 : 8'b10010100;
													assign node4529 = (inp[2]) ? 8'b10010100 : 8'b10000101;
												assign node4532 = (inp[2]) ? 8'b10010001 : node4533;
													assign node4533 = (inp[12]) ? 8'b10000100 : 8'b10010000;
											assign node4537 = (inp[1]) ? node4541 : node4538;
												assign node4538 = (inp[8]) ? 8'b10001101 : 8'b10101001;
												assign node4541 = (inp[8]) ? node4549 : node4542;
													assign node4542 = (inp[12]) ? node4546 : node4543;
														assign node4543 = (inp[2]) ? 8'b10000101 : 8'b10010101;
														assign node4546 = (inp[2]) ? 8'b10010101 : 8'b10100000;
													assign node4549 = (inp[12]) ? 8'b10010001 : node4550;
														assign node4550 = (inp[2]) ? 8'b10000001 : 8'b10010001;
										assign node4554 = (inp[8]) ? node4568 : node4555;
											assign node4555 = (inp[1]) ? node4563 : node4556;
												assign node4556 = (inp[3]) ? node4558 : 8'b10111000;
													assign node4558 = (inp[12]) ? node4560 : 8'b10111000;
														assign node4560 = (inp[2]) ? 8'b10101001 : 8'b10111001;
												assign node4563 = (inp[3]) ? node4565 : 8'b10010100;
													assign node4565 = (inp[2]) ? 8'b10100000 : 8'b10111000;
											assign node4568 = (inp[3]) ? node4570 : 8'b10010001;
												assign node4570 = (inp[2]) ? node4576 : node4571;
													assign node4571 = (inp[12]) ? node4573 : 8'b10001100;
														assign node4573 = (inp[1]) ? 8'b10011100 : 8'b10011101;
													assign node4576 = (inp[1]) ? node4578 : 8'b10011100;
														assign node4578 = (inp[12]) ? 8'b10000100 : 8'b10010001;
									assign node4581 = (inp[8]) ? node4615 : node4582;
										assign node4582 = (inp[1]) ? node4602 : node4583;
											assign node4583 = (inp[2]) ? node4595 : node4584;
												assign node4584 = (inp[12]) ? node4592 : node4585;
													assign node4585 = (inp[6]) ? node4589 : node4586;
														assign node4586 = (inp[3]) ? 8'b10111100 : 8'b10111001;
														assign node4589 = (inp[3]) ? 8'b10101101 : 8'b10101100;
													assign node4592 = (inp[3]) ? 8'b11111101 : 8'b10111100;
												assign node4595 = (inp[12]) ? node4599 : node4596;
													assign node4596 = (inp[6]) ? 8'b10111001 : 8'b10101001;
													assign node4599 = (inp[3]) ? 8'b10101101 : 8'b10101100;
											assign node4602 = (inp[2]) ? node4608 : node4603;
												assign node4603 = (inp[3]) ? node4605 : 8'b10101001;
													assign node4605 = (inp[12]) ? 8'b10101100 : 8'b10111001;
												assign node4608 = (inp[3]) ? 8'b10101001 : node4609;
													assign node4609 = (inp[6]) ? 8'b10111000 : node4610;
														assign node4610 = (inp[12]) ? 8'b10111000 : 8'b10101000;
										assign node4615 = (inp[3]) ? node4633 : node4616;
											assign node4616 = (inp[1]) ? node4626 : node4617;
												assign node4617 = (inp[12]) ? node4623 : node4618;
													assign node4618 = (inp[6]) ? 8'b10010101 : node4619;
														assign node4619 = (inp[2]) ? 8'b10000101 : 8'b10010101;
													assign node4623 = (inp[6]) ? 8'b10100000 : 8'b10010101;
												assign node4626 = (inp[2]) ? node4628 : 8'b10000101;
													assign node4628 = (inp[12]) ? 8'b10010100 : node4629;
														assign node4629 = (inp[6]) ? 8'b10010100 : 8'b10000100;
											assign node4633 = (inp[1]) ? node4641 : node4634;
												assign node4634 = (inp[12]) ? node4636 : 8'b10111000;
													assign node4636 = (inp[2]) ? node4638 : 8'b10101001;
														assign node4638 = (inp[6]) ? 8'b10101001 : 8'b10111000;
												assign node4641 = (inp[6]) ? node4643 : 8'b10100000;
													assign node4643 = (inp[12]) ? 8'b10111000 : 8'b10101000;
							assign node4646 = (inp[8]) ? node4764 : node4647;
								assign node4647 = (inp[10]) ? node4687 : node4648;
									assign node4648 = (inp[1]) ? node4666 : node4649;
										assign node4649 = (inp[3]) ? node4657 : node4650;
											assign node4650 = (inp[6]) ? node4654 : node4651;
												assign node4651 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node4654 = (inp[2]) ? 8'b00000010 : 8'b00011010;
											assign node4657 = (inp[11]) ? node4663 : node4658;
												assign node4658 = (inp[6]) ? node4660 : 8'b00001011;
													assign node4660 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node4663 = (inp[6]) ? 8'b00001011 : 8'b00011010;
										assign node4666 = (inp[2]) ? node4676 : node4667;
											assign node4667 = (inp[3]) ? node4673 : node4668;
												assign node4668 = (inp[11]) ? 8'b11111101 : node4669;
													assign node4669 = (inp[12]) ? 8'b10000001 : 8'b10011001;
												assign node4673 = (inp[6]) ? 8'b00011010 : 8'b00000010;
											assign node4676 = (inp[11]) ? node4678 : 8'b10000001;
												assign node4678 = (inp[3]) ? node4684 : node4679;
													assign node4679 = (inp[6]) ? node4681 : 8'b10110100;
														assign node4681 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node4684 = (inp[12]) ? 8'b11110101 : 8'b10100101;
									assign node4687 = (inp[11]) ? node4727 : node4688;
										assign node4688 = (inp[12]) ? node4708 : node4689;
											assign node4689 = (inp[3]) ? node4701 : node4690;
												assign node4690 = (inp[1]) ? node4696 : node4691;
													assign node4691 = (inp[2]) ? 8'b00001110 : node4692;
														assign node4692 = (inp[6]) ? 8'b00011110 : 8'b00001110;
													assign node4696 = (inp[2]) ? 8'b00001111 : node4697;
														assign node4697 = (inp[6]) ? 8'b00011111 : 8'b00001111;
												assign node4701 = (inp[2]) ? node4705 : node4702;
													assign node4702 = (inp[6]) ? 8'b00011111 : 8'b00001111;
													assign node4705 = (inp[6]) ? 8'b00001111 : 8'b00011111;
											assign node4708 = (inp[2]) ? node4720 : node4709;
												assign node4709 = (inp[6]) ? node4715 : node4710;
													assign node4710 = (inp[3]) ? node4712 : 8'b00001111;
														assign node4712 = (inp[1]) ? 8'b00001110 : 8'b00001111;
													assign node4715 = (inp[3]) ? 8'b00011110 : node4716;
														assign node4716 = (inp[1]) ? 8'b00011111 : 8'b00011110;
												assign node4720 = (inp[6]) ? 8'b00001111 : node4721;
													assign node4721 = (inp[1]) ? 8'b00011110 : node4722;
														assign node4722 = (inp[3]) ? 8'b00011111 : 8'b00011110;
										assign node4727 = (inp[3]) ? node4749 : node4728;
											assign node4728 = (inp[2]) ? node4736 : node4729;
												assign node4729 = (inp[6]) ? 8'b00001110 : node4730;
													assign node4730 = (inp[12]) ? node4732 : 8'b00011011;
														assign node4732 = (inp[1]) ? 8'b00001011 : 8'b00001110;
												assign node4736 = (inp[1]) ? node4744 : node4737;
													assign node4737 = (inp[6]) ? node4741 : node4738;
														assign node4738 = (inp[12]) ? 8'b00011011 : 8'b00001011;
														assign node4741 = (inp[12]) ? 8'b00001110 : 8'b00011011;
													assign node4744 = (inp[6]) ? node4746 : 8'b00011010;
														assign node4746 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node4749 = (inp[1]) ? node4755 : node4750;
												assign node4750 = (inp[12]) ? node4752 : 8'b00011110;
													assign node4752 = (inp[6]) ? 8'b00011111 : 8'b00011110;
												assign node4755 = (inp[2]) ? node4761 : node4756;
													assign node4756 = (inp[12]) ? node4758 : 8'b00001110;
														assign node4758 = (inp[6]) ? 8'b00011110 : 8'b00001110;
													assign node4761 = (inp[12]) ? 8'b00011011 : 8'b00001011;
								assign node4764 = (inp[10]) ? node4802 : node4765;
									assign node4765 = (inp[11]) ? node4791 : node4766;
										assign node4766 = (inp[2]) ? node4782 : node4767;
											assign node4767 = (inp[6]) ? node4771 : node4768;
												assign node4768 = (inp[12]) ? 8'b10001101 : 8'b10000100;
												assign node4771 = (inp[12]) ? node4777 : node4772;
													assign node4772 = (inp[1]) ? node4774 : 8'b10011100;
														assign node4774 = (inp[3]) ? 8'b10011100 : 8'b10011101;
													assign node4777 = (inp[1]) ? 8'b10011100 : node4778;
														assign node4778 = (inp[3]) ? 8'b10011101 : 8'b10011100;
											assign node4782 = (inp[6]) ? node4784 : 8'b10010101;
												assign node4784 = (inp[1]) ? node4788 : node4785;
													assign node4785 = (inp[3]) ? 8'b10001101 : 8'b10000100;
													assign node4788 = (inp[3]) ? 8'b10000100 : 8'b10000101;
										assign node4791 = (inp[1]) ? node4797 : node4792;
											assign node4792 = (inp[6]) ? node4794 : 8'b10111100;
												assign node4794 = (inp[3]) ? 8'b10101101 : 8'b10100100;
											assign node4797 = (inp[12]) ? node4799 : 8'b10110001;
												assign node4799 = (inp[3]) ? 8'b10100100 : 8'b10100001;
									assign node4802 = (inp[1]) ? node4832 : node4803;
										assign node4803 = (inp[3]) ? node4821 : node4804;
											assign node4804 = (inp[2]) ? node4812 : node4805;
												assign node4805 = (inp[6]) ? node4809 : node4806;
													assign node4806 = (inp[11]) ? 8'b00000010 : 8'b10000010;
													assign node4809 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node4812 = (inp[11]) ? node4818 : node4813;
													assign node4813 = (inp[6]) ? node4815 : 8'b10010000;
														assign node4815 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node4818 = (inp[12]) ? 8'b11110101 : 8'b11110111;
											assign node4821 = (inp[2]) ? node4829 : node4822;
												assign node4822 = (inp[12]) ? node4826 : node4823;
													assign node4823 = (inp[6]) ? 8'b00001011 : 8'b00011010;
													assign node4826 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node4829 = (inp[11]) ? 8'b00011010 : 8'b00011011;
										assign node4832 = (inp[11]) ? node4844 : node4833;
											assign node4833 = (inp[3]) ? node4839 : node4834;
												assign node4834 = (inp[2]) ? node4836 : 8'b10000001;
													assign node4836 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node4839 = (inp[12]) ? node4841 : 8'b10010000;
													assign node4841 = (inp[2]) ? 8'b00000010 : 8'b00011010;
											assign node4844 = (inp[3]) ? node4852 : node4845;
												assign node4845 = (inp[6]) ? node4847 : 8'b10110100;
													assign node4847 = (inp[2]) ? 8'b10100101 : node4848;
														assign node4848 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node4852 = (inp[12]) ? 8'b00000010 : 8'b11110111;
					assign node4855 = (inp[11]) ? node5017 : node4856;
						assign node4856 = (inp[10]) ? node4936 : node4857;
							assign node4857 = (inp[3]) ? node4893 : node4858;
								assign node4858 = (inp[0]) ? node4872 : node4859;
									assign node4859 = (inp[9]) ? node4867 : node4860;
										assign node4860 = (inp[6]) ? node4864 : node4861;
											assign node4861 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node4864 = (inp[2]) ? 8'b10010000 : 8'b00011010;
										assign node4867 = (inp[6]) ? node4869 : 8'b10100000;
											assign node4869 = (inp[2]) ? 8'b10110000 : 8'b10111000;
									assign node4872 = (inp[8]) ? node4884 : node4873;
										assign node4873 = (inp[1]) ? node4879 : node4874;
											assign node4874 = (inp[2]) ? 8'b10110000 : node4875;
												assign node4875 = (inp[6]) ? 8'b10111000 : 8'b10100000;
											assign node4879 = (inp[2]) ? 8'b10110001 : node4880;
												assign node4880 = (inp[6]) ? 8'b10111001 : 8'b10100001;
										assign node4884 = (inp[1]) ? node4890 : node4885;
											assign node4885 = (inp[2]) ? 8'b10110100 : node4886;
												assign node4886 = (inp[6]) ? 8'b10111100 : 8'b10100100;
											assign node4890 = (inp[2]) ? 8'b11110101 : 8'b11111101;
								assign node4893 = (inp[0]) ? node4913 : node4894;
									assign node4894 = (inp[9]) ? node4904 : node4895;
										assign node4895 = (inp[1]) ? node4899 : node4896;
											assign node4896 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node4899 = (inp[6]) ? node4901 : 8'b10000001;
												assign node4901 = (inp[2]) ? 8'b10010001 : 8'b10011001;
										assign node4904 = (inp[6]) ? node4908 : node4905;
											assign node4905 = (inp[1]) ? 8'b10100001 : 8'b10101001;
											assign node4908 = (inp[2]) ? node4910 : 8'b10111001;
												assign node4910 = (inp[1]) ? 8'b10110001 : 8'b10111001;
									assign node4913 = (inp[8]) ? node4927 : node4914;
										assign node4914 = (inp[1]) ? node4920 : node4915;
											assign node4915 = (inp[12]) ? 8'b10111001 : node4916;
												assign node4916 = (inp[6]) ? 8'b10111001 : 8'b10101001;
											assign node4920 = (inp[6]) ? node4924 : node4921;
												assign node4921 = (inp[2]) ? 8'b10110001 : 8'b10100001;
												assign node4924 = (inp[2]) ? 8'b10110001 : 8'b10111001;
										assign node4927 = (inp[6]) ? 8'b11111101 : node4928;
											assign node4928 = (inp[2]) ? node4932 : node4929;
												assign node4929 = (inp[1]) ? 8'b10100101 : 8'b10101101;
												assign node4932 = (inp[1]) ? 8'b11110101 : 8'b11111101;
							assign node4936 = (inp[3]) ? node4978 : node4937;
								assign node4937 = (inp[0]) ? node4957 : node4938;
									assign node4938 = (inp[9]) ? node4948 : node4939;
										assign node4939 = (inp[8]) ? node4943 : node4940;
											assign node4940 = (inp[6]) ? 8'b00011110 : 8'b00001110;
											assign node4943 = (inp[6]) ? node4945 : 8'b10000100;
												assign node4945 = (inp[2]) ? 8'b10010100 : 8'b10011100;
										assign node4948 = (inp[6]) ? node4952 : node4949;
											assign node4949 = (inp[8]) ? 8'b10100100 : 8'b10101100;
											assign node4952 = (inp[2]) ? node4954 : 8'b10111100;
												assign node4954 = (inp[1]) ? 8'b10110100 : 8'b10111100;
									assign node4957 = (inp[1]) ? node4969 : node4958;
										assign node4958 = (inp[8]) ? node4964 : node4959;
											assign node4959 = (inp[2]) ? 8'b10111100 : node4960;
												assign node4960 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node4964 = (inp[2]) ? 8'b10110100 : node4965;
												assign node4965 = (inp[6]) ? 8'b10111100 : 8'b10100100;
										assign node4969 = (inp[2]) ? node4975 : node4970;
											assign node4970 = (inp[9]) ? 8'b11111101 : node4971;
												assign node4971 = (inp[8]) ? 8'b10100101 : 8'b10101101;
											assign node4975 = (inp[8]) ? 8'b11110101 : 8'b11111101;
								assign node4978 = (inp[6]) ? node4998 : node4979;
									assign node4979 = (inp[0]) ? node4991 : node4980;
										assign node4980 = (inp[9]) ? node4986 : node4981;
											assign node4981 = (inp[8]) ? node4983 : 8'b00001111;
												assign node4983 = (inp[1]) ? 8'b10000101 : 8'b10001101;
											assign node4986 = (inp[8]) ? node4988 : 8'b10101101;
												assign node4988 = (inp[1]) ? 8'b10100101 : 8'b10101101;
										assign node4991 = (inp[2]) ? node4993 : 8'b10101101;
											assign node4993 = (inp[1]) ? node4995 : 8'b11111101;
												assign node4995 = (inp[12]) ? 8'b11111101 : 8'b11110101;
									assign node4998 = (inp[9]) ? node5010 : node4999;
										assign node4999 = (inp[0]) ? node5005 : node5000;
											assign node5000 = (inp[8]) ? node5002 : 8'b00011111;
												assign node5002 = (inp[1]) ? 8'b10010101 : 8'b10011101;
											assign node5005 = (inp[1]) ? node5007 : 8'b11111101;
												assign node5007 = (inp[2]) ? 8'b11110101 : 8'b11111101;
										assign node5010 = (inp[1]) ? node5012 : 8'b11111101;
											assign node5012 = (inp[8]) ? node5014 : 8'b11111101;
												assign node5014 = (inp[2]) ? 8'b11110101 : 8'b11111101;
						assign node5017 = (inp[8]) ? node5203 : node5018;
							assign node5018 = (inp[10]) ? node5110 : node5019;
								assign node5019 = (inp[1]) ? node5067 : node5020;
									assign node5020 = (inp[3]) ? node5044 : node5021;
										assign node5021 = (inp[2]) ? node5033 : node5022;
											assign node5022 = (inp[6]) ? node5028 : node5023;
												assign node5023 = (inp[12]) ? 8'b10100000 : node5024;
													assign node5024 = (inp[9]) ? 8'b10010101 : 8'b11110111;
												assign node5028 = (inp[0]) ? node5030 : 8'b00001010;
													assign node5030 = (inp[12]) ? 8'b10111000 : 8'b10101000;
											assign node5033 = (inp[6]) ? node5039 : node5034;
												assign node5034 = (inp[12]) ? node5036 : 8'b10000101;
													assign node5036 = (inp[9]) ? 8'b10100000 : 8'b00000010;
												assign node5039 = (inp[12]) ? node5041 : 8'b10000101;
													assign node5041 = (inp[0]) ? 8'b10010101 : 8'b11110101;
										assign node5044 = (inp[0]) ? node5058 : node5045;
											assign node5045 = (inp[9]) ? node5049 : node5046;
												assign node5046 = (inp[12]) ? 8'b00001011 : 8'b00001010;
												assign node5049 = (inp[2]) ? 8'b10111000 : node5050;
													assign node5050 = (inp[6]) ? node5054 : node5051;
														assign node5051 = (inp[12]) ? 8'b10101001 : 8'b10111000;
														assign node5054 = (inp[12]) ? 8'b10111001 : 8'b10101001;
											assign node5058 = (inp[2]) ? node5064 : node5059;
												assign node5059 = (inp[12]) ? 8'b10101001 : node5060;
													assign node5060 = (inp[6]) ? 8'b10101001 : 8'b10111000;
												assign node5064 = (inp[12]) ? 8'b10111000 : 8'b10101000;
									assign node5067 = (inp[0]) ? node5099 : node5068;
										assign node5068 = (inp[9]) ? node5090 : node5069;
											assign node5069 = (inp[3]) ? node5083 : node5070;
												assign node5070 = (inp[2]) ? node5076 : node5071;
													assign node5071 = (inp[6]) ? 8'b00001010 : node5072;
														assign node5072 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node5076 = (inp[6]) ? node5080 : node5077;
														assign node5077 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node5080 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node5083 = (inp[6]) ? node5087 : node5084;
													assign node5084 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node5087 = (inp[2]) ? 8'b10110100 : 8'b11111101;
											assign node5090 = (inp[2]) ? node5092 : 8'b10001101;
												assign node5092 = (inp[3]) ? 8'b10010100 : node5093;
													assign node5093 = (inp[6]) ? node5095 : 8'b10100000;
														assign node5095 = (inp[12]) ? 8'b10010101 : 8'b10000101;
										assign node5099 = (inp[2]) ? node5107 : node5100;
											assign node5100 = (inp[6]) ? node5104 : node5101;
												assign node5101 = (inp[12]) ? 8'b10000101 : 8'b10010100;
												assign node5104 = (inp[12]) ? 8'b10011101 : 8'b10001101;
											assign node5107 = (inp[12]) ? 8'b10010100 : 8'b10000100;
								assign node5110 = (inp[0]) ? node5172 : node5111;
									assign node5111 = (inp[9]) ? node5137 : node5112;
										assign node5112 = (inp[2]) ? node5128 : node5113;
											assign node5113 = (inp[3]) ? node5121 : node5114;
												assign node5114 = (inp[6]) ? node5118 : node5115;
													assign node5115 = (inp[12]) ? 8'b00001110 : 8'b00011011;
													assign node5118 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node5121 = (inp[1]) ? node5123 : 8'b00001111;
													assign node5123 = (inp[12]) ? 8'b00001011 : node5124;
														assign node5124 = (inp[6]) ? 8'b00001011 : 8'b00011010;
											assign node5128 = (inp[12]) ? node5130 : 8'b00011011;
												assign node5130 = (inp[6]) ? node5134 : node5131;
													assign node5131 = (inp[3]) ? 8'b00001011 : 8'b00001110;
													assign node5134 = (inp[3]) ? 8'b00011110 : 8'b00011011;
										assign node5137 = (inp[1]) ? node5153 : node5138;
											assign node5138 = (inp[3]) ? node5146 : node5139;
												assign node5139 = (inp[6]) ? node5141 : 8'b10111001;
													assign node5141 = (inp[2]) ? 8'b10101001 : node5142;
														assign node5142 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node5146 = (inp[2]) ? 8'b10101100 : node5147;
													assign node5147 = (inp[6]) ? 8'b10101101 : node5148;
														assign node5148 = (inp[12]) ? 8'b10101101 : 8'b10111100;
											assign node5153 = (inp[3]) ? node5165 : node5154;
												assign node5154 = (inp[2]) ? node5160 : node5155;
													assign node5155 = (inp[6]) ? node5157 : 8'b10111001;
														assign node5157 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node5160 = (inp[6]) ? 8'b10111001 : node5161;
														assign node5161 = (inp[12]) ? 8'b10101100 : 8'b10111001;
												assign node5165 = (inp[2]) ? 8'b10111000 : node5166;
													assign node5166 = (inp[6]) ? 8'b10101001 : node5167;
														assign node5167 = (inp[12]) ? 8'b10101001 : 8'b10111000;
									assign node5172 = (inp[1]) ? node5192 : node5173;
										assign node5173 = (inp[3]) ? node5185 : node5174;
											assign node5174 = (inp[2]) ? node5182 : node5175;
												assign node5175 = (inp[9]) ? 8'b10111001 : node5176;
													assign node5176 = (inp[6]) ? 8'b10101100 : node5177;
														assign node5177 = (inp[12]) ? 8'b10101100 : 8'b10111001;
												assign node5182 = (inp[12]) ? 8'b10111001 : 8'b10101001;
											assign node5185 = (inp[12]) ? node5189 : node5186;
												assign node5186 = (inp[6]) ? 8'b10101101 : 8'b10101100;
												assign node5189 = (inp[2]) ? 8'b10111100 : 8'b11111101;
										assign node5192 = (inp[2]) ? node5200 : node5193;
											assign node5193 = (inp[6]) ? node5197 : node5194;
												assign node5194 = (inp[12]) ? 8'b10101001 : 8'b10111000;
												assign node5197 = (inp[12]) ? 8'b10111001 : 8'b10101001;
											assign node5200 = (inp[12]) ? 8'b10111000 : 8'b10101000;
							assign node5203 = (inp[2]) ? node5297 : node5204;
								assign node5204 = (inp[6]) ? node5242 : node5205;
									assign node5205 = (inp[12]) ? node5219 : node5206;
										assign node5206 = (inp[3]) ? node5212 : node5207;
											assign node5207 = (inp[0]) ? 8'b10010001 : node5208;
												assign node5208 = (inp[10]) ? 8'b10010001 : 8'b10010101;
											assign node5212 = (inp[1]) ? node5216 : node5213;
												assign node5213 = (inp[0]) ? 8'b10011100 : 8'b10111000;
												assign node5216 = (inp[0]) ? 8'b10010000 : 8'b10110000;
										assign node5219 = (inp[1]) ? node5231 : node5220;
											assign node5220 = (inp[3]) ? node5226 : node5221;
												assign node5221 = (inp[10]) ? node5223 : 8'b10000100;
													assign node5223 = (inp[9]) ? 8'b10000100 : 8'b10100100;
												assign node5226 = (inp[0]) ? 8'b10001101 : node5227;
													assign node5227 = (inp[9]) ? 8'b10001101 : 8'b10101101;
											assign node5231 = (inp[0]) ? 8'b10000001 : node5232;
												assign node5232 = (inp[3]) ? node5238 : node5233;
													assign node5233 = (inp[10]) ? 8'b10100100 : node5234;
														assign node5234 = (inp[9]) ? 8'b10100000 : 8'b00000010;
													assign node5238 = (inp[9]) ? 8'b10000101 : 8'b10100101;
									assign node5242 = (inp[12]) ? node5268 : node5243;
										assign node5243 = (inp[3]) ? node5255 : node5244;
											assign node5244 = (inp[0]) ? node5252 : node5245;
												assign node5245 = (inp[10]) ? node5249 : node5246;
													assign node5246 = (inp[9]) ? 8'b10101000 : 8'b00001010;
													assign node5249 = (inp[9]) ? 8'b10001100 : 8'b10101100;
												assign node5252 = (inp[1]) ? 8'b10001001 : 8'b10001100;
											assign node5255 = (inp[0]) ? node5265 : node5256;
												assign node5256 = (inp[10]) ? node5262 : node5257;
													assign node5257 = (inp[1]) ? node5259 : 8'b10101001;
														assign node5259 = (inp[9]) ? 8'b10001101 : 8'b10101101;
													assign node5262 = (inp[9]) ? 8'b10001001 : 8'b10101001;
												assign node5265 = (inp[1]) ? 8'b10001001 : 8'b10001101;
										assign node5268 = (inp[3]) ? node5280 : node5269;
											assign node5269 = (inp[0]) ? node5277 : node5270;
												assign node5270 = (inp[10]) ? node5274 : node5271;
													assign node5271 = (inp[9]) ? 8'b10111000 : 8'b00011010;
													assign node5274 = (inp[9]) ? 8'b10011100 : 8'b10111100;
												assign node5277 = (inp[1]) ? 8'b10011001 : 8'b10011100;
											assign node5280 = (inp[1]) ? node5290 : node5281;
												assign node5281 = (inp[10]) ? node5285 : node5282;
													assign node5282 = (inp[9]) ? 8'b10011101 : 8'b00011011;
													assign node5285 = (inp[9]) ? 8'b10011101 : node5286;
														assign node5286 = (inp[0]) ? 8'b10011101 : 8'b11111101;
												assign node5290 = (inp[9]) ? node5294 : node5291;
													assign node5291 = (inp[0]) ? 8'b10011001 : 8'b10111001;
													assign node5294 = (inp[0]) ? 8'b10011001 : 8'b10011101;
								assign node5297 = (inp[3]) ? node5335 : node5298;
									assign node5298 = (inp[0]) ? node5328 : node5299;
										assign node5299 = (inp[9]) ? node5313 : node5300;
											assign node5300 = (inp[12]) ? node5308 : node5301;
												assign node5301 = (inp[6]) ? node5305 : node5302;
													assign node5302 = (inp[10]) ? 8'b10110001 : 8'b11110111;
													assign node5305 = (inp[10]) ? 8'b10100001 : 8'b10100101;
												assign node5308 = (inp[6]) ? 8'b11110101 : node5309;
													assign node5309 = (inp[10]) ? 8'b10100100 : 8'b00000010;
											assign node5313 = (inp[12]) ? node5321 : node5314;
												assign node5314 = (inp[10]) ? node5318 : node5315;
													assign node5315 = (inp[6]) ? 8'b10000101 : 8'b10010101;
													assign node5318 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node5321 = (inp[6]) ? node5325 : node5322;
													assign node5322 = (inp[10]) ? 8'b10000100 : 8'b10100000;
													assign node5325 = (inp[10]) ? 8'b10010001 : 8'b10010101;
										assign node5328 = (inp[12]) ? node5332 : node5329;
											assign node5329 = (inp[1]) ? 8'b10000000 : 8'b10000001;
											assign node5332 = (inp[1]) ? 8'b10010000 : 8'b10010001;
									assign node5335 = (inp[1]) ? node5345 : node5336;
										assign node5336 = (inp[0]) ? node5342 : node5337;
											assign node5337 = (inp[10]) ? node5339 : 8'b00011010;
												assign node5339 = (inp[9]) ? 8'b10011100 : 8'b10101100;
											assign node5342 = (inp[12]) ? 8'b10011100 : 8'b10001100;
										assign node5345 = (inp[12]) ? node5357 : node5346;
											assign node5346 = (inp[0]) ? 8'b10000000 : node5347;
												assign node5347 = (inp[9]) ? node5353 : node5348;
													assign node5348 = (inp[10]) ? node5350 : 8'b10110100;
														assign node5350 = (inp[6]) ? 8'b10100000 : 8'b10110000;
													assign node5353 = (inp[6]) ? 8'b10000000 : 8'b10010000;
											assign node5357 = (inp[0]) ? 8'b10010000 : node5358;
												assign node5358 = (inp[10]) ? 8'b10010000 : 8'b10010100;
			assign node5362 = (inp[12]) ? node5838 : node5363;
				assign node5363 = (inp[11]) ? node5589 : node5364;
					assign node5364 = (inp[5]) ? node5446 : node5365;
						assign node5365 = (inp[0]) ? node5367 : 8'b10000010;
							assign node5367 = (inp[9]) ? node5407 : node5368;
								assign node5368 = (inp[13]) ? node5382 : node5369;
									assign node5369 = (inp[6]) ? node5377 : node5370;
										assign node5370 = (inp[2]) ? 8'b10010000 : node5371;
											assign node5371 = (inp[8]) ? 8'b10000100 : node5372;
												assign node5372 = (inp[3]) ? 8'b10000010 : 8'b10000001;
										assign node5377 = (inp[1]) ? node5379 : 8'b10000010;
											assign node5379 = (inp[3]) ? 8'b10000010 : 8'b10000001;
									assign node5382 = (inp[2]) ? node5394 : node5383;
										assign node5383 = (inp[3]) ? node5389 : node5384;
											assign node5384 = (inp[1]) ? node5386 : 8'b10100000;
												assign node5386 = (inp[8]) ? 8'b10100101 : 8'b10100001;
											assign node5389 = (inp[8]) ? node5391 : 8'b10100000;
												assign node5391 = (inp[10]) ? 8'b10100000 : 8'b10100100;
										assign node5394 = (inp[6]) ? node5400 : node5395;
											assign node5395 = (inp[8]) ? node5397 : 8'b10110000;
												assign node5397 = (inp[10]) ? 8'b10110000 : 8'b10110100;
											assign node5400 = (inp[8]) ? 8'b10100100 : node5401;
												assign node5401 = (inp[1]) ? node5403 : 8'b10100000;
													assign node5403 = (inp[3]) ? 8'b10100000 : 8'b10100001;
								assign node5407 = (inp[10]) ? node5433 : node5408;
									assign node5408 = (inp[8]) ? node5422 : node5409;
										assign node5409 = (inp[13]) ? node5417 : node5410;
											assign node5410 = (inp[2]) ? node5414 : node5411;
												assign node5411 = (inp[1]) ? 8'b10000001 : 8'b10000010;
												assign node5414 = (inp[6]) ? 8'b10000001 : 8'b10010000;
											assign node5417 = (inp[1]) ? node5419 : 8'b10000010;
												assign node5419 = (inp[3]) ? 8'b10000010 : 8'b10000001;
										assign node5422 = (inp[1]) ? node5424 : 8'b10000100;
											assign node5424 = (inp[3]) ? node5430 : node5425;
												assign node5425 = (inp[13]) ? node5427 : 8'b10000101;
													assign node5427 = (inp[6]) ? 8'b10000101 : 8'b10010101;
												assign node5430 = (inp[13]) ? 8'b10000100 : 8'b10010100;
									assign node5433 = (inp[6]) ? node5441 : node5434;
										assign node5434 = (inp[2]) ? 8'b10010000 : node5435;
											assign node5435 = (inp[3]) ? 8'b10000010 : node5436;
												assign node5436 = (inp[1]) ? 8'b10000001 : 8'b10000010;
										assign node5441 = (inp[3]) ? 8'b10000010 : node5442;
											assign node5442 = (inp[1]) ? 8'b10000001 : 8'b10000010;
						assign node5446 = (inp[13]) ? node5502 : node5447;
							assign node5447 = (inp[2]) ? node5469 : node5448;
								assign node5448 = (inp[1]) ? node5456 : node5449;
									assign node5449 = (inp[8]) ? node5451 : 8'b10000010;
										assign node5451 = (inp[10]) ? 8'b10000100 : node5452;
											assign node5452 = (inp[0]) ? 8'b10000100 : 8'b10000010;
									assign node5456 = (inp[8]) ? node5462 : node5457;
										assign node5457 = (inp[3]) ? 8'b10000001 : node5458;
											assign node5458 = (inp[0]) ? 8'b10000001 : 8'b10000010;
										assign node5462 = (inp[10]) ? 8'b10000101 : node5463;
											assign node5463 = (inp[0]) ? 8'b10000101 : node5464;
												assign node5464 = (inp[3]) ? 8'b10000001 : 8'b10000010;
								assign node5469 = (inp[1]) ? node5485 : node5470;
									assign node5470 = (inp[8]) ? node5476 : node5471;
										assign node5471 = (inp[0]) ? 8'b10010000 : node5472;
											assign node5472 = (inp[6]) ? 8'b10010000 : 8'b10000010;
										assign node5476 = (inp[0]) ? 8'b10010100 : node5477;
											assign node5477 = (inp[6]) ? node5481 : node5478;
												assign node5478 = (inp[10]) ? 8'b10000100 : 8'b10000010;
												assign node5481 = (inp[10]) ? 8'b10010100 : 8'b10010000;
									assign node5485 = (inp[8]) ? node5495 : node5486;
										assign node5486 = (inp[0]) ? 8'b10010001 : node5487;
											assign node5487 = (inp[3]) ? node5491 : node5488;
												assign node5488 = (inp[6]) ? 8'b10010000 : 8'b10000010;
												assign node5491 = (inp[10]) ? 8'b10000001 : 8'b10010001;
										assign node5495 = (inp[0]) ? 8'b10010101 : node5496;
											assign node5496 = (inp[6]) ? node5498 : 8'b10000101;
												assign node5498 = (inp[3]) ? 8'b10010001 : 8'b10010000;
							assign node5502 = (inp[8]) ? node5538 : node5503;
								assign node5503 = (inp[1]) ? node5517 : node5504;
									assign node5504 = (inp[2]) ? node5510 : node5505;
										assign node5505 = (inp[0]) ? 8'b10100000 : node5506;
											assign node5506 = (inp[9]) ? 8'b10100000 : 8'b10000010;
										assign node5510 = (inp[0]) ? 8'b10110000 : node5511;
											assign node5511 = (inp[6]) ? node5513 : 8'b10100000;
												assign node5513 = (inp[9]) ? 8'b10110000 : 8'b10010000;
									assign node5517 = (inp[0]) ? node5535 : node5518;
										assign node5518 = (inp[3]) ? node5526 : node5519;
											assign node5519 = (inp[9]) ? node5523 : node5520;
												assign node5520 = (inp[10]) ? 8'b10000010 : 8'b10010000;
												assign node5523 = (inp[10]) ? 8'b10110000 : 8'b10100000;
											assign node5526 = (inp[9]) ? node5532 : node5527;
												assign node5527 = (inp[6]) ? node5529 : 8'b10000001;
													assign node5529 = (inp[2]) ? 8'b10010001 : 8'b10000001;
												assign node5532 = (inp[6]) ? 8'b10110001 : 8'b10100001;
										assign node5535 = (inp[2]) ? 8'b10110001 : 8'b10100001;
								assign node5538 = (inp[1]) ? node5562 : node5539;
									assign node5539 = (inp[2]) ? node5549 : node5540;
										assign node5540 = (inp[9]) ? node5544 : node5541;
											assign node5541 = (inp[0]) ? 8'b10100100 : 8'b10000100;
											assign node5544 = (inp[0]) ? 8'b10100100 : node5545;
												assign node5545 = (inp[10]) ? 8'b10100100 : 8'b10100000;
										assign node5549 = (inp[0]) ? 8'b10110100 : node5550;
											assign node5550 = (inp[9]) ? node5554 : node5551;
												assign node5551 = (inp[6]) ? 8'b10010100 : 8'b10000100;
												assign node5554 = (inp[10]) ? node5558 : node5555;
													assign node5555 = (inp[6]) ? 8'b10110000 : 8'b10100000;
													assign node5558 = (inp[6]) ? 8'b10110100 : 8'b10100100;
									assign node5562 = (inp[2]) ? node5574 : node5563;
										assign node5563 = (inp[0]) ? 8'b10100101 : node5564;
											assign node5564 = (inp[3]) ? node5568 : node5565;
												assign node5565 = (inp[6]) ? 8'b10100100 : 8'b10000010;
												assign node5568 = (inp[10]) ? 8'b10000101 : node5569;
													assign node5569 = (inp[9]) ? 8'b10100001 : 8'b10000001;
										assign node5574 = (inp[0]) ? 8'b11110101 : node5575;
											assign node5575 = (inp[6]) ? node5581 : node5576;
												assign node5576 = (inp[10]) ? node5578 : 8'b10100000;
													assign node5578 = (inp[3]) ? 8'b10100101 : 8'b10100100;
												assign node5581 = (inp[9]) ? node5585 : node5582;
													assign node5582 = (inp[10]) ? 8'b10010101 : 8'b10010000;
													assign node5585 = (inp[10]) ? 8'b11110101 : 8'b10110001;
					assign node5589 = (inp[0]) ? node5693 : node5590;
						assign node5590 = (inp[5]) ? node5592 : 8'b11110111;
							assign node5592 = (inp[10]) ? node5634 : node5593;
								assign node5593 = (inp[3]) ? node5611 : node5594;
									assign node5594 = (inp[6]) ? node5600 : node5595;
										assign node5595 = (inp[13]) ? node5597 : 8'b11110111;
											assign node5597 = (inp[9]) ? 8'b10010101 : 8'b11110111;
										assign node5600 = (inp[2]) ? node5606 : node5601;
											assign node5601 = (inp[9]) ? node5603 : 8'b11110111;
												assign node5603 = (inp[13]) ? 8'b10010101 : 8'b11110111;
											assign node5606 = (inp[13]) ? node5608 : 8'b10100101;
												assign node5608 = (inp[9]) ? 8'b10000101 : 8'b10100101;
									assign node5611 = (inp[1]) ? node5625 : node5612;
										assign node5612 = (inp[13]) ? node5614 : 8'b11110111;
											assign node5614 = (inp[9]) ? node5620 : node5615;
												assign node5615 = (inp[2]) ? node5617 : 8'b11110111;
													assign node5617 = (inp[6]) ? 8'b10100101 : 8'b11110111;
												assign node5620 = (inp[2]) ? node5622 : 8'b10010101;
													assign node5622 = (inp[6]) ? 8'b10000101 : 8'b10010101;
										assign node5625 = (inp[2]) ? node5631 : node5626;
											assign node5626 = (inp[13]) ? node5628 : 8'b10110100;
												assign node5628 = (inp[9]) ? 8'b10010100 : 8'b10110100;
											assign node5631 = (inp[6]) ? 8'b10100100 : 8'b10110100;
								assign node5634 = (inp[8]) ? node5666 : node5635;
									assign node5635 = (inp[9]) ? node5653 : node5636;
										assign node5636 = (inp[2]) ? node5642 : node5637;
											assign node5637 = (inp[1]) ? node5639 : 8'b11110111;
												assign node5639 = (inp[3]) ? 8'b10110100 : 8'b11110111;
											assign node5642 = (inp[6]) ? node5648 : node5643;
												assign node5643 = (inp[1]) ? node5645 : 8'b11110111;
													assign node5645 = (inp[3]) ? 8'b10110100 : 8'b11110111;
												assign node5648 = (inp[3]) ? node5650 : 8'b10100101;
													assign node5650 = (inp[13]) ? 8'b10100101 : 8'b10100100;
										assign node5653 = (inp[13]) ? node5657 : node5654;
											assign node5654 = (inp[6]) ? 8'b10100101 : 8'b11110111;
											assign node5657 = (inp[3]) ? node5663 : node5658;
												assign node5658 = (inp[6]) ? node5660 : 8'b10010101;
													assign node5660 = (inp[2]) ? 8'b10000101 : 8'b10010101;
												assign node5663 = (inp[6]) ? 8'b10010101 : 8'b10010100;
									assign node5666 = (inp[3]) ? node5676 : node5667;
										assign node5667 = (inp[13]) ? node5673 : node5668;
											assign node5668 = (inp[6]) ? node5670 : 8'b10110001;
												assign node5670 = (inp[2]) ? 8'b10100001 : 8'b10110001;
											assign node5673 = (inp[9]) ? 8'b10010001 : 8'b10110001;
										assign node5676 = (inp[1]) ? node5684 : node5677;
											assign node5677 = (inp[13]) ? 8'b10010001 : node5678;
												assign node5678 = (inp[6]) ? node5680 : 8'b10110001;
													assign node5680 = (inp[2]) ? 8'b10100001 : 8'b10110001;
											assign node5684 = (inp[2]) ? node5690 : node5685;
												assign node5685 = (inp[9]) ? node5687 : 8'b10110000;
													assign node5687 = (inp[13]) ? 8'b10010000 : 8'b10110000;
												assign node5690 = (inp[6]) ? 8'b10100000 : 8'b10110000;
						assign node5693 = (inp[2]) ? node5757 : node5694;
							assign node5694 = (inp[8]) ? node5720 : node5695;
								assign node5695 = (inp[1]) ? node5703 : node5696;
									assign node5696 = (inp[13]) ? node5698 : 8'b11110111;
										assign node5698 = (inp[9]) ? node5700 : 8'b10010101;
											assign node5700 = (inp[5]) ? 8'b10010101 : 8'b11110111;
									assign node5703 = (inp[3]) ? node5711 : node5704;
										assign node5704 = (inp[13]) ? node5706 : 8'b10110100;
											assign node5706 = (inp[5]) ? 8'b10010100 : node5707;
												assign node5707 = (inp[9]) ? 8'b10110100 : 8'b10010100;
										assign node5711 = (inp[5]) ? node5717 : node5712;
											assign node5712 = (inp[13]) ? node5714 : 8'b11110111;
												assign node5714 = (inp[9]) ? 8'b11110111 : 8'b10010101;
											assign node5717 = (inp[13]) ? 8'b10010100 : 8'b10110100;
								assign node5720 = (inp[1]) ? node5736 : node5721;
									assign node5721 = (inp[5]) ? node5733 : node5722;
										assign node5722 = (inp[10]) ? node5728 : node5723;
											assign node5723 = (inp[9]) ? 8'b10110001 : node5724;
												assign node5724 = (inp[13]) ? 8'b10010001 : 8'b10110001;
											assign node5728 = (inp[9]) ? 8'b11110111 : node5729;
												assign node5729 = (inp[13]) ? 8'b10010101 : 8'b11110111;
										assign node5733 = (inp[13]) ? 8'b10010001 : 8'b10110001;
									assign node5736 = (inp[5]) ? node5754 : node5737;
										assign node5737 = (inp[10]) ? node5745 : node5738;
											assign node5738 = (inp[3]) ? node5742 : node5739;
												assign node5739 = (inp[9]) ? 8'b10110000 : 8'b10010000;
												assign node5742 = (inp[9]) ? 8'b10110001 : 8'b10010001;
											assign node5745 = (inp[3]) ? node5751 : node5746;
												assign node5746 = (inp[6]) ? 8'b10110100 : node5747;
													assign node5747 = (inp[9]) ? 8'b10110100 : 8'b10010100;
												assign node5751 = (inp[9]) ? 8'b11110111 : 8'b10010101;
										assign node5754 = (inp[13]) ? 8'b10010000 : 8'b10110000;
							assign node5757 = (inp[1]) ? node5793 : node5758;
								assign node5758 = (inp[13]) ? node5776 : node5759;
									assign node5759 = (inp[8]) ? node5767 : node5760;
										assign node5760 = (inp[10]) ? 8'b10100101 : node5761;
											assign node5761 = (inp[5]) ? 8'b10100101 : node5762;
												assign node5762 = (inp[3]) ? 8'b10100101 : 8'b11110111;
										assign node5767 = (inp[5]) ? 8'b10100001 : node5768;
											assign node5768 = (inp[6]) ? node5772 : node5769;
												assign node5769 = (inp[10]) ? 8'b10100101 : 8'b10100001;
												assign node5772 = (inp[10]) ? 8'b11110111 : 8'b10110001;
									assign node5776 = (inp[5]) ? node5790 : node5777;
										assign node5777 = (inp[9]) ? node5785 : node5778;
											assign node5778 = (inp[6]) ? node5780 : 8'b10000101;
												assign node5780 = (inp[8]) ? node5782 : 8'b10010101;
													assign node5782 = (inp[10]) ? 8'b10010101 : 8'b10010001;
											assign node5785 = (inp[6]) ? 8'b11110111 : node5786;
												assign node5786 = (inp[8]) ? 8'b10100001 : 8'b10100101;
										assign node5790 = (inp[8]) ? 8'b10000001 : 8'b10000101;
								assign node5793 = (inp[5]) ? node5831 : node5794;
									assign node5794 = (inp[3]) ? node5814 : node5795;
										assign node5795 = (inp[6]) ? node5805 : node5796;
											assign node5796 = (inp[10]) ? 8'b10100100 : node5797;
												assign node5797 = (inp[8]) ? node5801 : node5798;
													assign node5798 = (inp[9]) ? 8'b10100100 : 8'b10000100;
													assign node5801 = (inp[9]) ? 8'b10100000 : 8'b10000000;
											assign node5805 = (inp[10]) ? node5809 : node5806;
												assign node5806 = (inp[8]) ? 8'b10110000 : 8'b10110100;
												assign node5809 = (inp[13]) ? node5811 : 8'b10110100;
													assign node5811 = (inp[9]) ? 8'b10110100 : 8'b10010100;
										assign node5814 = (inp[6]) ? node5824 : node5815;
											assign node5815 = (inp[9]) ? node5819 : node5816;
												assign node5816 = (inp[10]) ? 8'b10000101 : 8'b10000001;
												assign node5819 = (inp[10]) ? 8'b10100101 : node5820;
													assign node5820 = (inp[8]) ? 8'b10100001 : 8'b10100101;
											assign node5824 = (inp[8]) ? node5826 : 8'b11110111;
												assign node5826 = (inp[10]) ? 8'b11110111 : node5827;
													assign node5827 = (inp[13]) ? 8'b10010001 : 8'b10110001;
									assign node5831 = (inp[13]) ? node5835 : node5832;
										assign node5832 = (inp[8]) ? 8'b10100000 : 8'b10100100;
										assign node5835 = (inp[8]) ? 8'b10000000 : 8'b10000100;
				assign node5838 = (inp[0]) ? node6022 : node5839;
					assign node5839 = (inp[5]) ? node5841 : 8'b00000010;
						assign node5841 = (inp[6]) ? node5903 : node5842;
							assign node5842 = (inp[3]) ? node5862 : node5843;
								assign node5843 = (inp[10]) ? node5849 : node5844;
									assign node5844 = (inp[9]) ? node5846 : 8'b00000010;
										assign node5846 = (inp[13]) ? 8'b10100000 : 8'b00000010;
									assign node5849 = (inp[8]) ? node5855 : node5850;
										assign node5850 = (inp[13]) ? node5852 : 8'b00000010;
											assign node5852 = (inp[9]) ? 8'b10100000 : 8'b00000010;
										assign node5855 = (inp[11]) ? 8'b10100100 : node5856;
											assign node5856 = (inp[9]) ? node5858 : 8'b10000100;
												assign node5858 = (inp[13]) ? 8'b10100100 : 8'b10000100;
								assign node5862 = (inp[1]) ? node5882 : node5863;
									assign node5863 = (inp[9]) ? node5871 : node5864;
										assign node5864 = (inp[8]) ? node5866 : 8'b00000010;
											assign node5866 = (inp[10]) ? node5868 : 8'b00000010;
												assign node5868 = (inp[13]) ? 8'b10000100 : 8'b10100100;
										assign node5871 = (inp[8]) ? node5875 : node5872;
											assign node5872 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node5875 = (inp[10]) ? node5877 : 8'b10100000;
												assign node5877 = (inp[13]) ? node5879 : 8'b10100100;
													assign node5879 = (inp[11]) ? 8'b10000100 : 8'b10100100;
									assign node5882 = (inp[11]) ? node5890 : node5883;
										assign node5883 = (inp[13]) ? node5885 : 8'b10000001;
											assign node5885 = (inp[9]) ? 8'b10100001 : node5886;
												assign node5886 = (inp[2]) ? 8'b10000001 : 8'b10000101;
										assign node5890 = (inp[10]) ? node5896 : node5891;
											assign node5891 = (inp[9]) ? node5893 : 8'b10100101;
												assign node5893 = (inp[13]) ? 8'b10000101 : 8'b10100101;
											assign node5896 = (inp[8]) ? 8'b10100001 : node5897;
												assign node5897 = (inp[2]) ? 8'b10100101 : node5898;
													assign node5898 = (inp[9]) ? 8'b10000101 : 8'b10100101;
							assign node5903 = (inp[2]) ? node5959 : node5904;
								assign node5904 = (inp[8]) ? node5920 : node5905;
									assign node5905 = (inp[9]) ? node5911 : node5906;
										assign node5906 = (inp[3]) ? node5908 : 8'b00000010;
											assign node5908 = (inp[1]) ? 8'b10100101 : 8'b00000010;
										assign node5911 = (inp[13]) ? node5915 : node5912;
											assign node5912 = (inp[1]) ? 8'b10000001 : 8'b00000010;
											assign node5915 = (inp[1]) ? node5917 : 8'b10100000;
												assign node5917 = (inp[3]) ? 8'b10100001 : 8'b10100000;
									assign node5920 = (inp[10]) ? node5938 : node5921;
										assign node5921 = (inp[1]) ? node5927 : node5922;
											assign node5922 = (inp[9]) ? node5924 : 8'b00000010;
												assign node5924 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node5927 = (inp[3]) ? node5931 : node5928;
												assign node5928 = (inp[11]) ? 8'b10100000 : 8'b00000010;
												assign node5931 = (inp[11]) ? node5935 : node5932;
													assign node5932 = (inp[13]) ? 8'b10100001 : 8'b10000001;
													assign node5935 = (inp[13]) ? 8'b10000101 : 8'b10100101;
										assign node5938 = (inp[1]) ? node5950 : node5939;
											assign node5939 = (inp[11]) ? node5945 : node5940;
												assign node5940 = (inp[9]) ? node5942 : 8'b10000100;
													assign node5942 = (inp[13]) ? 8'b10100100 : 8'b10000100;
												assign node5945 = (inp[13]) ? node5947 : 8'b10100100;
													assign node5947 = (inp[9]) ? 8'b10000100 : 8'b10100100;
											assign node5950 = (inp[3]) ? node5954 : node5951;
												assign node5951 = (inp[11]) ? 8'b10100100 : 8'b10000100;
												assign node5954 = (inp[11]) ? 8'b10100001 : node5955;
													assign node5955 = (inp[9]) ? 8'b10100101 : 8'b10000101;
								assign node5959 = (inp[11]) ? node5989 : node5960;
									assign node5960 = (inp[3]) ? node5976 : node5961;
										assign node5961 = (inp[9]) ? node5967 : node5962;
											assign node5962 = (inp[8]) ? node5964 : 8'b10010000;
												assign node5964 = (inp[10]) ? 8'b10010100 : 8'b10010000;
											assign node5967 = (inp[13]) ? node5971 : node5968;
												assign node5968 = (inp[10]) ? 8'b10010100 : 8'b10010000;
												assign node5971 = (inp[10]) ? node5973 : 8'b10110000;
													assign node5973 = (inp[8]) ? 8'b10110100 : 8'b10110000;
										assign node5976 = (inp[1]) ? node5984 : node5977;
											assign node5977 = (inp[10]) ? node5979 : 8'b10010000;
												assign node5979 = (inp[8]) ? node5981 : 8'b10110000;
													assign node5981 = (inp[13]) ? 8'b10110100 : 8'b10010100;
											assign node5984 = (inp[10]) ? node5986 : 8'b10010001;
												assign node5986 = (inp[8]) ? 8'b10010101 : 8'b10010001;
									assign node5989 = (inp[10]) ? node6003 : node5990;
										assign node5990 = (inp[1]) ? node5996 : node5991;
											assign node5991 = (inp[13]) ? node5993 : 8'b11110101;
												assign node5993 = (inp[9]) ? 8'b10010101 : 8'b11110101;
											assign node5996 = (inp[3]) ? node5998 : 8'b11110101;
												assign node5998 = (inp[9]) ? node6000 : 8'b10110100;
													assign node6000 = (inp[13]) ? 8'b10010100 : 8'b10110100;
										assign node6003 = (inp[8]) ? node6009 : node6004;
											assign node6004 = (inp[9]) ? node6006 : 8'b11110101;
												assign node6006 = (inp[13]) ? 8'b10010101 : 8'b11110101;
											assign node6009 = (inp[3]) ? node6015 : node6010;
												assign node6010 = (inp[13]) ? node6012 : 8'b10110001;
													assign node6012 = (inp[9]) ? 8'b10010001 : 8'b10110001;
												assign node6015 = (inp[1]) ? node6017 : 8'b10110001;
													assign node6017 = (inp[13]) ? node6019 : 8'b10110000;
														assign node6019 = (inp[9]) ? 8'b10010000 : 8'b10110000;
					assign node6022 = (inp[2]) ? node6152 : node6023;
						assign node6023 = (inp[1]) ? node6061 : node6024;
							assign node6024 = (inp[13]) ? node6036 : node6025;
								assign node6025 = (inp[8]) ? node6027 : 8'b00000010;
									assign node6027 = (inp[5]) ? node6033 : node6028;
										assign node6028 = (inp[10]) ? 8'b00000010 : node6029;
											assign node6029 = (inp[11]) ? 8'b10100100 : 8'b10000100;
										assign node6033 = (inp[11]) ? 8'b10100100 : 8'b10000100;
								assign node6036 = (inp[8]) ? node6042 : node6037;
									assign node6037 = (inp[9]) ? node6039 : 8'b10100000;
										assign node6039 = (inp[5]) ? 8'b10100000 : 8'b00000010;
									assign node6042 = (inp[5]) ? node6058 : node6043;
										assign node6043 = (inp[10]) ? node6055 : node6044;
											assign node6044 = (inp[6]) ? 8'b10100100 : node6045;
												assign node6045 = (inp[3]) ? 8'b10100100 : node6046;
													assign node6046 = (inp[11]) ? node6050 : node6047;
														assign node6047 = (inp[9]) ? 8'b10000100 : 8'b10100100;
														assign node6050 = (inp[9]) ? 8'b10100100 : 8'b10000100;
											assign node6055 = (inp[9]) ? 8'b00000010 : 8'b10100000;
										assign node6058 = (inp[11]) ? 8'b10000100 : 8'b10100100;
							assign node6061 = (inp[3]) ? node6103 : node6062;
								assign node6062 = (inp[11]) ? node6082 : node6063;
									assign node6063 = (inp[13]) ? node6071 : node6064;
										assign node6064 = (inp[8]) ? node6066 : 8'b10000001;
											assign node6066 = (inp[10]) ? node6068 : 8'b10000101;
												assign node6068 = (inp[5]) ? 8'b10000101 : 8'b10000001;
										assign node6071 = (inp[8]) ? node6077 : node6072;
											assign node6072 = (inp[5]) ? 8'b10100001 : node6073;
												assign node6073 = (inp[9]) ? 8'b10000001 : 8'b10100001;
											assign node6077 = (inp[5]) ? 8'b10100101 : node6078;
												assign node6078 = (inp[10]) ? 8'b10000001 : 8'b10000101;
									assign node6082 = (inp[8]) ? node6090 : node6083;
										assign node6083 = (inp[13]) ? node6085 : 8'b10100101;
											assign node6085 = (inp[9]) ? node6087 : 8'b10000101;
												assign node6087 = (inp[5]) ? 8'b10000101 : 8'b10100101;
										assign node6090 = (inp[13]) ? node6096 : node6091;
											assign node6091 = (inp[5]) ? 8'b10100001 : node6092;
												assign node6092 = (inp[10]) ? 8'b10100101 : 8'b10100001;
											assign node6096 = (inp[5]) ? 8'b10000001 : node6097;
												assign node6097 = (inp[10]) ? node6099 : 8'b10000001;
													assign node6099 = (inp[9]) ? 8'b10100101 : 8'b10000101;
								assign node6103 = (inp[5]) ? node6121 : node6104;
									assign node6104 = (inp[8]) ? node6110 : node6105;
										assign node6105 = (inp[9]) ? 8'b00000010 : node6106;
											assign node6106 = (inp[13]) ? 8'b10100000 : 8'b00000010;
										assign node6110 = (inp[10]) ? node6118 : node6111;
											assign node6111 = (inp[11]) ? node6113 : 8'b10000100;
												assign node6113 = (inp[13]) ? node6115 : 8'b10100100;
													assign node6115 = (inp[9]) ? 8'b10100100 : 8'b10000100;
											assign node6118 = (inp[13]) ? 8'b10100000 : 8'b00000010;
									assign node6121 = (inp[10]) ? node6133 : node6122;
										assign node6122 = (inp[13]) ? node6130 : node6123;
											assign node6123 = (inp[11]) ? node6127 : node6124;
												assign node6124 = (inp[8]) ? 8'b10000101 : 8'b10000001;
												assign node6127 = (inp[8]) ? 8'b10100001 : 8'b10100101;
											assign node6130 = (inp[8]) ? 8'b10000001 : 8'b10000101;
										assign node6133 = (inp[9]) ? node6145 : node6134;
											assign node6134 = (inp[11]) ? node6138 : node6135;
												assign node6135 = (inp[13]) ? 8'b10100001 : 8'b10000001;
												assign node6138 = (inp[8]) ? node6142 : node6139;
													assign node6139 = (inp[13]) ? 8'b10000101 : 8'b10100101;
													assign node6142 = (inp[13]) ? 8'b10000001 : 8'b10100001;
											assign node6145 = (inp[11]) ? node6149 : node6146;
												assign node6146 = (inp[6]) ? 8'b10000001 : 8'b10000101;
												assign node6149 = (inp[13]) ? 8'b10000001 : 8'b10100001;
						assign node6152 = (inp[5]) ? node6262 : node6153;
							assign node6153 = (inp[6]) ? node6209 : node6154;
								assign node6154 = (inp[11]) ? node6178 : node6155;
									assign node6155 = (inp[10]) ? node6167 : node6156;
										assign node6156 = (inp[8]) ? node6158 : 8'b10010000;
											assign node6158 = (inp[1]) ? node6162 : node6159;
												assign node6159 = (inp[9]) ? 8'b10010100 : 8'b10110100;
												assign node6162 = (inp[3]) ? node6164 : 8'b10010101;
													assign node6164 = (inp[13]) ? 8'b10110100 : 8'b10010100;
										assign node6167 = (inp[13]) ? node6173 : node6168;
											assign node6168 = (inp[1]) ? node6170 : 8'b10010000;
												assign node6170 = (inp[3]) ? 8'b10010000 : 8'b10010001;
											assign node6173 = (inp[3]) ? node6175 : 8'b10110001;
												assign node6175 = (inp[9]) ? 8'b10010000 : 8'b10110000;
									assign node6178 = (inp[13]) ? node6194 : node6179;
										assign node6179 = (inp[10]) ? node6189 : node6180;
											assign node6180 = (inp[8]) ? node6184 : node6181;
												assign node6181 = (inp[1]) ? 8'b10110100 : 8'b11110101;
												assign node6184 = (inp[3]) ? 8'b10110001 : node6185;
													assign node6185 = (inp[1]) ? 8'b10110000 : 8'b10110001;
											assign node6189 = (inp[9]) ? node6191 : 8'b11110101;
												assign node6191 = (inp[3]) ? 8'b11110101 : 8'b10110100;
										assign node6194 = (inp[9]) ? node6204 : node6195;
											assign node6195 = (inp[8]) ? node6201 : node6196;
												assign node6196 = (inp[3]) ? 8'b10010101 : node6197;
													assign node6197 = (inp[1]) ? 8'b10010100 : 8'b10010101;
												assign node6201 = (inp[10]) ? 8'b10010101 : 8'b10010001;
											assign node6204 = (inp[3]) ? 8'b11110101 : node6205;
												assign node6205 = (inp[1]) ? 8'b10110100 : 8'b11110101;
								assign node6209 = (inp[3]) ? node6247 : node6210;
									assign node6210 = (inp[1]) ? node6224 : node6211;
										assign node6211 = (inp[11]) ? node6217 : node6212;
											assign node6212 = (inp[10]) ? 8'b00000010 : node6213;
												assign node6213 = (inp[8]) ? 8'b10000100 : 8'b00000010;
											assign node6217 = (inp[9]) ? node6221 : node6218;
												assign node6218 = (inp[13]) ? 8'b10100000 : 8'b00000010;
												assign node6221 = (inp[13]) ? 8'b00000010 : 8'b10100100;
										assign node6224 = (inp[11]) ? node6238 : node6225;
											assign node6225 = (inp[9]) ? node6233 : node6226;
												assign node6226 = (inp[13]) ? node6230 : node6227;
													assign node6227 = (inp[10]) ? 8'b10000001 : 8'b10000101;
													assign node6230 = (inp[8]) ? 8'b10100101 : 8'b10100001;
												assign node6233 = (inp[8]) ? node6235 : 8'b10000001;
													assign node6235 = (inp[10]) ? 8'b10000001 : 8'b10000101;
											assign node6238 = (inp[9]) ? node6244 : node6239;
												assign node6239 = (inp[10]) ? 8'b10000101 : node6240;
													assign node6240 = (inp[8]) ? 8'b10000001 : 8'b10000101;
												assign node6244 = (inp[10]) ? 8'b10100101 : 8'b10100001;
									assign node6247 = (inp[10]) ? node6257 : node6248;
										assign node6248 = (inp[8]) ? node6254 : node6249;
											assign node6249 = (inp[9]) ? 8'b00000010 : node6250;
												assign node6250 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node6254 = (inp[11]) ? 8'b10100100 : 8'b10000100;
										assign node6257 = (inp[9]) ? 8'b00000010 : node6258;
											assign node6258 = (inp[13]) ? 8'b10100000 : 8'b00000010;
							assign node6262 = (inp[6]) ? node6314 : node6263;
								assign node6263 = (inp[3]) ? node6289 : node6264;
									assign node6264 = (inp[11]) ? node6280 : node6265;
										assign node6265 = (inp[1]) ? node6273 : node6266;
											assign node6266 = (inp[8]) ? node6270 : node6267;
												assign node6267 = (inp[13]) ? 8'b10110000 : 8'b10010000;
												assign node6270 = (inp[13]) ? 8'b10110100 : 8'b10010100;
											assign node6273 = (inp[13]) ? node6277 : node6274;
												assign node6274 = (inp[8]) ? 8'b10010101 : 8'b10010001;
												assign node6277 = (inp[8]) ? 8'b11110101 : 8'b10110001;
										assign node6280 = (inp[8]) ? node6284 : node6281;
											assign node6281 = (inp[13]) ? 8'b10010101 : 8'b11110101;
											assign node6284 = (inp[13]) ? 8'b10010000 : node6285;
												assign node6285 = (inp[1]) ? 8'b10110000 : 8'b10110001;
									assign node6289 = (inp[11]) ? node6301 : node6290;
										assign node6290 = (inp[13]) ? node6298 : node6291;
											assign node6291 = (inp[1]) ? node6295 : node6292;
												assign node6292 = (inp[8]) ? 8'b10010100 : 8'b10010000;
												assign node6295 = (inp[8]) ? 8'b10010101 : 8'b10010001;
											assign node6298 = (inp[1]) ? 8'b11110101 : 8'b10110100;
										assign node6301 = (inp[1]) ? node6309 : node6302;
											assign node6302 = (inp[13]) ? node6306 : node6303;
												assign node6303 = (inp[8]) ? 8'b10110001 : 8'b11110101;
												assign node6306 = (inp[8]) ? 8'b10010001 : 8'b10010101;
											assign node6309 = (inp[8]) ? node6311 : 8'b10010100;
												assign node6311 = (inp[13]) ? 8'b10010000 : 8'b10110000;
								assign node6314 = (inp[8]) ? node6330 : node6315;
									assign node6315 = (inp[11]) ? node6323 : node6316;
										assign node6316 = (inp[1]) ? node6320 : node6317;
											assign node6317 = (inp[13]) ? 8'b10110000 : 8'b10010000;
											assign node6320 = (inp[13]) ? 8'b10110001 : 8'b10010001;
										assign node6323 = (inp[13]) ? node6327 : node6324;
											assign node6324 = (inp[1]) ? 8'b10110100 : 8'b11110101;
											assign node6327 = (inp[1]) ? 8'b10010100 : 8'b10010101;
									assign node6330 = (inp[11]) ? node6338 : node6331;
										assign node6331 = (inp[13]) ? node6335 : node6332;
											assign node6332 = (inp[1]) ? 8'b10010101 : 8'b10010100;
											assign node6335 = (inp[1]) ? 8'b11110101 : 8'b10110100;
										assign node6338 = (inp[13]) ? node6342 : node6339;
											assign node6339 = (inp[1]) ? 8'b10110000 : 8'b10110001;
											assign node6342 = (inp[1]) ? 8'b10010000 : 8'b10010001;

endmodule