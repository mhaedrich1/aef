module dtc_split875_bm49 (
	input  wire [7-1:0] inp,
	output wire [10-1:0] outp
);

	wire [10-1:0] node1;
	wire [10-1:0] node2;
	wire [10-1:0] node3;
	wire [10-1:0] node4;
	wire [10-1:0] node5;
	wire [10-1:0] node6;
	wire [10-1:0] node9;
	wire [10-1:0] node12;
	wire [10-1:0] node13;
	wire [10-1:0] node16;
	wire [10-1:0] node19;
	wire [10-1:0] node20;
	wire [10-1:0] node21;
	wire [10-1:0] node24;
	wire [10-1:0] node27;
	wire [10-1:0] node28;
	wire [10-1:0] node31;
	wire [10-1:0] node34;
	wire [10-1:0] node35;
	wire [10-1:0] node36;
	wire [10-1:0] node37;
	wire [10-1:0] node40;
	wire [10-1:0] node43;
	wire [10-1:0] node44;
	wire [10-1:0] node47;
	wire [10-1:0] node50;
	wire [10-1:0] node51;
	wire [10-1:0] node53;
	wire [10-1:0] node56;
	wire [10-1:0] node59;
	wire [10-1:0] node60;
	wire [10-1:0] node61;
	wire [10-1:0] node62;
	wire [10-1:0] node63;
	wire [10-1:0] node66;
	wire [10-1:0] node69;
	wire [10-1:0] node70;
	wire [10-1:0] node73;
	wire [10-1:0] node76;
	wire [10-1:0] node77;
	wire [10-1:0] node78;
	wire [10-1:0] node81;
	wire [10-1:0] node84;
	wire [10-1:0] node85;
	wire [10-1:0] node88;
	wire [10-1:0] node91;
	wire [10-1:0] node92;
	wire [10-1:0] node93;
	wire [10-1:0] node94;
	wire [10-1:0] node97;
	wire [10-1:0] node100;
	wire [10-1:0] node101;
	wire [10-1:0] node104;
	wire [10-1:0] node107;
	wire [10-1:0] node108;
	wire [10-1:0] node109;
	wire [10-1:0] node114;
	wire [10-1:0] node115;
	wire [10-1:0] node116;
	wire [10-1:0] node117;
	wire [10-1:0] node118;
	wire [10-1:0] node119;
	wire [10-1:0] node123;
	wire [10-1:0] node124;
	wire [10-1:0] node128;
	wire [10-1:0] node129;
	wire [10-1:0] node130;
	wire [10-1:0] node133;
	wire [10-1:0] node136;
	wire [10-1:0] node138;
	wire [10-1:0] node141;
	wire [10-1:0] node142;
	wire [10-1:0] node143;
	wire [10-1:0] node144;
	wire [10-1:0] node147;
	wire [10-1:0] node150;
	wire [10-1:0] node151;
	wire [10-1:0] node154;
	wire [10-1:0] node157;
	wire [10-1:0] node158;
	wire [10-1:0] node160;
	wire [10-1:0] node163;
	wire [10-1:0] node164;
	wire [10-1:0] node167;
	wire [10-1:0] node170;
	wire [10-1:0] node171;
	wire [10-1:0] node172;
	wire [10-1:0] node173;
	wire [10-1:0] node174;
	wire [10-1:0] node177;
	wire [10-1:0] node180;
	wire [10-1:0] node183;
	wire [10-1:0] node184;
	wire [10-1:0] node185;
	wire [10-1:0] node189;
	wire [10-1:0] node190;
	wire [10-1:0] node193;
	wire [10-1:0] node196;
	wire [10-1:0] node197;
	wire [10-1:0] node198;
	wire [10-1:0] node200;
	wire [10-1:0] node203;
	wire [10-1:0] node204;
	wire [10-1:0] node207;
	wire [10-1:0] node210;
	wire [10-1:0] node211;
	wire [10-1:0] node213;
	wire [10-1:0] node216;
	wire [10-1:0] node217;
	wire [10-1:0] node220;

	assign outp = (inp[3]) ? node114 : node1;
		assign node1 = (inp[1]) ? node59 : node2;
			assign node2 = (inp[2]) ? node34 : node3;
				assign node3 = (inp[0]) ? node19 : node4;
					assign node4 = (inp[6]) ? node12 : node5;
						assign node5 = (inp[4]) ? node9 : node6;
							assign node6 = (inp[5]) ? 10'b1000010111 : 10'b1101010011;
							assign node9 = (inp[5]) ? 10'b1100011001 : 10'b1001010001;
						assign node12 = (inp[5]) ? node16 : node13;
							assign node13 = (inp[4]) ? 10'b1000001101 : 10'b1100001111;
							assign node16 = (inp[4]) ? 10'b1100000001 : 10'b1000001011;
					assign node19 = (inp[4]) ? node27 : node20;
						assign node20 = (inp[6]) ? node24 : node21;
							assign node21 = (inp[5]) ? 10'b0000010101 : 10'b0101010001;
							assign node24 = (inp[5]) ? 10'b0000001001 : 10'b0100001101;
						assign node27 = (inp[6]) ? node31 : node28;
							assign node28 = (inp[5]) ? 10'b0100001011 : 10'b0001000011;
							assign node31 = (inp[5]) ? 10'b0000010011 : 10'b0100010111;
				assign node34 = (inp[0]) ? node50 : node35;
					assign node35 = (inp[6]) ? node43 : node36;
						assign node36 = (inp[4]) ? node40 : node37;
							assign node37 = (inp[5]) ? 10'b1000000110 : 10'b1101000010;
							assign node40 = (inp[5]) ? 10'b1100001000 : 10'b1001000000;
						assign node43 = (inp[4]) ? node47 : node44;
							assign node44 = (inp[5]) ? 10'b1100010010 : 10'b1000011110;
							assign node47 = (inp[5]) ? 10'b1000010000 : 10'b1100010100;
					assign node50 = (inp[4]) ? node56 : node51;
						assign node51 = (inp[6]) ? node53 : 10'b0101000000;
							assign node53 = (inp[5]) ? 10'b0100010000 : 10'b0000011100;
						assign node56 = (inp[6]) ? 10'b0000000010 : 10'b0100011110;
			assign node59 = (inp[0]) ? node91 : node60;
				assign node60 = (inp[2]) ? node76 : node61;
					assign node61 = (inp[6]) ? node69 : node62;
						assign node62 = (inp[4]) ? node66 : node63;
							assign node63 = (inp[5]) ? 10'b0000110110 : 10'b0101110010;
							assign node66 = (inp[5]) ? 10'b0100111000 : 10'b0001110000;
						assign node69 = (inp[5]) ? node73 : node70;
							assign node70 = (inp[4]) ? 10'b0000101100 : 10'b0100101110;
							assign node73 = (inp[4]) ? 10'b0100100000 : 10'b0000101010;
					assign node76 = (inp[4]) ? node84 : node77;
						assign node77 = (inp[6]) ? node81 : node78;
							assign node78 = (inp[5]) ? 10'b0000100101 : 10'b0101100001;
							assign node81 = (inp[5]) ? 10'b0100110001 : 10'b0000111101;
						assign node84 = (inp[5]) ? node88 : node85;
							assign node85 = (inp[6]) ? 10'b0100100111 : 10'b0100111111;
							assign node88 = (inp[6]) ? 10'b0000100011 : 10'b0000111011;
				assign node91 = (inp[2]) ? node107 : node92;
					assign node92 = (inp[6]) ? node100 : node93;
						assign node93 = (inp[4]) ? node97 : node94;
							assign node94 = (inp[5]) ? 10'b1000100111 : 10'b1101100011;
							assign node97 = (inp[5]) ? 10'b1100101001 : 10'b1001100001;
						assign node100 = (inp[4]) ? node104 : node101;
							assign node101 = (inp[5]) ? 10'b1100110011 : 10'b1000111111;
							assign node104 = (inp[5]) ? 10'b1000110001 : 10'b1100110101;
					assign node107 = (inp[4]) ? 10'b1100111100 : node108;
						assign node108 = (inp[6]) ? 10'b1000101110 : node109;
							assign node109 = (inp[5]) ? 10'b1100111010 : 10'b1001110010;
		assign node114 = (inp[1]) ? node170 : node115;
			assign node115 = (inp[2]) ? node141 : node116;
				assign node116 = (inp[0]) ? node128 : node117;
					assign node117 = (inp[6]) ? node123 : node118;
						assign node118 = (inp[5]) ? 10'b1110111000 : node119;
							assign node119 = (inp[4]) ? 10'b1011110000 : 10'b1111110010;
						assign node123 = (inp[4]) ? 10'b1010101100 : node124;
							assign node124 = (inp[5]) ? 10'b1010101010 : 10'b1110101110;
					assign node128 = (inp[4]) ? node136 : node129;
						assign node129 = (inp[6]) ? node133 : node130;
							assign node130 = (inp[5]) ? 10'b0010110100 : 10'b0111110000;
							assign node133 = (inp[5]) ? 10'b0010101000 : 10'b0110101100;
						assign node136 = (inp[6]) ? node138 : 10'b0110101010;
							assign node138 = (inp[5]) ? 10'b0010110010 : 10'b0110110110;
				assign node141 = (inp[0]) ? node157 : node142;
					assign node142 = (inp[4]) ? node150 : node143;
						assign node143 = (inp[6]) ? node147 : node144;
							assign node144 = (inp[5]) ? 10'b1010100101 : 10'b1111100001;
							assign node147 = (inp[5]) ? 10'b1110110001 : 10'b1010111101;
						assign node150 = (inp[6]) ? node154 : node151;
							assign node151 = (inp[5]) ? 10'b1010111011 : 10'b1110111111;
							assign node154 = (inp[5]) ? 10'b1010100011 : 10'b1110100111;
					assign node157 = (inp[6]) ? node163 : node158;
						assign node158 = (inp[4]) ? node160 : 10'b0110111011;
							assign node160 = (inp[5]) ? 10'b0010111001 : 10'b0110111101;
						assign node163 = (inp[4]) ? node167 : node164;
							assign node164 = (inp[5]) ? 10'b0110100011 : 10'b0010101111;
							assign node167 = (inp[5]) ? 10'b0010100001 : 10'b0110100101;
			assign node170 = (inp[2]) ? node196 : node171;
				assign node171 = (inp[0]) ? node183 : node172;
					assign node172 = (inp[4]) ? node180 : node173;
						assign node173 = (inp[6]) ? node177 : node174;
							assign node174 = (inp[5]) ? 10'b1010010101 : 10'b1111010001;
							assign node177 = (inp[5]) ? 10'b1010001001 : 10'b1110001101;
						assign node180 = (inp[6]) ? 10'b1010010011 : 10'b1011000011;
					assign node183 = (inp[6]) ? node189 : node184;
						assign node184 = (inp[5]) ? 10'b0110001001 : node185;
							assign node185 = (inp[4]) ? 10'b0011000001 : 10'b0111000011;
						assign node189 = (inp[5]) ? node193 : node190;
							assign node190 = (inp[4]) ? 10'b0110010101 : 10'b0010011111;
							assign node193 = (inp[4]) ? 10'b0010010001 : 10'b0110010011;
				assign node196 = (inp[0]) ? node210 : node197;
					assign node197 = (inp[4]) ? node203 : node198;
						assign node198 = (inp[6]) ? node200 : 10'b1111000000;
							assign node200 = (inp[5]) ? 10'b1110010000 : 10'b1010011100;
						assign node203 = (inp[6]) ? node207 : node204;
							assign node204 = (inp[5]) ? 10'b1010011010 : 10'b1110011110;
							assign node207 = (inp[5]) ? 10'b1010000010 : 10'b1110000110;
					assign node210 = (inp[6]) ? node216 : node211;
						assign node211 = (inp[4]) ? node213 : 10'b0011010010;
							assign node213 = (inp[5]) ? 10'b0010011000 : 10'b0110011100;
						assign node216 = (inp[4]) ? node220 : node217;
							assign node217 = (inp[5]) ? 10'b0110000010 : 10'b0010001110;
							assign node220 = (inp[5]) ? 10'b0010000000 : 10'b0110000100;

endmodule