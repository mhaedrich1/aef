module dtc_split5_bm66 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node9;
	wire [4-1:0] node11;
	wire [4-1:0] node13;
	wire [4-1:0] node15;
	wire [4-1:0] node16;
	wire [4-1:0] node18;
	wire [4-1:0] node22;
	wire [4-1:0] node23;
	wire [4-1:0] node24;
	wire [4-1:0] node25;
	wire [4-1:0] node27;
	wire [4-1:0] node29;
	wire [4-1:0] node31;
	wire [4-1:0] node34;
	wire [4-1:0] node37;
	wire [4-1:0] node38;
	wire [4-1:0] node39;
	wire [4-1:0] node45;
	wire [4-1:0] node46;
	wire [4-1:0] node48;
	wire [4-1:0] node50;
	wire [4-1:0] node52;
	wire [4-1:0] node54;
	wire [4-1:0] node57;
	wire [4-1:0] node58;
	wire [4-1:0] node60;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node65;
	wire [4-1:0] node67;
	wire [4-1:0] node71;
	wire [4-1:0] node72;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node76;
	wire [4-1:0] node78;
	wire [4-1:0] node84;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node88;
	wire [4-1:0] node90;
	wire [4-1:0] node91;
	wire [4-1:0] node93;
	wire [4-1:0] node94;
	wire [4-1:0] node96;
	wire [4-1:0] node98;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node104;
	wire [4-1:0] node105;
	wire [4-1:0] node107;
	wire [4-1:0] node113;
	wire [4-1:0] node114;
	wire [4-1:0] node115;
	wire [4-1:0] node117;
	wire [4-1:0] node118;
	wire [4-1:0] node120;
	wire [4-1:0] node122;
	wire [4-1:0] node124;
	wire [4-1:0] node126;
	wire [4-1:0] node130;
	wire [4-1:0] node131;
	wire [4-1:0] node132;
	wire [4-1:0] node134;
	wire [4-1:0] node135;
	wire [4-1:0] node137;
	wire [4-1:0] node144;
	wire [4-1:0] node145;
	wire [4-1:0] node147;
	wire [4-1:0] node149;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node153;
	wire [4-1:0] node155;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node162;
	wire [4-1:0] node163;
	wire [4-1:0] node165;
	wire [4-1:0] node167;
	wire [4-1:0] node169;
	wire [4-1:0] node174;
	wire [4-1:0] node176;
	wire [4-1:0] node178;
	wire [4-1:0] node179;
	wire [4-1:0] node181;
	wire [4-1:0] node183;
	wire [4-1:0] node184;
	wire [4-1:0] node186;
	wire [4-1:0] node191;
	wire [4-1:0] node192;
	wire [4-1:0] node193;
	wire [4-1:0] node194;
	wire [4-1:0] node195;
	wire [4-1:0] node196;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node201;
	wire [4-1:0] node203;
	wire [4-1:0] node207;
	wire [4-1:0] node209;
	wire [4-1:0] node211;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node218;
	wire [4-1:0] node220;
	wire [4-1:0] node222;
	wire [4-1:0] node224;
	wire [4-1:0] node228;
	wire [4-1:0] node229;
	wire [4-1:0] node231;
	wire [4-1:0] node233;
	wire [4-1:0] node235;
	wire [4-1:0] node241;
	wire [4-1:0] node243;
	wire [4-1:0] node244;
	wire [4-1:0] node246;
	wire [4-1:0] node248;
	wire [4-1:0] node250;
	wire [4-1:0] node252;
	wire [4-1:0] node255;
	wire [4-1:0] node258;
	wire [4-1:0] node259;
	wire [4-1:0] node260;
	wire [4-1:0] node261;
	wire [4-1:0] node263;
	wire [4-1:0] node264;
	wire [4-1:0] node266;
	wire [4-1:0] node268;
	wire [4-1:0] node270;
	wire [4-1:0] node272;
	wire [4-1:0] node275;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node282;
	wire [4-1:0] node283;
	wire [4-1:0] node285;
	wire [4-1:0] node287;
	wire [4-1:0] node289;
	wire [4-1:0] node291;
	wire [4-1:0] node296;
	wire [4-1:0] node297;
	wire [4-1:0] node298;
	wire [4-1:0] node299;
	wire [4-1:0] node300;
	wire [4-1:0] node302;
	wire [4-1:0] node304;
	wire [4-1:0] node309;
	wire [4-1:0] node311;
	wire [4-1:0] node312;
	wire [4-1:0] node313;
	wire [4-1:0] node314;
	wire [4-1:0] node316;
	wire [4-1:0] node318;
	wire [4-1:0] node324;
	wire [4-1:0] node326;
	wire [4-1:0] node327;
	wire [4-1:0] node328;
	wire [4-1:0] node330;
	wire [4-1:0] node332;
	wire [4-1:0] node334;
	wire [4-1:0] node336;
	wire [4-1:0] node341;
	wire [4-1:0] node342;
	wire [4-1:0] node343;
	wire [4-1:0] node344;
	wire [4-1:0] node345;
	wire [4-1:0] node346;
	wire [4-1:0] node348;
	wire [4-1:0] node350;
	wire [4-1:0] node352;
	wire [4-1:0] node356;
	wire [4-1:0] node358;
	wire [4-1:0] node359;
	wire [4-1:0] node361;
	wire [4-1:0] node362;
	wire [4-1:0] node364;
	wire [4-1:0] node366;
	wire [4-1:0] node371;
	wire [4-1:0] node372;
	wire [4-1:0] node374;
	wire [4-1:0] node375;
	wire [4-1:0] node376;
	wire [4-1:0] node378;
	wire [4-1:0] node380;
	wire [4-1:0] node385;
	wire [4-1:0] node387;
	wire [4-1:0] node388;
	wire [4-1:0] node390;
	wire [4-1:0] node392;
	wire [4-1:0] node396;
	wire [4-1:0] node397;
	wire [4-1:0] node398;
	wire [4-1:0] node400;
	wire [4-1:0] node402;
	wire [4-1:0] node405;
	wire [4-1:0] node407;
	wire [4-1:0] node409;
	wire [4-1:0] node410;
	wire [4-1:0] node411;
	wire [4-1:0] node413;
	wire [4-1:0] node415;
	wire [4-1:0] node420;
	wire [4-1:0] node422;
	wire [4-1:0] node424;
	wire [4-1:0] node426;
	wire [4-1:0] node429;
	wire [4-1:0] node430;
	wire [4-1:0] node431;
	wire [4-1:0] node432;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node436;
	wire [4-1:0] node438;
	wire [4-1:0] node440;
	wire [4-1:0] node446;
	wire [4-1:0] node448;
	wire [4-1:0] node449;
	wire [4-1:0] node451;
	wire [4-1:0] node453;
	wire [4-1:0] node455;
	wire [4-1:0] node460;
	wire [4-1:0] node462;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node467;
	wire [4-1:0] node469;
	wire [4-1:0] node471;
	wire [4-1:0] node472;
	wire [4-1:0] node476;
	wire [4-1:0] node478;
	wire [4-1:0] node480;
	wire [4-1:0] node482;
	wire [4-1:0] node485;
	wire [4-1:0] node486;
	wire [4-1:0] node487;
	wire [4-1:0] node488;
	wire [4-1:0] node489;
	wire [4-1:0] node491;
	wire [4-1:0] node493;
	wire [4-1:0] node498;
	wire [4-1:0] node501;
	wire [4-1:0] node503;
	wire [4-1:0] node505;
	wire [4-1:0] node507;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node516;
	wire [4-1:0] node517;
	wire [4-1:0] node518;
	wire [4-1:0] node519;
	wire [4-1:0] node520;
	wire [4-1:0] node522;
	wire [4-1:0] node524;
	wire [4-1:0] node525;
	wire [4-1:0] node526;
	wire [4-1:0] node528;
	wire [4-1:0] node530;
	wire [4-1:0] node536;
	wire [4-1:0] node537;
	wire [4-1:0] node539;
	wire [4-1:0] node540;
	wire [4-1:0] node542;
	wire [4-1:0] node544;
	wire [4-1:0] node548;
	wire [4-1:0] node550;
	wire [4-1:0] node552;
	wire [4-1:0] node555;
	wire [4-1:0] node556;
	wire [4-1:0] node558;
	wire [4-1:0] node559;
	wire [4-1:0] node560;
	wire [4-1:0] node562;
	wire [4-1:0] node563;
	wire [4-1:0] node565;
	wire [4-1:0] node567;
	wire [4-1:0] node573;
	wire [4-1:0] node575;
	wire [4-1:0] node576;
	wire [4-1:0] node578;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node584;
	wire [4-1:0] node590;
	wire [4-1:0] node591;
	wire [4-1:0] node592;
	wire [4-1:0] node593;
	wire [4-1:0] node595;
	wire [4-1:0] node597;
	wire [4-1:0] node600;
	wire [4-1:0] node602;
	wire [4-1:0] node604;
	wire [4-1:0] node606;
	wire [4-1:0] node608;
	wire [4-1:0] node612;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node616;
	wire [4-1:0] node618;
	wire [4-1:0] node620;
	wire [4-1:0] node622;
	wire [4-1:0] node624;
	wire [4-1:0] node627;
	wire [4-1:0] node628;
	wire [4-1:0] node629;
	wire [4-1:0] node630;
	wire [4-1:0] node631;
	wire [4-1:0] node633;
	wire [4-1:0] node641;
	wire [4-1:0] node642;
	wire [4-1:0] node643;
	wire [4-1:0] node644;
	wire [4-1:0] node645;
	wire [4-1:0] node646;
	wire [4-1:0] node647;
	wire [4-1:0] node649;
	wire [4-1:0] node651;
	wire [4-1:0] node656;
	wire [4-1:0] node658;
	wire [4-1:0] node660;
	wire [4-1:0] node661;
	wire [4-1:0] node663;
	wire [4-1:0] node665;
	wire [4-1:0] node669;
	wire [4-1:0] node671;
	wire [4-1:0] node674;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node681;
	wire [4-1:0] node682;
	wire [4-1:0] node684;
	wire [4-1:0] node686;
	wire [4-1:0] node688;
	wire [4-1:0] node694;
	wire [4-1:0] node695;
	wire [4-1:0] node696;
	wire [4-1:0] node698;
	wire [4-1:0] node700;
	wire [4-1:0] node702;
	wire [4-1:0] node706;
	wire [4-1:0] node709;
	wire [4-1:0] node710;
	wire [4-1:0] node711;
	wire [4-1:0] node713;
	wire [4-1:0] node714;
	wire [4-1:0] node716;
	wire [4-1:0] node718;
	wire [4-1:0] node720;
	wire [4-1:0] node722;
	wire [4-1:0] node724;
	wire [4-1:0] node728;
	wire [4-1:0] node729;
	wire [4-1:0] node731;
	wire [4-1:0] node733;
	wire [4-1:0] node735;
	wire [4-1:0] node737;
	wire [4-1:0] node741;
	wire [4-1:0] node742;
	wire [4-1:0] node743;
	wire [4-1:0] node744;
	wire [4-1:0] node746;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node751;
	wire [4-1:0] node756;
	wire [4-1:0] node758;
	wire [4-1:0] node760;
	wire [4-1:0] node763;
	wire [4-1:0] node765;
	wire [4-1:0] node766;
	wire [4-1:0] node768;
	wire [4-1:0] node769;
	wire [4-1:0] node770;
	wire [4-1:0] node772;
	wire [4-1:0] node774;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node782;
	wire [4-1:0] node783;
	wire [4-1:0] node784;
	wire [4-1:0] node786;
	wire [4-1:0] node788;
	wire [4-1:0] node790;
	wire [4-1:0] node791;
	wire [4-1:0] node793;
	wire [4-1:0] node795;
	wire [4-1:0] node797;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node803;
	wire [4-1:0] node807;
	wire [4-1:0] node808;
	wire [4-1:0] node809;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node814;
	wire [4-1:0] node816;
	wire [4-1:0] node818;
	wire [4-1:0] node822;
	wire [4-1:0] node823;
	wire [4-1:0] node824;
	wire [4-1:0] node825;
	wire [4-1:0] node827;
	wire [4-1:0] node829;
	wire [4-1:0] node835;
	wire [4-1:0] node837;
	wire [4-1:0] node839;
	wire [4-1:0] node842;
	wire [4-1:0] node843;
	wire [4-1:0] node845;
	wire [4-1:0] node847;
	wire [4-1:0] node849;
	wire [4-1:0] node850;
	wire [4-1:0] node852;
	wire [4-1:0] node856;
	wire [4-1:0] node857;
	wire [4-1:0] node858;
	wire [4-1:0] node859;
	wire [4-1:0] node861;
	wire [4-1:0] node863;
	wire [4-1:0] node868;
	wire [4-1:0] node870;
	wire [4-1:0] node871;
	wire [4-1:0] node873;
	wire [4-1:0] node874;
	wire [4-1:0] node876;
	wire [4-1:0] node878;
	wire [4-1:0] node883;
	wire [4-1:0] node884;
	wire [4-1:0] node885;
	wire [4-1:0] node886;
	wire [4-1:0] node888;
	wire [4-1:0] node890;
	wire [4-1:0] node892;
	wire [4-1:0] node894;
	wire [4-1:0] node897;
	wire [4-1:0] node898;
	wire [4-1:0] node900;
	wire [4-1:0] node901;
	wire [4-1:0] node902;
	wire [4-1:0] node904;
	wire [4-1:0] node906;
	wire [4-1:0] node912;
	wire [4-1:0] node913;
	wire [4-1:0] node915;
	wire [4-1:0] node916;
	wire [4-1:0] node918;
	wire [4-1:0] node920;
	wire [4-1:0] node922;
	wire [4-1:0] node924;
	wire [4-1:0] node928;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node932;
	wire [4-1:0] node934;
	wire [4-1:0] node939;
	wire [4-1:0] node940;
	wire [4-1:0] node941;
	wire [4-1:0] node943;
	wire [4-1:0] node944;
	wire [4-1:0] node945;
	wire [4-1:0] node947;
	wire [4-1:0] node949;
	wire [4-1:0] node951;
	wire [4-1:0] node956;
	wire [4-1:0] node959;
	wire [4-1:0] node960;
	wire [4-1:0] node962;
	wire [4-1:0] node963;
	wire [4-1:0] node965;
	wire [4-1:0] node967;
	wire [4-1:0] node969;
	wire [4-1:0] node973;
	wire [4-1:0] node974;
	wire [4-1:0] node976;
	wire [4-1:0] node978;
	wire [4-1:0] node980;
	wire [4-1:0] node984;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node987;
	wire [4-1:0] node988;
	wire [4-1:0] node989;
	wire [4-1:0] node990;
	wire [4-1:0] node994;
	wire [4-1:0] node995;
	wire [4-1:0] node996;
	wire [4-1:0] node997;
	wire [4-1:0] node999;
	wire [4-1:0] node1001;
	wire [4-1:0] node1006;
	wire [4-1:0] node1009;
	wire [4-1:0] node1011;
	wire [4-1:0] node1012;
	wire [4-1:0] node1013;
	wire [4-1:0] node1014;
	wire [4-1:0] node1016;
	wire [4-1:0] node1018;
	wire [4-1:0] node1024;
	wire [4-1:0] node1025;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1029;
	wire [4-1:0] node1031;
	wire [4-1:0] node1033;
	wire [4-1:0] node1035;
	wire [4-1:0] node1038;
	wire [4-1:0] node1040;
	wire [4-1:0] node1041;
	wire [4-1:0] node1043;
	wire [4-1:0] node1045;
	wire [4-1:0] node1049;
	wire [4-1:0] node1051;
	wire [4-1:0] node1054;
	wire [4-1:0] node1055;
	wire [4-1:0] node1056;
	wire [4-1:0] node1060;
	wire [4-1:0] node1061;
	wire [4-1:0] node1062;
	wire [4-1:0] node1064;
	wire [4-1:0] node1068;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1073;
	wire [4-1:0] node1074;
	wire [4-1:0] node1075;
	wire [4-1:0] node1077;
	wire [4-1:0] node1079;
	wire [4-1:0] node1084;
	wire [4-1:0] node1086;
	wire [4-1:0] node1088;
	wire [4-1:0] node1089;
	wire [4-1:0] node1090;
	wire [4-1:0] node1092;
	wire [4-1:0] node1094;
	wire [4-1:0] node1098;
	wire [4-1:0] node1100;
	wire [4-1:0] node1102;
	wire [4-1:0] node1104;
	wire [4-1:0] node1107;
	wire [4-1:0] node1108;
	wire [4-1:0] node1109;
	wire [4-1:0] node1111;
	wire [4-1:0] node1115;
	wire [4-1:0] node1117;
	wire [4-1:0] node1119;
	wire [4-1:0] node1121;
	wire [4-1:0] node1123;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1128;
	wire [4-1:0] node1129;
	wire [4-1:0] node1131;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1136;
	wire [4-1:0] node1138;
	wire [4-1:0] node1140;
	wire [4-1:0] node1143;
	wire [4-1:0] node1144;
	wire [4-1:0] node1146;
	wire [4-1:0] node1148;
	wire [4-1:0] node1152;
	wire [4-1:0] node1154;
	wire [4-1:0] node1156;
	wire [4-1:0] node1157;
	wire [4-1:0] node1159;
	wire [4-1:0] node1163;
	wire [4-1:0] node1164;
	wire [4-1:0] node1165;
	wire [4-1:0] node1166;
	wire [4-1:0] node1168;
	wire [4-1:0] node1169;
	wire [4-1:0] node1171;
	wire [4-1:0] node1173;
	wire [4-1:0] node1177;
	wire [4-1:0] node1179;
	wire [4-1:0] node1180;
	wire [4-1:0] node1184;
	wire [4-1:0] node1185;
	wire [4-1:0] node1188;
	wire [4-1:0] node1191;
	wire [4-1:0] node1192;
	wire [4-1:0] node1194;
	wire [4-1:0] node1195;
	wire [4-1:0] node1197;
	wire [4-1:0] node1199;
	wire [4-1:0] node1201;
	wire [4-1:0] node1203;
	wire [4-1:0] node1206;
	wire [4-1:0] node1208;
	wire [4-1:0] node1210;
	wire [4-1:0] node1212;
	wire [4-1:0] node1215;
	wire [4-1:0] node1217;
	wire [4-1:0] node1219;
	wire [4-1:0] node1221;
	wire [4-1:0] node1224;
	wire [4-1:0] node1225;
	wire [4-1:0] node1226;
	wire [4-1:0] node1227;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1232;
	wire [4-1:0] node1234;
	wire [4-1:0] node1236;
	wire [4-1:0] node1240;
	wire [4-1:0] node1241;
	wire [4-1:0] node1242;
	wire [4-1:0] node1243;
	wire [4-1:0] node1245;
	wire [4-1:0] node1247;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1257;
	wire [4-1:0] node1259;
	wire [4-1:0] node1263;
	wire [4-1:0] node1265;
	wire [4-1:0] node1266;
	wire [4-1:0] node1268;
	wire [4-1:0] node1270;
	wire [4-1:0] node1274;
	wire [4-1:0] node1275;
	wire [4-1:0] node1276;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1281;
	wire [4-1:0] node1283;
	wire [4-1:0] node1285;
	wire [4-1:0] node1288;
	wire [4-1:0] node1289;
	wire [4-1:0] node1291;
	wire [4-1:0] node1293;
	wire [4-1:0] node1297;
	wire [4-1:0] node1299;
	wire [4-1:0] node1300;
	wire [4-1:0] node1302;
	wire [4-1:0] node1306;
	wire [4-1:0] node1307;
	wire [4-1:0] node1308;
	wire [4-1:0] node1309;
	wire [4-1:0] node1311;
	wire [4-1:0] node1313;
	wire [4-1:0] node1315;
	wire [4-1:0] node1316;
	wire [4-1:0] node1320;
	wire [4-1:0] node1322;
	wire [4-1:0] node1324;
	wire [4-1:0] node1326;
	wire [4-1:0] node1328;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1334;
	wire [4-1:0] node1338;
	wire [4-1:0] node1339;
	wire [4-1:0] node1340;
	wire [4-1:0] node1342;
	wire [4-1:0] node1344;
	wire [4-1:0] node1346;
	wire [4-1:0] node1349;
	wire [4-1:0] node1350;
	wire [4-1:0] node1352;
	wire [4-1:0] node1356;
	wire [4-1:0] node1357;
	wire [4-1:0] node1359;
	wire [4-1:0] node1362;
	wire [4-1:0] node1363;
	wire [4-1:0] node1364;
	wire [4-1:0] node1366;
	wire [4-1:0] node1370;
	wire [4-1:0] node1372;

	assign outp = (inp[10]) ? node514 : node1;
		assign node1 = (inp[5]) ? node191 : node2;
			assign node2 = (inp[4]) ? node84 : node3;
				assign node3 = (inp[14]) ? node45 : node4;
					assign node4 = (inp[13]) ? node6 : 4'b1111;
						assign node6 = (inp[12]) ? node22 : node7;
							assign node7 = (inp[8]) ? node9 : 4'b1111;
								assign node9 = (inp[2]) ? node11 : 4'b1111;
									assign node11 = (inp[6]) ? node13 : 4'b1111;
										assign node13 = (inp[9]) ? node15 : 4'b1111;
											assign node15 = (inp[7]) ? 4'b1101 : node16;
												assign node16 = (inp[1]) ? node18 : 4'b1111;
													assign node18 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node22 = (inp[2]) ? 4'b1101 : node23;
								assign node23 = (inp[6]) ? node37 : node24;
									assign node24 = (inp[8]) ? node34 : node25;
										assign node25 = (inp[11]) ? node27 : 4'b1111;
											assign node27 = (inp[7]) ? node29 : 4'b1111;
												assign node29 = (inp[15]) ? node31 : 4'b1111;
													assign node31 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node34 = (inp[9]) ? 4'b1101 : 4'b1111;
									assign node37 = (inp[9]) ? 4'b1101 : node38;
										assign node38 = (inp[7]) ? 4'b1101 : node39;
											assign node39 = (inp[8]) ? 4'b1101 : 4'b1111;
					assign node45 = (inp[13]) ? node57 : node46;
						assign node46 = (inp[12]) ? node48 : 4'b1101;
							assign node48 = (inp[8]) ? node50 : 4'b1101;
								assign node50 = (inp[2]) ? node52 : 4'b1101;
									assign node52 = (inp[6]) ? node54 : 4'b1101;
										assign node54 = (inp[9]) ? 4'b1011 : 4'b1101;
						assign node57 = (inp[12]) ? node71 : node58;
							assign node58 = (inp[2]) ? node60 : 4'b1101;
								assign node60 = (inp[9]) ? node62 : 4'b1101;
									assign node62 = (inp[8]) ? node64 : 4'b1101;
										assign node64 = (inp[6]) ? 4'b1011 : node65;
											assign node65 = (inp[15]) ? node67 : 4'b1101;
												assign node67 = (inp[7]) ? 4'b1111 : 4'b1101;
							assign node71 = (inp[6]) ? 4'b1011 : node72;
								assign node72 = (inp[2]) ? 4'b1111 : node73;
									assign node73 = (inp[9]) ? 4'b1111 : node74;
										assign node74 = (inp[7]) ? node76 : 4'b1101;
											assign node76 = (inp[8]) ? node78 : 4'b1101;
												assign node78 = (inp[15]) ? 4'b1111 : 4'b1101;
				assign node84 = (inp[14]) ? node144 : node85;
					assign node85 = (inp[12]) ? node113 : node86;
						assign node86 = (inp[2]) ? node88 : 4'b1011;
							assign node88 = (inp[13]) ? node90 : 4'b1011;
								assign node90 = (inp[9]) ? node102 : node91;
									assign node91 = (inp[6]) ? node93 : 4'b1011;
										assign node93 = (inp[8]) ? 4'b1001 : node94;
											assign node94 = (inp[15]) ? node96 : 4'b1011;
												assign node96 = (inp[11]) ? node98 : 4'b1011;
													assign node98 = (inp[1]) ? 4'b1001 : 4'b1011;
									assign node102 = (inp[8]) ? 4'b1001 : node103;
										assign node103 = (inp[6]) ? 4'b1001 : node104;
											assign node104 = (inp[7]) ? 4'b1001 : node105;
												assign node105 = (inp[15]) ? node107 : 4'b1011;
													assign node107 = (inp[11]) ? 4'b1001 : 4'b1011;
						assign node113 = (inp[13]) ? 4'b1001 : node114;
							assign node114 = (inp[2]) ? node130 : node115;
								assign node115 = (inp[6]) ? node117 : 4'b1011;
									assign node117 = (inp[9]) ? 4'b1001 : node118;
										assign node118 = (inp[15]) ? node120 : 4'b1011;
											assign node120 = (inp[11]) ? node122 : 4'b1011;
												assign node122 = (inp[8]) ? node124 : 4'b1011;
													assign node124 = (inp[1]) ? node126 : 4'b1011;
														assign node126 = (inp[7]) ? 4'b1001 : 4'b1011;
								assign node130 = (inp[6]) ? 4'b1001 : node131;
									assign node131 = (inp[9]) ? 4'b1001 : node132;
										assign node132 = (inp[8]) ? node134 : 4'b1011;
											assign node134 = (inp[7]) ? 4'b1001 : node135;
												assign node135 = (inp[11]) ? node137 : 4'b1011;
													assign node137 = (inp[0]) ? 4'b1001 : 4'b1011;
					assign node144 = (inp[12]) ? node160 : node145;
						assign node145 = (inp[13]) ? node147 : 4'b1001;
							assign node147 = (inp[2]) ? node149 : 4'b1001;
								assign node149 = (inp[6]) ? 4'b1111 : node150;
									assign node150 = (inp[9]) ? 4'b1011 : node151;
										assign node151 = (inp[8]) ? node153 : 4'b1001;
											assign node153 = (inp[7]) ? node155 : 4'b1001;
												assign node155 = (inp[15]) ? 4'b1011 : 4'b1001;
						assign node160 = (inp[6]) ? node174 : node161;
							assign node161 = (inp[2]) ? 4'b1011 : node162;
								assign node162 = (inp[13]) ? 4'b1011 : node163;
									assign node163 = (inp[15]) ? node165 : 4'b1001;
										assign node165 = (inp[9]) ? node167 : 4'b1001;
											assign node167 = (inp[8]) ? node169 : 4'b1001;
												assign node169 = (inp[7]) ? 4'b1011 : 4'b1001;
							assign node174 = (inp[2]) ? node176 : 4'b1110;
								assign node176 = (inp[13]) ? node178 : 4'b1110;
									assign node178 = (inp[9]) ? 4'b1100 : node179;
										assign node179 = (inp[1]) ? node181 : 4'b1110;
											assign node181 = (inp[7]) ? node183 : 4'b1110;
												assign node183 = (inp[3]) ? 4'b1110 : node184;
													assign node184 = (inp[0]) ? node186 : 4'b1110;
														assign node186 = (inp[11]) ? 4'b1100 : 4'b1110;
			assign node191 = (inp[12]) ? node341 : node192;
				assign node192 = (inp[6]) ? node258 : node193;
					assign node193 = (inp[13]) ? node241 : node194;
						assign node194 = (inp[14]) ? node214 : node195;
							assign node195 = (inp[4]) ? node207 : node196;
								assign node196 = (inp[2]) ? node198 : 4'b1001;
									assign node198 = (inp[9]) ? 4'b1011 : node199;
										assign node199 = (inp[8]) ? node201 : 4'b1001;
											assign node201 = (inp[15]) ? node203 : 4'b1001;
												assign node203 = (inp[7]) ? 4'b1011 : 4'b1001;
								assign node207 = (inp[2]) ? node209 : 4'b1101;
									assign node209 = (inp[9]) ? node211 : 4'b1101;
										assign node211 = (inp[8]) ? 4'b1011 : 4'b1101;
							assign node214 = (inp[9]) ? 4'b1001 : node215;
								assign node215 = (inp[2]) ? 4'b1001 : node216;
									assign node216 = (inp[8]) ? node228 : node217;
										assign node217 = (inp[3]) ? 4'b1011 : node218;
											assign node218 = (inp[15]) ? node220 : 4'b1011;
												assign node220 = (inp[11]) ? node222 : 4'b1011;
													assign node222 = (inp[7]) ? node224 : 4'b1011;
														assign node224 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node228 = (inp[7]) ? 4'b1001 : node229;
											assign node229 = (inp[4]) ? node231 : 4'b1001;
												assign node231 = (inp[1]) ? node233 : 4'b1011;
													assign node233 = (inp[15]) ? node235 : 4'b1011;
														assign node235 = (inp[11]) ? 4'b1001 : 4'b1011;
						assign node241 = (inp[14]) ? node243 : 4'b1011;
							assign node243 = (inp[2]) ? node255 : node244;
								assign node244 = (inp[7]) ? node246 : 4'b1001;
									assign node246 = (inp[15]) ? node248 : 4'b1001;
										assign node248 = (inp[4]) ? node250 : 4'b1001;
											assign node250 = (inp[8]) ? node252 : 4'b1001;
												assign node252 = (inp[9]) ? 4'b1011 : 4'b1001;
								assign node255 = (inp[4]) ? 4'b1011 : 4'b1111;
					assign node258 = (inp[14]) ? node296 : node259;
						assign node259 = (inp[4]) ? node279 : node260;
							assign node260 = (inp[13]) ? 4'b1101 : node261;
								assign node261 = (inp[9]) ? node263 : 4'b1111;
									assign node263 = (inp[8]) ? node275 : node264;
										assign node264 = (inp[7]) ? node266 : 4'b1111;
											assign node266 = (inp[11]) ? node268 : 4'b1111;
												assign node268 = (inp[1]) ? node270 : 4'b1111;
													assign node270 = (inp[2]) ? node272 : 4'b1111;
														assign node272 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node275 = (inp[2]) ? 4'b1101 : 4'b1111;
							assign node279 = (inp[13]) ? 4'b1001 : node280;
								assign node280 = (inp[2]) ? node282 : 4'b1011;
									assign node282 = (inp[9]) ? 4'b1001 : node283;
										assign node283 = (inp[15]) ? node285 : 4'b1011;
											assign node285 = (inp[11]) ? node287 : 4'b1011;
												assign node287 = (inp[8]) ? node289 : 4'b1011;
													assign node289 = (inp[7]) ? node291 : 4'b1011;
														assign node291 = (inp[1]) ? 4'b1001 : 4'b1011;
						assign node296 = (inp[4]) ? node324 : node297;
							assign node297 = (inp[2]) ? node309 : node298;
								assign node298 = (inp[13]) ? 4'b1111 : node299;
									assign node299 = (inp[9]) ? 4'b1111 : node300;
										assign node300 = (inp[7]) ? node302 : 4'b1101;
											assign node302 = (inp[8]) ? node304 : 4'b1101;
												assign node304 = (inp[15]) ? 4'b1111 : 4'b1101;
								assign node309 = (inp[13]) ? node311 : 4'b1111;
									assign node311 = (inp[8]) ? 4'b1101 : node312;
										assign node312 = (inp[7]) ? 4'b1101 : node313;
											assign node313 = (inp[9]) ? 4'b1101 : node314;
												assign node314 = (inp[15]) ? node316 : 4'b1111;
													assign node316 = (inp[11]) ? node318 : 4'b1111;
														assign node318 = (inp[1]) ? 4'b1101 : 4'b1111;
							assign node324 = (inp[13]) ? node326 : 4'b1110;
								assign node326 = (inp[2]) ? 4'b1100 : node327;
									assign node327 = (inp[9]) ? 4'b1100 : node328;
										assign node328 = (inp[7]) ? node330 : 4'b1110;
											assign node330 = (inp[8]) ? node332 : 4'b1110;
												assign node332 = (inp[1]) ? node334 : 4'b1110;
													assign node334 = (inp[11]) ? node336 : 4'b1110;
														assign node336 = (inp[15]) ? 4'b1100 : 4'b1110;
				assign node341 = (inp[6]) ? node429 : node342;
					assign node342 = (inp[14]) ? node396 : node343;
						assign node343 = (inp[4]) ? node371 : node344;
							assign node344 = (inp[13]) ? node356 : node345;
								assign node345 = (inp[2]) ? 4'b1110 : node346;
									assign node346 = (inp[15]) ? node348 : 4'b1100;
										assign node348 = (inp[9]) ? node350 : 4'b1100;
											assign node350 = (inp[8]) ? node352 : 4'b1100;
												assign node352 = (inp[7]) ? 4'b1110 : 4'b1100;
								assign node356 = (inp[2]) ? node358 : 4'b1110;
									assign node358 = (inp[9]) ? 4'b1100 : node359;
										assign node359 = (inp[8]) ? node361 : 4'b1110;
											assign node361 = (inp[7]) ? 4'b1100 : node362;
												assign node362 = (inp[15]) ? node364 : 4'b1110;
													assign node364 = (inp[11]) ? node366 : 4'b1110;
														assign node366 = (inp[1]) ? 4'b1100 : 4'b1110;
							assign node371 = (inp[13]) ? node385 : node372;
								assign node372 = (inp[2]) ? node374 : 4'b1110;
									assign node374 = (inp[8]) ? 4'b1100 : node375;
										assign node375 = (inp[9]) ? 4'b1100 : node376;
											assign node376 = (inp[7]) ? node378 : 4'b1110;
												assign node378 = (inp[11]) ? node380 : 4'b1110;
													assign node380 = (inp[1]) ? 4'b1100 : 4'b1110;
								assign node385 = (inp[2]) ? node387 : 4'b1100;
									assign node387 = (inp[9]) ? 4'b1110 : node388;
										assign node388 = (inp[8]) ? node390 : 4'b1100;
											assign node390 = (inp[15]) ? node392 : 4'b1100;
												assign node392 = (inp[7]) ? 4'b1110 : 4'b1100;
						assign node396 = (inp[13]) ? node420 : node397;
							assign node397 = (inp[4]) ? node405 : node398;
								assign node398 = (inp[8]) ? node400 : 4'b1100;
									assign node400 = (inp[2]) ? node402 : 4'b1100;
										assign node402 = (inp[9]) ? 4'b1010 : 4'b1100;
								assign node405 = (inp[2]) ? node407 : 4'b1110;
									assign node407 = (inp[9]) ? node409 : 4'b1110;
										assign node409 = (inp[7]) ? 4'b1100 : node410;
											assign node410 = (inp[8]) ? 4'b1100 : node411;
												assign node411 = (inp[0]) ? node413 : 4'b1110;
													assign node413 = (inp[1]) ? node415 : 4'b1110;
														assign node415 = (inp[11]) ? 4'b1100 : 4'b1110;
							assign node420 = (inp[4]) ? node422 : 4'b1010;
								assign node422 = (inp[8]) ? node424 : 4'b1100;
									assign node424 = (inp[2]) ? node426 : 4'b1100;
										assign node426 = (inp[9]) ? 4'b1010 : 4'b1100;
					assign node429 = (inp[13]) ? node485 : node430;
						assign node430 = (inp[4]) ? node460 : node431;
							assign node431 = (inp[2]) ? 4'b1000 : node432;
								assign node432 = (inp[14]) ? node446 : node433;
									assign node433 = (inp[8]) ? 4'b1000 : node434;
										assign node434 = (inp[9]) ? 4'b1000 : node435;
											assign node435 = (inp[7]) ? 4'b1000 : node436;
												assign node436 = (inp[1]) ? node438 : 4'b1010;
													assign node438 = (inp[15]) ? node440 : 4'b1010;
														assign node440 = (inp[11]) ? 4'b1000 : 4'b1010;
									assign node446 = (inp[9]) ? node448 : 4'b1010;
										assign node448 = (inp[8]) ? 4'b1000 : node449;
											assign node449 = (inp[11]) ? node451 : 4'b1010;
												assign node451 = (inp[1]) ? node453 : 4'b1010;
													assign node453 = (inp[7]) ? node455 : 4'b1010;
														assign node455 = (inp[15]) ? 4'b1000 : 4'b1010;
							assign node460 = (inp[8]) ? node462 : 4'b1010;
								assign node462 = (inp[2]) ? node464 : 4'b1010;
									assign node464 = (inp[9]) ? node466 : 4'b1010;
										assign node466 = (inp[7]) ? node476 : node467;
											assign node467 = (inp[15]) ? node469 : 4'b1010;
												assign node469 = (inp[1]) ? node471 : 4'b1010;
													assign node471 = (inp[3]) ? 4'b1010 : node472;
														assign node472 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node476 = (inp[14]) ? node478 : 4'b1000;
												assign node478 = (inp[11]) ? node480 : 4'b1010;
													assign node480 = (inp[15]) ? node482 : 4'b1010;
														assign node482 = (inp[1]) ? 4'b1000 : 4'b1010;
						assign node485 = (inp[4]) ? node501 : node486;
							assign node486 = (inp[2]) ? node498 : node487;
								assign node487 = (inp[14]) ? 4'b1000 : node488;
									assign node488 = (inp[9]) ? 4'b1010 : node489;
										assign node489 = (inp[7]) ? node491 : 4'b1000;
											assign node491 = (inp[15]) ? node493 : 4'b1000;
												assign node493 = (inp[8]) ? 4'b1010 : 4'b1000;
								assign node498 = (inp[14]) ? 4'b1110 : 4'b1010;
							assign node501 = (inp[2]) ? node503 : 4'b1000;
								assign node503 = (inp[15]) ? node505 : 4'b1000;
									assign node505 = (inp[9]) ? node507 : 4'b1000;
										assign node507 = (inp[8]) ? node509 : 4'b1000;
											assign node509 = (inp[14]) ? 4'b1000 : node510;
												assign node510 = (inp[7]) ? 4'b1010 : 4'b1000;
		assign node514 = (inp[5]) ? node780 : node515;
			assign node515 = (inp[4]) ? node641 : node516;
				assign node516 = (inp[6]) ? node590 : node517;
					assign node517 = (inp[14]) ? node555 : node518;
						assign node518 = (inp[13]) ? node536 : node519;
							assign node519 = (inp[2]) ? 4'b1100 : node520;
								assign node520 = (inp[12]) ? node522 : 4'b1100;
									assign node522 = (inp[9]) ? node524 : 4'b1110;
										assign node524 = (inp[7]) ? 4'b1100 : node525;
											assign node525 = (inp[8]) ? 4'b1100 : node526;
												assign node526 = (inp[3]) ? node528 : 4'b1110;
													assign node528 = (inp[15]) ? node530 : 4'b1110;
														assign node530 = (inp[11]) ? 4'b1100 : 4'b1110;
							assign node536 = (inp[2]) ? node548 : node537;
								assign node537 = (inp[9]) ? node539 : 4'b1100;
									assign node539 = (inp[12]) ? 4'b1100 : node540;
										assign node540 = (inp[7]) ? node542 : 4'b1100;
											assign node542 = (inp[15]) ? node544 : 4'b1100;
												assign node544 = (inp[8]) ? 4'b1110 : 4'b1100;
								assign node548 = (inp[12]) ? node550 : 4'b1110;
									assign node550 = (inp[9]) ? node552 : 4'b1100;
										assign node552 = (inp[8]) ? 4'b1010 : 4'b1100;
						assign node555 = (inp[12]) ? node573 : node556;
							assign node556 = (inp[13]) ? node558 : 4'b1110;
								assign node558 = (inp[2]) ? 4'b1100 : node559;
									assign node559 = (inp[9]) ? 4'b1100 : node560;
										assign node560 = (inp[8]) ? node562 : 4'b1110;
											assign node562 = (inp[7]) ? 4'b1100 : node563;
												assign node563 = (inp[15]) ? node565 : 4'b1110;
													assign node565 = (inp[1]) ? node567 : 4'b1110;
														assign node567 = (inp[11]) ? 4'b1100 : 4'b1110;
							assign node573 = (inp[13]) ? node575 : 4'b1010;
								assign node575 = (inp[2]) ? 4'b1000 : node576;
									assign node576 = (inp[9]) ? node578 : 4'b1010;
										assign node578 = (inp[8]) ? node580 : 4'b1010;
											assign node580 = (inp[7]) ? 4'b1000 : node581;
												assign node581 = (inp[0]) ? 4'b1010 : node582;
													assign node582 = (inp[15]) ? node584 : 4'b1010;
														assign node584 = (inp[1]) ? 4'b1000 : 4'b1010;
					assign node590 = (inp[14]) ? node612 : node591;
						assign node591 = (inp[13]) ? 4'b1010 : node592;
							assign node592 = (inp[12]) ? node600 : node593;
								assign node593 = (inp[8]) ? node595 : 4'b1100;
									assign node595 = (inp[9]) ? node597 : 4'b1100;
										assign node597 = (inp[2]) ? 4'b1010 : 4'b1100;
								assign node600 = (inp[2]) ? node602 : 4'b1000;
									assign node602 = (inp[7]) ? node604 : 4'b1000;
										assign node604 = (inp[15]) ? node606 : 4'b1000;
											assign node606 = (inp[8]) ? node608 : 4'b1000;
												assign node608 = (inp[9]) ? 4'b1010 : 4'b1000;
						assign node612 = (inp[13]) ? 4'b1000 : node613;
							assign node613 = (inp[2]) ? node627 : node614;
								assign node614 = (inp[7]) ? node616 : 4'b1010;
									assign node616 = (inp[9]) ? node618 : 4'b1010;
										assign node618 = (inp[12]) ? node620 : 4'b1010;
											assign node620 = (inp[3]) ? node622 : 4'b1010;
												assign node622 = (inp[8]) ? node624 : 4'b1010;
													assign node624 = (inp[0]) ? 4'b1010 : 4'b1000;
								assign node627 = (inp[7]) ? 4'b1000 : node628;
									assign node628 = (inp[12]) ? 4'b1000 : node629;
										assign node629 = (inp[8]) ? 4'b1000 : node630;
											assign node630 = (inp[9]) ? 4'b1000 : node631;
												assign node631 = (inp[15]) ? node633 : 4'b1010;
													assign node633 = (inp[11]) ? 4'b1000 : 4'b1010;
				assign node641 = (inp[12]) ? node709 : node642;
					assign node642 = (inp[6]) ? node674 : node643;
						assign node643 = (inp[14]) ? node669 : node644;
							assign node644 = (inp[9]) ? node656 : node645;
								assign node645 = (inp[13]) ? 4'b1010 : node646;
									assign node646 = (inp[2]) ? 4'b1010 : node647;
										assign node647 = (inp[8]) ? node649 : 4'b1000;
											assign node649 = (inp[7]) ? node651 : 4'b1000;
												assign node651 = (inp[15]) ? 4'b1010 : 4'b1000;
								assign node656 = (inp[2]) ? node658 : 4'b1010;
									assign node658 = (inp[13]) ? node660 : 4'b1010;
										assign node660 = (inp[8]) ? 4'b1000 : node661;
											assign node661 = (inp[7]) ? node663 : 4'b1010;
												assign node663 = (inp[11]) ? node665 : 4'b1010;
													assign node665 = (inp[1]) ? 4'b1000 : 4'b1010;
							assign node669 = (inp[2]) ? node671 : 4'b1000;
								assign node671 = (inp[13]) ? 4'b1110 : 4'b1000;
						assign node674 = (inp[2]) ? node694 : node675;
							assign node675 = (inp[13]) ? node679 : node676;
								assign node676 = (inp[14]) ? 4'b1100 : 4'b1110;
								assign node679 = (inp[14]) ? 4'b1110 : node680;
									assign node680 = (inp[9]) ? 4'b1100 : node681;
										assign node681 = (inp[8]) ? 4'b1100 : node682;
											assign node682 = (inp[7]) ? node684 : 4'b1110;
												assign node684 = (inp[15]) ? node686 : 4'b1110;
													assign node686 = (inp[11]) ? node688 : 4'b1110;
														assign node688 = (inp[1]) ? 4'b1100 : 4'b1110;
							assign node694 = (inp[13]) ? node706 : node695;
								assign node695 = (inp[9]) ? 4'b1110 : node696;
									assign node696 = (inp[14]) ? node698 : 4'b1110;
										assign node698 = (inp[15]) ? node700 : 4'b1100;
											assign node700 = (inp[7]) ? node702 : 4'b1100;
												assign node702 = (inp[8]) ? 4'b1110 : 4'b1100;
								assign node706 = (inp[14]) ? 4'b1110 : 4'b1100;
					assign node709 = (inp[6]) ? node741 : node710;
						assign node710 = (inp[14]) ? node728 : node711;
							assign node711 = (inp[13]) ? node713 : 4'b1111;
								assign node713 = (inp[2]) ? 4'b1101 : node714;
									assign node714 = (inp[11]) ? node716 : 4'b1111;
										assign node716 = (inp[1]) ? node718 : 4'b1111;
											assign node718 = (inp[9]) ? node720 : 4'b1111;
												assign node720 = (inp[7]) ? node722 : 4'b1111;
													assign node722 = (inp[8]) ? node724 : 4'b1111;
														assign node724 = (inp[15]) ? 4'b1101 : 4'b1111;
							assign node728 = (inp[13]) ? 4'b1111 : node729;
								assign node729 = (inp[7]) ? node731 : 4'b1101;
									assign node731 = (inp[15]) ? node733 : 4'b1101;
										assign node733 = (inp[9]) ? node735 : 4'b1101;
											assign node735 = (inp[2]) ? node737 : 4'b1101;
												assign node737 = (inp[8]) ? 4'b1111 : 4'b1101;
						assign node741 = (inp[14]) ? node763 : node742;
							assign node742 = (inp[2]) ? node756 : node743;
								assign node743 = (inp[13]) ? 4'b1101 : node744;
									assign node744 = (inp[8]) ? node746 : 4'b1111;
										assign node746 = (inp[9]) ? node748 : 4'b1111;
											assign node748 = (inp[7]) ? 4'b1101 : node749;
												assign node749 = (inp[1]) ? node751 : 4'b1111;
													assign node751 = (inp[15]) ? 4'b1101 : 4'b1111;
								assign node756 = (inp[8]) ? node758 : 4'b1101;
									assign node758 = (inp[13]) ? node760 : 4'b1101;
										assign node760 = (inp[9]) ? 4'b1011 : 4'b1101;
							assign node763 = (inp[13]) ? node765 : 4'b1011;
								assign node765 = (inp[2]) ? 4'b1001 : node766;
									assign node766 = (inp[9]) ? node768 : 4'b1011;
										assign node768 = (inp[8]) ? 4'b1001 : node769;
											assign node769 = (inp[7]) ? 4'b1001 : node770;
												assign node770 = (inp[11]) ? node772 : 4'b1011;
													assign node772 = (inp[1]) ? node774 : 4'b1011;
														assign node774 = (inp[15]) ? 4'b1001 : 4'b1011;
			assign node780 = (inp[12]) ? node984 : node781;
				assign node781 = (inp[6]) ? node883 : node782;
					assign node782 = (inp[13]) ? node842 : node783;
						assign node783 = (inp[4]) ? node807 : node784;
							assign node784 = (inp[2]) ? node786 : 4'b0111;
								assign node786 = (inp[8]) ? node788 : 4'b0111;
									assign node788 = (inp[9]) ? node790 : 4'b0111;
										assign node790 = (inp[14]) ? node800 : node791;
											assign node791 = (inp[1]) ? node793 : 4'b0111;
												assign node793 = (inp[15]) ? node795 : 4'b0111;
													assign node795 = (inp[11]) ? node797 : 4'b0111;
														assign node797 = (inp[7]) ? 4'b0101 : 4'b0111;
											assign node800 = (inp[7]) ? 4'b0101 : node801;
												assign node801 = (inp[1]) ? node803 : 4'b0111;
													assign node803 = (inp[15]) ? 4'b0101 : 4'b0111;
							assign node807 = (inp[2]) ? node835 : node808;
								assign node808 = (inp[14]) ? node822 : node809;
									assign node809 = (inp[9]) ? node811 : 4'b0111;
										assign node811 = (inp[8]) ? 4'b0101 : node812;
											assign node812 = (inp[11]) ? node814 : 4'b0111;
												assign node814 = (inp[15]) ? node816 : 4'b0111;
													assign node816 = (inp[1]) ? node818 : 4'b0111;
														assign node818 = (inp[7]) ? 4'b0101 : 4'b0111;
									assign node822 = (inp[7]) ? 4'b0101 : node823;
										assign node823 = (inp[8]) ? 4'b0101 : node824;
											assign node824 = (inp[9]) ? 4'b0101 : node825;
												assign node825 = (inp[15]) ? node827 : 4'b0111;
													assign node827 = (inp[1]) ? node829 : 4'b0111;
														assign node829 = (inp[11]) ? 4'b0101 : 4'b0111;
								assign node835 = (inp[8]) ? node837 : 4'b0101;
									assign node837 = (inp[9]) ? node839 : 4'b0101;
										assign node839 = (inp[14]) ? 4'b0011 : 4'b0101;
						assign node842 = (inp[4]) ? node856 : node843;
							assign node843 = (inp[8]) ? node845 : 4'b0101;
								assign node845 = (inp[9]) ? node847 : 4'b0101;
									assign node847 = (inp[2]) ? node849 : 4'b0101;
										assign node849 = (inp[14]) ? 4'b0011 : node850;
											assign node850 = (inp[15]) ? node852 : 4'b0101;
												assign node852 = (inp[7]) ? 4'b0111 : 4'b0101;
							assign node856 = (inp[14]) ? node868 : node857;
								assign node857 = (inp[2]) ? 4'b0111 : node858;
									assign node858 = (inp[9]) ? 4'b0111 : node859;
										assign node859 = (inp[8]) ? node861 : 4'b0101;
											assign node861 = (inp[7]) ? node863 : 4'b0101;
												assign node863 = (inp[15]) ? 4'b0111 : 4'b0101;
								assign node868 = (inp[2]) ? node870 : 4'b0011;
									assign node870 = (inp[9]) ? 4'b0001 : node871;
										assign node871 = (inp[8]) ? node873 : 4'b0011;
											assign node873 = (inp[7]) ? 4'b0001 : node874;
												assign node874 = (inp[15]) ? node876 : 4'b0011;
													assign node876 = (inp[1]) ? node878 : 4'b0011;
														assign node878 = (inp[11]) ? 4'b0001 : 4'b0011;
					assign node883 = (inp[14]) ? node939 : node884;
						assign node884 = (inp[13]) ? node912 : node885;
							assign node885 = (inp[2]) ? node897 : node886;
								assign node886 = (inp[4]) ? node888 : 4'b0011;
									assign node888 = (inp[9]) ? node890 : 4'b0001;
										assign node890 = (inp[7]) ? node892 : 4'b0001;
											assign node892 = (inp[8]) ? node894 : 4'b0001;
												assign node894 = (inp[15]) ? 4'b0011 : 4'b0001;
								assign node897 = (inp[4]) ? 4'b0011 : node898;
									assign node898 = (inp[9]) ? node900 : 4'b0011;
										assign node900 = (inp[8]) ? 4'b0001 : node901;
											assign node901 = (inp[7]) ? 4'b0001 : node902;
												assign node902 = (inp[1]) ? node904 : 4'b0011;
													assign node904 = (inp[15]) ? node906 : 4'b0011;
														assign node906 = (inp[11]) ? 4'b0001 : 4'b0011;
							assign node912 = (inp[2]) ? node928 : node913;
								assign node913 = (inp[4]) ? node915 : 4'b0001;
									assign node915 = (inp[9]) ? 4'b0001 : node916;
										assign node916 = (inp[1]) ? node918 : 4'b0011;
											assign node918 = (inp[7]) ? node920 : 4'b0011;
												assign node920 = (inp[11]) ? node922 : 4'b0011;
													assign node922 = (inp[15]) ? node924 : 4'b0011;
														assign node924 = (inp[8]) ? 4'b0001 : 4'b0011;
								assign node928 = (inp[4]) ? 4'b0001 : node929;
									assign node929 = (inp[9]) ? 4'b0011 : node930;
										assign node930 = (inp[15]) ? node932 : 4'b0001;
											assign node932 = (inp[8]) ? node934 : 4'b0001;
												assign node934 = (inp[7]) ? 4'b0011 : 4'b0001;
						assign node939 = (inp[4]) ? node959 : node940;
							assign node940 = (inp[13]) ? node956 : node941;
								assign node941 = (inp[2]) ? node943 : 4'b0011;
									assign node943 = (inp[9]) ? 4'b0001 : node944;
										assign node944 = (inp[8]) ? 4'b0001 : node945;
											assign node945 = (inp[7]) ? node947 : 4'b0011;
												assign node947 = (inp[1]) ? node949 : 4'b0011;
													assign node949 = (inp[15]) ? node951 : 4'b0011;
														assign node951 = (inp[11]) ? 4'b0001 : 4'b0011;
								assign node956 = (inp[2]) ? 4'b0111 : 4'b0001;
							assign node959 = (inp[13]) ? node973 : node960;
								assign node960 = (inp[2]) ? node962 : 4'b0110;
									assign node962 = (inp[9]) ? 4'b0100 : node963;
										assign node963 = (inp[11]) ? node965 : 4'b0110;
											assign node965 = (inp[15]) ? node967 : 4'b0110;
												assign node967 = (inp[7]) ? node969 : 4'b0110;
													assign node969 = (inp[8]) ? 4'b0100 : 4'b0110;
								assign node973 = (inp[2]) ? 4'b0110 : node974;
									assign node974 = (inp[9]) ? node976 : 4'b0100;
										assign node976 = (inp[8]) ? node978 : 4'b0100;
											assign node978 = (inp[15]) ? node980 : 4'b0100;
												assign node980 = (inp[7]) ? 4'b0110 : 4'b0100;
				assign node984 = (inp[4]) ? node1126 : node985;
					assign node985 = (inp[14]) ? node1071 : node986;
						assign node986 = (inp[6]) ? node1024 : node987;
							assign node987 = (inp[13]) ? node1009 : node988;
								assign node988 = (inp[8]) ? node994 : node989;
									assign node989 = (inp[2]) ? 4'b0100 : node990;
										assign node990 = (inp[9]) ? 4'b0100 : 4'b0110;
									assign node994 = (inp[2]) ? node1006 : node995;
										assign node995 = (inp[9]) ? 4'b0100 : node996;
											assign node996 = (inp[7]) ? 4'b0100 : node997;
												assign node997 = (inp[11]) ? node999 : 4'b0110;
													assign node999 = (inp[15]) ? node1001 : 4'b0110;
														assign node1001 = (inp[1]) ? 4'b0100 : 4'b0110;
										assign node1006 = (inp[9]) ? 4'b0010 : 4'b0100;
								assign node1009 = (inp[2]) ? node1011 : 4'b0010;
									assign node1011 = (inp[7]) ? 4'b0000 : node1012;
										assign node1012 = (inp[9]) ? 4'b0000 : node1013;
											assign node1013 = (inp[8]) ? 4'b0000 : node1014;
												assign node1014 = (inp[15]) ? node1016 : 4'b0010;
													assign node1016 = (inp[11]) ? node1018 : 4'b0010;
														assign node1018 = (inp[1]) ? 4'b0000 : 4'b0010;
							assign node1024 = (inp[8]) ? node1054 : node1025;
								assign node1025 = (inp[2]) ? node1049 : node1026;
									assign node1026 = (inp[9]) ? node1038 : node1027;
										assign node1027 = (inp[11]) ? node1029 : 4'b0110;
											assign node1029 = (inp[3]) ? node1031 : 4'b0110;
												assign node1031 = (inp[0]) ? node1033 : 4'b0110;
													assign node1033 = (inp[15]) ? node1035 : 4'b0110;
														assign node1035 = (inp[13]) ? 4'b0110 : 4'b0100;
										assign node1038 = (inp[13]) ? node1040 : 4'b0100;
											assign node1040 = (inp[7]) ? 4'b0100 : node1041;
												assign node1041 = (inp[1]) ? node1043 : 4'b0110;
													assign node1043 = (inp[11]) ? node1045 : 4'b0110;
														assign node1045 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node1049 = (inp[9]) ? node1051 : 4'b0100;
										assign node1051 = (inp[13]) ? 4'b0100 : 4'b0110;
								assign node1054 = (inp[2]) ? node1060 : node1055;
									assign node1055 = (inp[9]) ? 4'b0100 : node1056;
										assign node1056 = (inp[13]) ? 4'b0110 : 4'b0100;
									assign node1060 = (inp[9]) ? node1068 : node1061;
										assign node1061 = (inp[13]) ? 4'b0100 : node1062;
											assign node1062 = (inp[7]) ? node1064 : 4'b0100;
												assign node1064 = (inp[15]) ? 4'b0110 : 4'b0100;
										assign node1068 = (inp[13]) ? 4'b0010 : 4'b0110;
						assign node1071 = (inp[2]) ? node1107 : node1072;
							assign node1072 = (inp[6]) ? node1084 : node1073;
								assign node1073 = (inp[13]) ? 4'b0000 : node1074;
									assign node1074 = (inp[9]) ? 4'b0010 : node1075;
										assign node1075 = (inp[8]) ? node1077 : 4'b0000;
											assign node1077 = (inp[15]) ? node1079 : 4'b0000;
												assign node1079 = (inp[7]) ? 4'b0010 : 4'b0000;
								assign node1084 = (inp[9]) ? node1086 : 4'b0010;
									assign node1086 = (inp[8]) ? node1088 : 4'b0010;
										assign node1088 = (inp[13]) ? node1098 : node1089;
											assign node1089 = (inp[7]) ? 4'b0000 : node1090;
												assign node1090 = (inp[15]) ? node1092 : 4'b0010;
													assign node1092 = (inp[1]) ? node1094 : 4'b0010;
														assign node1094 = (inp[11]) ? 4'b0000 : 4'b0010;
											assign node1098 = (inp[15]) ? node1100 : 4'b0010;
												assign node1100 = (inp[7]) ? node1102 : 4'b0010;
													assign node1102 = (inp[1]) ? node1104 : 4'b0010;
														assign node1104 = (inp[11]) ? 4'b0000 : 4'b0010;
							assign node1107 = (inp[6]) ? node1115 : node1108;
								assign node1108 = (inp[13]) ? 4'b0110 : node1109;
									assign node1109 = (inp[9]) ? node1111 : 4'b0010;
										assign node1111 = (inp[8]) ? 4'b0000 : 4'b0010;
								assign node1115 = (inp[8]) ? node1117 : 4'b0000;
									assign node1117 = (inp[15]) ? node1119 : 4'b0000;
										assign node1119 = (inp[9]) ? node1121 : 4'b0000;
											assign node1121 = (inp[7]) ? node1123 : 4'b0000;
												assign node1123 = (inp[13]) ? 4'b0000 : 4'b0010;
					assign node1126 = (inp[14]) ? node1224 : node1127;
						assign node1127 = (inp[6]) ? node1163 : node1128;
							assign node1128 = (inp[2]) ? node1152 : node1129;
								assign node1129 = (inp[9]) ? node1131 : 4'b0111;
									assign node1131 = (inp[8]) ? node1133 : 4'b0111;
										assign node1133 = (inp[7]) ? node1143 : node1134;
											assign node1134 = (inp[15]) ? node1136 : 4'b0111;
												assign node1136 = (inp[1]) ? node1138 : 4'b0111;
													assign node1138 = (inp[11]) ? node1140 : 4'b0111;
														assign node1140 = (inp[13]) ? 4'b0101 : 4'b0111;
											assign node1143 = (inp[13]) ? 4'b0101 : node1144;
												assign node1144 = (inp[11]) ? node1146 : 4'b0111;
													assign node1146 = (inp[15]) ? node1148 : 4'b0111;
														assign node1148 = (inp[1]) ? 4'b0101 : 4'b0111;
								assign node1152 = (inp[8]) ? node1154 : 4'b0101;
									assign node1154 = (inp[9]) ? node1156 : 4'b0101;
										assign node1156 = (inp[13]) ? 4'b0011 : node1157;
											assign node1157 = (inp[15]) ? node1159 : 4'b0101;
												assign node1159 = (inp[7]) ? 4'b0111 : 4'b0101;
							assign node1163 = (inp[13]) ? node1191 : node1164;
								assign node1164 = (inp[9]) ? node1184 : node1165;
									assign node1165 = (inp[8]) ? node1177 : node1166;
										assign node1166 = (inp[2]) ? node1168 : 4'b0101;
											assign node1168 = (inp[7]) ? 4'b0101 : node1169;
												assign node1169 = (inp[11]) ? node1171 : 4'b0111;
													assign node1171 = (inp[1]) ? node1173 : 4'b0111;
														assign node1173 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node1177 = (inp[15]) ? node1179 : 4'b0101;
											assign node1179 = (inp[2]) ? 4'b0101 : node1180;
												assign node1180 = (inp[7]) ? 4'b0111 : 4'b0101;
									assign node1184 = (inp[8]) ? node1188 : node1185;
										assign node1185 = (inp[2]) ? 4'b0101 : 4'b0111;
										assign node1188 = (inp[2]) ? 4'b0011 : 4'b0111;
								assign node1191 = (inp[9]) ? node1215 : node1192;
									assign node1192 = (inp[8]) ? node1194 : 4'b0011;
										assign node1194 = (inp[7]) ? node1206 : node1195;
											assign node1195 = (inp[0]) ? node1197 : 4'b0011;
												assign node1197 = (inp[15]) ? node1199 : 4'b0011;
													assign node1199 = (inp[11]) ? node1201 : 4'b0011;
														assign node1201 = (inp[1]) ? node1203 : 4'b0011;
															assign node1203 = (inp[2]) ? 4'b0011 : 4'b0001;
											assign node1206 = (inp[2]) ? node1208 : 4'b0001;
												assign node1208 = (inp[1]) ? node1210 : 4'b0011;
													assign node1210 = (inp[11]) ? node1212 : 4'b0011;
														assign node1212 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node1215 = (inp[8]) ? node1217 : 4'b0001;
										assign node1217 = (inp[7]) ? node1219 : 4'b0001;
											assign node1219 = (inp[15]) ? node1221 : 4'b0001;
												assign node1221 = (inp[2]) ? 4'b0001 : 4'b0011;
						assign node1224 = (inp[6]) ? node1274 : node1225;
							assign node1225 = (inp[2]) ? node1253 : node1226;
								assign node1226 = (inp[9]) ? node1240 : node1227;
									assign node1227 = (inp[13]) ? node1229 : 4'b0011;
										assign node1229 = (inp[8]) ? 4'b0001 : node1230;
											assign node1230 = (inp[1]) ? node1232 : 4'b0011;
												assign node1232 = (inp[15]) ? node1234 : 4'b0011;
													assign node1234 = (inp[7]) ? node1236 : 4'b0011;
														assign node1236 = (inp[0]) ? 4'b0011 : 4'b0001;
									assign node1240 = (inp[13]) ? 4'b0001 : node1241;
										assign node1241 = (inp[7]) ? 4'b0001 : node1242;
											assign node1242 = (inp[8]) ? 4'b0001 : node1243;
												assign node1243 = (inp[1]) ? node1245 : 4'b0011;
													assign node1245 = (inp[15]) ? node1247 : 4'b0011;
														assign node1247 = (inp[11]) ? 4'b0001 : 4'b0011;
								assign node1253 = (inp[13]) ? node1263 : node1254;
									assign node1254 = (inp[9]) ? 4'b0011 : node1255;
										assign node1255 = (inp[8]) ? node1257 : 4'b0001;
											assign node1257 = (inp[15]) ? node1259 : 4'b0001;
												assign node1259 = (inp[7]) ? 4'b0011 : 4'b0001;
									assign node1263 = (inp[9]) ? node1265 : 4'b0111;
										assign node1265 = (inp[8]) ? 4'b0101 : node1266;
											assign node1266 = (inp[11]) ? node1268 : 4'b0111;
												assign node1268 = (inp[1]) ? node1270 : 4'b0111;
													assign node1270 = (inp[15]) ? 4'b0101 : 4'b0111;
							assign node1274 = (inp[13]) ? node1306 : node1275;
								assign node1275 = (inp[9]) ? node1297 : node1276;
									assign node1276 = (inp[8]) ? node1278 : 4'b0110;
										assign node1278 = (inp[7]) ? node1288 : node1279;
											assign node1279 = (inp[2]) ? node1281 : 4'b0110;
												assign node1281 = (inp[11]) ? node1283 : 4'b0110;
													assign node1283 = (inp[1]) ? node1285 : 4'b0110;
														assign node1285 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node1288 = (inp[2]) ? 4'b0100 : node1289;
												assign node1289 = (inp[1]) ? node1291 : 4'b0110;
													assign node1291 = (inp[15]) ? node1293 : 4'b0110;
														assign node1293 = (inp[11]) ? 4'b0100 : 4'b0110;
									assign node1297 = (inp[8]) ? node1299 : 4'b0100;
										assign node1299 = (inp[2]) ? 4'b0010 : node1300;
											assign node1300 = (inp[15]) ? node1302 : 4'b0100;
												assign node1302 = (inp[7]) ? 4'b0110 : 4'b0100;
								assign node1306 = (inp[2]) ? node1338 : node1307;
									assign node1307 = (inp[8]) ? node1331 : node1308;
										assign node1308 = (inp[7]) ? node1320 : node1309;
											assign node1309 = (inp[0]) ? node1311 : 4'b0010;
												assign node1311 = (inp[15]) ? node1313 : 4'b0010;
													assign node1313 = (inp[11]) ? node1315 : 4'b0010;
														assign node1315 = (inp[9]) ? 4'b0010 : node1316;
															assign node1316 = (inp[1]) ? 4'b0000 : 4'b0010;
											assign node1320 = (inp[9]) ? node1322 : 4'b0000;
												assign node1322 = (inp[11]) ? node1324 : 4'b0010;
													assign node1324 = (inp[0]) ? node1326 : 4'b0010;
														assign node1326 = (inp[15]) ? node1328 : 4'b0010;
															assign node1328 = (inp[1]) ? 4'b0000 : 4'b0010;
										assign node1331 = (inp[9]) ? 4'b0000 : node1332;
											assign node1332 = (inp[15]) ? node1334 : 4'b0000;
												assign node1334 = (inp[7]) ? 4'b0010 : 4'b0000;
									assign node1338 = (inp[8]) ? node1356 : node1339;
										assign node1339 = (inp[9]) ? node1349 : node1340;
											assign node1340 = (inp[3]) ? node1342 : 4'b0110;
												assign node1342 = (inp[11]) ? node1344 : 4'b0110;
													assign node1344 = (inp[0]) ? node1346 : 4'b0110;
														assign node1346 = (inp[1]) ? 4'b0100 : 4'b0110;
											assign node1349 = (inp[7]) ? 4'b0100 : node1350;
												assign node1350 = (inp[1]) ? node1352 : 4'b0110;
													assign node1352 = (inp[11]) ? 4'b0100 : 4'b0110;
										assign node1356 = (inp[9]) ? node1362 : node1357;
											assign node1357 = (inp[7]) ? node1359 : 4'b0100;
												assign node1359 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node1362 = (inp[7]) ? node1370 : node1363;
												assign node1363 = (inp[3]) ? 4'b0010 : node1364;
													assign node1364 = (inp[15]) ? node1366 : 4'b0010;
														assign node1366 = (inp[11]) ? 4'b0000 : 4'b0010;
												assign node1370 = (inp[15]) ? node1372 : 4'b0000;
													assign node1372 = (inp[11]) ? 4'b0000 : 4'b0010;

endmodule