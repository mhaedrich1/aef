module dtc_split25_bm87 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node60;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node113;
	wire [3-1:0] node115;
	wire [3-1:0] node117;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node156;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node196;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node218;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node222;
	wire [3-1:0] node224;
	wire [3-1:0] node226;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node236;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node271;
	wire [3-1:0] node273;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node307;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node317;
	wire [3-1:0] node318;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node335;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node346;
	wire [3-1:0] node348;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node355;
	wire [3-1:0] node357;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node363;
	wire [3-1:0] node364;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node377;
	wire [3-1:0] node379;
	wire [3-1:0] node382;
	wire [3-1:0] node383;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node396;
	wire [3-1:0] node397;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node408;
	wire [3-1:0] node409;
	wire [3-1:0] node410;
	wire [3-1:0] node415;
	wire [3-1:0] node416;
	wire [3-1:0] node417;
	wire [3-1:0] node419;
	wire [3-1:0] node421;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node431;
	wire [3-1:0] node433;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node440;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node455;
	wire [3-1:0] node456;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node463;
	wire [3-1:0] node464;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node470;
	wire [3-1:0] node471;
	wire [3-1:0] node474;
	wire [3-1:0] node477;
	wire [3-1:0] node479;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node489;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node492;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node508;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node513;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node519;
	wire [3-1:0] node522;
	wire [3-1:0] node525;
	wire [3-1:0] node527;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node534;
	wire [3-1:0] node535;
	wire [3-1:0] node537;
	wire [3-1:0] node538;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node550;
	wire [3-1:0] node551;
	wire [3-1:0] node556;
	wire [3-1:0] node557;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node569;
	wire [3-1:0] node572;
	wire [3-1:0] node574;
	wire [3-1:0] node575;
	wire [3-1:0] node576;
	wire [3-1:0] node577;
	wire [3-1:0] node579;
	wire [3-1:0] node582;

	assign outp = (inp[6]) ? node122 : node1;
		assign node1 = (inp[7]) ? node19 : node2;
			assign node2 = (inp[10]) ? 3'b000 : node3;
				assign node3 = (inp[8]) ? node5 : 3'b000;
					assign node5 = (inp[0]) ? node7 : 3'b000;
						assign node7 = (inp[1]) ? 3'b000 : node8;
							assign node8 = (inp[9]) ? 3'b000 : node9;
								assign node9 = (inp[11]) ? node13 : node10;
									assign node10 = (inp[2]) ? 3'b000 : 3'b100;
									assign node13 = (inp[2]) ? 3'b100 : 3'b000;
			assign node19 = (inp[9]) ? node97 : node20;
				assign node20 = (inp[0]) ? node64 : node21;
					assign node21 = (inp[1]) ? node27 : node22;
						assign node22 = (inp[10]) ? 3'b110 : node23;
							assign node23 = (inp[11]) ? 3'b001 : 3'b101;
						assign node27 = (inp[10]) ? node53 : node28;
							assign node28 = (inp[8]) ? node44 : node29;
								assign node29 = (inp[5]) ? node35 : node30;
									assign node30 = (inp[11]) ? 3'b010 : node31;
										assign node31 = (inp[3]) ? 3'b110 : 3'b010;
									assign node35 = (inp[4]) ? 3'b110 : node36;
										assign node36 = (inp[3]) ? node40 : node37;
											assign node37 = (inp[11]) ? 3'b010 : 3'b110;
											assign node40 = (inp[11]) ? 3'b110 : 3'b010;
								assign node44 = (inp[11]) ? node48 : node45;
									assign node45 = (inp[4]) ? 3'b001 : 3'b101;
									assign node48 = (inp[4]) ? 3'b110 : node49;
										assign node49 = (inp[2]) ? 3'b010 : 3'b110;
							assign node53 = (inp[8]) ? node57 : node54;
								assign node54 = (inp[11]) ? 3'b000 : 3'b100;
								assign node57 = (inp[11]) ? 3'b000 : node58;
									assign node58 = (inp[2]) ? node60 : 3'b010;
										assign node60 = (inp[3]) ? 3'b100 : 3'b010;
					assign node64 = (inp[10]) ? node88 : node65;
						assign node65 = (inp[1]) ? node81 : node66;
							assign node66 = (inp[2]) ? node74 : node67;
								assign node67 = (inp[11]) ? node71 : node68;
									assign node68 = (inp[8]) ? 3'b110 : 3'b010;
									assign node71 = (inp[8]) ? 3'b010 : 3'b100;
								assign node74 = (inp[8]) ? node76 : 3'b100;
									assign node76 = (inp[11]) ? 3'b100 : node77;
										assign node77 = (inp[4]) ? 3'b010 : 3'b110;
							assign node81 = (inp[4]) ? 3'b000 : node82;
								assign node82 = (inp[8]) ? 3'b100 : node83;
									assign node83 = (inp[2]) ? 3'b000 : 3'b100;
						assign node88 = (inp[2]) ? 3'b000 : node89;
							assign node89 = (inp[1]) ? 3'b000 : node90;
								assign node90 = (inp[8]) ? node92 : 3'b000;
									assign node92 = (inp[11]) ? 3'b000 : 3'b100;
				assign node97 = (inp[0]) ? 3'b000 : node98;
					assign node98 = (inp[10]) ? 3'b000 : node99;
						assign node99 = (inp[2]) ? node109 : node100;
							assign node100 = (inp[1]) ? node104 : node101;
								assign node101 = (inp[11]) ? 3'b110 : 3'b010;
								assign node104 = (inp[4]) ? 3'b100 : node105;
									assign node105 = (inp[3]) ? 3'b000 : 3'b100;
							assign node109 = (inp[1]) ? node113 : node110;
								assign node110 = (inp[11]) ? 3'b000 : 3'b100;
								assign node113 = (inp[11]) ? node115 : 3'b000;
									assign node115 = (inp[8]) ? node117 : 3'b000;
										assign node117 = (inp[4]) ? 3'b000 : 3'b100;
		assign node122 = (inp[9]) ? node394 : node123;
			assign node123 = (inp[0]) ? node241 : node124;
				assign node124 = (inp[7]) ? node206 : node125;
					assign node125 = (inp[10]) ? node159 : node126;
						assign node126 = (inp[8]) ? node140 : node127;
							assign node127 = (inp[2]) ? node131 : node128;
								assign node128 = (inp[11]) ? 3'b001 : 3'b101;
								assign node131 = (inp[11]) ? 3'b101 : node132;
									assign node132 = (inp[1]) ? node134 : 3'b011;
										assign node134 = (inp[4]) ? 3'b101 : node135;
											assign node135 = (inp[5]) ? 3'b001 : 3'b101;
							assign node140 = (inp[1]) ? node146 : node141;
								assign node141 = (inp[11]) ? 3'b011 : node142;
									assign node142 = (inp[2]) ? 3'b111 : 3'b011;
								assign node146 = (inp[4]) ? node156 : node147;
									assign node147 = (inp[5]) ? 3'b101 : node148;
										assign node148 = (inp[3]) ? 3'b101 : node149;
											assign node149 = (inp[2]) ? 3'b011 : node150;
												assign node150 = (inp[11]) ? 3'b011 : 3'b101;
									assign node156 = (inp[5]) ? 3'b001 : 3'b011;
						assign node159 = (inp[1]) ? node185 : node160;
							assign node160 = (inp[11]) ? node170 : node161;
								assign node161 = (inp[2]) ? 3'b101 : node162;
									assign node162 = (inp[8]) ? 3'b011 : node163;
										assign node163 = (inp[5]) ? node165 : 3'b101;
											assign node165 = (inp[4]) ? 3'b101 : 3'b001;
								assign node170 = (inp[5]) ? node178 : node171;
									assign node171 = (inp[4]) ? node173 : 3'b001;
										assign node173 = (inp[2]) ? 3'b101 : node174;
											assign node174 = (inp[8]) ? 3'b101 : 3'b001;
									assign node178 = (inp[4]) ? node180 : 3'b010;
										assign node180 = (inp[3]) ? node182 : 3'b001;
											assign node182 = (inp[8]) ? 3'b001 : 3'b110;
							assign node185 = (inp[8]) ? node193 : node186;
								assign node186 = (inp[11]) ? node188 : 3'b110;
									assign node188 = (inp[5]) ? node190 : 3'b010;
										assign node190 = (inp[2]) ? 3'b010 : 3'b110;
								assign node193 = (inp[11]) ? node201 : node194;
									assign node194 = (inp[3]) ? node196 : 3'b001;
										assign node196 = (inp[4]) ? node198 : 3'b001;
											assign node198 = (inp[5]) ? 3'b110 : 3'b101;
									assign node201 = (inp[2]) ? 3'b001 : node202;
										assign node202 = (inp[3]) ? 3'b110 : 3'b010;
					assign node206 = (inp[10]) ? node218 : node207;
						assign node207 = (inp[1]) ? node209 : 3'b111;
							assign node209 = (inp[4]) ? node211 : 3'b111;
								assign node211 = (inp[8]) ? 3'b111 : node212;
									assign node212 = (inp[11]) ? 3'b011 : node213;
										assign node213 = (inp[5]) ? 3'b011 : 3'b111;
						assign node218 = (inp[1]) ? node230 : node219;
							assign node219 = (inp[8]) ? 3'b111 : node220;
								assign node220 = (inp[3]) ? node222 : 3'b011;
									assign node222 = (inp[5]) ? node224 : 3'b011;
										assign node224 = (inp[11]) ? node226 : 3'b111;
											assign node226 = (inp[4]) ? 3'b101 : 3'b001;
							assign node230 = (inp[5]) ? node236 : node231;
								assign node231 = (inp[11]) ? 3'b001 : node232;
									assign node232 = (inp[8]) ? 3'b011 : 3'b101;
								assign node236 = (inp[3]) ? node238 : 3'b101;
									assign node238 = (inp[8]) ? 3'b101 : 3'b001;
				assign node241 = (inp[7]) ? node307 : node242;
					assign node242 = (inp[10]) ? node278 : node243;
						assign node243 = (inp[1]) ? node269 : node244;
							assign node244 = (inp[8]) ? node254 : node245;
								assign node245 = (inp[2]) ? node249 : node246;
									assign node246 = (inp[11]) ? 3'b110 : 3'b001;
									assign node249 = (inp[5]) ? node251 : 3'b110;
										assign node251 = (inp[11]) ? 3'b010 : 3'b110;
								assign node254 = (inp[5]) ? node264 : node255;
									assign node255 = (inp[2]) ? node257 : 3'b101;
										assign node257 = (inp[11]) ? 3'b101 : node258;
											assign node258 = (inp[4]) ? 3'b001 : node259;
												assign node259 = (inp[3]) ? 3'b001 : 3'b101;
									assign node264 = (inp[3]) ? node266 : 3'b001;
										assign node266 = (inp[2]) ? 3'b110 : 3'b001;
							assign node269 = (inp[8]) ? 3'b110 : node270;
								assign node270 = (inp[3]) ? 3'b010 : node271;
									assign node271 = (inp[5]) ? node273 : 3'b010;
										assign node273 = (inp[2]) ? 3'b100 : 3'b010;
						assign node278 = (inp[4]) ? node286 : node279;
							assign node279 = (inp[1]) ? 3'b100 : node280;
								assign node280 = (inp[8]) ? 3'b100 : node281;
									assign node281 = (inp[11]) ? 3'b000 : 3'b010;
							assign node286 = (inp[1]) ? node300 : node287;
								assign node287 = (inp[5]) ? node291 : node288;
									assign node288 = (inp[8]) ? 3'b110 : 3'b100;
									assign node291 = (inp[3]) ? 3'b010 : node292;
										assign node292 = (inp[2]) ? 3'b100 : node293;
											assign node293 = (inp[11]) ? node295 : 3'b010;
												assign node295 = (inp[8]) ? 3'b010 : 3'b100;
								assign node300 = (inp[8]) ? node302 : 3'b000;
									assign node302 = (inp[3]) ? 3'b100 : node303;
										assign node303 = (inp[5]) ? 3'b010 : 3'b000;
					assign node307 = (inp[10]) ? node351 : node308;
						assign node308 = (inp[1]) ? node328 : node309;
							assign node309 = (inp[8]) ? node323 : node310;
								assign node310 = (inp[2]) ? 3'b001 : node311;
									assign node311 = (inp[11]) ? node317 : node312;
										assign node312 = (inp[4]) ? 3'b011 : node313;
											assign node313 = (inp[5]) ? 3'b001 : 3'b101;
										assign node317 = (inp[3]) ? 3'b101 : node318;
											assign node318 = (inp[4]) ? 3'b101 : 3'b111;
								assign node323 = (inp[2]) ? 3'b011 : node324;
									assign node324 = (inp[11]) ? 3'b011 : 3'b111;
							assign node328 = (inp[4]) ? node338 : node329;
								assign node329 = (inp[11]) ? node335 : node330;
									assign node330 = (inp[2]) ? 3'b101 : node331;
										assign node331 = (inp[8]) ? 3'b011 : 3'b101;
									assign node335 = (inp[8]) ? 3'b101 : 3'b111;
								assign node338 = (inp[5]) ? node346 : node339;
									assign node339 = (inp[11]) ? 3'b001 : node340;
										assign node340 = (inp[2]) ? node342 : 3'b101;
											assign node342 = (inp[8]) ? 3'b101 : 3'b001;
									assign node346 = (inp[8]) ? node348 : 3'b111;
										assign node348 = (inp[11]) ? 3'b001 : 3'b101;
						assign node351 = (inp[4]) ? node375 : node352;
							assign node352 = (inp[1]) ? node360 : node353;
								assign node353 = (inp[5]) ? node355 : 3'b001;
									assign node355 = (inp[11]) ? node357 : 3'b101;
										assign node357 = (inp[8]) ? 3'b010 : 3'b101;
								assign node360 = (inp[8]) ? node368 : node361;
									assign node361 = (inp[3]) ? node363 : 3'b010;
										assign node363 = (inp[11]) ? 3'b100 : node364;
											assign node364 = (inp[2]) ? 3'b010 : 3'b110;
									assign node368 = (inp[2]) ? node372 : node369;
										assign node369 = (inp[5]) ? 3'b000 : 3'b001;
										assign node372 = (inp[11]) ? 3'b010 : 3'b111;
							assign node375 = (inp[8]) ? node387 : node376;
								assign node376 = (inp[1]) ? node382 : node377;
									assign node377 = (inp[11]) ? node379 : 3'b110;
										assign node379 = (inp[3]) ? 3'b110 : 3'b010;
									assign node382 = (inp[5]) ? 3'b010 : node383;
										assign node383 = (inp[3]) ? 3'b010 : 3'b110;
								assign node387 = (inp[11]) ? node391 : node388;
									assign node388 = (inp[1]) ? 3'b111 : 3'b101;
									assign node391 = (inp[3]) ? 3'b010 : 3'b110;
			assign node394 = (inp[0]) ? node530 : node395;
				assign node395 = (inp[7]) ? node453 : node396;
					assign node396 = (inp[10]) ? node438 : node397;
						assign node397 = (inp[11]) ? node415 : node398;
							assign node398 = (inp[3]) ? node408 : node399;
								assign node399 = (inp[5]) ? node403 : node400;
									assign node400 = (inp[2]) ? 3'b100 : 3'b110;
									assign node403 = (inp[2]) ? 3'b010 : node404;
										assign node404 = (inp[1]) ? 3'b110 : 3'b010;
								assign node408 = (inp[5]) ? 3'b010 : node409;
									assign node409 = (inp[2]) ? 3'b010 : node410;
										assign node410 = (inp[8]) ? 3'b001 : 3'b000;
							assign node415 = (inp[8]) ? node429 : node416;
								assign node416 = (inp[5]) ? node424 : node417;
									assign node417 = (inp[4]) ? node419 : 3'b000;
										assign node419 = (inp[1]) ? node421 : 3'b100;
											assign node421 = (inp[2]) ? 3'b000 : 3'b100;
									assign node424 = (inp[4]) ? 3'b100 : node425;
										assign node425 = (inp[1]) ? 3'b100 : 3'b000;
								assign node429 = (inp[2]) ? 3'b010 : node430;
									assign node430 = (inp[4]) ? 3'b110 : node431;
										assign node431 = (inp[1]) ? node433 : 3'b101;
											assign node433 = (inp[3]) ? 3'b100 : 3'b010;
						assign node438 = (inp[1]) ? 3'b000 : node439;
							assign node439 = (inp[2]) ? node445 : node440;
								assign node440 = (inp[8]) ? node442 : 3'b100;
									assign node442 = (inp[11]) ? 3'b100 : 3'b010;
								assign node445 = (inp[11]) ? node449 : node446;
									assign node446 = (inp[8]) ? 3'b100 : 3'b000;
									assign node449 = (inp[8]) ? 3'b000 : 3'b100;
					assign node453 = (inp[10]) ? node489 : node454;
						assign node454 = (inp[8]) ? node468 : node455;
							assign node455 = (inp[11]) ? node463 : node456;
								assign node456 = (inp[1]) ? node458 : 3'b101;
									assign node458 = (inp[5]) ? 3'b110 : node459;
										assign node459 = (inp[2]) ? 3'b110 : 3'b001;
								assign node463 = (inp[5]) ? 3'b110 : node464;
									assign node464 = (inp[2]) ? 3'b010 : 3'b110;
							assign node468 = (inp[2]) ? node482 : node469;
								assign node469 = (inp[3]) ? node477 : node470;
									assign node470 = (inp[11]) ? node474 : node471;
										assign node471 = (inp[1]) ? 3'b101 : 3'b011;
										assign node474 = (inp[5]) ? 3'b010 : 3'b001;
									assign node477 = (inp[1]) ? node479 : 3'b101;
										assign node479 = (inp[5]) ? 3'b001 : 3'b101;
								assign node482 = (inp[3]) ? 3'b001 : node483;
									assign node483 = (inp[4]) ? 3'b101 : node484;
										assign node484 = (inp[11]) ? 3'b001 : 3'b011;
						assign node489 = (inp[11]) ? node511 : node490;
							assign node490 = (inp[2]) ? node500 : node491;
								assign node491 = (inp[8]) ? node497 : node492;
									assign node492 = (inp[3]) ? node494 : 3'b110;
										assign node494 = (inp[4]) ? 3'b100 : 3'b000;
									assign node497 = (inp[1]) ? 3'b010 : 3'b001;
								assign node500 = (inp[1]) ? node506 : node501;
									assign node501 = (inp[8]) ? node503 : 3'b010;
										assign node503 = (inp[3]) ? 3'b110 : 3'b111;
									assign node506 = (inp[4]) ? node508 : 3'b010;
										assign node508 = (inp[5]) ? 3'b010 : 3'b100;
							assign node511 = (inp[2]) ? node525 : node512;
								assign node512 = (inp[1]) ? node516 : node513;
									assign node513 = (inp[8]) ? 3'b110 : 3'b010;
									assign node516 = (inp[8]) ? node522 : node517;
										assign node517 = (inp[4]) ? node519 : 3'b100;
											assign node519 = (inp[3]) ? 3'b000 : 3'b100;
										assign node522 = (inp[3]) ? 3'b100 : 3'b010;
								assign node525 = (inp[4]) ? node527 : 3'b100;
									assign node527 = (inp[5]) ? 3'b000 : 3'b100;
				assign node530 = (inp[7]) ? node544 : node531;
					assign node531 = (inp[10]) ? 3'b000 : node532;
						assign node532 = (inp[8]) ? node534 : 3'b000;
							assign node534 = (inp[1]) ? 3'b000 : node535;
								assign node535 = (inp[4]) ? node537 : 3'b100;
									assign node537 = (inp[11]) ? 3'b000 : node538;
										assign node538 = (inp[2]) ? 3'b000 : 3'b100;
					assign node544 = (inp[10]) ? node572 : node545;
						assign node545 = (inp[1]) ? node561 : node546;
							assign node546 = (inp[8]) ? node556 : node547;
								assign node547 = (inp[3]) ? 3'b010 : node548;
									assign node548 = (inp[4]) ? node550 : 3'b010;
										assign node550 = (inp[11]) ? 3'b100 : node551;
											assign node551 = (inp[2]) ? 3'b100 : 3'b010;
								assign node556 = (inp[11]) ? 3'b100 : node557;
									assign node557 = (inp[4]) ? 3'b010 : 3'b110;
							assign node561 = (inp[8]) ? node565 : node562;
								assign node562 = (inp[11]) ? 3'b100 : 3'b000;
								assign node565 = (inp[11]) ? node569 : node566;
									assign node566 = (inp[4]) ? 3'b100 : 3'b110;
									assign node569 = (inp[2]) ? 3'b000 : 3'b100;
						assign node572 = (inp[8]) ? node574 : 3'b000;
							assign node574 = (inp[1]) ? 3'b000 : node575;
								assign node575 = (inp[3]) ? 3'b100 : node576;
									assign node576 = (inp[5]) ? node582 : node577;
										assign node577 = (inp[2]) ? node579 : 3'b100;
											assign node579 = (inp[11]) ? 3'b000 : 3'b100;
										assign node582 = (inp[2]) ? 3'b100 : 3'b010;

endmodule