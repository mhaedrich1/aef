module dtc_split33_bm48 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node2;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node6;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node11;
	wire [14-1:0] node12;
	wire [14-1:0] node14;
	wire [14-1:0] node20;
	wire [14-1:0] node21;
	wire [14-1:0] node22;
	wire [14-1:0] node23;
	wire [14-1:0] node24;
	wire [14-1:0] node29;
	wire [14-1:0] node30;
	wire [14-1:0] node32;
	wire [14-1:0] node36;
	wire [14-1:0] node37;
	wire [14-1:0] node39;
	wire [14-1:0] node40;
	wire [14-1:0] node45;
	wire [14-1:0] node47;
	wire [14-1:0] node48;
	wire [14-1:0] node49;
	wire [14-1:0] node51;
	wire [14-1:0] node53;
	wire [14-1:0] node55;
	wire [14-1:0] node57;
	wire [14-1:0] node60;
	wire [14-1:0] node61;
	wire [14-1:0] node64;
	wire [14-1:0] node65;
	wire [14-1:0] node66;
	wire [14-1:0] node71;
	wire [14-1:0] node73;
	wire [14-1:0] node75;
	wire [14-1:0] node77;
	wire [14-1:0] node78;
	wire [14-1:0] node80;
	wire [14-1:0] node83;
	wire [14-1:0] node86;
	wire [14-1:0] node87;
	wire [14-1:0] node89;
	wire [14-1:0] node90;
	wire [14-1:0] node91;
	wire [14-1:0] node92;
	wire [14-1:0] node94;
	wire [14-1:0] node96;
	wire [14-1:0] node99;
	wire [14-1:0] node101;
	wire [14-1:0] node102;
	wire [14-1:0] node107;
	wire [14-1:0] node109;
	wire [14-1:0] node111;
	wire [14-1:0] node112;
	wire [14-1:0] node114;
	wire [14-1:0] node118;
	wire [14-1:0] node119;
	wire [14-1:0] node120;
	wire [14-1:0] node122;
	wire [14-1:0] node123;
	wire [14-1:0] node124;
	wire [14-1:0] node126;
	wire [14-1:0] node127;
	wire [14-1:0] node131;
	wire [14-1:0] node132;
	wire [14-1:0] node133;
	wire [14-1:0] node137;
	wire [14-1:0] node142;
	wire [14-1:0] node143;
	wire [14-1:0] node144;
	wire [14-1:0] node145;
	wire [14-1:0] node146;
	wire [14-1:0] node150;
	wire [14-1:0] node152;
	wire [14-1:0] node154;
	wire [14-1:0] node157;
	wire [14-1:0] node158;
	wire [14-1:0] node159;
	wire [14-1:0] node160;
	wire [14-1:0] node162;
	wire [14-1:0] node168;
	wire [14-1:0] node169;
	wire [14-1:0] node171;
	wire [14-1:0] node174;
	wire [14-1:0] node176;
	wire [14-1:0] node177;
	wire [14-1:0] node178;
	wire [14-1:0] node180;
	wire [14-1:0] node184;
	wire [14-1:0] node185;
	wire [14-1:0] node189;
	wire [14-1:0] node190;
	wire [14-1:0] node191;
	wire [14-1:0] node192;
	wire [14-1:0] node194;
	wire [14-1:0] node195;
	wire [14-1:0] node197;
	wire [14-1:0] node199;
	wire [14-1:0] node200;
	wire [14-1:0] node206;
	wire [14-1:0] node207;
	wire [14-1:0] node208;
	wire [14-1:0] node209;
	wire [14-1:0] node210;
	wire [14-1:0] node212;
	wire [14-1:0] node214;
	wire [14-1:0] node217;
	wire [14-1:0] node218;
	wire [14-1:0] node219;
	wire [14-1:0] node224;
	wire [14-1:0] node226;
	wire [14-1:0] node228;
	wire [14-1:0] node230;
	wire [14-1:0] node231;
	wire [14-1:0] node235;
	wire [14-1:0] node237;
	wire [14-1:0] node238;
	wire [14-1:0] node239;
	wire [14-1:0] node241;
	wire [14-1:0] node246;
	wire [14-1:0] node247;
	wire [14-1:0] node248;
	wire [14-1:0] node249;
	wire [14-1:0] node252;
	wire [14-1:0] node253;
	wire [14-1:0] node254;
	wire [14-1:0] node259;
	wire [14-1:0] node260;
	wire [14-1:0] node261;
	wire [14-1:0] node266;
	wire [14-1:0] node268;
	wire [14-1:0] node269;
	wire [14-1:0] node270;
	wire [14-1:0] node271;
	wire [14-1:0] node272;
	wire [14-1:0] node277;
	wire [14-1:0] node279;
	wire [14-1:0] node282;
	wire [14-1:0] node283;
	wire [14-1:0] node284;
	wire [14-1:0] node289;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node293;
	wire [14-1:0] node294;
	wire [14-1:0] node295;
	wire [14-1:0] node296;
	wire [14-1:0] node297;
	wire [14-1:0] node300;
	wire [14-1:0] node301;
	wire [14-1:0] node307;
	wire [14-1:0] node309;
	wire [14-1:0] node310;
	wire [14-1:0] node314;
	wire [14-1:0] node315;
	wire [14-1:0] node317;
	wire [14-1:0] node318;
	wire [14-1:0] node319;
	wire [14-1:0] node320;
	wire [14-1:0] node322;
	wire [14-1:0] node328;
	wire [14-1:0] node330;
	wire [14-1:0] node331;
	wire [14-1:0] node334;
	wire [14-1:0] node336;
	wire [14-1:0] node338;
	wire [14-1:0] node341;
	wire [14-1:0] node342;
	wire [14-1:0] node343;
	wire [14-1:0] node344;
	wire [14-1:0] node346;
	wire [14-1:0] node347;
	wire [14-1:0] node348;
	wire [14-1:0] node350;
	wire [14-1:0] node354;
	wire [14-1:0] node355;
	wire [14-1:0] node360;
	wire [14-1:0] node361;
	wire [14-1:0] node362;
	wire [14-1:0] node364;
	wire [14-1:0] node365;
	wire [14-1:0] node367;
	wire [14-1:0] node370;
	wire [14-1:0] node374;
	wire [14-1:0] node376;
	wire [14-1:0] node378;
	wire [14-1:0] node379;
	wire [14-1:0] node381;
	wire [14-1:0] node386;
	wire [14-1:0] node387;
	wire [14-1:0] node388;
	wire [14-1:0] node389;
	wire [14-1:0] node390;
	wire [14-1:0] node391;
	wire [14-1:0] node392;
	wire [14-1:0] node393;
	wire [14-1:0] node398;
	wire [14-1:0] node400;
	wire [14-1:0] node402;
	wire [14-1:0] node405;
	wire [14-1:0] node406;
	wire [14-1:0] node407;
	wire [14-1:0] node408;
	wire [14-1:0] node409;
	wire [14-1:0] node414;
	wire [14-1:0] node416;
	wire [14-1:0] node418;
	wire [14-1:0] node421;
	wire [14-1:0] node422;
	wire [14-1:0] node423;
	wire [14-1:0] node425;
	wire [14-1:0] node426;
	wire [14-1:0] node428;
	wire [14-1:0] node432;
	wire [14-1:0] node433;
	wire [14-1:0] node434;
	wire [14-1:0] node438;
	wire [14-1:0] node440;
	wire [14-1:0] node443;
	wire [14-1:0] node444;
	wire [14-1:0] node445;
	wire [14-1:0] node446;
	wire [14-1:0] node451;
	wire [14-1:0] node453;
	wire [14-1:0] node455;
	wire [14-1:0] node458;
	wire [14-1:0] node459;
	wire [14-1:0] node460;
	wire [14-1:0] node461;
	wire [14-1:0] node462;
	wire [14-1:0] node463;
	wire [14-1:0] node464;
	wire [14-1:0] node469;
	wire [14-1:0] node471;
	wire [14-1:0] node473;
	wire [14-1:0] node476;
	wire [14-1:0] node478;
	wire [14-1:0] node480;
	wire [14-1:0] node482;
	wire [14-1:0] node485;
	wire [14-1:0] node486;
	wire [14-1:0] node487;
	wire [14-1:0] node488;
	wire [14-1:0] node489;
	wire [14-1:0] node494;
	wire [14-1:0] node496;
	wire [14-1:0] node498;
	wire [14-1:0] node502;
	wire [14-1:0] node503;
	wire [14-1:0] node504;
	wire [14-1:0] node506;
	wire [14-1:0] node508;
	wire [14-1:0] node510;
	wire [14-1:0] node513;
	wire [14-1:0] node514;
	wire [14-1:0] node515;
	wire [14-1:0] node516;
	wire [14-1:0] node521;
	wire [14-1:0] node523;
	wire [14-1:0] node524;
	wire [14-1:0] node528;
	wire [14-1:0] node529;
	wire [14-1:0] node530;
	wire [14-1:0] node531;
	wire [14-1:0] node536;
	wire [14-1:0] node538;
	wire [14-1:0] node540;
	wire [14-1:0] node543;
	wire [14-1:0] node544;
	wire [14-1:0] node545;
	wire [14-1:0] node546;
	wire [14-1:0] node547;
	wire [14-1:0] node552;
	wire [14-1:0] node554;
	wire [14-1:0] node556;
	wire [14-1:0] node559;
	wire [14-1:0] node560;
	wire [14-1:0] node561;
	wire [14-1:0] node562;
	wire [14-1:0] node566;
	wire [14-1:0] node567;
	wire [14-1:0] node569;
	wire [14-1:0] node570;
	wire [14-1:0] node571;
	wire [14-1:0] node573;
	wire [14-1:0] node579;
	wire [14-1:0] node580;
	wire [14-1:0] node581;
	wire [14-1:0] node582;
	wire [14-1:0] node583;
	wire [14-1:0] node584;
	wire [14-1:0] node589;
	wire [14-1:0] node592;
	wire [14-1:0] node593;
	wire [14-1:0] node597;
	wire [14-1:0] node598;
	wire [14-1:0] node599;
	wire [14-1:0] node600;
	wire [14-1:0] node604;
	wire [14-1:0] node607;
	wire [14-1:0] node608;
	wire [14-1:0] node612;
	wire [14-1:0] node613;
	wire [14-1:0] node614;
	wire [14-1:0] node615;
	wire [14-1:0] node616;
	wire [14-1:0] node617;
	wire [14-1:0] node618;
	wire [14-1:0] node621;
	wire [14-1:0] node622;
	wire [14-1:0] node624;
	wire [14-1:0] node628;
	wire [14-1:0] node630;
	wire [14-1:0] node631;
	wire [14-1:0] node632;
	wire [14-1:0] node633;
	wire [14-1:0] node636;
	wire [14-1:0] node639;
	wire [14-1:0] node643;
	wire [14-1:0] node644;
	wire [14-1:0] node645;
	wire [14-1:0] node646;
	wire [14-1:0] node648;
	wire [14-1:0] node649;
	wire [14-1:0] node652;
	wire [14-1:0] node656;
	wire [14-1:0] node657;
	wire [14-1:0] node658;
	wire [14-1:0] node659;
	wire [14-1:0] node662;
	wire [14-1:0] node665;
	wire [14-1:0] node667;
	wire [14-1:0] node670;
	wire [14-1:0] node673;
	wire [14-1:0] node674;
	wire [14-1:0] node675;
	wire [14-1:0] node676;
	wire [14-1:0] node677;
	wire [14-1:0] node681;
	wire [14-1:0] node682;
	wire [14-1:0] node685;
	wire [14-1:0] node689;
	wire [14-1:0] node690;
	wire [14-1:0] node691;
	wire [14-1:0] node693;
	wire [14-1:0] node698;
	wire [14-1:0] node699;
	wire [14-1:0] node700;
	wire [14-1:0] node701;
	wire [14-1:0] node702;
	wire [14-1:0] node703;
	wire [14-1:0] node706;
	wire [14-1:0] node708;
	wire [14-1:0] node711;
	wire [14-1:0] node712;
	wire [14-1:0] node713;
	wire [14-1:0] node717;
	wire [14-1:0] node720;
	wire [14-1:0] node721;
	wire [14-1:0] node723;
	wire [14-1:0] node724;
	wire [14-1:0] node728;
	wire [14-1:0] node729;
	wire [14-1:0] node730;
	wire [14-1:0] node734;
	wire [14-1:0] node737;
	wire [14-1:0] node738;
	wire [14-1:0] node739;
	wire [14-1:0] node740;
	wire [14-1:0] node745;
	wire [14-1:0] node747;
	wire [14-1:0] node749;
	wire [14-1:0] node752;
	wire [14-1:0] node753;
	wire [14-1:0] node754;
	wire [14-1:0] node755;
	wire [14-1:0] node760;
	wire [14-1:0] node762;
	wire [14-1:0] node764;
	wire [14-1:0] node767;
	wire [14-1:0] node768;
	wire [14-1:0] node769;
	wire [14-1:0] node770;
	wire [14-1:0] node771;
	wire [14-1:0] node772;
	wire [14-1:0] node773;
	wire [14-1:0] node774;
	wire [14-1:0] node780;
	wire [14-1:0] node781;
	wire [14-1:0] node782;
	wire [14-1:0] node783;
	wire [14-1:0] node787;
	wire [14-1:0] node789;
	wire [14-1:0] node793;
	wire [14-1:0] node794;
	wire [14-1:0] node795;
	wire [14-1:0] node796;
	wire [14-1:0] node800;
	wire [14-1:0] node802;
	wire [14-1:0] node804;
	wire [14-1:0] node807;
	wire [14-1:0] node808;
	wire [14-1:0] node809;
	wire [14-1:0] node810;
	wire [14-1:0] node814;
	wire [14-1:0] node815;
	wire [14-1:0] node819;
	wire [14-1:0] node821;
	wire [14-1:0] node824;
	wire [14-1:0] node825;
	wire [14-1:0] node826;
	wire [14-1:0] node827;
	wire [14-1:0] node828;
	wire [14-1:0] node832;
	wire [14-1:0] node833;
	wire [14-1:0] node836;
	wire [14-1:0] node838;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node843;
	wire [14-1:0] node844;
	wire [14-1:0] node848;
	wire [14-1:0] node850;
	wire [14-1:0] node853;
	wire [14-1:0] node855;
	wire [14-1:0] node857;
	wire [14-1:0] node860;
	wire [14-1:0] node861;
	wire [14-1:0] node862;
	wire [14-1:0] node863;
	wire [14-1:0] node868;
	wire [14-1:0] node870;
	wire [14-1:0] node872;
	wire [14-1:0] node875;
	wire [14-1:0] node876;
	wire [14-1:0] node877;
	wire [14-1:0] node878;
	wire [14-1:0] node879;
	wire [14-1:0] node884;
	wire [14-1:0] node886;
	wire [14-1:0] node888;
	wire [14-1:0] node891;
	wire [14-1:0] node892;
	wire [14-1:0] node893;
	wire [14-1:0] node894;
	wire [14-1:0] node899;
	wire [14-1:0] node901;
	wire [14-1:0] node903;
	wire [14-1:0] node906;
	wire [14-1:0] node907;
	wire [14-1:0] node908;
	wire [14-1:0] node909;
	wire [14-1:0] node910;
	wire [14-1:0] node911;
	wire [14-1:0] node914;
	wire [14-1:0] node916;
	wire [14-1:0] node917;
	wire [14-1:0] node918;
	wire [14-1:0] node924;
	wire [14-1:0] node926;
	wire [14-1:0] node927;
	wire [14-1:0] node928;
	wire [14-1:0] node929;
	wire [14-1:0] node930;
	wire [14-1:0] node933;
	wire [14-1:0] node938;
	wire [14-1:0] node941;
	wire [14-1:0] node942;
	wire [14-1:0] node943;
	wire [14-1:0] node944;
	wire [14-1:0] node945;
	wire [14-1:0] node950;
	wire [14-1:0] node952;
	wire [14-1:0] node954;
	wire [14-1:0] node957;
	wire [14-1:0] node958;
	wire [14-1:0] node959;
	wire [14-1:0] node960;
	wire [14-1:0] node965;
	wire [14-1:0] node967;
	wire [14-1:0] node969;
	wire [14-1:0] node972;
	wire [14-1:0] node973;
	wire [14-1:0] node974;
	wire [14-1:0] node975;
	wire [14-1:0] node976;
	wire [14-1:0] node981;
	wire [14-1:0] node983;
	wire [14-1:0] node985;
	wire [14-1:0] node988;
	wire [14-1:0] node989;
	wire [14-1:0] node990;
	wire [14-1:0] node991;
	wire [14-1:0] node993;
	wire [14-1:0] node995;
	wire [14-1:0] node996;
	wire [14-1:0] node1000;
	wire [14-1:0] node1001;
	wire [14-1:0] node1002;
	wire [14-1:0] node1004;
	wire [14-1:0] node1009;
	wire [14-1:0] node1011;
	wire [14-1:0] node1012;
	wire [14-1:0] node1014;
	wire [14-1:0] node1017;
	wire [14-1:0] node1018;
	wire [14-1:0] node1019;
	wire [14-1:0] node1023;
	wire [14-1:0] node1026;
	wire [14-1:0] node1027;
	wire [14-1:0] node1028;
	wire [14-1:0] node1030;
	wire [14-1:0] node1032;
	wire [14-1:0] node1035;
	wire [14-1:0] node1036;
	wire [14-1:0] node1040;
	wire [14-1:0] node1041;
	wire [14-1:0] node1043;
	wire [14-1:0] node1044;
	wire [14-1:0] node1045;
	wire [14-1:0] node1048;
	wire [14-1:0] node1051;
	wire [14-1:0] node1054;
	wire [14-1:0] node1055;
	wire [14-1:0] node1057;

	assign outp = (inp[10]) ? node386 : node1;
		assign node1 = (inp[8]) ? node189 : node2;
			assign node2 = (inp[13]) ? node86 : node3;
				assign node3 = (inp[12]) ? node45 : node4;
					assign node4 = (inp[11]) ? node6 : 14'b00000100000011;
						assign node6 = (inp[1]) ? node8 : 14'b00000000000000;
							assign node8 = (inp[7]) ? node20 : node9;
								assign node9 = (inp[3]) ? 14'b00000000000000 : node10;
									assign node10 = (inp[6]) ? 14'b00000000000000 : node11;
										assign node11 = (inp[9]) ? 14'b00000000000000 : node12;
											assign node12 = (inp[0]) ? node14 : 14'b00000000000000;
												assign node14 = (inp[4]) ? 14'b00000000000000 : 14'b00100000000011;
								assign node20 = (inp[6]) ? node36 : node21;
									assign node21 = (inp[2]) ? node29 : node22;
										assign node22 = (inp[0]) ? 14'b00000000000000 : node23;
											assign node23 = (inp[9]) ? 14'b10010000001101 : node24;
												assign node24 = (inp[3]) ? 14'b10010000001101 : 14'b00000000000000;
										assign node29 = (inp[9]) ? 14'b00000000000000 : node30;
											assign node30 = (inp[5]) ? node32 : 14'b00000000000000;
												assign node32 = (inp[3]) ? 14'b00000000000000 : 14'b00100000000011;
									assign node36 = (inp[5]) ? 14'b00000000000000 : node37;
										assign node37 = (inp[3]) ? node39 : 14'b00000000000000;
											assign node39 = (inp[0]) ? 14'b01001000000100 : node40;
												assign node40 = (inp[2]) ? 14'b00000000000000 : 14'b10100000101010;
					assign node45 = (inp[11]) ? node47 : 14'b00000000000000;
						assign node47 = (inp[9]) ? node71 : node48;
							assign node48 = (inp[3]) ? node60 : node49;
								assign node49 = (inp[1]) ? node51 : 14'b00000000000000;
									assign node51 = (inp[6]) ? node53 : 14'b10000100011000;
										assign node53 = (inp[7]) ? node55 : 14'b00000000000000;
											assign node55 = (inp[5]) ? node57 : 14'b00000000000000;
												assign node57 = (inp[0]) ? 14'b00000000000000 : 14'b10100000001000;
								assign node60 = (inp[1]) ? node64 : node61;
									assign node61 = (inp[6]) ? 14'b01100000001010 : 14'b00000000000000;
									assign node64 = (inp[0]) ? 14'b00000000000000 : node65;
										assign node65 = (inp[2]) ? 14'b00000000000000 : node66;
											assign node66 = (inp[6]) ? 14'b00000000000000 : 14'b01001000000100;
							assign node71 = (inp[5]) ? node73 : 14'b00000000000000;
								assign node73 = (inp[3]) ? node75 : 14'b00000000000000;
									assign node75 = (inp[1]) ? node77 : 14'b00000000000000;
										assign node77 = (inp[6]) ? node83 : node78;
											assign node78 = (inp[7]) ? node80 : 14'b00000000000000;
												assign node80 = (inp[2]) ? 14'b00000000000000 : 14'b01001000000100;
											assign node83 = (inp[7]) ? 14'b00000000000000 : 14'b01001000001100;
				assign node86 = (inp[3]) ? node118 : node87;
					assign node87 = (inp[1]) ? node89 : 14'b00000000000000;
						assign node89 = (inp[11]) ? node107 : node90;
							assign node90 = (inp[6]) ? 14'b00000000000000 : node91;
								assign node91 = (inp[9]) ? node99 : node92;
									assign node92 = (inp[12]) ? node94 : 14'b11000000000100;
										assign node94 = (inp[2]) ? node96 : 14'b00000000000000;
											assign node96 = (inp[0]) ? 14'b10000000101100 : 14'b00000000000000;
									assign node99 = (inp[12]) ? node101 : 14'b00000000000000;
										assign node101 = (inp[2]) ? 14'b00000000000000 : node102;
											assign node102 = (inp[0]) ? 14'b00000000000000 : 14'b11110111110010;
							assign node107 = (inp[7]) ? node109 : 14'b00000000000000;
								assign node109 = (inp[9]) ? node111 : 14'b00000000000000;
									assign node111 = (inp[6]) ? 14'b00000000000000 : node112;
										assign node112 = (inp[12]) ? node114 : 14'b00000000000000;
											assign node114 = (inp[2]) ? 14'b00000000000000 : 14'b10100010001100;
					assign node118 = (inp[6]) ? node142 : node119;
						assign node119 = (inp[2]) ? 14'b00000000000000 : node120;
							assign node120 = (inp[1]) ? node122 : 14'b00000000000000;
								assign node122 = (inp[0]) ? 14'b00000000000000 : node123;
									assign node123 = (inp[7]) ? node131 : node124;
										assign node124 = (inp[11]) ? node126 : 14'b00000000000000;
											assign node126 = (inp[12]) ? 14'b00000000000000 : node127;
												assign node127 = (inp[9]) ? 14'b10000100101010 : 14'b10000100111010;
										assign node131 = (inp[11]) ? node137 : node132;
											assign node132 = (inp[9]) ? 14'b11110111110010 : node133;
												assign node133 = (inp[5]) ? 14'b11110111110010 : 14'b00000000000000;
											assign node137 = (inp[12]) ? 14'b10100010001100 : 14'b10000100111010;
						assign node142 = (inp[11]) ? node168 : node143;
							assign node143 = (inp[12]) ? node157 : node144;
								assign node144 = (inp[7]) ? node150 : node145;
									assign node145 = (inp[1]) ? 14'b00000000000000 : node146;
										assign node146 = (inp[9]) ? 14'b00000000000000 : 14'b11000000000100;
									assign node150 = (inp[1]) ? node152 : 14'b00000000000000;
										assign node152 = (inp[0]) ? node154 : 14'b00000000000000;
											assign node154 = (inp[9]) ? 14'b01100000000110 : 14'b00000000000000;
								assign node157 = (inp[7]) ? 14'b00000000000000 : node158;
									assign node158 = (inp[0]) ? 14'b00000000000000 : node159;
										assign node159 = (inp[2]) ? 14'b00000000000000 : node160;
											assign node160 = (inp[4]) ? node162 : 14'b00000000000000;
												assign node162 = (inp[5]) ? 14'b00000000000000 : 14'b00000000000000;
							assign node168 = (inp[9]) ? node174 : node169;
								assign node169 = (inp[12]) ? node171 : 14'b00000000000000;
									assign node171 = (inp[1]) ? 14'b00000000000000 : 14'b00100100001101;
								assign node174 = (inp[1]) ? node176 : 14'b00000000000000;
									assign node176 = (inp[12]) ? node184 : node177;
										assign node177 = (inp[5]) ? 14'b01001000000101 : node178;
											assign node178 = (inp[7]) ? node180 : 14'b00000000000000;
												assign node180 = (inp[2]) ? 14'b10000010001100 : 14'b10000000001000;
										assign node184 = (inp[7]) ? 14'b00000000000000 : node185;
											assign node185 = (inp[5]) ? 14'b00000000011100 : 14'b00000000000000;
			assign node189 = (inp[12]) ? node289 : node190;
				assign node190 = (inp[1]) ? node206 : node191;
					assign node191 = (inp[9]) ? 14'b00000000000000 : node192;
						assign node192 = (inp[5]) ? node194 : 14'b00000000000000;
							assign node194 = (inp[0]) ? 14'b00000000000000 : node195;
								assign node195 = (inp[3]) ? node197 : 14'b00000000000000;
									assign node197 = (inp[13]) ? node199 : 14'b00000000000000;
										assign node199 = (inp[2]) ? 14'b00000000000000 : node200;
											assign node200 = (inp[11]) ? 14'b00100000000011 : 14'b00000000000000;
					assign node206 = (inp[11]) ? node246 : node207;
						assign node207 = (inp[13]) ? node235 : node208;
							assign node208 = (inp[6]) ? node224 : node209;
								assign node209 = (inp[3]) ? node217 : node210;
									assign node210 = (inp[0]) ? node212 : 14'b00000000000000;
										assign node212 = (inp[2]) ? node214 : 14'b00000000000000;
											assign node214 = (inp[9]) ? 14'b00000000000000 : 14'b10000000011010;
									assign node217 = (inp[2]) ? 14'b00000000000000 : node218;
										assign node218 = (inp[0]) ? 14'b00000000000000 : node219;
											assign node219 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
								assign node224 = (inp[9]) ? node226 : 14'b00000000000000;
									assign node226 = (inp[3]) ? node228 : 14'b00000000000000;
										assign node228 = (inp[7]) ? node230 : 14'b00000000000000;
											assign node230 = (inp[5]) ? 14'b00000000011100 : node231;
												assign node231 = (inp[2]) ? 14'b00000000000000 : 14'b01000000010000;
							assign node235 = (inp[6]) ? node237 : 14'b00000000000000;
								assign node237 = (inp[5]) ? 14'b00000000000000 : node238;
									assign node238 = (inp[2]) ? 14'b00000000000000 : node239;
										assign node239 = (inp[9]) ? node241 : 14'b00000000000000;
											assign node241 = (inp[0]) ? 14'b00000000000000 : 14'b00000000011100;
						assign node246 = (inp[9]) ? node266 : node247;
							assign node247 = (inp[3]) ? node259 : node248;
								assign node248 = (inp[6]) ? node252 : node249;
									assign node249 = (inp[13]) ? 14'b00000000011100 : 14'b01001000000100;
									assign node252 = (inp[7]) ? 14'b00000000000000 : node253;
										assign node253 = (inp[13]) ? 14'b00000000000000 : node254;
											assign node254 = (inp[5]) ? 14'b00000000000000 : 14'b11000000000100;
								assign node259 = (inp[7]) ? 14'b00000000000000 : node260;
									assign node260 = (inp[2]) ? 14'b00000000000000 : node261;
										assign node261 = (inp[13]) ? 14'b00000000000000 : 14'b00000100000001;
							assign node266 = (inp[3]) ? node268 : 14'b00000000000000;
								assign node268 = (inp[5]) ? node282 : node269;
									assign node269 = (inp[7]) ? node277 : node270;
										assign node270 = (inp[2]) ? 14'b00000000000000 : node271;
											assign node271 = (inp[6]) ? 14'b00000000000000 : node272;
												assign node272 = (inp[4]) ? 14'b00000000000000 : 14'b00000000011100;
										assign node277 = (inp[13]) ? node279 : 14'b01100000001010;
											assign node279 = (inp[6]) ? 14'b10100010001100 : 14'b00000000000000;
									assign node282 = (inp[2]) ? 14'b00000000000000 : node283;
										assign node283 = (inp[7]) ? 14'b00000000000000 : node284;
											assign node284 = (inp[4]) ? 14'b00000100000001 : 14'b00000000000000;
				assign node289 = (inp[13]) ? node341 : node290;
					assign node290 = (inp[6]) ? node314 : node291;
						assign node291 = (inp[1]) ? node293 : 14'b00000000000000;
							assign node293 = (inp[9]) ? node307 : node294;
								assign node294 = (inp[3]) ? 14'b00000000000000 : node295;
									assign node295 = (inp[11]) ? 14'b00100100011111 : node296;
										assign node296 = (inp[0]) ? node300 : node297;
											assign node297 = (inp[4]) ? 14'b00000000000000 : 14'b00100000000011;
											assign node300 = (inp[2]) ? 14'b00000000000000 : node301;
												assign node301 = (inp[4]) ? 14'b00000000000000 : 14'b00000000011100;
								assign node307 = (inp[3]) ? node309 : 14'b00000000000000;
									assign node309 = (inp[5]) ? 14'b00000000000000 : node310;
										assign node310 = (inp[2]) ? 14'b00000000000000 : 14'b00001000000101;
						assign node314 = (inp[9]) ? node328 : node315;
							assign node315 = (inp[1]) ? node317 : 14'b00000000000000;
								assign node317 = (inp[3]) ? 14'b00000000000000 : node318;
									assign node318 = (inp[11]) ? 14'b01000100000100 : node319;
										assign node319 = (inp[0]) ? 14'b00000000000000 : node320;
											assign node320 = (inp[7]) ? node322 : 14'b00000000000000;
												assign node322 = (inp[5]) ? 14'b10100100111111 : 14'b00000000000000;
							assign node328 = (inp[3]) ? node330 : 14'b00000000000000;
								assign node330 = (inp[1]) ? node334 : node331;
									assign node331 = (inp[11]) ? 14'b10100010001100 : 14'b11110111110010;
									assign node334 = (inp[7]) ? node336 : 14'b00000000000000;
										assign node336 = (inp[5]) ? node338 : 14'b00000000000000;
											assign node338 = (inp[11]) ? 14'b10000000011010 : 14'b00000000000000;
					assign node341 = (inp[11]) ? 14'b01000000010100 : node342;
						assign node342 = (inp[6]) ? node360 : node343;
							assign node343 = (inp[2]) ? 14'b00000000000000 : node344;
								assign node344 = (inp[1]) ? node346 : 14'b00000000000000;
									assign node346 = (inp[7]) ? node354 : node347;
										assign node347 = (inp[0]) ? 14'b00000000000000 : node348;
											assign node348 = (inp[3]) ? node350 : 14'b00000000000000;
												assign node350 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
										assign node354 = (inp[3]) ? 14'b00000000000000 : node355;
											assign node355 = (inp[9]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node360 = (inp[9]) ? node374 : node361;
								assign node361 = (inp[3]) ? 14'b00000000000000 : node362;
									assign node362 = (inp[1]) ? node364 : 14'b00000000000000;
										assign node364 = (inp[5]) ? node370 : node365;
											assign node365 = (inp[7]) ? node367 : 14'b10010100011100;
												assign node367 = (inp[0]) ? 14'b00000000000000 : 14'b10010010001100;
											assign node370 = (inp[7]) ? 14'b11100100010100 : 14'b11100100000100;
								assign node374 = (inp[3]) ? node376 : 14'b00000000000000;
									assign node376 = (inp[1]) ? node378 : 14'b01001000000100;
										assign node378 = (inp[0]) ? 14'b00000000000000 : node379;
											assign node379 = (inp[5]) ? node381 : 14'b00000000000000;
												assign node381 = (inp[7]) ? 14'b01001000001001 : 14'b00000000000000;
		assign node386 = (inp[1]) ? node612 : node387;
			assign node387 = (inp[3]) ? node543 : node388;
				assign node388 = (inp[6]) ? node458 : node389;
					assign node389 = (inp[5]) ? node405 : node390;
						assign node390 = (inp[8]) ? node398 : node391;
							assign node391 = (inp[11]) ? 14'b00000000000000 : node392;
								assign node392 = (inp[12]) ? 14'b00000000000000 : node393;
									assign node393 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
							assign node398 = (inp[11]) ? node400 : 14'b00000000000000;
								assign node400 = (inp[12]) ? node402 : 14'b00000000000000;
									assign node402 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node405 = (inp[0]) ? node421 : node406;
							assign node406 = (inp[11]) ? node414 : node407;
								assign node407 = (inp[13]) ? 14'b00000000000000 : node408;
									assign node408 = (inp[8]) ? 14'b00000000000000 : node409;
										assign node409 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node414 = (inp[8]) ? node416 : 14'b00000000000000;
									assign node416 = (inp[13]) ? node418 : 14'b00000000000000;
										assign node418 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node421 = (inp[9]) ? node443 : node422;
								assign node422 = (inp[4]) ? node432 : node423;
									assign node423 = (inp[8]) ? node425 : 14'b00000000000000;
										assign node425 = (inp[2]) ? 14'b00000000000000 : node426;
											assign node426 = (inp[11]) ? node428 : 14'b00000000000000;
												assign node428 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node432 = (inp[8]) ? node438 : node433;
										assign node433 = (inp[13]) ? 14'b00000000000000 : node434;
											assign node434 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node438 = (inp[11]) ? node440 : 14'b00000000000000;
											assign node440 = (inp[2]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node443 = (inp[11]) ? node451 : node444;
									assign node444 = (inp[12]) ? 14'b00000000000000 : node445;
										assign node445 = (inp[13]) ? 14'b00000000000000 : node446;
											assign node446 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node451 = (inp[12]) ? node453 : 14'b00000000000000;
										assign node453 = (inp[8]) ? node455 : 14'b00000000000000;
											assign node455 = (inp[2]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node458 = (inp[9]) ? node502 : node459;
						assign node459 = (inp[5]) ? node485 : node460;
							assign node460 = (inp[4]) ? node476 : node461;
								assign node461 = (inp[8]) ? node469 : node462;
									assign node462 = (inp[11]) ? 14'b00000000000000 : node463;
										assign node463 = (inp[12]) ? 14'b00000000000000 : node464;
											assign node464 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node469 = (inp[12]) ? node471 : 14'b00000000000000;
										assign node471 = (inp[11]) ? node473 : 14'b00000000000000;
											assign node473 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node476 = (inp[8]) ? node478 : 14'b00000000000000;
									assign node478 = (inp[12]) ? node480 : 14'b00000000000000;
										assign node480 = (inp[13]) ? node482 : 14'b00000000000000;
											assign node482 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node485 = (inp[0]) ? 14'b00000000000000 : node486;
								assign node486 = (inp[13]) ? node494 : node487;
									assign node487 = (inp[8]) ? 14'b00000000000000 : node488;
										assign node488 = (inp[12]) ? 14'b00000000000000 : node489;
											assign node489 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node494 = (inp[8]) ? node496 : 14'b00000000000000;
										assign node496 = (inp[12]) ? node498 : 14'b00000000000000;
											assign node498 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node502 = (inp[7]) ? node528 : node503;
							assign node503 = (inp[4]) ? node513 : node504;
								assign node504 = (inp[5]) ? node506 : 14'b00000000000000;
									assign node506 = (inp[13]) ? node508 : 14'b00000000000000;
										assign node508 = (inp[2]) ? node510 : 14'b00000000000000;
											assign node510 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node513 = (inp[11]) ? node521 : node514;
									assign node514 = (inp[12]) ? 14'b00000000000000 : node515;
										assign node515 = (inp[8]) ? 14'b00000000000000 : node516;
											assign node516 = (inp[0]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node521 = (inp[12]) ? node523 : 14'b00000000000000;
										assign node523 = (inp[2]) ? 14'b00000000000000 : node524;
											assign node524 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node528 = (inp[12]) ? node536 : node529;
								assign node529 = (inp[13]) ? 14'b00000000000000 : node530;
									assign node530 = (inp[11]) ? 14'b00000000000000 : node531;
										assign node531 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node536 = (inp[13]) ? node538 : 14'b00000000000000;
									assign node538 = (inp[11]) ? node540 : 14'b00000000000000;
										assign node540 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
				assign node543 = (inp[6]) ? node559 : node544;
					assign node544 = (inp[13]) ? node552 : node545;
						assign node545 = (inp[8]) ? 14'b00000000000000 : node546;
							assign node546 = (inp[12]) ? 14'b00000000000000 : node547;
								assign node547 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
						assign node552 = (inp[8]) ? node554 : 14'b00000000000000;
							assign node554 = (inp[12]) ? node556 : 14'b00000000000000;
								assign node556 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node559 = (inp[12]) ? node579 : node560;
						assign node560 = (inp[8]) ? node566 : node561;
							assign node561 = (inp[13]) ? 14'b00000000000000 : node562;
								assign node562 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
							assign node566 = (inp[7]) ? 14'b00000000000000 : node567;
								assign node567 = (inp[13]) ? node569 : 14'b00000000000000;
									assign node569 = (inp[2]) ? 14'b00000000000000 : node570;
										assign node570 = (inp[0]) ? 14'b00000000000000 : node571;
											assign node571 = (inp[11]) ? node573 : 14'b00000000000000;
												assign node573 = (inp[4]) ? 14'b10000100101010 : 14'b10000100111010;
						assign node579 = (inp[13]) ? node597 : node580;
							assign node580 = (inp[11]) ? node592 : node581;
								assign node581 = (inp[9]) ? node589 : node582;
									assign node582 = (inp[8]) ? 14'b00000000000000 : node583;
										assign node583 = (inp[7]) ? 14'b00000000000000 : node584;
											assign node584 = (inp[2]) ? 14'b00000000000000 : 14'b10100100111000;
									assign node589 = (inp[8]) ? 14'b01100000001010 : 14'b00000000000000;
								assign node592 = (inp[8]) ? 14'b00000000000000 : node593;
									assign node593 = (inp[9]) ? 14'b00000000000000 : 14'b01001000000101;
							assign node597 = (inp[11]) ? node607 : node598;
								assign node598 = (inp[8]) ? node604 : node599;
									assign node599 = (inp[9]) ? 14'b00000000000000 : node600;
										assign node600 = (inp[7]) ? 14'b00000000000000 : 14'b10000000111000;
									assign node604 = (inp[9]) ? 14'b00100100001101 : 14'b00000000000000;
								assign node607 = (inp[8]) ? 14'b10000100001000 : node608;
									assign node608 = (inp[9]) ? 14'b00000000000000 : 14'b10010101111110;
			assign node612 = (inp[6]) ? node906 : node613;
				assign node613 = (inp[9]) ? node767 : node614;
					assign node614 = (inp[3]) ? node698 : node615;
						assign node615 = (inp[8]) ? node643 : node616;
							assign node616 = (inp[11]) ? node628 : node617;
								assign node617 = (inp[12]) ? node621 : node618;
									assign node618 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node621 = (inp[13]) ? 14'b00000000011101 : node622;
										assign node622 = (inp[0]) ? node624 : 14'b00000000000000;
											assign node624 = (inp[4]) ? 14'b00000000000000 : 14'b01001000000100;
								assign node628 = (inp[0]) ? node630 : 14'b00000000000000;
									assign node630 = (inp[4]) ? 14'b00000000000000 : node631;
										assign node631 = (inp[5]) ? node639 : node632;
											assign node632 = (inp[13]) ? node636 : node633;
												assign node633 = (inp[12]) ? 14'b00001000000101 : 14'b01000000000000;
												assign node636 = (inp[2]) ? 14'b00000000000000 : 14'b10000000001101;
											assign node639 = (inp[12]) ? 14'b00000000000000 : 14'b00000000011100;
							assign node643 = (inp[11]) ? node673 : node644;
								assign node644 = (inp[12]) ? node656 : node645;
									assign node645 = (inp[13]) ? 14'b00000000000000 : node646;
										assign node646 = (inp[0]) ? node648 : 14'b00100000000011;
											assign node648 = (inp[2]) ? node652 : node649;
												assign node649 = (inp[7]) ? 14'b00000000000000 : 14'b00000000000000;
												assign node652 = (inp[4]) ? 14'b00000000000000 : 14'b00100000000011;
									assign node656 = (inp[2]) ? node670 : node657;
										assign node657 = (inp[0]) ? node665 : node658;
											assign node658 = (inp[13]) ? node662 : node659;
												assign node659 = (inp[4]) ? 14'b10100100101000 : 14'b10100100111000;
												assign node662 = (inp[4]) ? 14'b10000000101000 : 14'b10000000111000;
											assign node665 = (inp[7]) ? node667 : 14'b10000100011000;
												assign node667 = (inp[13]) ? 14'b00001000000100 : 14'b00000000000000;
										assign node670 = (inp[13]) ? 14'b00001000000100 : 14'b00000000000000;
								assign node673 = (inp[13]) ? node689 : node674;
									assign node674 = (inp[12]) ? 14'b00000000000000 : node675;
										assign node675 = (inp[2]) ? node681 : node676;
											assign node676 = (inp[7]) ? 14'b00000000000000 : node677;
												assign node677 = (inp[4]) ? 14'b10000000011101 : 14'b10000001001101;
											assign node681 = (inp[7]) ? node685 : node682;
												assign node682 = (inp[0]) ? 14'b00000000000000 : 14'b00000000000000;
												assign node685 = (inp[0]) ? 14'b00000000000000 : 14'b10000100001101;
									assign node689 = (inp[12]) ? 14'b10000100001000 : node690;
										assign node690 = (inp[0]) ? 14'b10100100011000 : node691;
											assign node691 = (inp[2]) ? node693 : 14'b10000000001010;
												assign node693 = (inp[4]) ? 14'b10100100011000 : 14'b00000000000000;
						assign node698 = (inp[2]) ? node752 : node699;
							assign node699 = (inp[0]) ? node737 : node700;
								assign node700 = (inp[11]) ? node720 : node701;
									assign node701 = (inp[8]) ? node711 : node702;
										assign node702 = (inp[13]) ? node706 : node703;
											assign node703 = (inp[7]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node706 = (inp[7]) ? node708 : 14'b00000000000000;
												assign node708 = (inp[5]) ? 14'b01100000001010 : 14'b00000000000000;
										assign node711 = (inp[4]) ? node717 : node712;
											assign node712 = (inp[13]) ? 14'b00000000000000 : node713;
												assign node713 = (inp[7]) ? 14'b00000000000000 : 14'b00000000000000;
											assign node717 = (inp[13]) ? 14'b00001000001001 : 14'b00000000000000;
									assign node720 = (inp[12]) ? node728 : node721;
										assign node721 = (inp[8]) ? node723 : 14'b00100000000011;
											assign node723 = (inp[7]) ? 14'b00000000000000 : node724;
												assign node724 = (inp[13]) ? 14'b10100100111000 : 14'b00100000001010;
										assign node728 = (inp[8]) ? node734 : node729;
											assign node729 = (inp[5]) ? 14'b00000000000000 : node730;
												assign node730 = (inp[13]) ? 14'b00000000000000 : 14'b00100100001101;
											assign node734 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node737 = (inp[13]) ? node745 : node738;
									assign node738 = (inp[12]) ? 14'b00000000000000 : node739;
										assign node739 = (inp[8]) ? 14'b00000000000000 : node740;
											assign node740 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node745 = (inp[12]) ? node747 : 14'b00000000000000;
										assign node747 = (inp[11]) ? node749 : 14'b00000000000000;
											assign node749 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node752 = (inp[8]) ? node760 : node753;
								assign node753 = (inp[13]) ? 14'b00000000000000 : node754;
									assign node754 = (inp[12]) ? 14'b00000000000000 : node755;
										assign node755 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node760 = (inp[13]) ? node762 : 14'b00000000000000;
									assign node762 = (inp[12]) ? node764 : 14'b00000000000000;
										assign node764 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node767 = (inp[0]) ? node875 : node768;
						assign node768 = (inp[3]) ? node824 : node769;
							assign node769 = (inp[5]) ? node793 : node770;
								assign node770 = (inp[2]) ? node780 : node771;
									assign node771 = (inp[11]) ? 14'b00000000000000 : node772;
										assign node772 = (inp[8]) ? 14'b00000000000000 : node773;
											assign node773 = (inp[12]) ? 14'b00000000000000 : node774;
												assign node774 = (inp[4]) ? 14'b00000000000000 : 14'b00001000000100;
									assign node780 = (inp[4]) ? 14'b00000000000000 : node781;
										assign node781 = (inp[13]) ? node787 : node782;
											assign node782 = (inp[8]) ? 14'b00000000000000 : node783;
												assign node783 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node787 = (inp[8]) ? node789 : 14'b00000000000000;
												assign node789 = (inp[7]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node793 = (inp[7]) ? node807 : node794;
									assign node794 = (inp[8]) ? node800 : node795;
										assign node795 = (inp[12]) ? 14'b00000000000000 : node796;
											assign node796 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
										assign node800 = (inp[2]) ? node802 : 14'b00000000000000;
											assign node802 = (inp[12]) ? node804 : 14'b00000000000000;
												assign node804 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
									assign node807 = (inp[11]) ? node819 : node808;
										assign node808 = (inp[13]) ? node814 : node809;
											assign node809 = (inp[8]) ? 14'b00000000000000 : node810;
												assign node810 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
											assign node814 = (inp[12]) ? 14'b01100000001010 : node815;
												assign node815 = (inp[4]) ? 14'b00001000000100 : 14'b00000000000000;
										assign node819 = (inp[12]) ? node821 : 14'b00000000000000;
											assign node821 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node824 = (inp[2]) ? node860 : node825;
								assign node825 = (inp[7]) ? node841 : node826;
									assign node826 = (inp[8]) ? node832 : node827;
										assign node827 = (inp[12]) ? 14'b00000000000000 : node828;
											assign node828 = (inp[11]) ? 14'b00100000000011 : 14'b00000000000000;
										assign node832 = (inp[11]) ? node836 : node833;
											assign node833 = (inp[13]) ? 14'b00000000000000 : 14'b00000000011100;
											assign node836 = (inp[13]) ? node838 : 14'b00100000001010;
												assign node838 = (inp[12]) ? 14'b10000100001000 : 14'b10100100101000;
									assign node841 = (inp[8]) ? node853 : node842;
										assign node842 = (inp[12]) ? node848 : node843;
											assign node843 = (inp[11]) ? 14'b00000000000000 : node844;
												assign node844 = (inp[13]) ? 14'b00001000000100 : 14'b10000100001000;
											assign node848 = (inp[11]) ? node850 : 14'b01100000001010;
												assign node850 = (inp[4]) ? 14'b00000000000000 : 14'b00100100001101;
										assign node853 = (inp[13]) ? node855 : 14'b00000000000000;
											assign node855 = (inp[12]) ? node857 : 14'b00000000000000;
												assign node857 = (inp[11]) ? 14'b10000100001000 : 14'b00000000000000;
								assign node860 = (inp[13]) ? node868 : node861;
									assign node861 = (inp[11]) ? 14'b00000000000000 : node862;
										assign node862 = (inp[12]) ? 14'b00000000000000 : node863;
											assign node863 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node868 = (inp[11]) ? node870 : 14'b00000000000000;
										assign node870 = (inp[12]) ? node872 : 14'b00000000000000;
											assign node872 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node875 = (inp[7]) ? node891 : node876;
							assign node876 = (inp[11]) ? node884 : node877;
								assign node877 = (inp[13]) ? 14'b00000000000000 : node878;
									assign node878 = (inp[8]) ? 14'b00000000000000 : node879;
										assign node879 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node884 = (inp[12]) ? node886 : 14'b00000000000000;
									assign node886 = (inp[13]) ? node888 : 14'b00000000000000;
										assign node888 = (inp[8]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node891 = (inp[8]) ? node899 : node892;
								assign node892 = (inp[11]) ? 14'b00000000000000 : node893;
									assign node893 = (inp[13]) ? 14'b00000000000000 : node894;
										assign node894 = (inp[12]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node899 = (inp[12]) ? node901 : 14'b00000000000000;
									assign node901 = (inp[11]) ? node903 : 14'b00000000000000;
										assign node903 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
				assign node906 = (inp[9]) ? node972 : node907;
					assign node907 = (inp[3]) ? node941 : node908;
						assign node908 = (inp[13]) ? node924 : node909;
							assign node909 = (inp[11]) ? 14'b00000000000000 : node910;
								assign node910 = (inp[12]) ? node914 : node911;
									assign node911 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
									assign node914 = (inp[5]) ? node916 : 14'b00000000000000;
										assign node916 = (inp[8]) ? 14'b00000000000000 : node917;
											assign node917 = (inp[2]) ? 14'b00000000000000 : node918;
												assign node918 = (inp[4]) ? 14'b00000000000000 : 14'b00000000000000;
							assign node924 = (inp[12]) ? node926 : 14'b00000000000000;
								assign node926 = (inp[8]) ? node938 : node927;
									assign node927 = (inp[2]) ? 14'b00000000000000 : node928;
										assign node928 = (inp[4]) ? 14'b00000000000000 : node929;
											assign node929 = (inp[11]) ? node933 : node930;
												assign node930 = (inp[5]) ? 14'b00000000011100 : 14'b00000000000000;
												assign node933 = (inp[0]) ? 14'b00000000000000 : 14'b01001000000101;
									assign node938 = (inp[11]) ? 14'b10000100001000 : 14'b00000100001110;
						assign node941 = (inp[7]) ? node957 : node942;
							assign node942 = (inp[11]) ? node950 : node943;
								assign node943 = (inp[13]) ? 14'b00000000000000 : node944;
									assign node944 = (inp[12]) ? 14'b00000000000000 : node945;
										assign node945 = (inp[8]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node950 = (inp[8]) ? node952 : 14'b00000000000000;
									assign node952 = (inp[12]) ? node954 : 14'b00000000000000;
										assign node954 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
							assign node957 = (inp[12]) ? node965 : node958;
								assign node958 = (inp[8]) ? 14'b00000000000000 : node959;
									assign node959 = (inp[11]) ? 14'b00000000000000 : node960;
										assign node960 = (inp[13]) ? 14'b00000000000000 : 14'b10000100001000;
								assign node965 = (inp[8]) ? node967 : 14'b00000000000000;
									assign node967 = (inp[11]) ? node969 : 14'b00000000000000;
										assign node969 = (inp[13]) ? 14'b10000100001000 : 14'b00000000000000;
					assign node972 = (inp[3]) ? node988 : node973;
						assign node973 = (inp[13]) ? node981 : node974;
							assign node974 = (inp[12]) ? 14'b00000000000000 : node975;
								assign node975 = (inp[8]) ? 14'b00000000000000 : node976;
									assign node976 = (inp[11]) ? 14'b00000000000000 : 14'b10000100001000;
							assign node981 = (inp[11]) ? node983 : 14'b00000000000000;
								assign node983 = (inp[8]) ? node985 : 14'b00000000000000;
									assign node985 = (inp[12]) ? 14'b10000100001000 : 14'b00000000000000;
						assign node988 = (inp[11]) ? node1026 : node989;
							assign node989 = (inp[12]) ? node1009 : node990;
								assign node990 = (inp[13]) ? node1000 : node991;
									assign node991 = (inp[8]) ? node993 : 14'b10000100001000;
										assign node993 = (inp[7]) ? node995 : 14'b00000000000000;
											assign node995 = (inp[0]) ? 14'b10100000001000 : node996;
												assign node996 = (inp[2]) ? 14'b10010010001101 : 14'b00100000001010;
									assign node1000 = (inp[0]) ? 14'b00000000000000 : node1001;
										assign node1001 = (inp[5]) ? 14'b00000000000000 : node1002;
											assign node1002 = (inp[8]) ? node1004 : 14'b00000000011101;
												assign node1004 = (inp[7]) ? 14'b10100000001000 : 14'b00000000000000;
								assign node1009 = (inp[5]) ? node1011 : 14'b00000000000000;
									assign node1011 = (inp[2]) ? node1017 : node1012;
										assign node1012 = (inp[7]) ? node1014 : 14'b00000000000000;
											assign node1014 = (inp[8]) ? 14'b00000000011100 : 14'b00000000000000;
										assign node1017 = (inp[8]) ? node1023 : node1018;
											assign node1018 = (inp[7]) ? 14'b00000000000000 : node1019;
												assign node1019 = (inp[13]) ? 14'b10100000001000 : 14'b00001000001100;
											assign node1023 = (inp[7]) ? 14'b01100000000110 : 14'b00000000000000;
							assign node1026 = (inp[13]) ? node1040 : node1027;
								assign node1027 = (inp[7]) ? node1035 : node1028;
									assign node1028 = (inp[12]) ? node1030 : 14'b00000000000000;
										assign node1030 = (inp[5]) ? node1032 : 14'b00000000000000;
											assign node1032 = (inp[8]) ? 14'b00000000000000 : 14'b00000100001111;
									assign node1035 = (inp[12]) ? 14'b00000000000000 : node1036;
										assign node1036 = (inp[5]) ? 14'b00000000000000 : 14'b01001000000100;
								assign node1040 = (inp[12]) ? node1054 : node1041;
									assign node1041 = (inp[7]) ? node1043 : 14'b00000000000000;
										assign node1043 = (inp[5]) ? node1051 : node1044;
											assign node1044 = (inp[0]) ? node1048 : node1045;
												assign node1045 = (inp[2]) ? 14'b00100100001101 : 14'b00001000001001;
												assign node1048 = (inp[8]) ? 14'b00100100001101 : 14'b01000100000010;
											assign node1051 = (inp[8]) ? 14'b00000000000000 : 14'b10100101111111;
									assign node1054 = (inp[8]) ? 14'b10000100001000 : node1055;
										assign node1055 = (inp[5]) ? node1057 : 14'b00000000000000;
											assign node1057 = (inp[7]) ? 14'b00000000000000 : 14'b10100100001000;

endmodule