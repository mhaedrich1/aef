module dtc_split875_bm90 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node50;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node70;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node89;
	wire [3-1:0] node92;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node110;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node115;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node131;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node189;
	wire [3-1:0] node190;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node226;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node251;
	wire [3-1:0] node252;
	wire [3-1:0] node253;
	wire [3-1:0] node254;
	wire [3-1:0] node258;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node266;
	wire [3-1:0] node267;
	wire [3-1:0] node270;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node281;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node288;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node310;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node324;
	wire [3-1:0] node327;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node332;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node346;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node354;
	wire [3-1:0] node357;
	wire [3-1:0] node358;
	wire [3-1:0] node360;
	wire [3-1:0] node364;
	wire [3-1:0] node365;
	wire [3-1:0] node366;
	wire [3-1:0] node367;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node375;
	wire [3-1:0] node378;
	wire [3-1:0] node379;
	wire [3-1:0] node380;
	wire [3-1:0] node383;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node390;

	assign outp = (inp[0]) ? node156 : node1;
		assign node1 = (inp[6]) ? node31 : node2;
			assign node2 = (inp[3]) ? node14 : node3;
				assign node3 = (inp[4]) ? node5 : 3'b011;
					assign node5 = (inp[7]) ? node7 : 3'b011;
						assign node7 = (inp[1]) ? node9 : 3'b111;
							assign node9 = (inp[8]) ? node11 : 3'b111;
								assign node11 = (inp[2]) ? 3'b011 : 3'b111;
				assign node14 = (inp[9]) ? 3'b111 : node15;
					assign node15 = (inp[7]) ? node17 : 3'b111;
						assign node17 = (inp[1]) ? node23 : node18;
							assign node18 = (inp[2]) ? node20 : 3'b111;
								assign node20 = (inp[4]) ? 3'b111 : 3'b011;
							assign node23 = (inp[4]) ? node27 : node24;
								assign node24 = (inp[8]) ? 3'b001 : 3'b101;
								assign node27 = (inp[8]) ? 3'b011 : 3'b111;
			assign node31 = (inp[7]) ? node95 : node32;
				assign node32 = (inp[3]) ? node64 : node33;
					assign node33 = (inp[4]) ? node49 : node34;
						assign node34 = (inp[2]) ? node42 : node35;
							assign node35 = (inp[9]) ? node39 : node36;
								assign node36 = (inp[10]) ? 3'b101 : 3'b001;
								assign node39 = (inp[5]) ? 3'b001 : 3'b001;
							assign node42 = (inp[1]) ? node46 : node43;
								assign node43 = (inp[10]) ? 3'b001 : 3'b101;
								assign node46 = (inp[8]) ? 3'b110 : 3'b101;
						assign node49 = (inp[9]) ? node57 : node50;
							assign node50 = (inp[1]) ? node54 : node51;
								assign node51 = (inp[2]) ? 3'b001 : 3'b101;
								assign node54 = (inp[10]) ? 3'b001 : 3'b111;
							assign node57 = (inp[1]) ? node61 : node58;
								assign node58 = (inp[2]) ? 3'b011 : 3'b111;
								assign node61 = (inp[2]) ? 3'b101 : 3'b011;
					assign node64 = (inp[1]) ? node80 : node65;
						assign node65 = (inp[5]) ? node73 : node66;
							assign node66 = (inp[8]) ? node70 : node67;
								assign node67 = (inp[11]) ? 3'b111 : 3'b111;
								assign node70 = (inp[4]) ? 3'b101 : 3'b111;
							assign node73 = (inp[9]) ? node77 : node74;
								assign node74 = (inp[4]) ? 3'b111 : 3'b011;
								assign node77 = (inp[11]) ? 3'b111 : 3'b111;
						assign node80 = (inp[9]) ? node88 : node81;
							assign node81 = (inp[4]) ? node85 : node82;
								assign node82 = (inp[5]) ? 3'b001 : 3'b100;
								assign node85 = (inp[2]) ? 3'b101 : 3'b001;
							assign node88 = (inp[4]) ? node92 : node89;
								assign node89 = (inp[2]) ? 3'b001 : 3'b111;
								assign node92 = (inp[2]) ? 3'b111 : 3'b111;
				assign node95 = (inp[3]) ? node125 : node96;
					assign node96 = (inp[9]) ? node110 : node97;
						assign node97 = (inp[4]) ? node103 : node98;
							assign node98 = (inp[1]) ? 3'b000 : node99;
								assign node99 = (inp[2]) ? 3'b000 : 3'b000;
							assign node103 = (inp[1]) ? node107 : node104;
								assign node104 = (inp[2]) ? 3'b010 : 3'b111;
								assign node107 = (inp[10]) ? 3'b000 : 3'b000;
						assign node110 = (inp[1]) ? node118 : node111;
							assign node111 = (inp[4]) ? node115 : node112;
								assign node112 = (inp[2]) ? 3'b000 : 3'b101;
								assign node115 = (inp[10]) ? 3'b011 : 3'b101;
							assign node118 = (inp[5]) ? node122 : node119;
								assign node119 = (inp[2]) ? 3'b100 : 3'b010;
								assign node122 = (inp[8]) ? 3'b110 : 3'b001;
					assign node125 = (inp[1]) ? node141 : node126;
						assign node126 = (inp[9]) ? node134 : node127;
							assign node127 = (inp[2]) ? node131 : node128;
								assign node128 = (inp[4]) ? 3'b111 : 3'b001;
								assign node131 = (inp[4]) ? 3'b001 : 3'b010;
							assign node134 = (inp[4]) ? node138 : node135;
								assign node135 = (inp[10]) ? 3'b111 : 3'b011;
								assign node138 = (inp[10]) ? 3'b111 : 3'b111;
						assign node141 = (inp[9]) ? node149 : node142;
							assign node142 = (inp[2]) ? node146 : node143;
								assign node143 = (inp[4]) ? 3'b001 : 3'b010;
								assign node146 = (inp[10]) ? 3'b010 : 3'b110;
							assign node149 = (inp[4]) ? node153 : node150;
								assign node150 = (inp[10]) ? 3'b001 : 3'b110;
								assign node153 = (inp[2]) ? 3'b101 : 3'b111;
		assign node156 = (inp[6]) ? node280 : node157;
			assign node157 = (inp[3]) ? node219 : node158;
				assign node158 = (inp[4]) ? node188 : node159;
					assign node159 = (inp[9]) ? node175 : node160;
						assign node160 = (inp[7]) ? node168 : node161;
							assign node161 = (inp[1]) ? node165 : node162;
								assign node162 = (inp[2]) ? 3'b110 : 3'b010;
								assign node165 = (inp[2]) ? 3'b110 : 3'b000;
							assign node168 = (inp[1]) ? node172 : node169;
								assign node169 = (inp[2]) ? 3'b000 : 3'b100;
								assign node172 = (inp[10]) ? 3'b010 : 3'b110;
						assign node175 = (inp[1]) ? node181 : node176;
							assign node176 = (inp[7]) ? node178 : 3'b110;
								assign node178 = (inp[2]) ? 3'b010 : 3'b110;
							assign node181 = (inp[7]) ? node185 : node182;
								assign node182 = (inp[5]) ? 3'b110 : 3'b010;
								assign node185 = (inp[2]) ? 3'b100 : 3'b110;
					assign node188 = (inp[1]) ? node204 : node189;
						assign node189 = (inp[7]) ? node197 : node190;
							assign node190 = (inp[5]) ? node194 : node191;
								assign node191 = (inp[9]) ? 3'b001 : 3'b000;
								assign node194 = (inp[11]) ? 3'b110 : 3'b110;
							assign node197 = (inp[2]) ? node201 : node198;
								assign node198 = (inp[8]) ? 3'b101 : 3'b111;
								assign node201 = (inp[5]) ? 3'b101 : 3'b001;
						assign node204 = (inp[9]) ? node212 : node205;
							assign node205 = (inp[7]) ? node209 : node206;
								assign node206 = (inp[2]) ? 3'b001 : 3'b001;
								assign node209 = (inp[2]) ? 3'b000 : 3'b000;
							assign node212 = (inp[7]) ? node216 : node213;
								assign node213 = (inp[11]) ? 3'b110 : 3'b001;
								assign node216 = (inp[2]) ? 3'b010 : 3'b110;
				assign node219 = (inp[9]) ? node251 : node220;
					assign node220 = (inp[1]) ? node236 : node221;
						assign node221 = (inp[7]) ? node229 : node222;
							assign node222 = (inp[4]) ? node226 : node223;
								assign node223 = (inp[10]) ? 3'b111 : 3'b111;
								assign node226 = (inp[2]) ? 3'b101 : 3'b111;
							assign node229 = (inp[4]) ? node233 : node230;
								assign node230 = (inp[2]) ? 3'b110 : 3'b000;
								assign node233 = (inp[8]) ? 3'b101 : 3'b001;
						assign node236 = (inp[4]) ? node244 : node237;
							assign node237 = (inp[8]) ? node241 : node238;
								assign node238 = (inp[7]) ? 3'b010 : 3'b010;
								assign node241 = (inp[5]) ? 3'b010 : 3'b000;
							assign node244 = (inp[7]) ? node248 : node245;
								assign node245 = (inp[2]) ? 3'b010 : 3'b001;
								assign node248 = (inp[10]) ? 3'b000 : 3'b110;
					assign node251 = (inp[7]) ? node265 : node252;
						assign node252 = (inp[1]) ? node258 : node253;
							assign node253 = (inp[4]) ? 3'b111 : node254;
								assign node254 = (inp[10]) ? 3'b111 : 3'b111;
							assign node258 = (inp[2]) ? node262 : node259;
								assign node259 = (inp[4]) ? 3'b111 : 3'b011;
								assign node262 = (inp[4]) ? 3'b011 : 3'b001;
						assign node265 = (inp[1]) ? node273 : node266;
							assign node266 = (inp[4]) ? node270 : node267;
								assign node267 = (inp[10]) ? 3'b011 : 3'b101;
								assign node270 = (inp[2]) ? 3'b011 : 3'b111;
							assign node273 = (inp[10]) ? node277 : node274;
								assign node274 = (inp[4]) ? 3'b101 : 3'b010;
								assign node277 = (inp[4]) ? 3'b001 : 3'b001;
			assign node280 = (inp[1]) ? node342 : node281;
				assign node281 = (inp[7]) ? node313 : node282;
					assign node282 = (inp[3]) ? node298 : node283;
						assign node283 = (inp[4]) ? node291 : node284;
							assign node284 = (inp[2]) ? node288 : node285;
								assign node285 = (inp[10]) ? 3'b010 : 3'b010;
								assign node288 = (inp[5]) ? 3'b000 : 3'b100;
							assign node291 = (inp[2]) ? node295 : node292;
								assign node292 = (inp[5]) ? 3'b100 : 3'b100;
								assign node295 = (inp[8]) ? 3'b110 : 3'b110;
						assign node298 = (inp[9]) ? node306 : node299;
							assign node299 = (inp[2]) ? node303 : node300;
								assign node300 = (inp[4]) ? 3'b010 : 3'b010;
								assign node303 = (inp[4]) ? 3'b010 : 3'b100;
							assign node306 = (inp[4]) ? node310 : node307;
								assign node307 = (inp[2]) ? 3'b100 : 3'b001;
								assign node310 = (inp[2]) ? 3'b101 : 3'b101;
					assign node313 = (inp[3]) ? node327 : node314;
						assign node314 = (inp[2]) ? node322 : node315;
							assign node315 = (inp[9]) ? node319 : node316;
								assign node316 = (inp[10]) ? 3'b000 : 3'b000;
								assign node319 = (inp[4]) ? 3'b100 : 3'b000;
							assign node322 = (inp[9]) ? node324 : 3'b000;
								assign node324 = (inp[8]) ? 3'b000 : 3'b000;
						assign node327 = (inp[9]) ? node335 : node328;
							assign node328 = (inp[4]) ? node332 : node329;
								assign node329 = (inp[10]) ? 3'b000 : 3'b000;
								assign node332 = (inp[10]) ? 3'b010 : 3'b100;
							assign node335 = (inp[2]) ? node339 : node336;
								assign node336 = (inp[8]) ? 3'b110 : 3'b101;
								assign node339 = (inp[4]) ? 3'b010 : 3'b100;
				assign node342 = (inp[3]) ? node364 : node343;
					assign node343 = (inp[7]) ? node357 : node344;
						assign node344 = (inp[2]) ? node352 : node345;
							assign node345 = (inp[4]) ? node349 : node346;
								assign node346 = (inp[8]) ? 3'b000 : 3'b000;
								assign node349 = (inp[10]) ? 3'b000 : 3'b000;
							assign node352 = (inp[4]) ? node354 : 3'b000;
								assign node354 = (inp[8]) ? 3'b000 : 3'b000;
						assign node357 = (inp[2]) ? 3'b000 : node358;
							assign node358 = (inp[9]) ? node360 : 3'b000;
								assign node360 = (inp[5]) ? 3'b000 : 3'b000;
					assign node364 = (inp[9]) ? node378 : node365;
						assign node365 = (inp[4]) ? node371 : node366;
							assign node366 = (inp[8]) ? 3'b000 : node367;
								assign node367 = (inp[2]) ? 3'b000 : 3'b000;
							assign node371 = (inp[7]) ? node375 : node372;
								assign node372 = (inp[8]) ? 3'b000 : 3'b010;
								assign node375 = (inp[10]) ? 3'b000 : 3'b000;
						assign node378 = (inp[7]) ? node386 : node379;
							assign node379 = (inp[2]) ? node383 : node380;
								assign node380 = (inp[4]) ? 3'b001 : 3'b010;
								assign node383 = (inp[4]) ? 3'b110 : 3'b100;
							assign node386 = (inp[4]) ? node390 : node387;
								assign node387 = (inp[10]) ? 3'b000 : 3'b000;
								assign node390 = (inp[10]) ? 3'b010 : 3'b000;

endmodule