module dtc_split875_bm75 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node12;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node20;
	wire [3-1:0] node21;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node38;
	wire [3-1:0] node41;
	wire [3-1:0] node44;
	wire [3-1:0] node45;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node56;
	wire [3-1:0] node59;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node88;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node96;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node101;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node117;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node144;
	wire [3-1:0] node147;
	wire [3-1:0] node148;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node153;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node174;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node201;
	wire [3-1:0] node202;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node213;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node233;
	wire [3-1:0] node234;
	wire [3-1:0] node237;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node242;
	wire [3-1:0] node245;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node257;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node271;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node316;
	wire [3-1:0] node319;
	wire [3-1:0] node320;
	wire [3-1:0] node321;
	wire [3-1:0] node322;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node329;
	wire [3-1:0] node332;
	wire [3-1:0] node335;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node340;
	wire [3-1:0] node343;
	wire [3-1:0] node344;
	wire [3-1:0] node347;
	wire [3-1:0] node350;
	wire [3-1:0] node351;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node354;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node364;
	wire [3-1:0] node367;
	wire [3-1:0] node369;
	wire [3-1:0] node372;
	wire [3-1:0] node373;
	wire [3-1:0] node374;
	wire [3-1:0] node375;
	wire [3-1:0] node378;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node388;
	wire [3-1:0] node391;
	wire [3-1:0] node394;
	wire [3-1:0] node395;
	wire [3-1:0] node398;
	wire [3-1:0] node401;
	wire [3-1:0] node402;
	wire [3-1:0] node403;
	wire [3-1:0] node404;
	wire [3-1:0] node405;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node426;
	wire [3-1:0] node429;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node436;
	wire [3-1:0] node437;
	wire [3-1:0] node438;
	wire [3-1:0] node439;
	wire [3-1:0] node442;
	wire [3-1:0] node445;
	wire [3-1:0] node446;
	wire [3-1:0] node449;
	wire [3-1:0] node452;
	wire [3-1:0] node453;
	wire [3-1:0] node454;
	wire [3-1:0] node457;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node467;
	wire [3-1:0] node468;
	wire [3-1:0] node469;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node479;
	wire [3-1:0] node482;
	wire [3-1:0] node483;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node490;
	wire [3-1:0] node491;
	wire [3-1:0] node494;
	wire [3-1:0] node497;
	wire [3-1:0] node498;
	wire [3-1:0] node499;
	wire [3-1:0] node500;
	wire [3-1:0] node503;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node510;
	wire [3-1:0] node513;
	wire [3-1:0] node514;
	wire [3-1:0] node515;
	wire [3-1:0] node518;
	wire [3-1:0] node521;
	wire [3-1:0] node522;
	wire [3-1:0] node525;
	wire [3-1:0] node528;
	wire [3-1:0] node529;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node533;
	wire [3-1:0] node536;
	wire [3-1:0] node539;
	wire [3-1:0] node540;
	wire [3-1:0] node543;
	wire [3-1:0] node546;
	wire [3-1:0] node547;
	wire [3-1:0] node548;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node558;
	wire [3-1:0] node561;
	wire [3-1:0] node562;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node567;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node582;
	wire [3-1:0] node585;
	wire [3-1:0] node586;
	wire [3-1:0] node589;
	wire [3-1:0] node592;
	wire [3-1:0] node593;
	wire [3-1:0] node594;
	wire [3-1:0] node595;
	wire [3-1:0] node596;
	wire [3-1:0] node601;
	wire [3-1:0] node602;
	wire [3-1:0] node603;
	wire [3-1:0] node606;
	wire [3-1:0] node609;
	wire [3-1:0] node610;
	wire [3-1:0] node614;
	wire [3-1:0] node615;
	wire [3-1:0] node616;
	wire [3-1:0] node617;
	wire [3-1:0] node620;
	wire [3-1:0] node623;
	wire [3-1:0] node624;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node637;
	wire [3-1:0] node640;
	wire [3-1:0] node643;
	wire [3-1:0] node644;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node647;
	wire [3-1:0] node648;
	wire [3-1:0] node649;
	wire [3-1:0] node652;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node663;
	wire [3-1:0] node664;
	wire [3-1:0] node667;
	wire [3-1:0] node670;
	wire [3-1:0] node672;
	wire [3-1:0] node675;
	wire [3-1:0] node676;
	wire [3-1:0] node677;
	wire [3-1:0] node678;
	wire [3-1:0] node681;
	wire [3-1:0] node684;
	wire [3-1:0] node685;
	wire [3-1:0] node688;
	wire [3-1:0] node691;
	wire [3-1:0] node692;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node701;
	wire [3-1:0] node704;
	wire [3-1:0] node705;
	wire [3-1:0] node706;
	wire [3-1:0] node707;
	wire [3-1:0] node708;
	wire [3-1:0] node711;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node718;
	wire [3-1:0] node721;
	wire [3-1:0] node722;
	wire [3-1:0] node723;
	wire [3-1:0] node726;
	wire [3-1:0] node729;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node736;
	wire [3-1:0] node737;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node743;
	wire [3-1:0] node744;
	wire [3-1:0] node747;
	wire [3-1:0] node750;
	wire [3-1:0] node751;
	wire [3-1:0] node752;
	wire [3-1:0] node755;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node766;
	wire [3-1:0] node767;
	wire [3-1:0] node768;
	wire [3-1:0] node769;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node776;
	wire [3-1:0] node777;
	wire [3-1:0] node780;
	wire [3-1:0] node783;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node788;
	wire [3-1:0] node791;
	wire [3-1:0] node792;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node800;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node807;
	wire [3-1:0] node808;
	wire [3-1:0] node811;
	wire [3-1:0] node814;
	wire [3-1:0] node815;
	wire [3-1:0] node816;
	wire [3-1:0] node819;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node826;
	wire [3-1:0] node829;
	wire [3-1:0] node830;
	wire [3-1:0] node831;
	wire [3-1:0] node832;
	wire [3-1:0] node833;
	wire [3-1:0] node836;
	wire [3-1:0] node839;
	wire [3-1:0] node840;
	wire [3-1:0] node843;
	wire [3-1:0] node846;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node851;
	wire [3-1:0] node854;
	wire [3-1:0] node855;
	wire [3-1:0] node858;
	wire [3-1:0] node861;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node867;
	wire [3-1:0] node870;
	wire [3-1:0] node871;
	wire [3-1:0] node874;
	wire [3-1:0] node877;
	wire [3-1:0] node878;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node885;
	wire [3-1:0] node886;
	wire [3-1:0] node889;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node895;
	wire [3-1:0] node896;
	wire [3-1:0] node897;
	wire [3-1:0] node898;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node903;
	wire [3-1:0] node906;
	wire [3-1:0] node907;
	wire [3-1:0] node910;
	wire [3-1:0] node913;
	wire [3-1:0] node914;
	wire [3-1:0] node915;
	wire [3-1:0] node918;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node925;
	wire [3-1:0] node928;
	wire [3-1:0] node929;
	wire [3-1:0] node930;
	wire [3-1:0] node931;
	wire [3-1:0] node934;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node942;
	wire [3-1:0] node943;
	wire [3-1:0] node944;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node952;
	wire [3-1:0] node955;
	wire [3-1:0] node956;
	wire [3-1:0] node957;
	wire [3-1:0] node958;
	wire [3-1:0] node959;
	wire [3-1:0] node962;
	wire [3-1:0] node965;
	wire [3-1:0] node966;
	wire [3-1:0] node969;
	wire [3-1:0] node972;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node977;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node984;
	wire [3-1:0] node987;
	wire [3-1:0] node988;
	wire [3-1:0] node989;
	wire [3-1:0] node990;
	wire [3-1:0] node993;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1005;
	wire [3-1:0] node1008;
	wire [3-1:0] node1011;
	wire [3-1:0] node1012;
	wire [3-1:0] node1015;
	wire [3-1:0] node1018;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1026;
	wire [3-1:0] node1029;
	wire [3-1:0] node1030;
	wire [3-1:0] node1033;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1038;
	wire [3-1:0] node1041;
	wire [3-1:0] node1044;
	wire [3-1:0] node1045;
	wire [3-1:0] node1048;
	wire [3-1:0] node1051;
	wire [3-1:0] node1052;
	wire [3-1:0] node1053;
	wire [3-1:0] node1054;
	wire [3-1:0] node1057;
	wire [3-1:0] node1060;
	wire [3-1:0] node1061;
	wire [3-1:0] node1064;
	wire [3-1:0] node1067;
	wire [3-1:0] node1068;
	wire [3-1:0] node1069;
	wire [3-1:0] node1072;
	wire [3-1:0] node1075;
	wire [3-1:0] node1076;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1082;
	wire [3-1:0] node1083;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1090;
	wire [3-1:0] node1091;
	wire [3-1:0] node1094;
	wire [3-1:0] node1097;
	wire [3-1:0] node1098;
	wire [3-1:0] node1099;
	wire [3-1:0] node1102;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1109;
	wire [3-1:0] node1112;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1115;
	wire [3-1:0] node1118;
	wire [3-1:0] node1121;
	wire [3-1:0] node1122;
	wire [3-1:0] node1125;
	wire [3-1:0] node1128;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1133;
	wire [3-1:0] node1136;
	wire [3-1:0] node1137;
	wire [3-1:0] node1140;
	wire [3-1:0] node1143;
	wire [3-1:0] node1144;
	wire [3-1:0] node1145;
	wire [3-1:0] node1146;
	wire [3-1:0] node1147;
	wire [3-1:0] node1148;
	wire [3-1:0] node1150;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1157;
	wire [3-1:0] node1160;
	wire [3-1:0] node1161;
	wire [3-1:0] node1163;
	wire [3-1:0] node1168;
	wire [3-1:0] node1169;
	wire [3-1:0] node1170;
	wire [3-1:0] node1171;
	wire [3-1:0] node1172;
	wire [3-1:0] node1175;
	wire [3-1:0] node1178;
	wire [3-1:0] node1179;
	wire [3-1:0] node1182;
	wire [3-1:0] node1185;
	wire [3-1:0] node1186;
	wire [3-1:0] node1188;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1195;
	wire [3-1:0] node1198;
	wire [3-1:0] node1199;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1204;
	wire [3-1:0] node1207;
	wire [3-1:0] node1209;
	wire [3-1:0] node1212;
	wire [3-1:0] node1214;
	wire [3-1:0] node1216;
	wire [3-1:0] node1219;
	wire [3-1:0] node1220;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1224;
	wire [3-1:0] node1227;
	wire [3-1:0] node1230;
	wire [3-1:0] node1231;
	wire [3-1:0] node1235;
	wire [3-1:0] node1236;
	wire [3-1:0] node1237;
	wire [3-1:0] node1240;
	wire [3-1:0] node1243;
	wire [3-1:0] node1244;
	wire [3-1:0] node1247;
	wire [3-1:0] node1250;
	wire [3-1:0] node1251;
	wire [3-1:0] node1252;
	wire [3-1:0] node1254;
	wire [3-1:0] node1257;
	wire [3-1:0] node1258;
	wire [3-1:0] node1261;
	wire [3-1:0] node1264;
	wire [3-1:0] node1266;
	wire [3-1:0] node1268;
	wire [3-1:0] node1271;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1275;
	wire [3-1:0] node1278;
	wire [3-1:0] node1281;
	wire [3-1:0] node1282;
	wire [3-1:0] node1285;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1293;
	wire [3-1:0] node1296;
	wire [3-1:0] node1297;
	wire [3-1:0] node1300;
	wire [3-1:0] node1303;
	wire [3-1:0] node1304;
	wire [3-1:0] node1305;
	wire [3-1:0] node1306;
	wire [3-1:0] node1310;
	wire [3-1:0] node1311;
	wire [3-1:0] node1314;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1319;
	wire [3-1:0] node1322;
	wire [3-1:0] node1325;
	wire [3-1:0] node1326;
	wire [3-1:0] node1329;
	wire [3-1:0] node1332;
	wire [3-1:0] node1333;
	wire [3-1:0] node1334;
	wire [3-1:0] node1335;
	wire [3-1:0] node1336;
	wire [3-1:0] node1337;
	wire [3-1:0] node1339;
	wire [3-1:0] node1341;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1346;
	wire [3-1:0] node1349;
	wire [3-1:0] node1352;
	wire [3-1:0] node1354;
	wire [3-1:0] node1357;
	wire [3-1:0] node1358;
	wire [3-1:0] node1359;
	wire [3-1:0] node1361;
	wire [3-1:0] node1366;
	wire [3-1:0] node1367;
	wire [3-1:0] node1368;
	wire [3-1:0] node1369;
	wire [3-1:0] node1370;
	wire [3-1:0] node1373;
	wire [3-1:0] node1376;
	wire [3-1:0] node1377;
	wire [3-1:0] node1380;
	wire [3-1:0] node1383;
	wire [3-1:0] node1384;
	wire [3-1:0] node1386;
	wire [3-1:0] node1389;
	wire [3-1:0] node1390;
	wire [3-1:0] node1393;
	wire [3-1:0] node1396;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1400;
	wire [3-1:0] node1403;
	wire [3-1:0] node1404;
	wire [3-1:0] node1407;
	wire [3-1:0] node1410;
	wire [3-1:0] node1412;
	wire [3-1:0] node1414;
	wire [3-1:0] node1417;
	wire [3-1:0] node1418;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1421;
	wire [3-1:0] node1422;
	wire [3-1:0] node1425;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1432;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1440;
	wire [3-1:0] node1443;
	wire [3-1:0] node1444;
	wire [3-1:0] node1447;
	wire [3-1:0] node1450;
	wire [3-1:0] node1451;
	wire [3-1:0] node1452;
	wire [3-1:0] node1453;
	wire [3-1:0] node1456;
	wire [3-1:0] node1459;
	wire [3-1:0] node1460;
	wire [3-1:0] node1463;
	wire [3-1:0] node1466;
	wire [3-1:0] node1468;
	wire [3-1:0] node1470;
	wire [3-1:0] node1473;
	wire [3-1:0] node1474;
	wire [3-1:0] node1475;
	wire [3-1:0] node1476;
	wire [3-1:0] node1477;
	wire [3-1:0] node1480;
	wire [3-1:0] node1483;
	wire [3-1:0] node1484;
	wire [3-1:0] node1487;
	wire [3-1:0] node1490;
	wire [3-1:0] node1491;
	wire [3-1:0] node1492;
	wire [3-1:0] node1495;
	wire [3-1:0] node1498;
	wire [3-1:0] node1499;
	wire [3-1:0] node1502;
	wire [3-1:0] node1505;
	wire [3-1:0] node1506;
	wire [3-1:0] node1507;
	wire [3-1:0] node1508;
	wire [3-1:0] node1511;
	wire [3-1:0] node1514;
	wire [3-1:0] node1515;
	wire [3-1:0] node1518;
	wire [3-1:0] node1521;
	wire [3-1:0] node1522;
	wire [3-1:0] node1523;
	wire [3-1:0] node1526;
	wire [3-1:0] node1529;
	wire [3-1:0] node1530;
	wire [3-1:0] node1533;
	wire [3-1:0] node1536;
	wire [3-1:0] node1537;
	wire [3-1:0] node1538;
	wire [3-1:0] node1539;
	wire [3-1:0] node1541;
	wire [3-1:0] node1543;
	wire [3-1:0] node1545;
	wire [3-1:0] node1550;
	wire [3-1:0] node1551;
	wire [3-1:0] node1552;
	wire [3-1:0] node1554;
	wire [3-1:0] node1556;
	wire [3-1:0] node1557;
	wire [3-1:0] node1562;
	wire [3-1:0] node1563;
	wire [3-1:0] node1564;
	wire [3-1:0] node1565;
	wire [3-1:0] node1566;
	wire [3-1:0] node1569;
	wire [3-1:0] node1572;
	wire [3-1:0] node1573;
	wire [3-1:0] node1576;
	wire [3-1:0] node1579;
	wire [3-1:0] node1580;
	wire [3-1:0] node1581;
	wire [3-1:0] node1585;
	wire [3-1:0] node1586;
	wire [3-1:0] node1589;
	wire [3-1:0] node1592;
	wire [3-1:0] node1593;
	wire [3-1:0] node1595;
	wire [3-1:0] node1597;
	wire [3-1:0] node1600;
	wire [3-1:0] node1601;
	wire [3-1:0] node1602;
	wire [3-1:0] node1606;
	wire [3-1:0] node1607;
	wire [3-1:0] node1610;

	assign outp = (inp[3]) ? node892 : node1;
		assign node1 = (inp[9]) ? node401 : node2;
			assign node2 = (inp[4]) ? node158 : node3;
				assign node3 = (inp[6]) ? node111 : node4;
					assign node4 = (inp[0]) ? node66 : node5;
						assign node5 = (inp[10]) ? node35 : node6;
							assign node6 = (inp[5]) ? node20 : node7;
								assign node7 = (inp[7]) ? node15 : node8;
									assign node8 = (inp[1]) ? node12 : node9;
										assign node9 = (inp[11]) ? 3'b011 : 3'b011;
										assign node12 = (inp[2]) ? 3'b111 : 3'b011;
									assign node15 = (inp[1]) ? 3'b111 : node16;
										assign node16 = (inp[11]) ? 3'b011 : 3'b111;
								assign node20 = (inp[7]) ? node28 : node21;
									assign node21 = (inp[1]) ? node25 : node22;
										assign node22 = (inp[11]) ? 3'b001 : 3'b101;
										assign node25 = (inp[11]) ? 3'b101 : 3'b011;
									assign node28 = (inp[1]) ? node32 : node29;
										assign node29 = (inp[2]) ? 3'b011 : 3'b101;
										assign node32 = (inp[11]) ? 3'b011 : 3'b111;
							assign node35 = (inp[5]) ? node51 : node36;
								assign node36 = (inp[1]) ? node44 : node37;
									assign node37 = (inp[8]) ? node41 : node38;
										assign node38 = (inp[11]) ? 3'b101 : 3'b101;
										assign node41 = (inp[7]) ? 3'b011 : 3'b101;
									assign node44 = (inp[8]) ? node48 : node45;
										assign node45 = (inp[7]) ? 3'b011 : 3'b101;
										assign node48 = (inp[7]) ? 3'b111 : 3'b011;
								assign node51 = (inp[1]) ? node59 : node52;
									assign node52 = (inp[11]) ? node56 : node53;
										assign node53 = (inp[7]) ? 3'b101 : 3'b001;
										assign node56 = (inp[7]) ? 3'b001 : 3'b110;
									assign node59 = (inp[7]) ? node63 : node60;
										assign node60 = (inp[8]) ? 3'b101 : 3'b001;
										assign node63 = (inp[8]) ? 3'b001 : 3'b101;
						assign node66 = (inp[10]) ? node82 : node67;
							assign node67 = (inp[5]) ? node69 : 3'b111;
								assign node69 = (inp[1]) ? node77 : node70;
									assign node70 = (inp[7]) ? node74 : node71;
										assign node71 = (inp[11]) ? 3'b011 : 3'b111;
										assign node74 = (inp[8]) ? 3'b111 : 3'b111;
									assign node77 = (inp[2]) ? 3'b111 : node78;
										assign node78 = (inp[8]) ? 3'b111 : 3'b111;
							assign node82 = (inp[5]) ? node96 : node83;
								assign node83 = (inp[1]) ? node91 : node84;
									assign node84 = (inp[7]) ? node88 : node85;
										assign node85 = (inp[11]) ? 3'b011 : 3'b011;
										assign node88 = (inp[2]) ? 3'b111 : 3'b111;
									assign node91 = (inp[8]) ? 3'b111 : node92;
										assign node92 = (inp[2]) ? 3'b111 : 3'b011;
								assign node96 = (inp[7]) ? node104 : node97;
									assign node97 = (inp[1]) ? node101 : node98;
										assign node98 = (inp[11]) ? 3'b101 : 3'b101;
										assign node101 = (inp[2]) ? 3'b011 : 3'b011;
									assign node104 = (inp[11]) ? node108 : node105;
										assign node105 = (inp[1]) ? 3'b111 : 3'b011;
										assign node108 = (inp[2]) ? 3'b011 : 3'b011;
					assign node111 = (inp[0]) ? node147 : node112;
						assign node112 = (inp[10]) ? node122 : node113;
							assign node113 = (inp[7]) ? 3'b111 : node114;
								assign node114 = (inp[5]) ? node116 : 3'b111;
									assign node116 = (inp[1]) ? 3'b111 : node117;
										assign node117 = (inp[8]) ? 3'b111 : 3'b011;
							assign node122 = (inp[5]) ? node132 : node123;
								assign node123 = (inp[7]) ? 3'b111 : node124;
									assign node124 = (inp[2]) ? node128 : node125;
										assign node125 = (inp[11]) ? 3'b011 : 3'b111;
										assign node128 = (inp[1]) ? 3'b111 : 3'b111;
								assign node132 = (inp[7]) ? node140 : node133;
									assign node133 = (inp[1]) ? node137 : node134;
										assign node134 = (inp[11]) ? 3'b101 : 3'b011;
										assign node137 = (inp[11]) ? 3'b011 : 3'b011;
									assign node140 = (inp[1]) ? node144 : node141;
										assign node141 = (inp[11]) ? 3'b011 : 3'b011;
										assign node144 = (inp[8]) ? 3'b111 : 3'b111;
						assign node147 = (inp[7]) ? 3'b111 : node148;
							assign node148 = (inp[11]) ? node150 : 3'b111;
								assign node150 = (inp[2]) ? 3'b111 : node151;
									assign node151 = (inp[10]) ? node153 : 3'b111;
										assign node153 = (inp[8]) ? 3'b111 : 3'b111;
				assign node158 = (inp[6]) ? node286 : node159;
					assign node159 = (inp[0]) ? node223 : node160;
						assign node160 = (inp[10]) ? node192 : node161;
							assign node161 = (inp[1]) ? node177 : node162;
								assign node162 = (inp[5]) ? node170 : node163;
									assign node163 = (inp[11]) ? node167 : node164;
										assign node164 = (inp[7]) ? 3'b101 : 3'b001;
										assign node167 = (inp[2]) ? 3'b001 : 3'b110;
									assign node170 = (inp[7]) ? node174 : node171;
										assign node171 = (inp[11]) ? 3'b010 : 3'b110;
										assign node174 = (inp[2]) ? 3'b001 : 3'b110;
								assign node177 = (inp[5]) ? node185 : node178;
									assign node178 = (inp[11]) ? node182 : node179;
										assign node179 = (inp[7]) ? 3'b011 : 3'b101;
										assign node182 = (inp[7]) ? 3'b101 : 3'b001;
									assign node185 = (inp[7]) ? node189 : node186;
										assign node186 = (inp[11]) ? 3'b110 : 3'b001;
										assign node189 = (inp[11]) ? 3'b001 : 3'b001;
							assign node192 = (inp[5]) ? node208 : node193;
								assign node193 = (inp[7]) ? node201 : node194;
									assign node194 = (inp[1]) ? node198 : node195;
										assign node195 = (inp[8]) ? 3'b110 : 3'b010;
										assign node198 = (inp[11]) ? 3'b110 : 3'b001;
									assign node201 = (inp[1]) ? node205 : node202;
										assign node202 = (inp[11]) ? 3'b110 : 3'b001;
										assign node205 = (inp[11]) ? 3'b001 : 3'b001;
								assign node208 = (inp[11]) ? node216 : node209;
									assign node209 = (inp[1]) ? node213 : node210;
										assign node210 = (inp[7]) ? 3'b110 : 3'b010;
										assign node213 = (inp[2]) ? 3'b110 : 3'b110;
									assign node216 = (inp[7]) ? node220 : node217;
										assign node217 = (inp[1]) ? 3'b010 : 3'b100;
										assign node220 = (inp[1]) ? 3'b010 : 3'b010;
						assign node223 = (inp[10]) ? node255 : node224;
							assign node224 = (inp[5]) ? node240 : node225;
								assign node225 = (inp[7]) ? node233 : node226;
									assign node226 = (inp[1]) ? node230 : node227;
										assign node227 = (inp[8]) ? 3'b101 : 3'b101;
										assign node230 = (inp[2]) ? 3'b011 : 3'b001;
									assign node233 = (inp[1]) ? node237 : node234;
										assign node234 = (inp[8]) ? 3'b011 : 3'b011;
										assign node237 = (inp[11]) ? 3'b011 : 3'b111;
								assign node240 = (inp[11]) ? node248 : node241;
									assign node241 = (inp[1]) ? node245 : node242;
										assign node242 = (inp[7]) ? 3'b101 : 3'b001;
										assign node245 = (inp[7]) ? 3'b011 : 3'b101;
									assign node248 = (inp[7]) ? node252 : node249;
										assign node249 = (inp[1]) ? 3'b101 : 3'b001;
										assign node252 = (inp[8]) ? 3'b101 : 3'b101;
							assign node255 = (inp[7]) ? node271 : node256;
								assign node256 = (inp[5]) ? node264 : node257;
									assign node257 = (inp[1]) ? node261 : node258;
										assign node258 = (inp[11]) ? 3'b001 : 3'b001;
										assign node261 = (inp[8]) ? 3'b101 : 3'b101;
									assign node264 = (inp[1]) ? node268 : node265;
										assign node265 = (inp[2]) ? 3'b110 : 3'b110;
										assign node268 = (inp[8]) ? 3'b001 : 3'b000;
								assign node271 = (inp[11]) ? node279 : node272;
									assign node272 = (inp[5]) ? node276 : node273;
										assign node273 = (inp[1]) ? 3'b011 : 3'b101;
										assign node276 = (inp[1]) ? 3'b101 : 3'b001;
									assign node279 = (inp[5]) ? node283 : node280;
										assign node280 = (inp[8]) ? 3'b101 : 3'b101;
										assign node283 = (inp[2]) ? 3'b001 : 3'b000;
					assign node286 = (inp[0]) ? node350 : node287;
						assign node287 = (inp[5]) ? node319 : node288;
							assign node288 = (inp[10]) ? node304 : node289;
								assign node289 = (inp[7]) ? node297 : node290;
									assign node290 = (inp[11]) ? node294 : node291;
										assign node291 = (inp[2]) ? 3'b011 : 3'b011;
										assign node294 = (inp[1]) ? 3'b011 : 3'b101;
									assign node297 = (inp[1]) ? node301 : node298;
										assign node298 = (inp[11]) ? 3'b011 : 3'b011;
										assign node301 = (inp[11]) ? 3'b111 : 3'b111;
								assign node304 = (inp[1]) ? node312 : node305;
									assign node305 = (inp[11]) ? node309 : node306;
										assign node306 = (inp[7]) ? 3'b101 : 3'b101;
										assign node309 = (inp[7]) ? 3'b101 : 3'b001;
									assign node312 = (inp[7]) ? node316 : node313;
										assign node313 = (inp[8]) ? 3'b001 : 3'b101;
										assign node316 = (inp[11]) ? 3'b011 : 3'b011;
							assign node319 = (inp[10]) ? node335 : node320;
								assign node320 = (inp[7]) ? node328 : node321;
									assign node321 = (inp[1]) ? node325 : node322;
										assign node322 = (inp[11]) ? 3'b001 : 3'b101;
										assign node325 = (inp[8]) ? 3'b101 : 3'b101;
									assign node328 = (inp[1]) ? node332 : node329;
										assign node329 = (inp[11]) ? 3'b101 : 3'b101;
										assign node332 = (inp[2]) ? 3'b011 : 3'b011;
								assign node335 = (inp[8]) ? node343 : node336;
									assign node336 = (inp[7]) ? node340 : node337;
										assign node337 = (inp[1]) ? 3'b001 : 3'b110;
										assign node340 = (inp[1]) ? 3'b101 : 3'b001;
									assign node343 = (inp[2]) ? node347 : node344;
										assign node344 = (inp[1]) ? 3'b001 : 3'b001;
										assign node347 = (inp[7]) ? 3'b101 : 3'b001;
						assign node350 = (inp[10]) ? node372 : node351;
							assign node351 = (inp[5]) ? node359 : node352;
								assign node352 = (inp[7]) ? 3'b111 : node353;
									assign node353 = (inp[8]) ? 3'b111 : node354;
										assign node354 = (inp[11]) ? 3'b111 : 3'b111;
								assign node359 = (inp[7]) ? node367 : node360;
									assign node360 = (inp[1]) ? node364 : node361;
										assign node361 = (inp[2]) ? 3'b011 : 3'b011;
										assign node364 = (inp[8]) ? 3'b111 : 3'b011;
									assign node367 = (inp[11]) ? node369 : 3'b111;
										assign node369 = (inp[1]) ? 3'b111 : 3'b011;
							assign node372 = (inp[5]) ? node386 : node373;
								assign node373 = (inp[1]) ? node381 : node374;
									assign node374 = (inp[7]) ? node378 : node375;
										assign node375 = (inp[8]) ? 3'b011 : 3'b001;
										assign node378 = (inp[2]) ? 3'b111 : 3'b011;
									assign node381 = (inp[7]) ? 3'b111 : node382;
										assign node382 = (inp[2]) ? 3'b111 : 3'b011;
								assign node386 = (inp[1]) ? node394 : node387;
									assign node387 = (inp[7]) ? node391 : node388;
										assign node388 = (inp[11]) ? 3'b001 : 3'b101;
										assign node391 = (inp[8]) ? 3'b011 : 3'b101;
									assign node394 = (inp[7]) ? node398 : node395;
										assign node395 = (inp[8]) ? 3'b011 : 3'b101;
										assign node398 = (inp[11]) ? 3'b011 : 3'b111;
			assign node401 = (inp[4]) ? node643 : node402;
				assign node402 = (inp[6]) ? node528 : node403;
					assign node403 = (inp[0]) ? node465 : node404;
						assign node404 = (inp[5]) ? node436 : node405;
							assign node405 = (inp[10]) ? node421 : node406;
								assign node406 = (inp[1]) ? node414 : node407;
									assign node407 = (inp[7]) ? node411 : node408;
										assign node408 = (inp[8]) ? 3'b001 : 3'b110;
										assign node411 = (inp[11]) ? 3'b001 : 3'b101;
									assign node414 = (inp[7]) ? node418 : node415;
										assign node415 = (inp[11]) ? 3'b001 : 3'b101;
										assign node418 = (inp[11]) ? 3'b101 : 3'b101;
								assign node421 = (inp[1]) ? node429 : node422;
									assign node422 = (inp[7]) ? node426 : node423;
										assign node423 = (inp[8]) ? 3'b110 : 3'b010;
										assign node426 = (inp[11]) ? 3'b110 : 3'b001;
									assign node429 = (inp[2]) ? node433 : node430;
										assign node430 = (inp[8]) ? 3'b001 : 3'b110;
										assign node433 = (inp[7]) ? 3'b001 : 3'b001;
							assign node436 = (inp[10]) ? node452 : node437;
								assign node437 = (inp[7]) ? node445 : node438;
									assign node438 = (inp[1]) ? node442 : node439;
										assign node439 = (inp[11]) ? 3'b010 : 3'b110;
										assign node442 = (inp[11]) ? 3'b110 : 3'b001;
									assign node445 = (inp[8]) ? node449 : node446;
										assign node446 = (inp[11]) ? 3'b110 : 3'b001;
										assign node449 = (inp[2]) ? 3'b001 : 3'b001;
								assign node452 = (inp[7]) ? node460 : node453;
									assign node453 = (inp[1]) ? node457 : node454;
										assign node454 = (inp[2]) ? 3'b010 : 3'b100;
										assign node457 = (inp[2]) ? 3'b010 : 3'b010;
									assign node460 = (inp[11]) ? node462 : 3'b110;
										assign node462 = (inp[1]) ? 3'b110 : 3'b010;
						assign node465 = (inp[5]) ? node497 : node466;
							assign node466 = (inp[10]) ? node482 : node467;
								assign node467 = (inp[7]) ? node475 : node468;
									assign node468 = (inp[1]) ? node472 : node469;
										assign node469 = (inp[2]) ? 3'b101 : 3'b101;
										assign node472 = (inp[11]) ? 3'b011 : 3'b011;
									assign node475 = (inp[11]) ? node479 : node476;
										assign node476 = (inp[1]) ? 3'b111 : 3'b011;
										assign node479 = (inp[8]) ? 3'b011 : 3'b011;
								assign node482 = (inp[7]) ? node490 : node483;
									assign node483 = (inp[8]) ? node487 : node484;
										assign node484 = (inp[2]) ? 3'b001 : 3'b001;
										assign node487 = (inp[1]) ? 3'b101 : 3'b001;
									assign node490 = (inp[1]) ? node494 : node491;
										assign node491 = (inp[2]) ? 3'b101 : 3'b101;
										assign node494 = (inp[8]) ? 3'b011 : 3'b101;
							assign node497 = (inp[10]) ? node513 : node498;
								assign node498 = (inp[11]) ? node506 : node499;
									assign node499 = (inp[7]) ? node503 : node500;
										assign node500 = (inp[1]) ? 3'b101 : 3'b001;
										assign node503 = (inp[1]) ? 3'b011 : 3'b101;
									assign node506 = (inp[1]) ? node510 : node507;
										assign node507 = (inp[7]) ? 3'b101 : 3'b001;
										assign node510 = (inp[2]) ? 3'b101 : 3'b101;
								assign node513 = (inp[7]) ? node521 : node514;
									assign node514 = (inp[11]) ? node518 : node515;
										assign node515 = (inp[1]) ? 3'b001 : 3'b110;
										assign node518 = (inp[2]) ? 3'b110 : 3'b110;
									assign node521 = (inp[8]) ? node525 : node522;
										assign node522 = (inp[11]) ? 3'b000 : 3'b001;
										assign node525 = (inp[1]) ? 3'b101 : 3'b001;
					assign node528 = (inp[0]) ? node592 : node529;
						assign node529 = (inp[10]) ? node561 : node530;
							assign node530 = (inp[5]) ? node546 : node531;
								assign node531 = (inp[11]) ? node539 : node532;
									assign node532 = (inp[7]) ? node536 : node533;
										assign node533 = (inp[2]) ? 3'b011 : 3'b011;
										assign node536 = (inp[1]) ? 3'b111 : 3'b011;
									assign node539 = (inp[7]) ? node543 : node540;
										assign node540 = (inp[1]) ? 3'b011 : 3'b101;
										assign node543 = (inp[1]) ? 3'b111 : 3'b011;
								assign node546 = (inp[7]) ? node554 : node547;
									assign node547 = (inp[1]) ? node551 : node548;
										assign node548 = (inp[11]) ? 3'b001 : 3'b101;
										assign node551 = (inp[11]) ? 3'b101 : 3'b101;
									assign node554 = (inp[1]) ? node558 : node555;
										assign node555 = (inp[8]) ? 3'b101 : 3'b101;
										assign node558 = (inp[2]) ? 3'b011 : 3'b011;
							assign node561 = (inp[5]) ? node577 : node562;
								assign node562 = (inp[1]) ? node570 : node563;
									assign node563 = (inp[7]) ? node567 : node564;
										assign node564 = (inp[11]) ? 3'b001 : 3'b001;
										assign node567 = (inp[8]) ? 3'b101 : 3'b101;
									assign node570 = (inp[7]) ? node574 : node571;
										assign node571 = (inp[11]) ? 3'b101 : 3'b001;
										assign node574 = (inp[11]) ? 3'b001 : 3'b011;
								assign node577 = (inp[7]) ? node585 : node578;
									assign node578 = (inp[1]) ? node582 : node579;
										assign node579 = (inp[8]) ? 3'b110 : 3'b110;
										assign node582 = (inp[11]) ? 3'b110 : 3'b001;
									assign node585 = (inp[2]) ? node589 : node586;
										assign node586 = (inp[8]) ? 3'b001 : 3'b001;
										assign node589 = (inp[8]) ? 3'b101 : 3'b001;
						assign node592 = (inp[10]) ? node614 : node593;
							assign node593 = (inp[5]) ? node601 : node594;
								assign node594 = (inp[7]) ? 3'b111 : node595;
									assign node595 = (inp[1]) ? 3'b111 : node596;
										assign node596 = (inp[11]) ? 3'b011 : 3'b111;
								assign node601 = (inp[1]) ? node609 : node602;
									assign node602 = (inp[11]) ? node606 : node603;
										assign node603 = (inp[7]) ? 3'b111 : 3'b011;
										assign node606 = (inp[7]) ? 3'b011 : 3'b101;
									assign node609 = (inp[7]) ? 3'b111 : node610;
										assign node610 = (inp[11]) ? 3'b011 : 3'b111;
							assign node614 = (inp[5]) ? node628 : node615;
								assign node615 = (inp[7]) ? node623 : node616;
									assign node616 = (inp[11]) ? node620 : node617;
										assign node617 = (inp[1]) ? 3'b111 : 3'b011;
										assign node620 = (inp[1]) ? 3'b011 : 3'b101;
									assign node623 = (inp[1]) ? 3'b111 : node624;
										assign node624 = (inp[8]) ? 3'b111 : 3'b011;
								assign node628 = (inp[7]) ? node636 : node629;
									assign node629 = (inp[1]) ? node633 : node630;
										assign node630 = (inp[11]) ? 3'b001 : 3'b101;
										assign node633 = (inp[8]) ? 3'b011 : 3'b101;
									assign node636 = (inp[1]) ? node640 : node637;
										assign node637 = (inp[8]) ? 3'b011 : 3'b101;
										assign node640 = (inp[8]) ? 3'b011 : 3'b011;
				assign node643 = (inp[6]) ? node765 : node644;
					assign node644 = (inp[0]) ? node704 : node645;
						assign node645 = (inp[10]) ? node675 : node646;
							assign node646 = (inp[5]) ? node662 : node647;
								assign node647 = (inp[7]) ? node655 : node648;
									assign node648 = (inp[1]) ? node652 : node649;
										assign node649 = (inp[2]) ? 3'b010 : 3'b100;
										assign node652 = (inp[11]) ? 3'b010 : 3'b010;
									assign node655 = (inp[8]) ? node659 : node656;
										assign node656 = (inp[1]) ? 3'b110 : 3'b010;
										assign node659 = (inp[2]) ? 3'b110 : 3'b110;
								assign node662 = (inp[7]) ? node670 : node663;
									assign node663 = (inp[1]) ? node667 : node664;
										assign node664 = (inp[8]) ? 3'b100 : 3'b000;
										assign node667 = (inp[11]) ? 3'b100 : 3'b100;
									assign node670 = (inp[11]) ? node672 : 3'b010;
										assign node672 = (inp[1]) ? 3'b010 : 3'b100;
							assign node675 = (inp[5]) ? node691 : node676;
								assign node676 = (inp[7]) ? node684 : node677;
									assign node677 = (inp[8]) ? node681 : node678;
										assign node678 = (inp[2]) ? 3'b100 : 3'b000;
										assign node681 = (inp[11]) ? 3'b100 : 3'b100;
									assign node684 = (inp[1]) ? node688 : node685;
										assign node685 = (inp[8]) ? 3'b000 : 3'b100;
										assign node688 = (inp[8]) ? 3'b010 : 3'b010;
								assign node691 = (inp[1]) ? node697 : node692;
									assign node692 = (inp[7]) ? node694 : 3'b000;
										assign node694 = (inp[8]) ? 3'b000 : 3'b000;
									assign node697 = (inp[7]) ? node701 : node698;
										assign node698 = (inp[2]) ? 3'b000 : 3'b000;
										assign node701 = (inp[11]) ? 3'b100 : 3'b100;
						assign node704 = (inp[10]) ? node736 : node705;
							assign node705 = (inp[5]) ? node721 : node706;
								assign node706 = (inp[7]) ? node714 : node707;
									assign node707 = (inp[1]) ? node711 : node708;
										assign node708 = (inp[2]) ? 3'b110 : 3'b110;
										assign node711 = (inp[11]) ? 3'b110 : 3'b001;
									assign node714 = (inp[11]) ? node718 : node715;
										assign node715 = (inp[8]) ? 3'b101 : 3'b001;
										assign node718 = (inp[2]) ? 3'b001 : 3'b001;
								assign node721 = (inp[7]) ? node729 : node722;
									assign node722 = (inp[11]) ? node726 : node723;
										assign node723 = (inp[1]) ? 3'b110 : 3'b010;
										assign node726 = (inp[2]) ? 3'b010 : 3'b010;
									assign node729 = (inp[1]) ? node733 : node730;
										assign node730 = (inp[11]) ? 3'b010 : 3'b110;
										assign node733 = (inp[8]) ? 3'b001 : 3'b110;
							assign node736 = (inp[5]) ? node750 : node737;
								assign node737 = (inp[11]) ? node743 : node738;
									assign node738 = (inp[7]) ? 3'b110 : node739;
										assign node739 = (inp[1]) ? 3'b110 : 3'b010;
									assign node743 = (inp[7]) ? node747 : node744;
										assign node744 = (inp[2]) ? 3'b010 : 3'b010;
										assign node747 = (inp[1]) ? 3'b110 : 3'b010;
								assign node750 = (inp[7]) ? node758 : node751;
									assign node751 = (inp[1]) ? node755 : node752;
										assign node752 = (inp[2]) ? 3'b100 : 3'b100;
										assign node755 = (inp[8]) ? 3'b010 : 3'b100;
									assign node758 = (inp[11]) ? node762 : node759;
										assign node759 = (inp[1]) ? 3'b110 : 3'b010;
										assign node762 = (inp[1]) ? 3'b010 : 3'b100;
					assign node765 = (inp[0]) ? node829 : node766;
						assign node766 = (inp[10]) ? node798 : node767;
							assign node767 = (inp[5]) ? node783 : node768;
								assign node768 = (inp[1]) ? node776 : node769;
									assign node769 = (inp[7]) ? node773 : node770;
										assign node770 = (inp[11]) ? 3'b110 : 3'b110;
										assign node773 = (inp[8]) ? 3'b001 : 3'b000;
									assign node776 = (inp[7]) ? node780 : node777;
										assign node777 = (inp[8]) ? 3'b001 : 3'b001;
										assign node780 = (inp[8]) ? 3'b101 : 3'b001;
								assign node783 = (inp[11]) ? node791 : node784;
									assign node784 = (inp[7]) ? node788 : node785;
										assign node785 = (inp[1]) ? 3'b110 : 3'b010;
										assign node788 = (inp[1]) ? 3'b001 : 3'b110;
									assign node791 = (inp[1]) ? node795 : node792;
										assign node792 = (inp[7]) ? 3'b110 : 3'b010;
										assign node795 = (inp[7]) ? 3'b110 : 3'b110;
							assign node798 = (inp[7]) ? node814 : node799;
								assign node799 = (inp[5]) ? node807 : node800;
									assign node800 = (inp[1]) ? node804 : node801;
										assign node801 = (inp[8]) ? 3'b010 : 3'b010;
										assign node804 = (inp[2]) ? 3'b110 : 3'b110;
									assign node807 = (inp[1]) ? node811 : node808;
										assign node808 = (inp[8]) ? 3'b100 : 3'b100;
										assign node811 = (inp[11]) ? 3'b100 : 3'b010;
								assign node814 = (inp[5]) ? node822 : node815;
									assign node815 = (inp[11]) ? node819 : node816;
										assign node816 = (inp[1]) ? 3'b001 : 3'b110;
										assign node819 = (inp[2]) ? 3'b110 : 3'b110;
									assign node822 = (inp[2]) ? node826 : node823;
										assign node823 = (inp[1]) ? 3'b010 : 3'b010;
										assign node826 = (inp[1]) ? 3'b110 : 3'b010;
						assign node829 = (inp[5]) ? node861 : node830;
							assign node830 = (inp[10]) ? node846 : node831;
								assign node831 = (inp[7]) ? node839 : node832;
									assign node832 = (inp[11]) ? node836 : node833;
										assign node833 = (inp[1]) ? 3'b011 : 3'b101;
										assign node836 = (inp[1]) ? 3'b101 : 3'b001;
									assign node839 = (inp[1]) ? node843 : node840;
										assign node840 = (inp[11]) ? 3'b101 : 3'b011;
										assign node843 = (inp[11]) ? 3'b011 : 3'b111;
								assign node846 = (inp[7]) ? node854 : node847;
									assign node847 = (inp[1]) ? node851 : node848;
										assign node848 = (inp[11]) ? 3'b110 : 3'b001;
										assign node851 = (inp[11]) ? 3'b001 : 3'b101;
									assign node854 = (inp[8]) ? node858 : node855;
										assign node855 = (inp[2]) ? 3'b101 : 3'b001;
										assign node858 = (inp[1]) ? 3'b101 : 3'b101;
							assign node861 = (inp[10]) ? node877 : node862;
								assign node862 = (inp[7]) ? node870 : node863;
									assign node863 = (inp[1]) ? node867 : node864;
										assign node864 = (inp[11]) ? 3'b110 : 3'b001;
										assign node867 = (inp[11]) ? 3'b001 : 3'b101;
									assign node870 = (inp[2]) ? node874 : node871;
										assign node871 = (inp[1]) ? 3'b101 : 3'b001;
										assign node874 = (inp[11]) ? 3'b101 : 3'b101;
								assign node877 = (inp[11]) ? node885 : node878;
									assign node878 = (inp[7]) ? node882 : node879;
										assign node879 = (inp[1]) ? 3'b001 : 3'b110;
										assign node882 = (inp[8]) ? 3'b001 : 3'b001;
									assign node885 = (inp[7]) ? node889 : node886;
										assign node886 = (inp[1]) ? 3'b110 : 3'b010;
										assign node889 = (inp[1]) ? 3'b001 : 3'b110;
		assign node892 = (inp[9]) ? node1332 : node893;
			assign node893 = (inp[4]) ? node1143 : node894;
				assign node894 = (inp[6]) ? node1018 : node895;
					assign node895 = (inp[0]) ? node955 : node896;
						assign node896 = (inp[5]) ? node928 : node897;
							assign node897 = (inp[10]) ? node913 : node898;
								assign node898 = (inp[7]) ? node906 : node899;
									assign node899 = (inp[1]) ? node903 : node900;
										assign node900 = (inp[2]) ? 3'b010 : 3'b100;
										assign node903 = (inp[11]) ? 3'b010 : 3'b110;
									assign node906 = (inp[8]) ? node910 : node907;
										assign node907 = (inp[11]) ? 3'b010 : 3'b110;
										assign node910 = (inp[2]) ? 3'b110 : 3'b110;
								assign node913 = (inp[7]) ? node921 : node914;
									assign node914 = (inp[1]) ? node918 : node915;
										assign node915 = (inp[8]) ? 3'b100 : 3'b000;
										assign node918 = (inp[11]) ? 3'b100 : 3'b010;
									assign node921 = (inp[1]) ? node925 : node922;
										assign node922 = (inp[11]) ? 3'b100 : 3'b010;
										assign node925 = (inp[2]) ? 3'b010 : 3'b010;
							assign node928 = (inp[10]) ? node942 : node929;
								assign node929 = (inp[7]) ? node937 : node930;
									assign node930 = (inp[1]) ? node934 : node931;
										assign node931 = (inp[11]) ? 3'b000 : 3'b100;
										assign node934 = (inp[11]) ? 3'b100 : 3'b010;
									assign node937 = (inp[2]) ? 3'b010 : node938;
										assign node938 = (inp[8]) ? 3'b010 : 3'b100;
								assign node942 = (inp[7]) ? node948 : node943;
									assign node943 = (inp[11]) ? 3'b000 : node944;
										assign node944 = (inp[8]) ? 3'b000 : 3'b000;
									assign node948 = (inp[1]) ? node952 : node949;
										assign node949 = (inp[11]) ? 3'b000 : 3'b100;
										assign node952 = (inp[11]) ? 3'b100 : 3'b100;
						assign node955 = (inp[10]) ? node987 : node956;
							assign node956 = (inp[5]) ? node972 : node957;
								assign node957 = (inp[7]) ? node965 : node958;
									assign node958 = (inp[1]) ? node962 : node959;
										assign node959 = (inp[11]) ? 3'b110 : 3'b110;
										assign node962 = (inp[11]) ? 3'b000 : 3'b001;
									assign node965 = (inp[1]) ? node969 : node966;
										assign node966 = (inp[11]) ? 3'b001 : 3'b001;
										assign node969 = (inp[11]) ? 3'b001 : 3'b101;
								assign node972 = (inp[7]) ? node980 : node973;
									assign node973 = (inp[11]) ? node977 : node974;
										assign node974 = (inp[1]) ? 3'b110 : 3'b010;
										assign node977 = (inp[2]) ? 3'b010 : 3'b110;
									assign node980 = (inp[8]) ? node984 : node981;
										assign node981 = (inp[11]) ? 3'b110 : 3'b110;
										assign node984 = (inp[11]) ? 3'b110 : 3'b001;
							assign node987 = (inp[5]) ? node1003 : node988;
								assign node988 = (inp[7]) ? node996 : node989;
									assign node989 = (inp[11]) ? node993 : node990;
										assign node990 = (inp[1]) ? 3'b110 : 3'b010;
										assign node993 = (inp[1]) ? 3'b010 : 3'b010;
									assign node996 = (inp[1]) ? node1000 : node997;
										assign node997 = (inp[2]) ? 3'b110 : 3'b110;
										assign node1000 = (inp[8]) ? 3'b001 : 3'b110;
								assign node1003 = (inp[7]) ? node1011 : node1004;
									assign node1004 = (inp[11]) ? node1008 : node1005;
										assign node1005 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1008 = (inp[8]) ? 3'b100 : 3'b100;
									assign node1011 = (inp[1]) ? node1015 : node1012;
										assign node1012 = (inp[11]) ? 3'b100 : 3'b010;
										assign node1015 = (inp[11]) ? 3'b010 : 3'b110;
					assign node1018 = (inp[0]) ? node1080 : node1019;
						assign node1019 = (inp[10]) ? node1051 : node1020;
							assign node1020 = (inp[5]) ? node1036 : node1021;
								assign node1021 = (inp[1]) ? node1029 : node1022;
									assign node1022 = (inp[7]) ? node1026 : node1023;
										assign node1023 = (inp[11]) ? 3'b110 : 3'b001;
										assign node1026 = (inp[8]) ? 3'b001 : 3'b001;
									assign node1029 = (inp[7]) ? node1033 : node1030;
										assign node1030 = (inp[8]) ? 3'b001 : 3'b001;
										assign node1033 = (inp[8]) ? 3'b101 : 3'b101;
								assign node1036 = (inp[11]) ? node1044 : node1037;
									assign node1037 = (inp[7]) ? node1041 : node1038;
										assign node1038 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1041 = (inp[1]) ? 3'b001 : 3'b110;
									assign node1044 = (inp[7]) ? node1048 : node1045;
										assign node1045 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1048 = (inp[1]) ? 3'b110 : 3'b110;
							assign node1051 = (inp[5]) ? node1067 : node1052;
								assign node1052 = (inp[11]) ? node1060 : node1053;
									assign node1053 = (inp[7]) ? node1057 : node1054;
										assign node1054 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1057 = (inp[1]) ? 3'b001 : 3'b110;
									assign node1060 = (inp[7]) ? node1064 : node1061;
										assign node1061 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1064 = (inp[1]) ? 3'b110 : 3'b110;
								assign node1067 = (inp[1]) ? node1075 : node1068;
									assign node1068 = (inp[7]) ? node1072 : node1069;
										assign node1069 = (inp[11]) ? 3'b100 : 3'b100;
										assign node1072 = (inp[8]) ? 3'b010 : 3'b010;
									assign node1075 = (inp[11]) ? 3'b010 : node1076;
										assign node1076 = (inp[7]) ? 3'b110 : 3'b010;
						assign node1080 = (inp[10]) ? node1112 : node1081;
							assign node1081 = (inp[7]) ? node1097 : node1082;
								assign node1082 = (inp[5]) ? node1090 : node1083;
									assign node1083 = (inp[2]) ? node1087 : node1084;
										assign node1084 = (inp[1]) ? 3'b101 : 3'b101;
										assign node1087 = (inp[1]) ? 3'b011 : 3'b101;
									assign node1090 = (inp[1]) ? node1094 : node1091;
										assign node1091 = (inp[11]) ? 3'b000 : 3'b001;
										assign node1094 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1097 = (inp[5]) ? node1105 : node1098;
									assign node1098 = (inp[2]) ? node1102 : node1099;
										assign node1099 = (inp[1]) ? 3'b011 : 3'b101;
										assign node1102 = (inp[1]) ? 3'b011 : 3'b011;
									assign node1105 = (inp[1]) ? node1109 : node1106;
										assign node1106 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1109 = (inp[11]) ? 3'b101 : 3'b011;
							assign node1112 = (inp[5]) ? node1128 : node1113;
								assign node1113 = (inp[7]) ? node1121 : node1114;
									assign node1114 = (inp[11]) ? node1118 : node1115;
										assign node1115 = (inp[1]) ? 3'b101 : 3'b001;
										assign node1118 = (inp[1]) ? 3'b001 : 3'b110;
									assign node1121 = (inp[1]) ? node1125 : node1122;
										assign node1122 = (inp[11]) ? 3'b001 : 3'b101;
										assign node1125 = (inp[11]) ? 3'b101 : 3'b011;
								assign node1128 = (inp[7]) ? node1136 : node1129;
									assign node1129 = (inp[1]) ? node1133 : node1130;
										assign node1130 = (inp[2]) ? 3'b110 : 3'b010;
										assign node1133 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1136 = (inp[1]) ? node1140 : node1137;
										assign node1137 = (inp[2]) ? 3'b001 : 3'b110;
										assign node1140 = (inp[8]) ? 3'b001 : 3'b001;
				assign node1143 = (inp[6]) ? node1219 : node1144;
					assign node1144 = (inp[0]) ? node1168 : node1145;
						assign node1145 = (inp[5]) ? 3'b000 : node1146;
							assign node1146 = (inp[10]) ? node1160 : node1147;
								assign node1147 = (inp[7]) ? node1153 : node1148;
									assign node1148 = (inp[8]) ? node1150 : 3'b000;
										assign node1150 = (inp[11]) ? 3'b000 : 3'b000;
									assign node1153 = (inp[2]) ? node1157 : node1154;
										assign node1154 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1157 = (inp[8]) ? 3'b100 : 3'b100;
								assign node1160 = (inp[11]) ? 3'b000 : node1161;
									assign node1161 = (inp[2]) ? node1163 : 3'b000;
										assign node1163 = (inp[1]) ? 3'b000 : 3'b000;
						assign node1168 = (inp[5]) ? node1198 : node1169;
							assign node1169 = (inp[10]) ? node1185 : node1170;
								assign node1170 = (inp[7]) ? node1178 : node1171;
									assign node1171 = (inp[11]) ? node1175 : node1172;
										assign node1172 = (inp[1]) ? 3'b010 : 3'b100;
										assign node1175 = (inp[1]) ? 3'b100 : 3'b100;
									assign node1178 = (inp[1]) ? node1182 : node1179;
										assign node1179 = (inp[8]) ? 3'b010 : 3'b000;
										assign node1182 = (inp[11]) ? 3'b010 : 3'b110;
								assign node1185 = (inp[7]) ? node1191 : node1186;
									assign node1186 = (inp[2]) ? node1188 : 3'b000;
										assign node1188 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1191 = (inp[1]) ? node1195 : node1192;
										assign node1192 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1195 = (inp[11]) ? 3'b100 : 3'b010;
							assign node1198 = (inp[10]) ? node1212 : node1199;
								assign node1199 = (inp[11]) ? node1207 : node1200;
									assign node1200 = (inp[2]) ? node1204 : node1201;
										assign node1201 = (inp[7]) ? 3'b100 : 3'b000;
										assign node1204 = (inp[7]) ? 3'b000 : 3'b100;
									assign node1207 = (inp[7]) ? node1209 : 3'b000;
										assign node1209 = (inp[1]) ? 3'b100 : 3'b000;
								assign node1212 = (inp[1]) ? node1214 : 3'b000;
									assign node1214 = (inp[7]) ? node1216 : 3'b000;
										assign node1216 = (inp[2]) ? 3'b100 : 3'b000;
					assign node1219 = (inp[0]) ? node1271 : node1220;
						assign node1220 = (inp[10]) ? node1250 : node1221;
							assign node1221 = (inp[5]) ? node1235 : node1222;
								assign node1222 = (inp[7]) ? node1230 : node1223;
									assign node1223 = (inp[1]) ? node1227 : node1224;
										assign node1224 = (inp[2]) ? 3'b100 : 3'b100;
										assign node1227 = (inp[11]) ? 3'b010 : 3'b010;
									assign node1230 = (inp[11]) ? 3'b010 : node1231;
										assign node1231 = (inp[1]) ? 3'b110 : 3'b010;
								assign node1235 = (inp[7]) ? node1243 : node1236;
									assign node1236 = (inp[1]) ? node1240 : node1237;
										assign node1237 = (inp[2]) ? 3'b000 : 3'b000;
										assign node1240 = (inp[8]) ? 3'b100 : 3'b100;
									assign node1243 = (inp[1]) ? node1247 : node1244;
										assign node1244 = (inp[11]) ? 3'b100 : 3'b100;
										assign node1247 = (inp[11]) ? 3'b100 : 3'b010;
							assign node1250 = (inp[5]) ? node1264 : node1251;
								assign node1251 = (inp[7]) ? node1257 : node1252;
									assign node1252 = (inp[1]) ? node1254 : 3'b000;
										assign node1254 = (inp[2]) ? 3'b100 : 3'b100;
									assign node1257 = (inp[2]) ? node1261 : node1258;
										assign node1258 = (inp[11]) ? 3'b100 : 3'b100;
										assign node1261 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1264 = (inp[1]) ? node1266 : 3'b000;
									assign node1266 = (inp[7]) ? node1268 : 3'b000;
										assign node1268 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1271 = (inp[10]) ? node1303 : node1272;
							assign node1272 = (inp[5]) ? node1288 : node1273;
								assign node1273 = (inp[7]) ? node1281 : node1274;
									assign node1274 = (inp[1]) ? node1278 : node1275;
										assign node1275 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1278 = (inp[8]) ? 3'b001 : 3'b110;
									assign node1281 = (inp[1]) ? node1285 : node1282;
										assign node1282 = (inp[2]) ? 3'b001 : 3'b110;
										assign node1285 = (inp[11]) ? 3'b001 : 3'b101;
								assign node1288 = (inp[7]) ? node1296 : node1289;
									assign node1289 = (inp[2]) ? node1293 : node1290;
										assign node1290 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1293 = (inp[8]) ? 3'b010 : 3'b010;
									assign node1296 = (inp[2]) ? node1300 : node1297;
										assign node1297 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1300 = (inp[11]) ? 3'b110 : 3'b110;
							assign node1303 = (inp[5]) ? node1317 : node1304;
								assign node1304 = (inp[11]) ? node1310 : node1305;
									assign node1305 = (inp[1]) ? 3'b110 : node1306;
										assign node1306 = (inp[7]) ? 3'b110 : 3'b010;
									assign node1310 = (inp[1]) ? node1314 : node1311;
										assign node1311 = (inp[7]) ? 3'b010 : 3'b100;
										assign node1314 = (inp[7]) ? 3'b110 : 3'b010;
								assign node1317 = (inp[1]) ? node1325 : node1318;
									assign node1318 = (inp[7]) ? node1322 : node1319;
										assign node1319 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1322 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1325 = (inp[7]) ? node1329 : node1326;
										assign node1326 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1329 = (inp[11]) ? 3'b010 : 3'b010;
			assign node1332 = (inp[4]) ? node1536 : node1333;
				assign node1333 = (inp[6]) ? node1417 : node1334;
					assign node1334 = (inp[0]) ? node1366 : node1335;
						assign node1335 = (inp[5]) ? node1357 : node1336;
							assign node1336 = (inp[7]) ? node1344 : node1337;
								assign node1337 = (inp[2]) ? node1339 : 3'b000;
									assign node1339 = (inp[8]) ? node1341 : 3'b000;
										assign node1341 = (inp[11]) ? 3'b000 : 3'b000;
								assign node1344 = (inp[10]) ? node1352 : node1345;
									assign node1345 = (inp[1]) ? node1349 : node1346;
										assign node1346 = (inp[8]) ? 3'b000 : 3'b000;
										assign node1349 = (inp[8]) ? 3'b100 : 3'b100;
									assign node1352 = (inp[8]) ? node1354 : 3'b000;
										assign node1354 = (inp[11]) ? 3'b000 : 3'b000;
							assign node1357 = (inp[10]) ? 3'b000 : node1358;
								assign node1358 = (inp[11]) ? 3'b000 : node1359;
									assign node1359 = (inp[7]) ? node1361 : 3'b000;
										assign node1361 = (inp[8]) ? 3'b000 : 3'b000;
						assign node1366 = (inp[10]) ? node1396 : node1367;
							assign node1367 = (inp[5]) ? node1383 : node1368;
								assign node1368 = (inp[7]) ? node1376 : node1369;
									assign node1369 = (inp[2]) ? node1373 : node1370;
										assign node1370 = (inp[11]) ? 3'b100 : 3'b100;
										assign node1373 = (inp[11]) ? 3'b100 : 3'b010;
									assign node1376 = (inp[11]) ? node1380 : node1377;
										assign node1377 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1380 = (inp[1]) ? 3'b010 : 3'b100;
								assign node1383 = (inp[7]) ? node1389 : node1384;
									assign node1384 = (inp[1]) ? node1386 : 3'b000;
										assign node1386 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1389 = (inp[1]) ? node1393 : node1390;
										assign node1390 = (inp[11]) ? 3'b000 : 3'b100;
										assign node1393 = (inp[8]) ? 3'b010 : 3'b100;
							assign node1396 = (inp[5]) ? node1410 : node1397;
								assign node1397 = (inp[1]) ? node1403 : node1398;
									assign node1398 = (inp[2]) ? node1400 : 3'b000;
										assign node1400 = (inp[7]) ? 3'b100 : 3'b000;
									assign node1403 = (inp[7]) ? node1407 : node1404;
										assign node1404 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1407 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1410 = (inp[7]) ? node1412 : 3'b000;
									assign node1412 = (inp[1]) ? node1414 : 3'b000;
										assign node1414 = (inp[11]) ? 3'b000 : 3'b100;
					assign node1417 = (inp[0]) ? node1473 : node1418;
						assign node1418 = (inp[10]) ? node1450 : node1419;
							assign node1419 = (inp[5]) ? node1435 : node1420;
								assign node1420 = (inp[7]) ? node1428 : node1421;
									assign node1421 = (inp[1]) ? node1425 : node1422;
										assign node1422 = (inp[2]) ? 3'b100 : 3'b100;
										assign node1425 = (inp[8]) ? 3'b010 : 3'b000;
									assign node1428 = (inp[11]) ? node1432 : node1429;
										assign node1429 = (inp[1]) ? 3'b110 : 3'b010;
										assign node1432 = (inp[8]) ? 3'b010 : 3'b010;
								assign node1435 = (inp[7]) ? node1443 : node1436;
									assign node1436 = (inp[11]) ? node1440 : node1437;
										assign node1437 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1440 = (inp[2]) ? 3'b000 : 3'b000;
									assign node1443 = (inp[1]) ? node1447 : node1444;
										assign node1444 = (inp[8]) ? 3'b100 : 3'b100;
										assign node1447 = (inp[2]) ? 3'b010 : 3'b100;
							assign node1450 = (inp[5]) ? node1466 : node1451;
								assign node1451 = (inp[7]) ? node1459 : node1452;
									assign node1452 = (inp[1]) ? node1456 : node1453;
										assign node1453 = (inp[2]) ? 3'b000 : 3'b000;
										assign node1456 = (inp[11]) ? 3'b000 : 3'b100;
									assign node1459 = (inp[1]) ? node1463 : node1460;
										assign node1460 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1463 = (inp[11]) ? 3'b100 : 3'b010;
								assign node1466 = (inp[1]) ? node1468 : 3'b000;
									assign node1468 = (inp[7]) ? node1470 : 3'b000;
										assign node1470 = (inp[8]) ? 3'b100 : 3'b000;
						assign node1473 = (inp[5]) ? node1505 : node1474;
							assign node1474 = (inp[10]) ? node1490 : node1475;
								assign node1475 = (inp[7]) ? node1483 : node1476;
									assign node1476 = (inp[1]) ? node1480 : node1477;
										assign node1477 = (inp[8]) ? 3'b110 : 3'b010;
										assign node1480 = (inp[11]) ? 3'b110 : 3'b001;
									assign node1483 = (inp[11]) ? node1487 : node1484;
										assign node1484 = (inp[8]) ? 3'b001 : 3'b001;
										assign node1487 = (inp[8]) ? 3'b001 : 3'b110;
								assign node1490 = (inp[7]) ? node1498 : node1491;
									assign node1491 = (inp[1]) ? node1495 : node1492;
										assign node1492 = (inp[2]) ? 3'b010 : 3'b100;
										assign node1495 = (inp[8]) ? 3'b010 : 3'b010;
									assign node1498 = (inp[11]) ? node1502 : node1499;
										assign node1499 = (inp[1]) ? 3'b110 : 3'b110;
										assign node1502 = (inp[1]) ? 3'b110 : 3'b010;
							assign node1505 = (inp[10]) ? node1521 : node1506;
								assign node1506 = (inp[7]) ? node1514 : node1507;
									assign node1507 = (inp[1]) ? node1511 : node1508;
										assign node1508 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1511 = (inp[8]) ? 3'b110 : 3'b010;
									assign node1514 = (inp[1]) ? node1518 : node1515;
										assign node1515 = (inp[11]) ? 3'b010 : 3'b110;
										assign node1518 = (inp[2]) ? 3'b110 : 3'b110;
								assign node1521 = (inp[7]) ? node1529 : node1522;
									assign node1522 = (inp[11]) ? node1526 : node1523;
										assign node1523 = (inp[1]) ? 3'b100 : 3'b100;
										assign node1526 = (inp[8]) ? 3'b100 : 3'b000;
									assign node1529 = (inp[1]) ? node1533 : node1530;
										assign node1530 = (inp[8]) ? 3'b010 : 3'b100;
										assign node1533 = (inp[8]) ? 3'b010 : 3'b010;
				assign node1536 = (inp[0]) ? node1550 : node1537;
					assign node1537 = (inp[5]) ? 3'b000 : node1538;
						assign node1538 = (inp[10]) ? 3'b000 : node1539;
							assign node1539 = (inp[1]) ? node1541 : 3'b000;
								assign node1541 = (inp[7]) ? node1543 : 3'b000;
									assign node1543 = (inp[6]) ? node1545 : 3'b000;
										assign node1545 = (inp[2]) ? 3'b100 : 3'b000;
					assign node1550 = (inp[6]) ? node1562 : node1551;
						assign node1551 = (inp[11]) ? 3'b000 : node1552;
							assign node1552 = (inp[7]) ? node1554 : 3'b000;
								assign node1554 = (inp[1]) ? node1556 : 3'b000;
									assign node1556 = (inp[10]) ? 3'b000 : node1557;
										assign node1557 = (inp[5]) ? 3'b000 : 3'b100;
						assign node1562 = (inp[10]) ? node1592 : node1563;
							assign node1563 = (inp[5]) ? node1579 : node1564;
								assign node1564 = (inp[7]) ? node1572 : node1565;
									assign node1565 = (inp[1]) ? node1569 : node1566;
										assign node1566 = (inp[8]) ? 3'b100 : 3'b000;
										assign node1569 = (inp[11]) ? 3'b100 : 3'b100;
									assign node1572 = (inp[11]) ? node1576 : node1573;
										assign node1573 = (inp[2]) ? 3'b010 : 3'b010;
										assign node1576 = (inp[1]) ? 3'b000 : 3'b100;
								assign node1579 = (inp[7]) ? node1585 : node1580;
									assign node1580 = (inp[11]) ? 3'b000 : node1581;
										assign node1581 = (inp[8]) ? 3'b000 : 3'b000;
									assign node1585 = (inp[1]) ? node1589 : node1586;
										assign node1586 = (inp[11]) ? 3'b000 : 3'b000;
										assign node1589 = (inp[2]) ? 3'b100 : 3'b100;
							assign node1592 = (inp[7]) ? node1600 : node1593;
								assign node1593 = (inp[8]) ? node1595 : 3'b000;
									assign node1595 = (inp[1]) ? node1597 : 3'b000;
										assign node1597 = (inp[11]) ? 3'b000 : 3'b000;
								assign node1600 = (inp[1]) ? node1606 : node1601;
									assign node1601 = (inp[5]) ? 3'b000 : node1602;
										assign node1602 = (inp[11]) ? 3'b000 : 3'b000;
									assign node1606 = (inp[5]) ? node1610 : node1607;
										assign node1607 = (inp[11]) ? 3'b100 : 3'b100;
										assign node1610 = (inp[2]) ? 3'b000 : 3'b000;

endmodule