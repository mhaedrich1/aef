module dtc_split125_bm24 (
	input  wire [13-1:0] inp,
	output wire [13-1:0] outp
);

	wire [13-1:0] node1;
	wire [13-1:0] node2;
	wire [13-1:0] node3;
	wire [13-1:0] node4;
	wire [13-1:0] node5;
	wire [13-1:0] node6;
	wire [13-1:0] node7;
	wire [13-1:0] node8;
	wire [13-1:0] node11;
	wire [13-1:0] node12;
	wire [13-1:0] node13;
	wire [13-1:0] node15;
	wire [13-1:0] node18;
	wire [13-1:0] node19;
	wire [13-1:0] node24;
	wire [13-1:0] node25;
	wire [13-1:0] node26;
	wire [13-1:0] node27;
	wire [13-1:0] node29;
	wire [13-1:0] node35;
	wire [13-1:0] node36;
	wire [13-1:0] node37;
	wire [13-1:0] node38;
	wire [13-1:0] node40;
	wire [13-1:0] node44;
	wire [13-1:0] node46;
	wire [13-1:0] node47;
	wire [13-1:0] node51;
	wire [13-1:0] node52;
	wire [13-1:0] node53;
	wire [13-1:0] node57;
	wire [13-1:0] node60;
	wire [13-1:0] node61;
	wire [13-1:0] node62;
	wire [13-1:0] node63;
	wire [13-1:0] node65;
	wire [13-1:0] node68;
	wire [13-1:0] node71;
	wire [13-1:0] node72;
	wire [13-1:0] node76;
	wire [13-1:0] node77;
	wire [13-1:0] node78;
	wire [13-1:0] node80;
	wire [13-1:0] node83;
	wire [13-1:0] node85;
	wire [13-1:0] node86;
	wire [13-1:0] node90;
	wire [13-1:0] node91;
	wire [13-1:0] node93;
	wire [13-1:0] node96;
	wire [13-1:0] node97;
	wire [13-1:0] node101;
	wire [13-1:0] node102;
	wire [13-1:0] node103;
	wire [13-1:0] node104;
	wire [13-1:0] node105;
	wire [13-1:0] node106;
	wire [13-1:0] node108;
	wire [13-1:0] node112;
	wire [13-1:0] node115;
	wire [13-1:0] node117;
	wire [13-1:0] node119;
	wire [13-1:0] node122;
	wire [13-1:0] node123;
	wire [13-1:0] node124;
	wire [13-1:0] node125;
	wire [13-1:0] node129;
	wire [13-1:0] node130;
	wire [13-1:0] node131;
	wire [13-1:0] node136;
	wire [13-1:0] node137;
	wire [13-1:0] node138;
	wire [13-1:0] node143;
	wire [13-1:0] node144;
	wire [13-1:0] node145;
	wire [13-1:0] node146;
	wire [13-1:0] node147;
	wire [13-1:0] node150;
	wire [13-1:0] node153;
	wire [13-1:0] node156;
	wire [13-1:0] node157;
	wire [13-1:0] node159;
	wire [13-1:0] node162;
	wire [13-1:0] node164;
	wire [13-1:0] node167;
	wire [13-1:0] node168;
	wire [13-1:0] node170;
	wire [13-1:0] node172;
	wire [13-1:0] node173;
	wire [13-1:0] node177;
	wire [13-1:0] node178;
	wire [13-1:0] node180;
	wire [13-1:0] node183;
	wire [13-1:0] node186;
	wire [13-1:0] node187;
	wire [13-1:0] node188;
	wire [13-1:0] node189;
	wire [13-1:0] node190;
	wire [13-1:0] node191;
	wire [13-1:0] node192;
	wire [13-1:0] node193;
	wire [13-1:0] node197;
	wire [13-1:0] node201;
	wire [13-1:0] node202;
	wire [13-1:0] node204;
	wire [13-1:0] node206;
	wire [13-1:0] node209;
	wire [13-1:0] node212;
	wire [13-1:0] node213;
	wire [13-1:0] node214;
	wire [13-1:0] node216;
	wire [13-1:0] node217;
	wire [13-1:0] node221;
	wire [13-1:0] node222;
	wire [13-1:0] node224;
	wire [13-1:0] node228;
	wire [13-1:0] node231;
	wire [13-1:0] node232;
	wire [13-1:0] node233;
	wire [13-1:0] node234;
	wire [13-1:0] node236;
	wire [13-1:0] node240;
	wire [13-1:0] node241;
	wire [13-1:0] node242;
	wire [13-1:0] node243;
	wire [13-1:0] node246;
	wire [13-1:0] node250;
	wire [13-1:0] node251;
	wire [13-1:0] node253;
	wire [13-1:0] node257;
	wire [13-1:0] node258;
	wire [13-1:0] node259;
	wire [13-1:0] node261;
	wire [13-1:0] node262;
	wire [13-1:0] node266;
	wire [13-1:0] node268;
	wire [13-1:0] node271;
	wire [13-1:0] node272;
	wire [13-1:0] node275;
	wire [13-1:0] node276;
	wire [13-1:0] node279;
	wire [13-1:0] node280;
	wire [13-1:0] node284;
	wire [13-1:0] node285;
	wire [13-1:0] node286;
	wire [13-1:0] node287;
	wire [13-1:0] node288;
	wire [13-1:0] node289;
	wire [13-1:0] node293;
	wire [13-1:0] node294;
	wire [13-1:0] node295;
	wire [13-1:0] node300;
	wire [13-1:0] node301;
	wire [13-1:0] node302;
	wire [13-1:0] node306;
	wire [13-1:0] node308;
	wire [13-1:0] node309;
	wire [13-1:0] node313;
	wire [13-1:0] node314;
	wire [13-1:0] node315;
	wire [13-1:0] node317;
	wire [13-1:0] node319;
	wire [13-1:0] node322;
	wire [13-1:0] node324;
	wire [13-1:0] node327;
	wire [13-1:0] node328;
	wire [13-1:0] node331;
	wire [13-1:0] node334;
	wire [13-1:0] node335;
	wire [13-1:0] node336;
	wire [13-1:0] node337;
	wire [13-1:0] node339;
	wire [13-1:0] node342;
	wire [13-1:0] node343;
	wire [13-1:0] node345;
	wire [13-1:0] node349;
	wire [13-1:0] node350;
	wire [13-1:0] node351;
	wire [13-1:0] node356;
	wire [13-1:0] node357;
	wire [13-1:0] node358;
	wire [13-1:0] node359;
	wire [13-1:0] node361;
	wire [13-1:0] node365;
	wire [13-1:0] node367;
	wire [13-1:0] node370;
	wire [13-1:0] node371;
	wire [13-1:0] node375;
	wire [13-1:0] node376;
	wire [13-1:0] node377;
	wire [13-1:0] node378;
	wire [13-1:0] node379;
	wire [13-1:0] node380;
	wire [13-1:0] node381;
	wire [13-1:0] node383;
	wire [13-1:0] node384;
	wire [13-1:0] node389;
	wire [13-1:0] node390;
	wire [13-1:0] node392;
	wire [13-1:0] node396;
	wire [13-1:0] node397;
	wire [13-1:0] node398;
	wire [13-1:0] node401;
	wire [13-1:0] node403;
	wire [13-1:0] node406;
	wire [13-1:0] node409;
	wire [13-1:0] node410;
	wire [13-1:0] node411;
	wire [13-1:0] node412;
	wire [13-1:0] node413;
	wire [13-1:0] node417;
	wire [13-1:0] node419;
	wire [13-1:0] node421;
	wire [13-1:0] node424;
	wire [13-1:0] node425;
	wire [13-1:0] node427;
	wire [13-1:0] node430;
	wire [13-1:0] node431;
	wire [13-1:0] node435;
	wire [13-1:0] node436;
	wire [13-1:0] node437;
	wire [13-1:0] node440;
	wire [13-1:0] node443;
	wire [13-1:0] node445;
	wire [13-1:0] node447;
	wire [13-1:0] node450;
	wire [13-1:0] node451;
	wire [13-1:0] node452;
	wire [13-1:0] node453;
	wire [13-1:0] node454;
	wire [13-1:0] node456;
	wire [13-1:0] node460;
	wire [13-1:0] node461;
	wire [13-1:0] node462;
	wire [13-1:0] node464;
	wire [13-1:0] node468;
	wire [13-1:0] node471;
	wire [13-1:0] node472;
	wire [13-1:0] node473;
	wire [13-1:0] node477;
	wire [13-1:0] node478;
	wire [13-1:0] node481;
	wire [13-1:0] node483;
	wire [13-1:0] node484;
	wire [13-1:0] node488;
	wire [13-1:0] node489;
	wire [13-1:0] node490;
	wire [13-1:0] node491;
	wire [13-1:0] node492;
	wire [13-1:0] node495;
	wire [13-1:0] node496;
	wire [13-1:0] node500;
	wire [13-1:0] node503;
	wire [13-1:0] node504;
	wire [13-1:0] node505;
	wire [13-1:0] node509;
	wire [13-1:0] node512;
	wire [13-1:0] node513;
	wire [13-1:0] node514;
	wire [13-1:0] node515;
	wire [13-1:0] node519;
	wire [13-1:0] node521;
	wire [13-1:0] node523;
	wire [13-1:0] node526;
	wire [13-1:0] node527;
	wire [13-1:0] node529;
	wire [13-1:0] node532;
	wire [13-1:0] node535;
	wire [13-1:0] node536;
	wire [13-1:0] node537;
	wire [13-1:0] node538;
	wire [13-1:0] node539;
	wire [13-1:0] node540;
	wire [13-1:0] node541;
	wire [13-1:0] node544;
	wire [13-1:0] node545;
	wire [13-1:0] node550;
	wire [13-1:0] node551;
	wire [13-1:0] node552;
	wire [13-1:0] node553;
	wire [13-1:0] node556;
	wire [13-1:0] node559;
	wire [13-1:0] node561;
	wire [13-1:0] node564;
	wire [13-1:0] node567;
	wire [13-1:0] node568;
	wire [13-1:0] node569;
	wire [13-1:0] node573;
	wire [13-1:0] node574;
	wire [13-1:0] node575;
	wire [13-1:0] node579;
	wire [13-1:0] node581;
	wire [13-1:0] node582;
	wire [13-1:0] node586;
	wire [13-1:0] node587;
	wire [13-1:0] node588;
	wire [13-1:0] node589;
	wire [13-1:0] node591;
	wire [13-1:0] node592;
	wire [13-1:0] node596;
	wire [13-1:0] node597;
	wire [13-1:0] node601;
	wire [13-1:0] node603;
	wire [13-1:0] node604;
	wire [13-1:0] node605;
	wire [13-1:0] node610;
	wire [13-1:0] node611;
	wire [13-1:0] node612;
	wire [13-1:0] node613;
	wire [13-1:0] node617;
	wire [13-1:0] node619;
	wire [13-1:0] node622;
	wire [13-1:0] node623;
	wire [13-1:0] node625;
	wire [13-1:0] node628;
	wire [13-1:0] node629;
	wire [13-1:0] node632;
	wire [13-1:0] node634;
	wire [13-1:0] node637;
	wire [13-1:0] node638;
	wire [13-1:0] node639;
	wire [13-1:0] node640;
	wire [13-1:0] node643;
	wire [13-1:0] node644;
	wire [13-1:0] node647;
	wire [13-1:0] node648;
	wire [13-1:0] node649;
	wire [13-1:0] node654;
	wire [13-1:0] node655;
	wire [13-1:0] node656;
	wire [13-1:0] node657;
	wire [13-1:0] node661;
	wire [13-1:0] node663;
	wire [13-1:0] node665;
	wire [13-1:0] node668;
	wire [13-1:0] node669;
	wire [13-1:0] node670;
	wire [13-1:0] node674;
	wire [13-1:0] node675;
	wire [13-1:0] node679;
	wire [13-1:0] node680;
	wire [13-1:0] node681;
	wire [13-1:0] node683;
	wire [13-1:0] node686;
	wire [13-1:0] node687;
	wire [13-1:0] node688;
	wire [13-1:0] node692;
	wire [13-1:0] node694;
	wire [13-1:0] node695;
	wire [13-1:0] node699;
	wire [13-1:0] node700;
	wire [13-1:0] node702;
	wire [13-1:0] node705;
	wire [13-1:0] node706;
	wire [13-1:0] node708;
	wire [13-1:0] node710;
	wire [13-1:0] node711;
	wire [13-1:0] node715;
	wire [13-1:0] node716;
	wire [13-1:0] node720;
	wire [13-1:0] node721;
	wire [13-1:0] node722;
	wire [13-1:0] node723;
	wire [13-1:0] node724;
	wire [13-1:0] node725;
	wire [13-1:0] node726;
	wire [13-1:0] node727;
	wire [13-1:0] node728;
	wire [13-1:0] node730;
	wire [13-1:0] node731;
	wire [13-1:0] node736;
	wire [13-1:0] node737;
	wire [13-1:0] node741;
	wire [13-1:0] node742;
	wire [13-1:0] node744;
	wire [13-1:0] node747;
	wire [13-1:0] node748;
	wire [13-1:0] node752;
	wire [13-1:0] node753;
	wire [13-1:0] node754;
	wire [13-1:0] node755;
	wire [13-1:0] node757;
	wire [13-1:0] node761;
	wire [13-1:0] node762;
	wire [13-1:0] node763;
	wire [13-1:0] node764;
	wire [13-1:0] node769;
	wire [13-1:0] node772;
	wire [13-1:0] node773;
	wire [13-1:0] node775;
	wire [13-1:0] node778;
	wire [13-1:0] node781;
	wire [13-1:0] node782;
	wire [13-1:0] node783;
	wire [13-1:0] node784;
	wire [13-1:0] node785;
	wire [13-1:0] node786;
	wire [13-1:0] node789;
	wire [13-1:0] node792;
	wire [13-1:0] node795;
	wire [13-1:0] node798;
	wire [13-1:0] node801;
	wire [13-1:0] node802;
	wire [13-1:0] node803;
	wire [13-1:0] node805;
	wire [13-1:0] node808;
	wire [13-1:0] node811;
	wire [13-1:0] node812;
	wire [13-1:0] node813;
	wire [13-1:0] node817;
	wire [13-1:0] node820;
	wire [13-1:0] node821;
	wire [13-1:0] node822;
	wire [13-1:0] node823;
	wire [13-1:0] node824;
	wire [13-1:0] node825;
	wire [13-1:0] node826;
	wire [13-1:0] node831;
	wire [13-1:0] node832;
	wire [13-1:0] node833;
	wire [13-1:0] node838;
	wire [13-1:0] node839;
	wire [13-1:0] node840;
	wire [13-1:0] node842;
	wire [13-1:0] node846;
	wire [13-1:0] node849;
	wire [13-1:0] node850;
	wire [13-1:0] node851;
	wire [13-1:0] node852;
	wire [13-1:0] node854;
	wire [13-1:0] node857;
	wire [13-1:0] node858;
	wire [13-1:0] node860;
	wire [13-1:0] node864;
	wire [13-1:0] node867;
	wire [13-1:0] node868;
	wire [13-1:0] node870;
	wire [13-1:0] node873;
	wire [13-1:0] node876;
	wire [13-1:0] node877;
	wire [13-1:0] node878;
	wire [13-1:0] node879;
	wire [13-1:0] node881;
	wire [13-1:0] node882;
	wire [13-1:0] node886;
	wire [13-1:0] node887;
	wire [13-1:0] node889;
	wire [13-1:0] node893;
	wire [13-1:0] node894;
	wire [13-1:0] node896;
	wire [13-1:0] node897;
	wire [13-1:0] node901;
	wire [13-1:0] node902;
	wire [13-1:0] node903;
	wire [13-1:0] node905;
	wire [13-1:0] node909;
	wire [13-1:0] node912;
	wire [13-1:0] node913;
	wire [13-1:0] node914;
	wire [13-1:0] node916;
	wire [13-1:0] node919;
	wire [13-1:0] node922;
	wire [13-1:0] node923;
	wire [13-1:0] node924;
	wire [13-1:0] node926;
	wire [13-1:0] node930;
	wire [13-1:0] node931;
	wire [13-1:0] node933;
	wire [13-1:0] node934;
	wire [13-1:0] node939;
	wire [13-1:0] node940;
	wire [13-1:0] node941;
	wire [13-1:0] node942;
	wire [13-1:0] node943;
	wire [13-1:0] node944;
	wire [13-1:0] node946;
	wire [13-1:0] node949;
	wire [13-1:0] node951;
	wire [13-1:0] node954;
	wire [13-1:0] node955;
	wire [13-1:0] node958;
	wire [13-1:0] node961;
	wire [13-1:0] node962;
	wire [13-1:0] node963;
	wire [13-1:0] node966;
	wire [13-1:0] node968;
	wire [13-1:0] node971;
	wire [13-1:0] node973;
	wire [13-1:0] node975;
	wire [13-1:0] node977;
	wire [13-1:0] node978;
	wire [13-1:0] node982;
	wire [13-1:0] node983;
	wire [13-1:0] node984;
	wire [13-1:0] node985;
	wire [13-1:0] node986;
	wire [13-1:0] node988;
	wire [13-1:0] node992;
	wire [13-1:0] node994;
	wire [13-1:0] node997;
	wire [13-1:0] node1000;
	wire [13-1:0] node1001;
	wire [13-1:0] node1002;
	wire [13-1:0] node1006;
	wire [13-1:0] node1007;
	wire [13-1:0] node1010;
	wire [13-1:0] node1011;
	wire [13-1:0] node1013;
	wire [13-1:0] node1014;
	wire [13-1:0] node1017;
	wire [13-1:0] node1021;
	wire [13-1:0] node1022;
	wire [13-1:0] node1023;
	wire [13-1:0] node1024;
	wire [13-1:0] node1025;
	wire [13-1:0] node1029;
	wire [13-1:0] node1030;
	wire [13-1:0] node1032;
	wire [13-1:0] node1035;
	wire [13-1:0] node1036;
	wire [13-1:0] node1040;
	wire [13-1:0] node1041;
	wire [13-1:0] node1042;
	wire [13-1:0] node1043;
	wire [13-1:0] node1047;
	wire [13-1:0] node1049;
	wire [13-1:0] node1052;
	wire [13-1:0] node1053;
	wire [13-1:0] node1055;
	wire [13-1:0] node1057;
	wire [13-1:0] node1060;
	wire [13-1:0] node1062;
	wire [13-1:0] node1065;
	wire [13-1:0] node1066;
	wire [13-1:0] node1069;
	wire [13-1:0] node1070;
	wire [13-1:0] node1071;
	wire [13-1:0] node1072;
	wire [13-1:0] node1074;
	wire [13-1:0] node1078;
	wire [13-1:0] node1079;
	wire [13-1:0] node1083;
	wire [13-1:0] node1084;
	wire [13-1:0] node1088;
	wire [13-1:0] node1089;
	wire [13-1:0] node1090;
	wire [13-1:0] node1091;
	wire [13-1:0] node1092;
	wire [13-1:0] node1093;
	wire [13-1:0] node1094;
	wire [13-1:0] node1096;
	wire [13-1:0] node1097;
	wire [13-1:0] node1099;
	wire [13-1:0] node1103;
	wire [13-1:0] node1104;
	wire [13-1:0] node1108;
	wire [13-1:0] node1109;
	wire [13-1:0] node1111;
	wire [13-1:0] node1114;
	wire [13-1:0] node1117;
	wire [13-1:0] node1118;
	wire [13-1:0] node1119;
	wire [13-1:0] node1120;
	wire [13-1:0] node1121;
	wire [13-1:0] node1126;
	wire [13-1:0] node1127;
	wire [13-1:0] node1128;
	wire [13-1:0] node1133;
	wire [13-1:0] node1134;
	wire [13-1:0] node1138;
	wire [13-1:0] node1139;
	wire [13-1:0] node1140;
	wire [13-1:0] node1142;
	wire [13-1:0] node1145;
	wire [13-1:0] node1146;
	wire [13-1:0] node1148;
	wire [13-1:0] node1149;
	wire [13-1:0] node1153;
	wire [13-1:0] node1155;
	wire [13-1:0] node1157;
	wire [13-1:0] node1160;
	wire [13-1:0] node1161;
	wire [13-1:0] node1162;
	wire [13-1:0] node1163;
	wire [13-1:0] node1166;
	wire [13-1:0] node1168;
	wire [13-1:0] node1172;
	wire [13-1:0] node1173;
	wire [13-1:0] node1174;
	wire [13-1:0] node1177;
	wire [13-1:0] node1178;
	wire [13-1:0] node1183;
	wire [13-1:0] node1184;
	wire [13-1:0] node1185;
	wire [13-1:0] node1186;
	wire [13-1:0] node1187;
	wire [13-1:0] node1188;
	wire [13-1:0] node1192;
	wire [13-1:0] node1193;
	wire [13-1:0] node1195;
	wire [13-1:0] node1199;
	wire [13-1:0] node1202;
	wire [13-1:0] node1203;
	wire [13-1:0] node1205;
	wire [13-1:0] node1206;
	wire [13-1:0] node1210;
	wire [13-1:0] node1211;
	wire [13-1:0] node1212;
	wire [13-1:0] node1216;
	wire [13-1:0] node1218;
	wire [13-1:0] node1221;
	wire [13-1:0] node1222;
	wire [13-1:0] node1223;
	wire [13-1:0] node1224;
	wire [13-1:0] node1227;
	wire [13-1:0] node1229;
	wire [13-1:0] node1230;
	wire [13-1:0] node1233;
	wire [13-1:0] node1236;
	wire [13-1:0] node1238;
	wire [13-1:0] node1239;
	wire [13-1:0] node1243;
	wire [13-1:0] node1244;
	wire [13-1:0] node1247;
	wire [13-1:0] node1248;
	wire [13-1:0] node1250;
	wire [13-1:0] node1252;
	wire [13-1:0] node1255;
	wire [13-1:0] node1256;
	wire [13-1:0] node1259;
	wire [13-1:0] node1260;
	wire [13-1:0] node1262;
	wire [13-1:0] node1266;
	wire [13-1:0] node1267;
	wire [13-1:0] node1268;
	wire [13-1:0] node1269;
	wire [13-1:0] node1270;
	wire [13-1:0] node1271;
	wire [13-1:0] node1272;
	wire [13-1:0] node1276;
	wire [13-1:0] node1277;
	wire [13-1:0] node1278;
	wire [13-1:0] node1283;
	wire [13-1:0] node1284;
	wire [13-1:0] node1286;
	wire [13-1:0] node1287;
	wire [13-1:0] node1291;
	wire [13-1:0] node1293;
	wire [13-1:0] node1296;
	wire [13-1:0] node1297;
	wire [13-1:0] node1298;
	wire [13-1:0] node1299;
	wire [13-1:0] node1302;
	wire [13-1:0] node1305;
	wire [13-1:0] node1307;
	wire [13-1:0] node1309;
	wire [13-1:0] node1313;
	wire [13-1:0] node1314;
	wire [13-1:0] node1315;
	wire [13-1:0] node1317;
	wire [13-1:0] node1320;
	wire [13-1:0] node1321;
	wire [13-1:0] node1322;
	wire [13-1:0] node1323;
	wire [13-1:0] node1326;
	wire [13-1:0] node1329;
	wire [13-1:0] node1332;
	wire [13-1:0] node1333;
	wire [13-1:0] node1336;
	wire [13-1:0] node1339;
	wire [13-1:0] node1341;
	wire [13-1:0] node1342;
	wire [13-1:0] node1343;
	wire [13-1:0] node1344;
	wire [13-1:0] node1346;
	wire [13-1:0] node1351;
	wire [13-1:0] node1352;
	wire [13-1:0] node1356;
	wire [13-1:0] node1357;
	wire [13-1:0] node1358;
	wire [13-1:0] node1359;
	wire [13-1:0] node1360;
	wire [13-1:0] node1364;
	wire [13-1:0] node1365;
	wire [13-1:0] node1366;
	wire [13-1:0] node1369;
	wire [13-1:0] node1372;
	wire [13-1:0] node1373;
	wire [13-1:0] node1377;
	wire [13-1:0] node1378;
	wire [13-1:0] node1379;
	wire [13-1:0] node1382;
	wire [13-1:0] node1384;
	wire [13-1:0] node1386;
	wire [13-1:0] node1389;
	wire [13-1:0] node1390;
	wire [13-1:0] node1392;
	wire [13-1:0] node1394;
	wire [13-1:0] node1397;
	wire [13-1:0] node1400;
	wire [13-1:0] node1401;
	wire [13-1:0] node1402;
	wire [13-1:0] node1403;
	wire [13-1:0] node1404;
	wire [13-1:0] node1408;
	wire [13-1:0] node1409;
	wire [13-1:0] node1411;
	wire [13-1:0] node1415;
	wire [13-1:0] node1416;
	wire [13-1:0] node1417;
	wire [13-1:0] node1421;
	wire [13-1:0] node1424;
	wire [13-1:0] node1425;
	wire [13-1:0] node1428;
	wire [13-1:0] node1429;
	wire [13-1:0] node1430;
	wire [13-1:0] node1434;
	wire [13-1:0] node1435;

	assign outp = (inp[4]) ? node720 : node1;
		assign node1 = (inp[5]) ? node375 : node2;
			assign node2 = (inp[6]) ? node186 : node3;
				assign node3 = (inp[8]) ? node101 : node4;
					assign node4 = (inp[2]) ? node60 : node5;
						assign node5 = (inp[12]) ? node35 : node6;
							assign node6 = (inp[7]) ? node24 : node7;
								assign node7 = (inp[9]) ? node11 : node8;
									assign node8 = (inp[3]) ? 13'b0001111111111 : 13'b0011111111111;
									assign node11 = (inp[0]) ? 13'b0000111111111 : node12;
										assign node12 = (inp[10]) ? node18 : node13;
											assign node13 = (inp[11]) ? node15 : 13'b0001111111111;
												assign node15 = (inp[3]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node18 = (inp[3]) ? 13'b0001111111111 : node19;
												assign node19 = (inp[11]) ? 13'b0001111111111 : 13'b0011111111111;
								assign node24 = (inp[10]) ? 13'b0000111111111 : node25;
									assign node25 = (inp[9]) ? 13'b0000111111111 : node26;
										assign node26 = (inp[3]) ? 13'b0001111111111 : node27;
											assign node27 = (inp[0]) ? node29 : 13'b0011111111111;
												assign node29 = (inp[11]) ? 13'b0001111111111 : 13'b0011111111111;
							assign node35 = (inp[3]) ? node51 : node36;
								assign node36 = (inp[0]) ? node44 : node37;
									assign node37 = (inp[10]) ? 13'b0000111111111 : node38;
										assign node38 = (inp[11]) ? node40 : 13'b0001111111111;
											assign node40 = (inp[7]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node44 = (inp[7]) ? node46 : 13'b0000111111111;
										assign node46 = (inp[9]) ? 13'b0000011111111 : node47;
											assign node47 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node51 = (inp[10]) ? node57 : node52;
									assign node52 = (inp[11]) ? 13'b0000011111111 : node53;
										assign node53 = (inp[7]) ? 13'b0001111111111 : 13'b0000111111111;
									assign node57 = (inp[1]) ? 13'b0000001111111 : 13'b0000011111111;
						assign node60 = (inp[11]) ? node76 : node61;
							assign node61 = (inp[7]) ? node71 : node62;
								assign node62 = (inp[0]) ? node68 : node63;
									assign node63 = (inp[9]) ? node65 : 13'b0001111111111;
										assign node65 = (inp[3]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node68 = (inp[9]) ? 13'b0000111111111 : 13'b0000011111111;
								assign node71 = (inp[9]) ? 13'b0000011111111 : node72;
									assign node72 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node76 = (inp[12]) ? node90 : node77;
								assign node77 = (inp[1]) ? node83 : node78;
									assign node78 = (inp[9]) ? node80 : 13'b0000111111111;
										assign node80 = (inp[0]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node83 = (inp[0]) ? node85 : 13'b0000011111111;
										assign node85 = (inp[3]) ? 13'b0000001111111 : node86;
											assign node86 = (inp[9]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node90 = (inp[7]) ? node96 : node91;
									assign node91 = (inp[9]) ? node93 : 13'b0000111111111;
										assign node93 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node96 = (inp[0]) ? 13'b0000000011111 : node97;
										assign node97 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
					assign node101 = (inp[10]) ? node143 : node102;
						assign node102 = (inp[1]) ? node122 : node103;
							assign node103 = (inp[0]) ? node115 : node104;
								assign node104 = (inp[3]) ? node112 : node105;
									assign node105 = (inp[2]) ? 13'b0000111111111 : node106;
										assign node106 = (inp[7]) ? node108 : 13'b0011111111111;
											assign node108 = (inp[9]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node112 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node115 = (inp[7]) ? node117 : 13'b0000111111111;
									assign node117 = (inp[12]) ? node119 : 13'b0000011111111;
										assign node119 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node122 = (inp[3]) ? node136 : node123;
								assign node123 = (inp[7]) ? node129 : node124;
									assign node124 = (inp[9]) ? 13'b0000011111111 : node125;
										assign node125 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node129 = (inp[0]) ? 13'b0000011111111 : node130;
										assign node130 = (inp[12]) ? 13'b0000001111111 : node131;
											assign node131 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node136 = (inp[7]) ? 13'b0000000111111 : node137;
									assign node137 = (inp[9]) ? 13'b0000001111111 : node138;
										assign node138 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
						assign node143 = (inp[7]) ? node167 : node144;
							assign node144 = (inp[1]) ? node156 : node145;
								assign node145 = (inp[0]) ? node153 : node146;
									assign node146 = (inp[2]) ? node150 : node147;
										assign node147 = (inp[12]) ? 13'b0000111111111 : 13'b0001111111111;
										assign node150 = (inp[9]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node153 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node156 = (inp[2]) ? node162 : node157;
									assign node157 = (inp[11]) ? node159 : 13'b0000011111111;
										assign node159 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node162 = (inp[3]) ? node164 : 13'b0000001111111;
										assign node164 = (inp[0]) ? 13'b0000000111111 : 13'b0000000011111;
							assign node167 = (inp[1]) ? node177 : node168;
								assign node168 = (inp[3]) ? node170 : 13'b0000001111111;
									assign node170 = (inp[12]) ? node172 : 13'b0000001111111;
										assign node172 = (inp[9]) ? 13'b0000000111111 : node173;
											assign node173 = (inp[0]) ? 13'b0000000111111 : 13'b0000011111111;
								assign node177 = (inp[0]) ? node183 : node178;
									assign node178 = (inp[2]) ? node180 : 13'b0000011111111;
										assign node180 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node183 = (inp[3]) ? 13'b0000000111111 : 13'b0000000011111;
				assign node186 = (inp[1]) ? node284 : node187;
					assign node187 = (inp[12]) ? node231 : node188;
						assign node188 = (inp[9]) ? node212 : node189;
							assign node189 = (inp[2]) ? node201 : node190;
								assign node190 = (inp[8]) ? 13'b0000011111111 : node191;
									assign node191 = (inp[3]) ? node197 : node192;
										assign node192 = (inp[0]) ? 13'b0001111111111 : node193;
											assign node193 = (inp[7]) ? 13'b0001111111111 : 13'b0011111111111;
										assign node197 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
								assign node201 = (inp[7]) ? node209 : node202;
									assign node202 = (inp[3]) ? node204 : 13'b0000111111111;
										assign node204 = (inp[11]) ? node206 : 13'b0000011111111;
											assign node206 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node209 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node212 = (inp[7]) ? node228 : node213;
								assign node213 = (inp[11]) ? node221 : node214;
									assign node214 = (inp[0]) ? node216 : 13'b0000111111111;
										assign node216 = (inp[3]) ? 13'b0000011111111 : node217;
											assign node217 = (inp[10]) ? 13'b0000011111111 : 13'b0001111111111;
									assign node221 = (inp[8]) ? 13'b0000001111111 : node222;
										assign node222 = (inp[0]) ? node224 : 13'b0000011111111;
											assign node224 = (inp[3]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node228 = (inp[2]) ? 13'b0000000111111 : 13'b0000001111111;
						assign node231 = (inp[9]) ? node257 : node232;
							assign node232 = (inp[8]) ? node240 : node233;
								assign node233 = (inp[10]) ? 13'b0000011111111 : node234;
									assign node234 = (inp[2]) ? node236 : 13'b0000111111111;
										assign node236 = (inp[3]) ? 13'b0000011111111 : 13'b0001111111111;
								assign node240 = (inp[0]) ? node250 : node241;
									assign node241 = (inp[2]) ? 13'b0000001111111 : node242;
										assign node242 = (inp[11]) ? node246 : node243;
											assign node243 = (inp[3]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node246 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node250 = (inp[3]) ? 13'b0000000111111 : node251;
										assign node251 = (inp[7]) ? node253 : 13'b0000001111111;
											assign node253 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node257 = (inp[2]) ? node271 : node258;
								assign node258 = (inp[8]) ? node266 : node259;
									assign node259 = (inp[10]) ? node261 : 13'b0000011111111;
										assign node261 = (inp[11]) ? 13'b0000001111111 : node262;
											assign node262 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node266 = (inp[3]) ? node268 : 13'b0000011111111;
										assign node268 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node271 = (inp[3]) ? node275 : node272;
									assign node272 = (inp[10]) ? 13'b0000001111111 : 13'b0000000111111;
									assign node275 = (inp[10]) ? node279 : node276;
										assign node276 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node279 = (inp[7]) ? 13'b0000000011111 : node280;
											assign node280 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node284 = (inp[2]) ? node334 : node285;
						assign node285 = (inp[0]) ? node313 : node286;
							assign node286 = (inp[3]) ? node300 : node287;
								assign node287 = (inp[9]) ? node293 : node288;
									assign node288 = (inp[11]) ? 13'b0000011111111 : node289;
										assign node289 = (inp[7]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node293 = (inp[12]) ? 13'b0000001111111 : node294;
										assign node294 = (inp[10]) ? 13'b0000011111111 : node295;
											assign node295 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node300 = (inp[12]) ? node306 : node301;
									assign node301 = (inp[8]) ? 13'b0000001111111 : node302;
										assign node302 = (inp[7]) ? 13'b0000001111111 : 13'b0000111111111;
									assign node306 = (inp[11]) ? node308 : 13'b0000011111111;
										assign node308 = (inp[7]) ? 13'b0000000111111 : node309;
											assign node309 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node313 = (inp[8]) ? node327 : node314;
								assign node314 = (inp[7]) ? node322 : node315;
									assign node315 = (inp[3]) ? node317 : 13'b0000001111111;
										assign node317 = (inp[10]) ? node319 : 13'b0000111111111;
											assign node319 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node322 = (inp[10]) ? node324 : 13'b0000001111111;
										assign node324 = (inp[3]) ? 13'b0000001111111 : 13'b0000000111111;
								assign node327 = (inp[9]) ? node331 : node328;
									assign node328 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node331 = (inp[7]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node334 = (inp[10]) ? node356 : node335;
							assign node335 = (inp[7]) ? node349 : node336;
								assign node336 = (inp[8]) ? node342 : node337;
									assign node337 = (inp[3]) ? node339 : 13'b0000011111111;
										assign node339 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node342 = (inp[9]) ? 13'b0000000001111 : node343;
										assign node343 = (inp[11]) ? node345 : 13'b0000001111111;
											assign node345 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node349 = (inp[3]) ? 13'b0000000111111 : node350;
									assign node350 = (inp[0]) ? 13'b0000000111111 : node351;
										assign node351 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node356 = (inp[9]) ? node370 : node357;
								assign node357 = (inp[12]) ? node365 : node358;
									assign node358 = (inp[3]) ? 13'b0000000111111 : node359;
										assign node359 = (inp[0]) ? node361 : 13'b0000001111111;
											assign node361 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node365 = (inp[11]) ? node367 : 13'b0000000111111;
										assign node367 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node370 = (inp[0]) ? 13'b0000000011111 : node371;
									assign node371 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
			assign node375 = (inp[11]) ? node535 : node376;
				assign node376 = (inp[6]) ? node450 : node377;
					assign node377 = (inp[3]) ? node409 : node378;
						assign node378 = (inp[9]) ? node396 : node379;
							assign node379 = (inp[0]) ? node389 : node380;
								assign node380 = (inp[1]) ? 13'b0000111111111 : node381;
									assign node381 = (inp[8]) ? node383 : 13'b0111111111111;
										assign node383 = (inp[7]) ? 13'b0000111111111 : node384;
											assign node384 = (inp[10]) ? 13'b0000111111111 : 13'b0001111111111;
								assign node389 = (inp[8]) ? 13'b0000011111111 : node390;
									assign node390 = (inp[10]) ? node392 : 13'b0001111111111;
										assign node392 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
							assign node396 = (inp[7]) ? node406 : node397;
								assign node397 = (inp[10]) ? node401 : node398;
									assign node398 = (inp[0]) ? 13'b0000111111111 : 13'b0000011111111;
									assign node401 = (inp[2]) ? node403 : 13'b0000011111111;
										assign node403 = (inp[12]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node406 = (inp[10]) ? 13'b0000001111111 : 13'b0000011111111;
						assign node409 = (inp[12]) ? node435 : node410;
							assign node410 = (inp[1]) ? node424 : node411;
								assign node411 = (inp[2]) ? node417 : node412;
									assign node412 = (inp[10]) ? 13'b0000111111111 : node413;
										assign node413 = (inp[9]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node417 = (inp[8]) ? node419 : 13'b0000111111111;
										assign node419 = (inp[7]) ? node421 : 13'b0000011111111;
											assign node421 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node424 = (inp[0]) ? node430 : node425;
									assign node425 = (inp[8]) ? node427 : 13'b0000011111111;
										assign node427 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node430 = (inp[10]) ? 13'b0000001111111 : node431;
										assign node431 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node435 = (inp[2]) ? node443 : node436;
								assign node436 = (inp[0]) ? node440 : node437;
									assign node437 = (inp[7]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node440 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node443 = (inp[7]) ? node445 : 13'b0000000111111;
									assign node445 = (inp[8]) ? node447 : 13'b0000000011111;
										assign node447 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node450 = (inp[3]) ? node488 : node451;
						assign node451 = (inp[7]) ? node471 : node452;
							assign node452 = (inp[2]) ? node460 : node453;
								assign node453 = (inp[9]) ? 13'b0000011111111 : node454;
									assign node454 = (inp[10]) ? node456 : 13'b0000111111111;
										assign node456 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node460 = (inp[8]) ? node468 : node461;
									assign node461 = (inp[9]) ? 13'b0000001111111 : node462;
										assign node462 = (inp[0]) ? node464 : 13'b0000011111111;
											assign node464 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node468 = (inp[10]) ? 13'b0000000001111 : 13'b0000001111111;
							assign node471 = (inp[12]) ? node477 : node472;
								assign node472 = (inp[8]) ? 13'b0000001111111 : node473;
									assign node473 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node477 = (inp[0]) ? node481 : node478;
									assign node478 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node481 = (inp[9]) ? node483 : 13'b0000000111111;
										assign node483 = (inp[8]) ? 13'b0000000001111 : node484;
											assign node484 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node488 = (inp[1]) ? node512 : node489;
							assign node489 = (inp[8]) ? node503 : node490;
								assign node490 = (inp[0]) ? node500 : node491;
									assign node491 = (inp[9]) ? node495 : node492;
										assign node492 = (inp[2]) ? 13'b0000111111111 : 13'b0000011111111;
										assign node495 = (inp[7]) ? 13'b0000001111111 : node496;
											assign node496 = (inp[2]) ? 13'b0000011111111 : 13'b0000001111111;
									assign node500 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node503 = (inp[10]) ? node509 : node504;
									assign node504 = (inp[9]) ? 13'b0000000111111 : node505;
										assign node505 = (inp[7]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node509 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node512 = (inp[0]) ? node526 : node513;
								assign node513 = (inp[12]) ? node519 : node514;
									assign node514 = (inp[2]) ? 13'b0000000111111 : node515;
										assign node515 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node519 = (inp[8]) ? node521 : 13'b0000011111111;
										assign node521 = (inp[7]) ? node523 : 13'b0000000011111;
											assign node523 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node526 = (inp[7]) ? node532 : node527;
									assign node527 = (inp[10]) ? node529 : 13'b0000000111111;
										assign node529 = (inp[8]) ? 13'b0000000001111 : 13'b0000000111111;
									assign node532 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
				assign node535 = (inp[3]) ? node637 : node536;
					assign node536 = (inp[1]) ? node586 : node537;
						assign node537 = (inp[9]) ? node567 : node538;
							assign node538 = (inp[12]) ? node550 : node539;
								assign node539 = (inp[2]) ? 13'b0000011111111 : node540;
									assign node540 = (inp[6]) ? node544 : node541;
										assign node541 = (inp[8]) ? 13'b0001111111111 : 13'b0000111111111;
										assign node544 = (inp[10]) ? 13'b0000001111111 : node545;
											assign node545 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node550 = (inp[6]) ? node564 : node551;
									assign node551 = (inp[10]) ? node559 : node552;
										assign node552 = (inp[2]) ? node556 : node553;
											assign node553 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
											assign node556 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node559 = (inp[2]) ? node561 : 13'b0000001111111;
											assign node561 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node564 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node567 = (inp[8]) ? node573 : node568;
								assign node568 = (inp[7]) ? 13'b0000000111111 : node569;
									assign node569 = (inp[12]) ? 13'b0000001111111 : 13'b0000111111111;
								assign node573 = (inp[6]) ? node579 : node574;
									assign node574 = (inp[0]) ? 13'b0000000111111 : node575;
										assign node575 = (inp[2]) ? 13'b0000000111111 : 13'b0000011111111;
									assign node579 = (inp[2]) ? node581 : 13'b0000000111111;
										assign node581 = (inp[10]) ? 13'b0000000001111 : node582;
											assign node582 = (inp[7]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node586 = (inp[9]) ? node610 : node587;
							assign node587 = (inp[7]) ? node601 : node588;
								assign node588 = (inp[0]) ? node596 : node589;
									assign node589 = (inp[12]) ? node591 : 13'b0000111111111;
										assign node591 = (inp[6]) ? 13'b0000001111111 : node592;
											assign node592 = (inp[2]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node596 = (inp[10]) ? 13'b0000001111111 : node597;
										assign node597 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node601 = (inp[2]) ? node603 : 13'b0000000111111;
									assign node603 = (inp[10]) ? 13'b0000000011111 : node604;
										assign node604 = (inp[6]) ? 13'b0000000111111 : node605;
											assign node605 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node610 = (inp[12]) ? node622 : node611;
								assign node611 = (inp[10]) ? node617 : node612;
									assign node612 = (inp[6]) ? 13'b0000000111111 : node613;
										assign node613 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node617 = (inp[0]) ? node619 : 13'b0000000111111;
										assign node619 = (inp[2]) ? 13'b0000000011111 : 13'b0000000001111;
								assign node622 = (inp[0]) ? node628 : node623;
									assign node623 = (inp[7]) ? node625 : 13'b0000000111111;
										assign node625 = (inp[8]) ? 13'b0000000001111 : 13'b0000000111111;
									assign node628 = (inp[6]) ? node632 : node629;
										assign node629 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node632 = (inp[10]) ? node634 : 13'b0000000001111;
											assign node634 = (inp[8]) ? 13'b0000000000111 : 13'b0000000001111;
					assign node637 = (inp[12]) ? node679 : node638;
						assign node638 = (inp[1]) ? node654 : node639;
							assign node639 = (inp[7]) ? node643 : node640;
								assign node640 = (inp[6]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node643 = (inp[0]) ? node647 : node644;
									assign node644 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node647 = (inp[6]) ? 13'b0000000011111 : node648;
										assign node648 = (inp[10]) ? 13'b0000000111111 : node649;
											assign node649 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node654 = (inp[6]) ? node668 : node655;
								assign node655 = (inp[10]) ? node661 : node656;
									assign node656 = (inp[2]) ? 13'b0000000111111 : node657;
										assign node657 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node661 = (inp[0]) ? node663 : 13'b0000000111111;
										assign node663 = (inp[9]) ? node665 : 13'b0000000111111;
											assign node665 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node668 = (inp[8]) ? node674 : node669;
									assign node669 = (inp[7]) ? 13'b0000000001111 : node670;
										assign node670 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node674 = (inp[9]) ? 13'b0000000000111 : node675;
										assign node675 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node679 = (inp[6]) ? node699 : node680;
							assign node680 = (inp[9]) ? node686 : node681;
								assign node681 = (inp[1]) ? node683 : 13'b0000000111111;
									assign node683 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node686 = (inp[7]) ? node692 : node687;
									assign node687 = (inp[10]) ? 13'b0000000011111 : node688;
										assign node688 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node692 = (inp[8]) ? node694 : 13'b0000000011111;
										assign node694 = (inp[1]) ? 13'b0000000001111 : node695;
											assign node695 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node699 = (inp[7]) ? node705 : node700;
								assign node700 = (inp[8]) ? node702 : 13'b0000001111111;
									assign node702 = (inp[2]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node705 = (inp[1]) ? node715 : node706;
									assign node706 = (inp[8]) ? node708 : 13'b0000000001111;
										assign node708 = (inp[0]) ? node710 : 13'b0000000001111;
											assign node710 = (inp[9]) ? 13'b0000000000111 : node711;
												assign node711 = (inp[10]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node715 = (inp[9]) ? 13'b0000000000111 : node716;
										assign node716 = (inp[0]) ? 13'b0000000000111 : 13'b0000000001111;
		assign node720 = (inp[7]) ? node1088 : node721;
			assign node721 = (inp[5]) ? node939 : node722;
				assign node722 = (inp[11]) ? node820 : node723;
					assign node723 = (inp[3]) ? node781 : node724;
						assign node724 = (inp[0]) ? node752 : node725;
							assign node725 = (inp[9]) ? node741 : node726;
								assign node726 = (inp[8]) ? node736 : node727;
									assign node727 = (inp[2]) ? 13'b0001111111111 : node728;
										assign node728 = (inp[6]) ? node730 : 13'b0011111111111;
											assign node730 = (inp[12]) ? 13'b0001111111111 : node731;
												assign node731 = (inp[1]) ? 13'b0001111111111 : 13'b0011111111111;
									assign node736 = (inp[12]) ? 13'b0000011111111 : node737;
										assign node737 = (inp[2]) ? 13'b0000111111111 : 13'b0001111111111;
								assign node741 = (inp[6]) ? node747 : node742;
									assign node742 = (inp[10]) ? node744 : 13'b0001111111111;
										assign node744 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node747 = (inp[1]) ? 13'b0000000111111 : node748;
										assign node748 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node752 = (inp[6]) ? node772 : node753;
								assign node753 = (inp[1]) ? node761 : node754;
									assign node754 = (inp[10]) ? 13'b0000011111111 : node755;
										assign node755 = (inp[9]) ? node757 : 13'b0001111111111;
											assign node757 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node761 = (inp[10]) ? node769 : node762;
										assign node762 = (inp[8]) ? 13'b0000001111111 : node763;
											assign node763 = (inp[9]) ? 13'b0000011111111 : node764;
												assign node764 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node769 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node772 = (inp[12]) ? node778 : node773;
									assign node773 = (inp[1]) ? node775 : 13'b0000001111111;
										assign node775 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node778 = (inp[10]) ? 13'b0000001111111 : 13'b0000000111111;
						assign node781 = (inp[12]) ? node801 : node782;
							assign node782 = (inp[9]) ? node798 : node783;
								assign node783 = (inp[6]) ? node795 : node784;
									assign node784 = (inp[10]) ? node792 : node785;
										assign node785 = (inp[1]) ? node789 : node786;
											assign node786 = (inp[0]) ? 13'b0000111111111 : 13'b0001111111111;
											assign node789 = (inp[8]) ? 13'b0000011111111 : 13'b0000111111111;
										assign node792 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node795 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node798 = (inp[1]) ? 13'b0000001111111 : 13'b0000000111111;
							assign node801 = (inp[8]) ? node811 : node802;
								assign node802 = (inp[2]) ? node808 : node803;
									assign node803 = (inp[1]) ? node805 : 13'b0000011111111;
										assign node805 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node808 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node811 = (inp[6]) ? node817 : node812;
									assign node812 = (inp[9]) ? 13'b0000000111111 : node813;
										assign node813 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node817 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node820 = (inp[6]) ? node876 : node821;
						assign node821 = (inp[3]) ? node849 : node822;
							assign node822 = (inp[10]) ? node838 : node823;
								assign node823 = (inp[8]) ? node831 : node824;
									assign node824 = (inp[2]) ? 13'b0000111111111 : node825;
										assign node825 = (inp[12]) ? 13'b0000111111111 : node826;
											assign node826 = (inp[1]) ? 13'b0000111111111 : 13'b0011111111111;
									assign node831 = (inp[9]) ? 13'b0000001111111 : node832;
										assign node832 = (inp[12]) ? 13'b0000001111111 : node833;
											assign node833 = (inp[2]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node838 = (inp[12]) ? node846 : node839;
									assign node839 = (inp[2]) ? 13'b0000001111111 : node840;
										assign node840 = (inp[1]) ? node842 : 13'b0000011111111;
											assign node842 = (inp[0]) ? 13'b0000000111111 : 13'b0000011111111;
									assign node846 = (inp[0]) ? 13'b0000000011111 : 13'b0000001111111;
							assign node849 = (inp[2]) ? node867 : node850;
								assign node850 = (inp[0]) ? node864 : node851;
									assign node851 = (inp[12]) ? node857 : node852;
										assign node852 = (inp[1]) ? node854 : 13'b0001111111111;
											assign node854 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
										assign node857 = (inp[1]) ? 13'b0000001111111 : node858;
											assign node858 = (inp[8]) ? node860 : 13'b0000001111111;
												assign node860 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node864 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node867 = (inp[10]) ? node873 : node868;
									assign node868 = (inp[0]) ? node870 : 13'b0000000111111;
										assign node870 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node873 = (inp[9]) ? 13'b0000000000111 : 13'b0000000111111;
						assign node876 = (inp[2]) ? node912 : node877;
							assign node877 = (inp[1]) ? node893 : node878;
								assign node878 = (inp[3]) ? node886 : node879;
									assign node879 = (inp[12]) ? node881 : 13'b0000011111111;
										assign node881 = (inp[8]) ? 13'b0000001111111 : node882;
											assign node882 = (inp[9]) ? 13'b0000001111111 : 13'b0000111111111;
									assign node886 = (inp[0]) ? 13'b0000000111111 : node887;
										assign node887 = (inp[8]) ? node889 : 13'b0000011111111;
											assign node889 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node893 = (inp[8]) ? node901 : node894;
									assign node894 = (inp[0]) ? node896 : 13'b0000001111111;
										assign node896 = (inp[12]) ? 13'b0000000111111 : node897;
											assign node897 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node901 = (inp[0]) ? node909 : node902;
										assign node902 = (inp[9]) ? 13'b0000000111111 : node903;
											assign node903 = (inp[12]) ? node905 : 13'b0000000111111;
												assign node905 = (inp[3]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node909 = (inp[9]) ? 13'b0000000000111 : 13'b0000000111111;
							assign node912 = (inp[0]) ? node922 : node913;
								assign node913 = (inp[8]) ? node919 : node914;
									assign node914 = (inp[9]) ? node916 : 13'b0000001111111;
										assign node916 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node919 = (inp[10]) ? 13'b0000000111111 : 13'b0000000011111;
								assign node922 = (inp[10]) ? node930 : node923;
									assign node923 = (inp[1]) ? 13'b0000000011111 : node924;
										assign node924 = (inp[12]) ? node926 : 13'b0000000111111;
											assign node926 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node930 = (inp[9]) ? 13'b0000000001111 : node931;
										assign node931 = (inp[8]) ? node933 : 13'b0000000011111;
											assign node933 = (inp[3]) ? 13'b0000000001111 : node934;
												assign node934 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
				assign node939 = (inp[12]) ? node1021 : node940;
					assign node940 = (inp[0]) ? node982 : node941;
						assign node941 = (inp[1]) ? node961 : node942;
							assign node942 = (inp[2]) ? node954 : node943;
								assign node943 = (inp[10]) ? node949 : node944;
									assign node944 = (inp[3]) ? node946 : 13'b0000111111111;
										assign node946 = (inp[11]) ? 13'b0000111111111 : 13'b0001111111111;
									assign node949 = (inp[3]) ? node951 : 13'b0000111111111;
										assign node951 = (inp[6]) ? 13'b0000011111111 : 13'b0000001111111;
								assign node954 = (inp[3]) ? node958 : node955;
									assign node955 = (inp[8]) ? 13'b0000000111111 : 13'b0000011111111;
									assign node958 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
							assign node961 = (inp[3]) ? node971 : node962;
								assign node962 = (inp[9]) ? node966 : node963;
									assign node963 = (inp[11]) ? 13'b0000111111111 : 13'b0000011111111;
									assign node966 = (inp[10]) ? node968 : 13'b0000001111111;
										assign node968 = (inp[6]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node971 = (inp[6]) ? node973 : 13'b0000001111111;
									assign node973 = (inp[11]) ? node975 : 13'b0000000111111;
										assign node975 = (inp[2]) ? node977 : 13'b0000000001111;
											assign node977 = (inp[8]) ? 13'b0000000011111 : node978;
												assign node978 = (inp[10]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node982 = (inp[10]) ? node1000 : node983;
							assign node983 = (inp[8]) ? node997 : node984;
								assign node984 = (inp[1]) ? node992 : node985;
									assign node985 = (inp[6]) ? 13'b0000001111111 : node986;
										assign node986 = (inp[3]) ? node988 : 13'b0000011111111;
											assign node988 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node992 = (inp[6]) ? node994 : 13'b0000001111111;
										assign node994 = (inp[3]) ? 13'b0000000011111 : 13'b0000001111111;
								assign node997 = (inp[9]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node1000 = (inp[3]) ? node1006 : node1001;
								assign node1001 = (inp[2]) ? 13'b0000000111111 : node1002;
									assign node1002 = (inp[11]) ? 13'b0000000111111 : 13'b0000011111111;
								assign node1006 = (inp[1]) ? node1010 : node1007;
									assign node1007 = (inp[2]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1010 = (inp[2]) ? 13'b0000000001111 : node1011;
										assign node1011 = (inp[8]) ? node1013 : 13'b0000000011111;
											assign node1013 = (inp[11]) ? node1017 : node1014;
												assign node1014 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
												assign node1017 = (inp[6]) ? 13'b0000000000111 : 13'b0000000001111;
					assign node1021 = (inp[2]) ? node1065 : node1022;
						assign node1022 = (inp[8]) ? node1040 : node1023;
							assign node1023 = (inp[1]) ? node1029 : node1024;
								assign node1024 = (inp[9]) ? 13'b0000001111111 : node1025;
									assign node1025 = (inp[0]) ? 13'b0000011111111 : 13'b0000001111111;
								assign node1029 = (inp[11]) ? node1035 : node1030;
									assign node1030 = (inp[6]) ? node1032 : 13'b0000001111111;
										assign node1032 = (inp[10]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1035 = (inp[6]) ? 13'b0000000111111 : node1036;
										assign node1036 = (inp[9]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1040 = (inp[10]) ? node1052 : node1041;
								assign node1041 = (inp[1]) ? node1047 : node1042;
									assign node1042 = (inp[6]) ? 13'b0000000111111 : node1043;
										assign node1043 = (inp[0]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1047 = (inp[3]) ? node1049 : 13'b0000000011111;
										assign node1049 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1052 = (inp[11]) ? node1060 : node1053;
									assign node1053 = (inp[0]) ? node1055 : 13'b0000000111111;
										assign node1055 = (inp[6]) ? node1057 : 13'b0000000011111;
											assign node1057 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1060 = (inp[0]) ? node1062 : 13'b0000000001111;
										assign node1062 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node1065 = (inp[1]) ? node1069 : node1066;
							assign node1066 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1069 = (inp[11]) ? node1083 : node1070;
								assign node1070 = (inp[8]) ? node1078 : node1071;
									assign node1071 = (inp[6]) ? 13'b0000000011111 : node1072;
										assign node1072 = (inp[10]) ? node1074 : 13'b0000000011111;
											assign node1074 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1078 = (inp[6]) ? 13'b0000000001111 : node1079;
										assign node1079 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1083 = (inp[9]) ? 13'b0000000000011 : node1084;
									assign node1084 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
			assign node1088 = (inp[2]) ? node1266 : node1089;
				assign node1089 = (inp[9]) ? node1183 : node1090;
					assign node1090 = (inp[6]) ? node1138 : node1091;
						assign node1091 = (inp[3]) ? node1117 : node1092;
							assign node1092 = (inp[5]) ? node1108 : node1093;
								assign node1093 = (inp[11]) ? node1103 : node1094;
									assign node1094 = (inp[10]) ? node1096 : 13'b0000111111111;
										assign node1096 = (inp[8]) ? 13'b0000011111111 : node1097;
											assign node1097 = (inp[0]) ? node1099 : 13'b0000111111111;
												assign node1099 = (inp[12]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1103 = (inp[8]) ? 13'b0000001111111 : node1104;
										assign node1104 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
								assign node1108 = (inp[12]) ? node1114 : node1109;
									assign node1109 = (inp[1]) ? node1111 : 13'b0000111111111;
										assign node1111 = (inp[11]) ? 13'b0000001111111 : 13'b0000011111111;
									assign node1114 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
							assign node1117 = (inp[10]) ? node1133 : node1118;
								assign node1118 = (inp[8]) ? node1126 : node1119;
									assign node1119 = (inp[0]) ? 13'b0000001111111 : node1120;
										assign node1120 = (inp[12]) ? 13'b0000011111111 : node1121;
											assign node1121 = (inp[1]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1126 = (inp[0]) ? 13'b0000000111111 : node1127;
										assign node1127 = (inp[11]) ? 13'b0000000111111 : node1128;
											assign node1128 = (inp[5]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1133 = (inp[12]) ? 13'b0000000111111 : node1134;
									assign node1134 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
						assign node1138 = (inp[10]) ? node1160 : node1139;
							assign node1139 = (inp[11]) ? node1145 : node1140;
								assign node1140 = (inp[3]) ? node1142 : 13'b0000111111111;
									assign node1142 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1145 = (inp[3]) ? node1153 : node1146;
									assign node1146 = (inp[1]) ? node1148 : 13'b0000001111111;
										assign node1148 = (inp[8]) ? 13'b0000000111111 : node1149;
											assign node1149 = (inp[0]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1153 = (inp[12]) ? node1155 : 13'b0000000111111;
										assign node1155 = (inp[5]) ? node1157 : 13'b0000000011111;
											assign node1157 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node1160 = (inp[8]) ? node1172 : node1161;
								assign node1161 = (inp[5]) ? 13'b0000000011111 : node1162;
									assign node1162 = (inp[1]) ? node1166 : node1163;
										assign node1163 = (inp[11]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1166 = (inp[11]) ? node1168 : 13'b0000000111111;
											assign node1168 = (inp[12]) ? 13'b0000000011111 : 13'b0000000111111;
								assign node1172 = (inp[5]) ? 13'b0000000001111 : node1173;
									assign node1173 = (inp[12]) ? node1177 : node1174;
										assign node1174 = (inp[1]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1177 = (inp[1]) ? 13'b0000000011111 : node1178;
											assign node1178 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
					assign node1183 = (inp[3]) ? node1221 : node1184;
						assign node1184 = (inp[8]) ? node1202 : node1185;
							assign node1185 = (inp[5]) ? node1199 : node1186;
								assign node1186 = (inp[6]) ? node1192 : node1187;
									assign node1187 = (inp[0]) ? 13'b0000001111111 : node1188;
										assign node1188 = (inp[10]) ? 13'b0000011111111 : 13'b0000111111111;
									assign node1192 = (inp[11]) ? 13'b0000000111111 : node1193;
										assign node1193 = (inp[10]) ? node1195 : 13'b0000001111111;
											assign node1195 = (inp[1]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1199 = (inp[6]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1202 = (inp[1]) ? node1210 : node1203;
								assign node1203 = (inp[11]) ? node1205 : 13'b0000001111111;
									assign node1205 = (inp[0]) ? 13'b0000000111111 : node1206;
										assign node1206 = (inp[12]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1210 = (inp[5]) ? node1216 : node1211;
									assign node1211 = (inp[0]) ? 13'b0000000011111 : node1212;
										assign node1212 = (inp[11]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1216 = (inp[6]) ? node1218 : 13'b0000000011111;
										assign node1218 = (inp[12]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node1221 = (inp[1]) ? node1243 : node1222;
							assign node1222 = (inp[10]) ? node1236 : node1223;
								assign node1223 = (inp[0]) ? node1227 : node1224;
									assign node1224 = (inp[8]) ? 13'b0000001111111 : 13'b0000000111111;
									assign node1227 = (inp[12]) ? node1229 : 13'b0000000111111;
										assign node1229 = (inp[6]) ? node1233 : node1230;
											assign node1230 = (inp[8]) ? 13'b0000000011111 : 13'b0000000111111;
											assign node1233 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1236 = (inp[6]) ? node1238 : 13'b0000000011111;
									assign node1238 = (inp[12]) ? 13'b0000000000111 : node1239;
										assign node1239 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
							assign node1243 = (inp[0]) ? node1247 : node1244;
								assign node1244 = (inp[8]) ? 13'b0000000001111 : 13'b0000000011111;
								assign node1247 = (inp[5]) ? node1255 : node1248;
									assign node1248 = (inp[8]) ? node1250 : 13'b0000000111111;
										assign node1250 = (inp[11]) ? node1252 : 13'b0000000001111;
											assign node1252 = (inp[10]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1255 = (inp[6]) ? node1259 : node1256;
										assign node1256 = (inp[11]) ? 13'b0000000001111 : 13'b0000000011111;
										assign node1259 = (inp[8]) ? 13'b0000000000111 : node1260;
											assign node1260 = (inp[10]) ? node1262 : 13'b0000000001111;
												assign node1262 = (inp[11]) ? 13'b0000000000111 : 13'b0000000001111;
				assign node1266 = (inp[12]) ? node1356 : node1267;
					assign node1267 = (inp[11]) ? node1313 : node1268;
						assign node1268 = (inp[3]) ? node1296 : node1269;
							assign node1269 = (inp[5]) ? node1283 : node1270;
								assign node1270 = (inp[0]) ? node1276 : node1271;
									assign node1271 = (inp[8]) ? 13'b0000001111111 : node1272;
										assign node1272 = (inp[1]) ? 13'b0000111111111 : 13'b0000011111111;
									assign node1276 = (inp[10]) ? 13'b0000000111111 : node1277;
										assign node1277 = (inp[1]) ? 13'b0000001111111 : node1278;
											assign node1278 = (inp[8]) ? 13'b0000001111111 : 13'b0000011111111;
								assign node1283 = (inp[10]) ? node1291 : node1284;
									assign node1284 = (inp[0]) ? node1286 : 13'b0000001111111;
										assign node1286 = (inp[9]) ? 13'b0000000111111 : node1287;
											assign node1287 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
									assign node1291 = (inp[8]) ? node1293 : 13'b0000000111111;
										assign node1293 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
							assign node1296 = (inp[0]) ? 13'b0000000001111 : node1297;
								assign node1297 = (inp[8]) ? node1305 : node1298;
									assign node1298 = (inp[9]) ? node1302 : node1299;
										assign node1299 = (inp[1]) ? 13'b0000011111111 : 13'b0000001111111;
										assign node1302 = (inp[5]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1305 = (inp[1]) ? node1307 : 13'b0000000111111;
										assign node1307 = (inp[9]) ? node1309 : 13'b0000000011111;
											assign node1309 = (inp[6]) ? 13'b0000000001111 : 13'b0000000011111;
						assign node1313 = (inp[1]) ? node1339 : node1314;
							assign node1314 = (inp[10]) ? node1320 : node1315;
								assign node1315 = (inp[9]) ? node1317 : 13'b0000000111111;
									assign node1317 = (inp[6]) ? 13'b0000000011111 : 13'b0000001111111;
								assign node1320 = (inp[3]) ? node1332 : node1321;
									assign node1321 = (inp[6]) ? node1329 : node1322;
										assign node1322 = (inp[5]) ? node1326 : node1323;
											assign node1323 = (inp[9]) ? 13'b0000000111111 : 13'b0000011111111;
											assign node1326 = (inp[0]) ? 13'b0000000011111 : 13'b0000000111111;
										assign node1329 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1332 = (inp[6]) ? node1336 : node1333;
										assign node1333 = (inp[5]) ? 13'b0000000011111 : 13'b0000000001111;
										assign node1336 = (inp[9]) ? 13'b0000000000011 : 13'b0000000001111;
							assign node1339 = (inp[6]) ? node1341 : 13'b0000000011111;
								assign node1341 = (inp[9]) ? node1351 : node1342;
									assign node1342 = (inp[3]) ? 13'b0000000001111 : node1343;
										assign node1343 = (inp[8]) ? 13'b0000000001111 : node1344;
											assign node1344 = (inp[10]) ? node1346 : 13'b0000000011111;
												assign node1346 = (inp[0]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1351 = (inp[5]) ? 13'b0000000000111 : node1352;
										assign node1352 = (inp[3]) ? 13'b0000000001111 : 13'b0000000011111;
					assign node1356 = (inp[10]) ? node1400 : node1357;
						assign node1357 = (inp[0]) ? node1377 : node1358;
							assign node1358 = (inp[9]) ? node1364 : node1359;
								assign node1359 = (inp[5]) ? 13'b0000000111111 : node1360;
									assign node1360 = (inp[3]) ? 13'b0000000111111 : 13'b0000001111111;
								assign node1364 = (inp[3]) ? node1372 : node1365;
									assign node1365 = (inp[5]) ? node1369 : node1366;
										assign node1366 = (inp[8]) ? 13'b0000000111111 : 13'b0000001111111;
										assign node1369 = (inp[1]) ? 13'b0000000011111 : 13'b0000000111111;
									assign node1372 = (inp[8]) ? 13'b0000000001111 : node1373;
										assign node1373 = (inp[6]) ? 13'b0000000000111 : 13'b0000000011111;
							assign node1377 = (inp[3]) ? node1389 : node1378;
								assign node1378 = (inp[11]) ? node1382 : node1379;
									assign node1379 = (inp[1]) ? 13'b0000000011111 : 13'b0000001111111;
									assign node1382 = (inp[1]) ? node1384 : 13'b0000000011111;
										assign node1384 = (inp[8]) ? node1386 : 13'b0000000001111;
											assign node1386 = (inp[6]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node1389 = (inp[5]) ? node1397 : node1390;
									assign node1390 = (inp[11]) ? node1392 : 13'b0000000011111;
										assign node1392 = (inp[8]) ? node1394 : 13'b0000000001111;
											assign node1394 = (inp[9]) ? 13'b0000000000111 : 13'b0000000001111;
									assign node1397 = (inp[1]) ? 13'b0000000000111 : 13'b0000000001111;
						assign node1400 = (inp[9]) ? node1424 : node1401;
							assign node1401 = (inp[0]) ? node1415 : node1402;
								assign node1402 = (inp[1]) ? node1408 : node1403;
									assign node1403 = (inp[6]) ? 13'b0000000011111 : node1404;
										assign node1404 = (inp[5]) ? 13'b0000000001111 : 13'b0000000011111;
									assign node1408 = (inp[5]) ? 13'b0000000001111 : node1409;
										assign node1409 = (inp[11]) ? node1411 : 13'b0000000001111;
											assign node1411 = (inp[8]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node1415 = (inp[8]) ? node1421 : node1416;
									assign node1416 = (inp[11]) ? 13'b0000000000111 : node1417;
										assign node1417 = (inp[5]) ? 13'b0000000001111 : 13'b0000000111111;
									assign node1421 = (inp[1]) ? 13'b0000000000011 : 13'b0000000000111;
							assign node1424 = (inp[6]) ? node1428 : node1425;
								assign node1425 = (inp[3]) ? 13'b0000000000111 : 13'b0000000001111;
								assign node1428 = (inp[0]) ? node1434 : node1429;
									assign node1429 = (inp[11]) ? 13'b0000000000111 : node1430;
										assign node1430 = (inp[3]) ? 13'b0000000001111 : 13'b0000000000111;
									assign node1434 = (inp[1]) ? 13'b0000000000111 : node1435;
										assign node1435 = (inp[5]) ? 13'b0000000000011 : 13'b0000000000111;

endmodule