module dtc_split5_bm56 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node40;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node51;
	wire [3-1:0] node52;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node114;
	wire [3-1:0] node118;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node127;
	wire [3-1:0] node130;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node145;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node153;
	wire [3-1:0] node156;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node160;
	wire [3-1:0] node163;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node172;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node177;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node182;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node212;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node218;
	wire [3-1:0] node221;
	wire [3-1:0] node224;
	wire [3-1:0] node225;
	wire [3-1:0] node226;
	wire [3-1:0] node228;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node242;
	wire [3-1:0] node243;
	wire [3-1:0] node247;
	wire [3-1:0] node248;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node253;
	wire [3-1:0] node257;
	wire [3-1:0] node259;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node264;
	wire [3-1:0] node266;
	wire [3-1:0] node269;
	wire [3-1:0] node270;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node277;
	wire [3-1:0] node280;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node286;
	wire [3-1:0] node287;
	wire [3-1:0] node290;
	wire [3-1:0] node293;
	wire [3-1:0] node295;
	wire [3-1:0] node298;
	wire [3-1:0] node299;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node305;
	wire [3-1:0] node308;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node313;
	wire [3-1:0] node314;
	wire [3-1:0] node317;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node324;
	wire [3-1:0] node325;
	wire [3-1:0] node328;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node338;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node341;
	wire [3-1:0] node342;
	wire [3-1:0] node343;
	wire [3-1:0] node347;
	wire [3-1:0] node349;
	wire [3-1:0] node352;
	wire [3-1:0] node353;
	wire [3-1:0] node356;
	wire [3-1:0] node359;
	wire [3-1:0] node360;
	wire [3-1:0] node361;
	wire [3-1:0] node362;
	wire [3-1:0] node365;
	wire [3-1:0] node368;
	wire [3-1:0] node369;
	wire [3-1:0] node373;
	wire [3-1:0] node375;
	wire [3-1:0] node376;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node382;
	wire [3-1:0] node385;
	wire [3-1:0] node386;
	wire [3-1:0] node387;
	wire [3-1:0] node390;
	wire [3-1:0] node393;
	wire [3-1:0] node395;
	wire [3-1:0] node398;
	wire [3-1:0] node399;
	wire [3-1:0] node400;
	wire [3-1:0] node402;
	wire [3-1:0] node406;
	wire [3-1:0] node407;
	wire [3-1:0] node408;
	wire [3-1:0] node411;
	wire [3-1:0] node414;
	wire [3-1:0] node415;
	wire [3-1:0] node418;
	wire [3-1:0] node421;
	wire [3-1:0] node422;
	wire [3-1:0] node423;
	wire [3-1:0] node424;
	wire [3-1:0] node425;
	wire [3-1:0] node427;
	wire [3-1:0] node430;
	wire [3-1:0] node433;
	wire [3-1:0] node434;
	wire [3-1:0] node437;
	wire [3-1:0] node440;
	wire [3-1:0] node441;
	wire [3-1:0] node442;
	wire [3-1:0] node443;
	wire [3-1:0] node447;
	wire [3-1:0] node450;
	wire [3-1:0] node451;
	wire [3-1:0] node453;
	wire [3-1:0] node457;
	wire [3-1:0] node458;
	wire [3-1:0] node459;
	wire [3-1:0] node460;
	wire [3-1:0] node462;
	wire [3-1:0] node465;
	wire [3-1:0] node466;
	wire [3-1:0] node470;
	wire [3-1:0] node472;
	wire [3-1:0] node475;
	wire [3-1:0] node476;
	wire [3-1:0] node477;
	wire [3-1:0] node481;
	wire [3-1:0] node482;
	wire [3-1:0] node484;
	wire [3-1:0] node487;
	wire [3-1:0] node489;
	wire [3-1:0] node492;
	wire [3-1:0] node493;
	wire [3-1:0] node494;
	wire [3-1:0] node495;
	wire [3-1:0] node496;
	wire [3-1:0] node497;
	wire [3-1:0] node500;
	wire [3-1:0] node501;
	wire [3-1:0] node505;
	wire [3-1:0] node506;
	wire [3-1:0] node507;
	wire [3-1:0] node511;
	wire [3-1:0] node512;
	wire [3-1:0] node516;
	wire [3-1:0] node517;
	wire [3-1:0] node518;
	wire [3-1:0] node520;
	wire [3-1:0] node523;
	wire [3-1:0] node524;
	wire [3-1:0] node527;
	wire [3-1:0] node530;
	wire [3-1:0] node531;
	wire [3-1:0] node532;
	wire [3-1:0] node536;
	wire [3-1:0] node538;
	wire [3-1:0] node541;
	wire [3-1:0] node542;
	wire [3-1:0] node543;
	wire [3-1:0] node544;
	wire [3-1:0] node545;
	wire [3-1:0] node549;
	wire [3-1:0] node551;
	wire [3-1:0] node554;
	wire [3-1:0] node555;
	wire [3-1:0] node556;
	wire [3-1:0] node560;
	wire [3-1:0] node563;
	wire [3-1:0] node564;
	wire [3-1:0] node565;
	wire [3-1:0] node566;
	wire [3-1:0] node570;
	wire [3-1:0] node571;
	wire [3-1:0] node574;
	wire [3-1:0] node577;
	wire [3-1:0] node578;
	wire [3-1:0] node579;
	wire [3-1:0] node583;
	wire [3-1:0] node586;
	wire [3-1:0] node587;
	wire [3-1:0] node588;
	wire [3-1:0] node589;
	wire [3-1:0] node590;
	wire [3-1:0] node592;
	wire [3-1:0] node596;
	wire [3-1:0] node597;
	wire [3-1:0] node599;
	wire [3-1:0] node602;
	wire [3-1:0] node604;
	wire [3-1:0] node607;
	wire [3-1:0] node608;
	wire [3-1:0] node609;
	wire [3-1:0] node611;
	wire [3-1:0] node614;
	wire [3-1:0] node617;
	wire [3-1:0] node619;
	wire [3-1:0] node620;
	wire [3-1:0] node623;
	wire [3-1:0] node626;
	wire [3-1:0] node627;
	wire [3-1:0] node628;
	wire [3-1:0] node629;
	wire [3-1:0] node630;
	wire [3-1:0] node633;
	wire [3-1:0] node636;
	wire [3-1:0] node638;
	wire [3-1:0] node641;
	wire [3-1:0] node642;
	wire [3-1:0] node645;
	wire [3-1:0] node646;
	wire [3-1:0] node650;
	wire [3-1:0] node651;
	wire [3-1:0] node654;
	wire [3-1:0] node655;
	wire [3-1:0] node656;
	wire [3-1:0] node659;
	wire [3-1:0] node662;
	wire [3-1:0] node665;
	wire [3-1:0] node666;
	wire [3-1:0] node667;
	wire [3-1:0] node668;
	wire [3-1:0] node669;
	wire [3-1:0] node670;
	wire [3-1:0] node671;
	wire [3-1:0] node672;
	wire [3-1:0] node673;
	wire [3-1:0] node677;
	wire [3-1:0] node679;
	wire [3-1:0] node682;
	wire [3-1:0] node683;
	wire [3-1:0] node684;
	wire [3-1:0] node687;
	wire [3-1:0] node690;
	wire [3-1:0] node691;
	wire [3-1:0] node694;
	wire [3-1:0] node697;
	wire [3-1:0] node698;
	wire [3-1:0] node699;
	wire [3-1:0] node702;
	wire [3-1:0] node705;
	wire [3-1:0] node707;
	wire [3-1:0] node709;
	wire [3-1:0] node712;
	wire [3-1:0] node713;
	wire [3-1:0] node714;
	wire [3-1:0] node715;
	wire [3-1:0] node717;
	wire [3-1:0] node720;
	wire [3-1:0] node722;
	wire [3-1:0] node725;
	wire [3-1:0] node726;
	wire [3-1:0] node727;
	wire [3-1:0] node730;
	wire [3-1:0] node733;
	wire [3-1:0] node734;
	wire [3-1:0] node738;
	wire [3-1:0] node739;
	wire [3-1:0] node740;
	wire [3-1:0] node743;
	wire [3-1:0] node746;
	wire [3-1:0] node747;
	wire [3-1:0] node748;
	wire [3-1:0] node752;
	wire [3-1:0] node754;
	wire [3-1:0] node757;
	wire [3-1:0] node758;
	wire [3-1:0] node759;
	wire [3-1:0] node760;
	wire [3-1:0] node761;
	wire [3-1:0] node762;
	wire [3-1:0] node765;
	wire [3-1:0] node768;
	wire [3-1:0] node770;
	wire [3-1:0] node773;
	wire [3-1:0] node774;
	wire [3-1:0] node776;
	wire [3-1:0] node779;
	wire [3-1:0] node781;
	wire [3-1:0] node784;
	wire [3-1:0] node785;
	wire [3-1:0] node786;
	wire [3-1:0] node787;
	wire [3-1:0] node790;
	wire [3-1:0] node793;
	wire [3-1:0] node795;
	wire [3-1:0] node798;
	wire [3-1:0] node799;
	wire [3-1:0] node801;
	wire [3-1:0] node804;
	wire [3-1:0] node805;
	wire [3-1:0] node809;
	wire [3-1:0] node810;
	wire [3-1:0] node811;
	wire [3-1:0] node812;
	wire [3-1:0] node813;
	wire [3-1:0] node817;
	wire [3-1:0] node818;
	wire [3-1:0] node822;
	wire [3-1:0] node823;
	wire [3-1:0] node825;
	wire [3-1:0] node828;
	wire [3-1:0] node829;
	wire [3-1:0] node832;
	wire [3-1:0] node835;
	wire [3-1:0] node836;
	wire [3-1:0] node837;
	wire [3-1:0] node838;
	wire [3-1:0] node842;
	wire [3-1:0] node844;
	wire [3-1:0] node847;
	wire [3-1:0] node848;
	wire [3-1:0] node849;
	wire [3-1:0] node852;
	wire [3-1:0] node855;
	wire [3-1:0] node856;
	wire [3-1:0] node859;
	wire [3-1:0] node862;
	wire [3-1:0] node863;
	wire [3-1:0] node864;
	wire [3-1:0] node865;
	wire [3-1:0] node866;
	wire [3-1:0] node867;
	wire [3-1:0] node869;
	wire [3-1:0] node872;
	wire [3-1:0] node875;
	wire [3-1:0] node876;
	wire [3-1:0] node879;
	wire [3-1:0] node882;
	wire [3-1:0] node883;
	wire [3-1:0] node884;
	wire [3-1:0] node885;
	wire [3-1:0] node889;
	wire [3-1:0] node892;
	wire [3-1:0] node893;
	wire [3-1:0] node894;
	wire [3-1:0] node899;
	wire [3-1:0] node900;
	wire [3-1:0] node901;
	wire [3-1:0] node903;
	wire [3-1:0] node905;
	wire [3-1:0] node908;
	wire [3-1:0] node909;
	wire [3-1:0] node911;
	wire [3-1:0] node914;
	wire [3-1:0] node916;
	wire [3-1:0] node919;
	wire [3-1:0] node920;
	wire [3-1:0] node921;
	wire [3-1:0] node922;
	wire [3-1:0] node925;
	wire [3-1:0] node929;
	wire [3-1:0] node931;
	wire [3-1:0] node932;
	wire [3-1:0] node936;
	wire [3-1:0] node937;
	wire [3-1:0] node938;
	wire [3-1:0] node939;
	wire [3-1:0] node940;
	wire [3-1:0] node943;
	wire [3-1:0] node945;
	wire [3-1:0] node948;
	wire [3-1:0] node949;
	wire [3-1:0] node950;
	wire [3-1:0] node954;
	wire [3-1:0] node955;
	wire [3-1:0] node958;
	wire [3-1:0] node961;
	wire [3-1:0] node962;
	wire [3-1:0] node963;
	wire [3-1:0] node967;
	wire [3-1:0] node968;
	wire [3-1:0] node969;
	wire [3-1:0] node973;
	wire [3-1:0] node974;
	wire [3-1:0] node978;
	wire [3-1:0] node979;
	wire [3-1:0] node980;
	wire [3-1:0] node981;
	wire [3-1:0] node985;
	wire [3-1:0] node986;
	wire [3-1:0] node987;
	wire [3-1:0] node990;
	wire [3-1:0] node994;
	wire [3-1:0] node995;
	wire [3-1:0] node996;
	wire [3-1:0] node997;
	wire [3-1:0] node1000;
	wire [3-1:0] node1003;
	wire [3-1:0] node1004;
	wire [3-1:0] node1008;
	wire [3-1:0] node1009;
	wire [3-1:0] node1011;
	wire [3-1:0] node1014;
	wire [3-1:0] node1016;
	wire [3-1:0] node1019;
	wire [3-1:0] node1020;
	wire [3-1:0] node1021;
	wire [3-1:0] node1022;
	wire [3-1:0] node1023;
	wire [3-1:0] node1024;
	wire [3-1:0] node1025;
	wire [3-1:0] node1028;
	wire [3-1:0] node1029;
	wire [3-1:0] node1032;
	wire [3-1:0] node1035;
	wire [3-1:0] node1036;
	wire [3-1:0] node1037;
	wire [3-1:0] node1041;
	wire [3-1:0] node1042;
	wire [3-1:0] node1046;
	wire [3-1:0] node1047;
	wire [3-1:0] node1049;
	wire [3-1:0] node1051;
	wire [3-1:0] node1054;
	wire [3-1:0] node1056;
	wire [3-1:0] node1057;
	wire [3-1:0] node1061;
	wire [3-1:0] node1062;
	wire [3-1:0] node1063;
	wire [3-1:0] node1064;
	wire [3-1:0] node1065;
	wire [3-1:0] node1069;
	wire [3-1:0] node1070;
	wire [3-1:0] node1073;
	wire [3-1:0] node1076;
	wire [3-1:0] node1077;
	wire [3-1:0] node1080;
	wire [3-1:0] node1081;
	wire [3-1:0] node1084;
	wire [3-1:0] node1087;
	wire [3-1:0] node1088;
	wire [3-1:0] node1089;
	wire [3-1:0] node1092;
	wire [3-1:0] node1095;
	wire [3-1:0] node1096;
	wire [3-1:0] node1099;
	wire [3-1:0] node1102;
	wire [3-1:0] node1103;
	wire [3-1:0] node1104;
	wire [3-1:0] node1105;
	wire [3-1:0] node1106;
	wire [3-1:0] node1107;
	wire [3-1:0] node1110;
	wire [3-1:0] node1113;
	wire [3-1:0] node1114;
	wire [3-1:0] node1118;
	wire [3-1:0] node1119;
	wire [3-1:0] node1121;
	wire [3-1:0] node1124;
	wire [3-1:0] node1126;
	wire [3-1:0] node1129;
	wire [3-1:0] node1130;
	wire [3-1:0] node1131;
	wire [3-1:0] node1132;
	wire [3-1:0] node1136;
	wire [3-1:0] node1139;
	wire [3-1:0] node1140;
	wire [3-1:0] node1141;
	wire [3-1:0] node1145;
	wire [3-1:0] node1147;
	wire [3-1:0] node1150;
	wire [3-1:0] node1151;
	wire [3-1:0] node1152;
	wire [3-1:0] node1153;
	wire [3-1:0] node1154;
	wire [3-1:0] node1159;
	wire [3-1:0] node1160;
	wire [3-1:0] node1162;
	wire [3-1:0] node1165;
	wire [3-1:0] node1166;
	wire [3-1:0] node1169;
	wire [3-1:0] node1172;
	wire [3-1:0] node1173;
	wire [3-1:0] node1174;
	wire [3-1:0] node1177;
	wire [3-1:0] node1180;
	wire [3-1:0] node1181;
	wire [3-1:0] node1182;
	wire [3-1:0] node1187;
	wire [3-1:0] node1188;
	wire [3-1:0] node1189;
	wire [3-1:0] node1190;
	wire [3-1:0] node1191;
	wire [3-1:0] node1192;
	wire [3-1:0] node1193;
	wire [3-1:0] node1197;
	wire [3-1:0] node1200;
	wire [3-1:0] node1201;
	wire [3-1:0] node1202;
	wire [3-1:0] node1205;
	wire [3-1:0] node1209;
	wire [3-1:0] node1210;
	wire [3-1:0] node1211;
	wire [3-1:0] node1212;
	wire [3-1:0] node1216;
	wire [3-1:0] node1218;
	wire [3-1:0] node1221;
	wire [3-1:0] node1222;
	wire [3-1:0] node1223;
	wire [3-1:0] node1227;
	wire [3-1:0] node1228;
	wire [3-1:0] node1232;
	wire [3-1:0] node1233;
	wire [3-1:0] node1234;
	wire [3-1:0] node1235;
	wire [3-1:0] node1237;
	wire [3-1:0] node1240;
	wire [3-1:0] node1241;
	wire [3-1:0] node1245;
	wire [3-1:0] node1246;
	wire [3-1:0] node1247;
	wire [3-1:0] node1250;
	wire [3-1:0] node1253;
	wire [3-1:0] node1254;
	wire [3-1:0] node1257;
	wire [3-1:0] node1260;
	wire [3-1:0] node1261;
	wire [3-1:0] node1262;
	wire [3-1:0] node1264;
	wire [3-1:0] node1267;
	wire [3-1:0] node1269;
	wire [3-1:0] node1272;
	wire [3-1:0] node1273;
	wire [3-1:0] node1274;
	wire [3-1:0] node1277;
	wire [3-1:0] node1280;
	wire [3-1:0] node1281;
	wire [3-1:0] node1284;
	wire [3-1:0] node1287;
	wire [3-1:0] node1288;
	wire [3-1:0] node1289;
	wire [3-1:0] node1290;
	wire [3-1:0] node1291;
	wire [3-1:0] node1293;
	wire [3-1:0] node1297;
	wire [3-1:0] node1298;
	wire [3-1:0] node1301;
	wire [3-1:0] node1303;
	wire [3-1:0] node1306;
	wire [3-1:0] node1307;
	wire [3-1:0] node1308;
	wire [3-1:0] node1309;
	wire [3-1:0] node1313;
	wire [3-1:0] node1316;
	wire [3-1:0] node1317;
	wire [3-1:0] node1318;
	wire [3-1:0] node1322;
	wire [3-1:0] node1323;
	wire [3-1:0] node1326;
	wire [3-1:0] node1329;
	wire [3-1:0] node1330;
	wire [3-1:0] node1331;
	wire [3-1:0] node1332;
	wire [3-1:0] node1333;
	wire [3-1:0] node1336;
	wire [3-1:0] node1339;
	wire [3-1:0] node1340;
	wire [3-1:0] node1344;
	wire [3-1:0] node1345;
	wire [3-1:0] node1348;
	wire [3-1:0] node1351;
	wire [3-1:0] node1352;
	wire [3-1:0] node1353;
	wire [3-1:0] node1355;
	wire [3-1:0] node1358;
	wire [3-1:0] node1361;
	wire [3-1:0] node1362;
	wire [3-1:0] node1363;
	wire [3-1:0] node1366;
	wire [3-1:0] node1369;
	wire [3-1:0] node1370;
	wire [3-1:0] node1374;
	wire [3-1:0] node1375;
	wire [3-1:0] node1376;
	wire [3-1:0] node1377;
	wire [3-1:0] node1378;
	wire [3-1:0] node1379;
	wire [3-1:0] node1380;
	wire [3-1:0] node1381;
	wire [3-1:0] node1382;
	wire [3-1:0] node1383;
	wire [3-1:0] node1386;
	wire [3-1:0] node1389;
	wire [3-1:0] node1390;
	wire [3-1:0] node1393;
	wire [3-1:0] node1396;
	wire [3-1:0] node1397;
	wire [3-1:0] node1398;
	wire [3-1:0] node1402;
	wire [3-1:0] node1403;
	wire [3-1:0] node1407;
	wire [3-1:0] node1408;
	wire [3-1:0] node1409;
	wire [3-1:0] node1410;
	wire [3-1:0] node1414;
	wire [3-1:0] node1415;
	wire [3-1:0] node1419;
	wire [3-1:0] node1420;
	wire [3-1:0] node1423;
	wire [3-1:0] node1425;
	wire [3-1:0] node1428;
	wire [3-1:0] node1429;
	wire [3-1:0] node1430;
	wire [3-1:0] node1432;
	wire [3-1:0] node1435;
	wire [3-1:0] node1436;
	wire [3-1:0] node1437;
	wire [3-1:0] node1441;
	wire [3-1:0] node1442;
	wire [3-1:0] node1445;
	wire [3-1:0] node1448;
	wire [3-1:0] node1449;
	wire [3-1:0] node1450;
	wire [3-1:0] node1453;
	wire [3-1:0] node1454;
	wire [3-1:0] node1458;
	wire [3-1:0] node1459;
	wire [3-1:0] node1460;
	wire [3-1:0] node1465;
	wire [3-1:0] node1466;
	wire [3-1:0] node1467;
	wire [3-1:0] node1468;
	wire [3-1:0] node1469;
	wire [3-1:0] node1470;
	wire [3-1:0] node1474;
	wire [3-1:0] node1476;
	wire [3-1:0] node1479;
	wire [3-1:0] node1480;
	wire [3-1:0] node1482;
	wire [3-1:0] node1486;
	wire [3-1:0] node1487;
	wire [3-1:0] node1488;
	wire [3-1:0] node1489;
	wire [3-1:0] node1493;
	wire [3-1:0] node1496;
	wire [3-1:0] node1497;
	wire [3-1:0] node1501;
	wire [3-1:0] node1502;
	wire [3-1:0] node1503;
	wire [3-1:0] node1504;
	wire [3-1:0] node1506;
	wire [3-1:0] node1509;
	wire [3-1:0] node1510;
	wire [3-1:0] node1514;
	wire [3-1:0] node1515;
	wire [3-1:0] node1516;
	wire [3-1:0] node1519;
	wire [3-1:0] node1522;
	wire [3-1:0] node1524;
	wire [3-1:0] node1527;
	wire [3-1:0] node1528;
	wire [3-1:0] node1529;
	wire [3-1:0] node1531;
	wire [3-1:0] node1534;
	wire [3-1:0] node1535;
	wire [3-1:0] node1539;
	wire [3-1:0] node1540;
	wire [3-1:0] node1542;
	wire [3-1:0] node1545;
	wire [3-1:0] node1546;
	wire [3-1:0] node1550;
	wire [3-1:0] node1551;
	wire [3-1:0] node1552;
	wire [3-1:0] node1553;
	wire [3-1:0] node1554;
	wire [3-1:0] node1555;
	wire [3-1:0] node1556;
	wire [3-1:0] node1559;
	wire [3-1:0] node1562;
	wire [3-1:0] node1565;
	wire [3-1:0] node1566;
	wire [3-1:0] node1568;
	wire [3-1:0] node1572;
	wire [3-1:0] node1573;
	wire [3-1:0] node1574;
	wire [3-1:0] node1576;
	wire [3-1:0] node1579;
	wire [3-1:0] node1581;
	wire [3-1:0] node1584;
	wire [3-1:0] node1585;
	wire [3-1:0] node1588;
	wire [3-1:0] node1590;
	wire [3-1:0] node1593;
	wire [3-1:0] node1594;
	wire [3-1:0] node1595;
	wire [3-1:0] node1596;
	wire [3-1:0] node1597;
	wire [3-1:0] node1601;
	wire [3-1:0] node1602;
	wire [3-1:0] node1606;
	wire [3-1:0] node1607;
	wire [3-1:0] node1608;
	wire [3-1:0] node1611;
	wire [3-1:0] node1615;
	wire [3-1:0] node1616;
	wire [3-1:0] node1617;
	wire [3-1:0] node1620;
	wire [3-1:0] node1622;
	wire [3-1:0] node1625;
	wire [3-1:0] node1626;
	wire [3-1:0] node1627;
	wire [3-1:0] node1631;
	wire [3-1:0] node1632;
	wire [3-1:0] node1635;
	wire [3-1:0] node1638;
	wire [3-1:0] node1639;
	wire [3-1:0] node1640;
	wire [3-1:0] node1641;
	wire [3-1:0] node1642;
	wire [3-1:0] node1645;
	wire [3-1:0] node1648;
	wire [3-1:0] node1649;
	wire [3-1:0] node1650;
	wire [3-1:0] node1653;
	wire [3-1:0] node1656;
	wire [3-1:0] node1658;
	wire [3-1:0] node1661;
	wire [3-1:0] node1662;
	wire [3-1:0] node1664;
	wire [3-1:0] node1665;
	wire [3-1:0] node1668;
	wire [3-1:0] node1671;
	wire [3-1:0] node1672;
	wire [3-1:0] node1674;
	wire [3-1:0] node1677;
	wire [3-1:0] node1678;
	wire [3-1:0] node1682;
	wire [3-1:0] node1683;
	wire [3-1:0] node1684;
	wire [3-1:0] node1685;
	wire [3-1:0] node1687;
	wire [3-1:0] node1690;
	wire [3-1:0] node1692;
	wire [3-1:0] node1695;
	wire [3-1:0] node1696;
	wire [3-1:0] node1697;
	wire [3-1:0] node1702;
	wire [3-1:0] node1703;
	wire [3-1:0] node1704;
	wire [3-1:0] node1705;
	wire [3-1:0] node1708;
	wire [3-1:0] node1711;
	wire [3-1:0] node1712;
	wire [3-1:0] node1715;
	wire [3-1:0] node1718;
	wire [3-1:0] node1719;
	wire [3-1:0] node1721;
	wire [3-1:0] node1724;
	wire [3-1:0] node1725;
	wire [3-1:0] node1729;
	wire [3-1:0] node1730;
	wire [3-1:0] node1731;
	wire [3-1:0] node1732;
	wire [3-1:0] node1733;
	wire [3-1:0] node1734;
	wire [3-1:0] node1735;
	wire [3-1:0] node1736;
	wire [3-1:0] node1740;
	wire [3-1:0] node1741;
	wire [3-1:0] node1744;
	wire [3-1:0] node1747;
	wire [3-1:0] node1748;
	wire [3-1:0] node1750;
	wire [3-1:0] node1753;
	wire [3-1:0] node1754;
	wire [3-1:0] node1758;
	wire [3-1:0] node1759;
	wire [3-1:0] node1761;
	wire [3-1:0] node1764;
	wire [3-1:0] node1765;
	wire [3-1:0] node1766;
	wire [3-1:0] node1769;
	wire [3-1:0] node1772;
	wire [3-1:0] node1773;
	wire [3-1:0] node1777;
	wire [3-1:0] node1778;
	wire [3-1:0] node1779;
	wire [3-1:0] node1781;
	wire [3-1:0] node1782;
	wire [3-1:0] node1785;
	wire [3-1:0] node1788;
	wire [3-1:0] node1789;
	wire [3-1:0] node1792;
	wire [3-1:0] node1795;
	wire [3-1:0] node1796;
	wire [3-1:0] node1797;
	wire [3-1:0] node1799;
	wire [3-1:0] node1802;
	wire [3-1:0] node1805;
	wire [3-1:0] node1806;
	wire [3-1:0] node1807;
	wire [3-1:0] node1811;
	wire [3-1:0] node1812;
	wire [3-1:0] node1816;
	wire [3-1:0] node1817;
	wire [3-1:0] node1818;
	wire [3-1:0] node1819;
	wire [3-1:0] node1820;
	wire [3-1:0] node1823;
	wire [3-1:0] node1824;
	wire [3-1:0] node1828;
	wire [3-1:0] node1829;
	wire [3-1:0] node1830;
	wire [3-1:0] node1834;
	wire [3-1:0] node1835;
	wire [3-1:0] node1839;
	wire [3-1:0] node1840;
	wire [3-1:0] node1841;
	wire [3-1:0] node1842;
	wire [3-1:0] node1845;
	wire [3-1:0] node1848;
	wire [3-1:0] node1849;
	wire [3-1:0] node1853;
	wire [3-1:0] node1854;
	wire [3-1:0] node1857;
	wire [3-1:0] node1860;
	wire [3-1:0] node1861;
	wire [3-1:0] node1862;
	wire [3-1:0] node1864;
	wire [3-1:0] node1865;
	wire [3-1:0] node1869;
	wire [3-1:0] node1872;
	wire [3-1:0] node1873;
	wire [3-1:0] node1874;
	wire [3-1:0] node1875;
	wire [3-1:0] node1880;
	wire [3-1:0] node1881;
	wire [3-1:0] node1884;
	wire [3-1:0] node1887;
	wire [3-1:0] node1888;
	wire [3-1:0] node1889;
	wire [3-1:0] node1890;
	wire [3-1:0] node1891;
	wire [3-1:0] node1892;
	wire [3-1:0] node1893;
	wire [3-1:0] node1897;
	wire [3-1:0] node1898;
	wire [3-1:0] node1902;
	wire [3-1:0] node1903;
	wire [3-1:0] node1905;
	wire [3-1:0] node1908;
	wire [3-1:0] node1910;
	wire [3-1:0] node1913;
	wire [3-1:0] node1914;
	wire [3-1:0] node1915;
	wire [3-1:0] node1917;
	wire [3-1:0] node1920;
	wire [3-1:0] node1921;
	wire [3-1:0] node1925;
	wire [3-1:0] node1926;
	wire [3-1:0] node1927;
	wire [3-1:0] node1931;
	wire [3-1:0] node1932;
	wire [3-1:0] node1936;
	wire [3-1:0] node1937;
	wire [3-1:0] node1938;
	wire [3-1:0] node1939;
	wire [3-1:0] node1942;
	wire [3-1:0] node1943;
	wire [3-1:0] node1947;
	wire [3-1:0] node1948;
	wire [3-1:0] node1951;
	wire [3-1:0] node1954;
	wire [3-1:0] node1955;
	wire [3-1:0] node1956;
	wire [3-1:0] node1958;
	wire [3-1:0] node1961;
	wire [3-1:0] node1962;
	wire [3-1:0] node1966;
	wire [3-1:0] node1967;
	wire [3-1:0] node1970;
	wire [3-1:0] node1973;
	wire [3-1:0] node1974;
	wire [3-1:0] node1975;
	wire [3-1:0] node1976;
	wire [3-1:0] node1977;
	wire [3-1:0] node1979;
	wire [3-1:0] node1982;
	wire [3-1:0] node1983;
	wire [3-1:0] node1987;
	wire [3-1:0] node1988;
	wire [3-1:0] node1991;
	wire [3-1:0] node1994;
	wire [3-1:0] node1995;
	wire [3-1:0] node1996;
	wire [3-1:0] node2000;
	wire [3-1:0] node2001;
	wire [3-1:0] node2002;
	wire [3-1:0] node2006;
	wire [3-1:0] node2007;
	wire [3-1:0] node2011;
	wire [3-1:0] node2012;
	wire [3-1:0] node2013;
	wire [3-1:0] node2014;
	wire [3-1:0] node2019;
	wire [3-1:0] node2020;
	wire [3-1:0] node2021;
	wire [3-1:0] node2022;
	wire [3-1:0] node2026;
	wire [3-1:0] node2029;
	wire [3-1:0] node2032;
	wire [3-1:0] node2033;
	wire [3-1:0] node2034;
	wire [3-1:0] node2035;
	wire [3-1:0] node2036;
	wire [3-1:0] node2037;
	wire [3-1:0] node2038;
	wire [3-1:0] node2039;
	wire [3-1:0] node2043;
	wire [3-1:0] node2044;
	wire [3-1:0] node2046;
	wire [3-1:0] node2050;
	wire [3-1:0] node2051;
	wire [3-1:0] node2052;
	wire [3-1:0] node2053;
	wire [3-1:0] node2057;
	wire [3-1:0] node2058;
	wire [3-1:0] node2062;
	wire [3-1:0] node2063;
	wire [3-1:0] node2064;
	wire [3-1:0] node2067;
	wire [3-1:0] node2070;
	wire [3-1:0] node2071;
	wire [3-1:0] node2074;
	wire [3-1:0] node2077;
	wire [3-1:0] node2078;
	wire [3-1:0] node2079;
	wire [3-1:0] node2080;
	wire [3-1:0] node2081;
	wire [3-1:0] node2085;
	wire [3-1:0] node2086;
	wire [3-1:0] node2089;
	wire [3-1:0] node2092;
	wire [3-1:0] node2093;
	wire [3-1:0] node2095;
	wire [3-1:0] node2098;
	wire [3-1:0] node2099;
	wire [3-1:0] node2103;
	wire [3-1:0] node2104;
	wire [3-1:0] node2105;
	wire [3-1:0] node2107;
	wire [3-1:0] node2111;
	wire [3-1:0] node2112;
	wire [3-1:0] node2113;
	wire [3-1:0] node2117;
	wire [3-1:0] node2120;
	wire [3-1:0] node2121;
	wire [3-1:0] node2122;
	wire [3-1:0] node2123;
	wire [3-1:0] node2124;
	wire [3-1:0] node2125;
	wire [3-1:0] node2128;
	wire [3-1:0] node2131;
	wire [3-1:0] node2134;
	wire [3-1:0] node2136;
	wire [3-1:0] node2138;
	wire [3-1:0] node2141;
	wire [3-1:0] node2142;
	wire [3-1:0] node2143;
	wire [3-1:0] node2144;
	wire [3-1:0] node2148;
	wire [3-1:0] node2150;
	wire [3-1:0] node2153;
	wire [3-1:0] node2154;
	wire [3-1:0] node2155;
	wire [3-1:0] node2158;
	wire [3-1:0] node2161;
	wire [3-1:0] node2162;
	wire [3-1:0] node2166;
	wire [3-1:0] node2167;
	wire [3-1:0] node2168;
	wire [3-1:0] node2169;
	wire [3-1:0] node2171;
	wire [3-1:0] node2174;
	wire [3-1:0] node2175;
	wire [3-1:0] node2179;
	wire [3-1:0] node2180;
	wire [3-1:0] node2183;
	wire [3-1:0] node2186;
	wire [3-1:0] node2187;
	wire [3-1:0] node2188;
	wire [3-1:0] node2190;
	wire [3-1:0] node2193;
	wire [3-1:0] node2195;
	wire [3-1:0] node2198;
	wire [3-1:0] node2199;
	wire [3-1:0] node2202;
	wire [3-1:0] node2205;
	wire [3-1:0] node2206;
	wire [3-1:0] node2207;
	wire [3-1:0] node2208;
	wire [3-1:0] node2209;
	wire [3-1:0] node2210;
	wire [3-1:0] node2211;
	wire [3-1:0] node2215;
	wire [3-1:0] node2216;
	wire [3-1:0] node2220;
	wire [3-1:0] node2221;
	wire [3-1:0] node2222;
	wire [3-1:0] node2225;
	wire [3-1:0] node2229;
	wire [3-1:0] node2230;
	wire [3-1:0] node2231;
	wire [3-1:0] node2233;
	wire [3-1:0] node2236;
	wire [3-1:0] node2237;
	wire [3-1:0] node2241;
	wire [3-1:0] node2242;
	wire [3-1:0] node2243;
	wire [3-1:0] node2246;
	wire [3-1:0] node2249;
	wire [3-1:0] node2251;
	wire [3-1:0] node2254;
	wire [3-1:0] node2255;
	wire [3-1:0] node2256;
	wire [3-1:0] node2258;
	wire [3-1:0] node2259;
	wire [3-1:0] node2262;
	wire [3-1:0] node2265;
	wire [3-1:0] node2266;
	wire [3-1:0] node2269;
	wire [3-1:0] node2272;
	wire [3-1:0] node2273;
	wire [3-1:0] node2274;
	wire [3-1:0] node2277;
	wire [3-1:0] node2279;
	wire [3-1:0] node2282;
	wire [3-1:0] node2283;
	wire [3-1:0] node2286;
	wire [3-1:0] node2289;
	wire [3-1:0] node2290;
	wire [3-1:0] node2291;
	wire [3-1:0] node2292;
	wire [3-1:0] node2293;
	wire [3-1:0] node2295;
	wire [3-1:0] node2298;
	wire [3-1:0] node2299;
	wire [3-1:0] node2303;
	wire [3-1:0] node2304;
	wire [3-1:0] node2305;
	wire [3-1:0] node2309;
	wire [3-1:0] node2311;
	wire [3-1:0] node2314;
	wire [3-1:0] node2315;
	wire [3-1:0] node2316;
	wire [3-1:0] node2317;
	wire [3-1:0] node2322;
	wire [3-1:0] node2323;
	wire [3-1:0] node2326;
	wire [3-1:0] node2329;
	wire [3-1:0] node2330;
	wire [3-1:0] node2331;
	wire [3-1:0] node2332;
	wire [3-1:0] node2333;
	wire [3-1:0] node2336;
	wire [3-1:0] node2339;
	wire [3-1:0] node2342;
	wire [3-1:0] node2343;
	wire [3-1:0] node2345;
	wire [3-1:0] node2348;
	wire [3-1:0] node2349;
	wire [3-1:0] node2353;
	wire [3-1:0] node2354;
	wire [3-1:0] node2355;
	wire [3-1:0] node2357;
	wire [3-1:0] node2360;
	wire [3-1:0] node2362;
	wire [3-1:0] node2365;
	wire [3-1:0] node2366;
	wire [3-1:0] node2369;
	wire [3-1:0] node2372;
	wire [3-1:0] node2373;
	wire [3-1:0] node2374;
	wire [3-1:0] node2375;
	wire [3-1:0] node2376;
	wire [3-1:0] node2377;
	wire [3-1:0] node2378;
	wire [3-1:0] node2380;
	wire [3-1:0] node2383;
	wire [3-1:0] node2384;
	wire [3-1:0] node2387;
	wire [3-1:0] node2390;
	wire [3-1:0] node2391;
	wire [3-1:0] node2392;
	wire [3-1:0] node2395;
	wire [3-1:0] node2398;
	wire [3-1:0] node2401;
	wire [3-1:0] node2402;
	wire [3-1:0] node2403;
	wire [3-1:0] node2404;
	wire [3-1:0] node2408;
	wire [3-1:0] node2409;
	wire [3-1:0] node2412;
	wire [3-1:0] node2415;
	wire [3-1:0] node2416;
	wire [3-1:0] node2418;
	wire [3-1:0] node2421;
	wire [3-1:0] node2422;
	wire [3-1:0] node2426;
	wire [3-1:0] node2427;
	wire [3-1:0] node2428;
	wire [3-1:0] node2429;
	wire [3-1:0] node2432;
	wire [3-1:0] node2435;
	wire [3-1:0] node2436;
	wire [3-1:0] node2437;
	wire [3-1:0] node2442;
	wire [3-1:0] node2443;
	wire [3-1:0] node2444;
	wire [3-1:0] node2445;
	wire [3-1:0] node2448;
	wire [3-1:0] node2452;
	wire [3-1:0] node2453;
	wire [3-1:0] node2454;
	wire [3-1:0] node2457;
	wire [3-1:0] node2461;
	wire [3-1:0] node2462;
	wire [3-1:0] node2463;
	wire [3-1:0] node2464;
	wire [3-1:0] node2465;
	wire [3-1:0] node2466;
	wire [3-1:0] node2469;
	wire [3-1:0] node2472;
	wire [3-1:0] node2475;
	wire [3-1:0] node2476;
	wire [3-1:0] node2477;
	wire [3-1:0] node2481;
	wire [3-1:0] node2483;
	wire [3-1:0] node2486;
	wire [3-1:0] node2487;
	wire [3-1:0] node2488;
	wire [3-1:0] node2490;
	wire [3-1:0] node2493;
	wire [3-1:0] node2494;
	wire [3-1:0] node2498;
	wire [3-1:0] node2499;
	wire [3-1:0] node2502;
	wire [3-1:0] node2505;
	wire [3-1:0] node2506;
	wire [3-1:0] node2507;
	wire [3-1:0] node2508;
	wire [3-1:0] node2511;
	wire [3-1:0] node2512;
	wire [3-1:0] node2516;
	wire [3-1:0] node2517;
	wire [3-1:0] node2520;
	wire [3-1:0] node2523;
	wire [3-1:0] node2524;
	wire [3-1:0] node2525;
	wire [3-1:0] node2526;
	wire [3-1:0] node2530;
	wire [3-1:0] node2531;
	wire [3-1:0] node2534;
	wire [3-1:0] node2537;
	wire [3-1:0] node2538;
	wire [3-1:0] node2539;
	wire [3-1:0] node2542;
	wire [3-1:0] node2545;
	wire [3-1:0] node2547;
	wire [3-1:0] node2550;
	wire [3-1:0] node2551;
	wire [3-1:0] node2552;
	wire [3-1:0] node2553;
	wire [3-1:0] node2554;
	wire [3-1:0] node2555;
	wire [3-1:0] node2556;
	wire [3-1:0] node2559;
	wire [3-1:0] node2562;
	wire [3-1:0] node2565;
	wire [3-1:0] node2566;
	wire [3-1:0] node2569;
	wire [3-1:0] node2572;
	wire [3-1:0] node2573;
	wire [3-1:0] node2574;
	wire [3-1:0] node2576;
	wire [3-1:0] node2579;
	wire [3-1:0] node2582;
	wire [3-1:0] node2583;
	wire [3-1:0] node2584;
	wire [3-1:0] node2588;
	wire [3-1:0] node2590;
	wire [3-1:0] node2593;
	wire [3-1:0] node2594;
	wire [3-1:0] node2595;
	wire [3-1:0] node2597;
	wire [3-1:0] node2598;
	wire [3-1:0] node2601;
	wire [3-1:0] node2604;
	wire [3-1:0] node2605;
	wire [3-1:0] node2606;
	wire [3-1:0] node2609;
	wire [3-1:0] node2612;
	wire [3-1:0] node2613;
	wire [3-1:0] node2617;
	wire [3-1:0] node2618;
	wire [3-1:0] node2619;
	wire [3-1:0] node2623;
	wire [3-1:0] node2625;
	wire [3-1:0] node2626;
	wire [3-1:0] node2630;
	wire [3-1:0] node2631;
	wire [3-1:0] node2632;
	wire [3-1:0] node2633;
	wire [3-1:0] node2634;
	wire [3-1:0] node2636;
	wire [3-1:0] node2639;
	wire [3-1:0] node2641;
	wire [3-1:0] node2644;
	wire [3-1:0] node2645;
	wire [3-1:0] node2646;
	wire [3-1:0] node2650;
	wire [3-1:0] node2652;
	wire [3-1:0] node2655;
	wire [3-1:0] node2656;
	wire [3-1:0] node2657;
	wire [3-1:0] node2658;
	wire [3-1:0] node2662;
	wire [3-1:0] node2664;
	wire [3-1:0] node2667;
	wire [3-1:0] node2668;
	wire [3-1:0] node2671;
	wire [3-1:0] node2674;
	wire [3-1:0] node2675;
	wire [3-1:0] node2676;
	wire [3-1:0] node2677;
	wire [3-1:0] node2679;
	wire [3-1:0] node2682;
	wire [3-1:0] node2684;
	wire [3-1:0] node2687;
	wire [3-1:0] node2688;
	wire [3-1:0] node2691;
	wire [3-1:0] node2694;
	wire [3-1:0] node2695;
	wire [3-1:0] node2696;
	wire [3-1:0] node2697;
	wire [3-1:0] node2700;
	wire [3-1:0] node2703;
	wire [3-1:0] node2704;
	wire [3-1:0] node2708;
	wire [3-1:0] node2710;

	assign outp = (inp[2]) ? node1374 : node1;
		assign node1 = (inp[4]) ? node665 : node2;
			assign node2 = (inp[8]) ? node336 : node3;
				assign node3 = (inp[5]) ? node175 : node4;
					assign node4 = (inp[3]) ? node98 : node5;
						assign node5 = (inp[0]) ? node51 : node6;
							assign node6 = (inp[6]) ? node26 : node7;
								assign node7 = (inp[10]) ? node13 : node8;
									assign node8 = (inp[7]) ? node10 : 3'b010;
										assign node10 = (inp[9]) ? 3'b011 : 3'b010;
									assign node13 = (inp[1]) ? node19 : node14;
										assign node14 = (inp[11]) ? 3'b110 : node15;
											assign node15 = (inp[9]) ? 3'b010 : 3'b010;
										assign node19 = (inp[9]) ? node23 : node20;
											assign node20 = (inp[7]) ? 3'b110 : 3'b111;
											assign node23 = (inp[11]) ? 3'b110 : 3'b111;
								assign node26 = (inp[10]) ? node40 : node27;
									assign node27 = (inp[1]) ? node35 : node28;
										assign node28 = (inp[11]) ? node32 : node29;
											assign node29 = (inp[7]) ? 3'b010 : 3'b011;
											assign node32 = (inp[9]) ? 3'b110 : 3'b111;
										assign node35 = (inp[11]) ? 3'b110 : node36;
											assign node36 = (inp[9]) ? 3'b111 : 3'b110;
									assign node40 = (inp[1]) ? node46 : node41;
										assign node41 = (inp[11]) ? 3'b011 : node42;
											assign node42 = (inp[7]) ? 3'b111 : 3'b110;
										assign node46 = (inp[7]) ? 3'b011 : node47;
											assign node47 = (inp[9]) ? 3'b010 : 3'b011;
							assign node51 = (inp[10]) ? node73 : node52;
								assign node52 = (inp[6]) ? node62 : node53;
									assign node53 = (inp[7]) ? node57 : node54;
										assign node54 = (inp[9]) ? 3'b010 : 3'b011;
										assign node57 = (inp[11]) ? 3'b011 : node58;
											assign node58 = (inp[1]) ? 3'b011 : 3'b111;
									assign node62 = (inp[9]) ? node68 : node63;
										assign node63 = (inp[7]) ? 3'b110 : node64;
											assign node64 = (inp[1]) ? 3'b111 : 3'b011;
										assign node68 = (inp[7]) ? 3'b111 : node69;
											assign node69 = (inp[11]) ? 3'b110 : 3'b010;
								assign node73 = (inp[6]) ? node87 : node74;
									assign node74 = (inp[1]) ? node80 : node75;
										assign node75 = (inp[11]) ? node77 : 3'b010;
											assign node77 = (inp[7]) ? 3'b110 : 3'b110;
										assign node80 = (inp[11]) ? node84 : node81;
											assign node81 = (inp[9]) ? 3'b111 : 3'b110;
											assign node84 = (inp[7]) ? 3'b110 : 3'b110;
									assign node87 = (inp[1]) ? node93 : node88;
										assign node88 = (inp[11]) ? node90 : 3'b110;
											assign node90 = (inp[7]) ? 3'b010 : 3'b011;
										assign node93 = (inp[9]) ? node95 : 3'b010;
											assign node95 = (inp[7]) ? 3'b011 : 3'b010;
						assign node98 = (inp[10]) ? node140 : node99;
							assign node99 = (inp[6]) ? node121 : node100;
								assign node100 = (inp[1]) ? node112 : node101;
									assign node101 = (inp[11]) ? node107 : node102;
										assign node102 = (inp[9]) ? 3'b110 : node103;
											assign node103 = (inp[7]) ? 3'b110 : 3'b111;
										assign node107 = (inp[9]) ? node109 : 3'b010;
											assign node109 = (inp[7]) ? 3'b011 : 3'b010;
									assign node112 = (inp[0]) ? node118 : node113;
										assign node113 = (inp[11]) ? 3'b011 : node114;
											assign node114 = (inp[9]) ? 3'b010 : 3'b011;
										assign node118 = (inp[7]) ? 3'b010 : 3'b011;
								assign node121 = (inp[1]) ? node133 : node122;
									assign node122 = (inp[11]) ? node130 : node123;
										assign node123 = (inp[0]) ? node127 : node124;
											assign node124 = (inp[7]) ? 3'b011 : 3'b010;
											assign node127 = (inp[7]) ? 3'b010 : 3'b011;
										assign node130 = (inp[9]) ? 3'b101 : 3'b100;
									assign node133 = (inp[7]) ? node137 : node134;
										assign node134 = (inp[9]) ? 3'b100 : 3'b101;
										assign node137 = (inp[9]) ? 3'b101 : 3'b100;
							assign node140 = (inp[6]) ? node156 : node141;
								assign node141 = (inp[1]) ? node149 : node142;
									assign node142 = (inp[11]) ? node144 : 3'b010;
										assign node144 = (inp[7]) ? 3'b100 : node145;
											assign node145 = (inp[9]) ? 3'b100 : 3'b101;
									assign node149 = (inp[7]) ? node153 : node150;
										assign node150 = (inp[9]) ? 3'b100 : 3'b101;
										assign node153 = (inp[9]) ? 3'b101 : 3'b100;
								assign node156 = (inp[1]) ? node168 : node157;
									assign node157 = (inp[11]) ? node163 : node158;
										assign node158 = (inp[0]) ? node160 : 3'b100;
											assign node160 = (inp[7]) ? 3'b101 : 3'b100;
										assign node163 = (inp[9]) ? node165 : 3'b000;
											assign node165 = (inp[7]) ? 3'b001 : 3'b000;
									assign node168 = (inp[7]) ? node172 : node169;
										assign node169 = (inp[11]) ? 3'b000 : 3'b001;
										assign node172 = (inp[9]) ? 3'b001 : 3'b000;
					assign node175 = (inp[3]) ? node247 : node176;
						assign node176 = (inp[10]) ? node204 : node177;
							assign node177 = (inp[11]) ? node191 : node178;
								assign node178 = (inp[1]) ? node188 : node179;
									assign node179 = (inp[6]) ? node181 : 3'b111;
										assign node181 = (inp[9]) ? node185 : node182;
											assign node182 = (inp[7]) ? 3'b010 : 3'b011;
											assign node185 = (inp[7]) ? 3'b011 : 3'b010;
									assign node188 = (inp[6]) ? 3'b101 : 3'b011;
								assign node191 = (inp[6]) ? node197 : node192;
									assign node192 = (inp[7]) ? node194 : 3'b011;
										assign node194 = (inp[9]) ? 3'b011 : 3'b010;
									assign node197 = (inp[0]) ? 3'b101 : node198;
										assign node198 = (inp[7]) ? 3'b100 : node199;
											assign node199 = (inp[9]) ? 3'b100 : 3'b101;
							assign node204 = (inp[6]) ? node224 : node205;
								assign node205 = (inp[11]) ? node217 : node206;
									assign node206 = (inp[1]) ? node212 : node207;
										assign node207 = (inp[0]) ? node209 : 3'b011;
											assign node209 = (inp[7]) ? 3'b011 : 3'b010;
										assign node212 = (inp[9]) ? node214 : 3'b100;
											assign node214 = (inp[7]) ? 3'b101 : 3'b100;
									assign node217 = (inp[7]) ? node221 : node218;
										assign node218 = (inp[9]) ? 3'b100 : 3'b101;
										assign node221 = (inp[9]) ? 3'b101 : 3'b100;
								assign node224 = (inp[1]) ? node236 : node225;
									assign node225 = (inp[11]) ? node231 : node226;
										assign node226 = (inp[9]) ? node228 : 3'b101;
											assign node228 = (inp[7]) ? 3'b101 : 3'b100;
										assign node231 = (inp[7]) ? 3'b001 : node232;
											assign node232 = (inp[0]) ? 3'b001 : 3'b000;
									assign node236 = (inp[0]) ? node242 : node237;
										assign node237 = (inp[9]) ? 3'b001 : node238;
											assign node238 = (inp[7]) ? 3'b000 : 3'b001;
										assign node242 = (inp[11]) ? 3'b000 : node243;
											assign node243 = (inp[9]) ? 3'b000 : 3'b001;
						assign node247 = (inp[6]) ? node283 : node248;
							assign node248 = (inp[10]) ? node262 : node249;
								assign node249 = (inp[11]) ? node257 : node250;
									assign node250 = (inp[1]) ? 3'b001 : node251;
										assign node251 = (inp[9]) ? node253 : 3'b101;
											assign node253 = (inp[7]) ? 3'b101 : 3'b100;
									assign node257 = (inp[7]) ? node259 : 3'b001;
										assign node259 = (inp[9]) ? 3'b001 : 3'b000;
								assign node262 = (inp[1]) ? node274 : node263;
									assign node263 = (inp[11]) ? node269 : node264;
										assign node264 = (inp[7]) ? node266 : 3'b001;
											assign node266 = (inp[9]) ? 3'b001 : 3'b000;
										assign node269 = (inp[0]) ? 3'b101 : node270;
											assign node270 = (inp[9]) ? 3'b101 : 3'b100;
									assign node274 = (inp[0]) ? node276 : 3'b101;
										assign node276 = (inp[11]) ? node280 : node277;
											assign node277 = (inp[7]) ? 3'b101 : 3'b100;
											assign node280 = (inp[9]) ? 3'b100 : 3'b100;
							assign node283 = (inp[10]) ? node311 : node284;
								assign node284 = (inp[11]) ? node298 : node285;
									assign node285 = (inp[1]) ? node293 : node286;
										assign node286 = (inp[9]) ? node290 : node287;
											assign node287 = (inp[0]) ? 3'b000 : 3'b001;
											assign node290 = (inp[7]) ? 3'b001 : 3'b000;
										assign node293 = (inp[9]) ? node295 : 3'b101;
											assign node295 = (inp[7]) ? 3'b101 : 3'b100;
									assign node298 = (inp[1]) ? node304 : node299;
										assign node299 = (inp[7]) ? node301 : 3'b101;
											assign node301 = (inp[0]) ? 3'b101 : 3'b100;
										assign node304 = (inp[9]) ? node308 : node305;
											assign node305 = (inp[7]) ? 3'b100 : 3'b101;
											assign node308 = (inp[7]) ? 3'b101 : 3'b100;
								assign node311 = (inp[11]) ? node323 : node312;
									assign node312 = (inp[1]) ? node320 : node313;
										assign node313 = (inp[7]) ? node317 : node314;
											assign node314 = (inp[9]) ? 3'b100 : 3'b101;
											assign node317 = (inp[9]) ? 3'b101 : 3'b100;
										assign node320 = (inp[0]) ? 3'b000 : 3'b001;
									assign node323 = (inp[1]) ? node331 : node324;
										assign node324 = (inp[9]) ? node328 : node325;
											assign node325 = (inp[7]) ? 3'b000 : 3'b001;
											assign node328 = (inp[7]) ? 3'b001 : 3'b000;
										assign node331 = (inp[0]) ? 3'b000 : node332;
											assign node332 = (inp[9]) ? 3'b000 : 3'b000;
				assign node336 = (inp[5]) ? node492 : node337;
					assign node337 = (inp[3]) ? node421 : node338;
						assign node338 = (inp[6]) ? node380 : node339;
							assign node339 = (inp[10]) ? node359 : node340;
								assign node340 = (inp[1]) ? node352 : node341;
									assign node341 = (inp[11]) ? node347 : node342;
										assign node342 = (inp[9]) ? 3'b100 : node343;
											assign node343 = (inp[7]) ? 3'b100 : 3'b101;
										assign node347 = (inp[7]) ? node349 : 3'b000;
											assign node349 = (inp[9]) ? 3'b001 : 3'b000;
									assign node352 = (inp[9]) ? node356 : node353;
										assign node353 = (inp[7]) ? 3'b000 : 3'b001;
										assign node356 = (inp[7]) ? 3'b001 : 3'b000;
								assign node359 = (inp[1]) ? node373 : node360;
									assign node360 = (inp[11]) ? node368 : node361;
										assign node361 = (inp[7]) ? node365 : node362;
											assign node362 = (inp[9]) ? 3'b000 : 3'b001;
											assign node365 = (inp[9]) ? 3'b001 : 3'b000;
										assign node368 = (inp[9]) ? 3'b101 : node369;
											assign node369 = (inp[7]) ? 3'b100 : 3'b101;
									assign node373 = (inp[0]) ? node375 : 3'b101;
										assign node375 = (inp[7]) ? 3'b100 : node376;
											assign node376 = (inp[9]) ? 3'b100 : 3'b101;
							assign node380 = (inp[10]) ? node398 : node381;
								assign node381 = (inp[1]) ? node385 : node382;
									assign node382 = (inp[11]) ? 3'b101 : 3'b001;
									assign node385 = (inp[0]) ? node393 : node386;
										assign node386 = (inp[9]) ? node390 : node387;
											assign node387 = (inp[7]) ? 3'b100 : 3'b101;
											assign node390 = (inp[7]) ? 3'b101 : 3'b100;
										assign node393 = (inp[7]) ? node395 : 3'b100;
											assign node395 = (inp[9]) ? 3'b101 : 3'b100;
								assign node398 = (inp[1]) ? node406 : node399;
									assign node399 = (inp[11]) ? 3'b001 : node400;
										assign node400 = (inp[7]) ? node402 : 3'b101;
											assign node402 = (inp[9]) ? 3'b101 : 3'b100;
									assign node406 = (inp[0]) ? node414 : node407;
										assign node407 = (inp[9]) ? node411 : node408;
											assign node408 = (inp[7]) ? 3'b000 : 3'b001;
											assign node411 = (inp[7]) ? 3'b001 : 3'b000;
										assign node414 = (inp[7]) ? node418 : node415;
											assign node415 = (inp[9]) ? 3'b000 : 3'b001;
											assign node418 = (inp[9]) ? 3'b001 : 3'b000;
						assign node421 = (inp[10]) ? node457 : node422;
							assign node422 = (inp[6]) ? node440 : node423;
								assign node423 = (inp[1]) ? node433 : node424;
									assign node424 = (inp[11]) ? node430 : node425;
										assign node425 = (inp[0]) ? node427 : 3'b100;
											assign node427 = (inp[7]) ? 3'b101 : 3'b100;
										assign node430 = (inp[0]) ? 3'b000 : 3'b001;
									assign node433 = (inp[7]) ? node437 : node434;
										assign node434 = (inp[9]) ? 3'b000 : 3'b001;
										assign node437 = (inp[9]) ? 3'b001 : 3'b000;
								assign node440 = (inp[1]) ? node450 : node441;
									assign node441 = (inp[11]) ? node447 : node442;
										assign node442 = (inp[7]) ? 3'b001 : node443;
											assign node443 = (inp[9]) ? 3'b000 : 3'b001;
										assign node447 = (inp[0]) ? 3'b110 : 3'b111;
									assign node450 = (inp[9]) ? 3'b111 : node451;
										assign node451 = (inp[0]) ? node453 : 3'b110;
											assign node453 = (inp[7]) ? 3'b111 : 3'b110;
							assign node457 = (inp[6]) ? node475 : node458;
								assign node458 = (inp[1]) ? node470 : node459;
									assign node459 = (inp[11]) ? node465 : node460;
										assign node460 = (inp[0]) ? node462 : 3'b000;
											assign node462 = (inp[9]) ? 3'b000 : 3'b001;
										assign node465 = (inp[7]) ? 3'b111 : node466;
											assign node466 = (inp[9]) ? 3'b110 : 3'b111;
									assign node470 = (inp[11]) ? node472 : 3'b111;
										assign node472 = (inp[7]) ? 3'b110 : 3'b111;
								assign node475 = (inp[1]) ? node481 : node476;
									assign node476 = (inp[11]) ? 3'b010 : node477;
										assign node477 = (inp[7]) ? 3'b111 : 3'b110;
									assign node481 = (inp[11]) ? node487 : node482;
										assign node482 = (inp[9]) ? node484 : 3'b010;
											assign node484 = (inp[0]) ? 3'b010 : 3'b011;
										assign node487 = (inp[9]) ? node489 : 3'b011;
											assign node489 = (inp[7]) ? 3'b010 : 3'b011;
					assign node492 = (inp[3]) ? node586 : node493;
						assign node493 = (inp[10]) ? node541 : node494;
							assign node494 = (inp[6]) ? node516 : node495;
								assign node495 = (inp[1]) ? node505 : node496;
									assign node496 = (inp[11]) ? node500 : node497;
										assign node497 = (inp[7]) ? 3'b100 : 3'b101;
										assign node500 = (inp[9]) ? 3'b001 : node501;
											assign node501 = (inp[7]) ? 3'b000 : 3'b001;
									assign node505 = (inp[11]) ? node511 : node506;
										assign node506 = (inp[9]) ? 3'b001 : node507;
											assign node507 = (inp[7]) ? 3'b000 : 3'b001;
										assign node511 = (inp[9]) ? 3'b000 : node512;
											assign node512 = (inp[7]) ? 3'b000 : 3'b001;
								assign node516 = (inp[1]) ? node530 : node517;
									assign node517 = (inp[11]) ? node523 : node518;
										assign node518 = (inp[0]) ? node520 : 3'b000;
											assign node520 = (inp[9]) ? 3'b000 : 3'b000;
										assign node523 = (inp[7]) ? node527 : node524;
											assign node524 = (inp[0]) ? 3'b110 : 3'b110;
											assign node527 = (inp[0]) ? 3'b111 : 3'b110;
									assign node530 = (inp[9]) ? node536 : node531;
										assign node531 = (inp[7]) ? 3'b110 : node532;
											assign node532 = (inp[0]) ? 3'b110 : 3'b111;
										assign node536 = (inp[7]) ? node538 : 3'b111;
											assign node538 = (inp[0]) ? 3'b110 : 3'b111;
							assign node541 = (inp[6]) ? node563 : node542;
								assign node542 = (inp[11]) ? node554 : node543;
									assign node543 = (inp[1]) ? node549 : node544;
										assign node544 = (inp[7]) ? 3'b001 : node545;
											assign node545 = (inp[9]) ? 3'b000 : 3'b001;
										assign node549 = (inp[0]) ? node551 : 3'b111;
											assign node551 = (inp[7]) ? 3'b110 : 3'b111;
									assign node554 = (inp[0]) ? node560 : node555;
										assign node555 = (inp[1]) ? 3'b110 : node556;
											assign node556 = (inp[7]) ? 3'b110 : 3'b111;
										assign node560 = (inp[1]) ? 3'b111 : 3'b110;
								assign node563 = (inp[1]) ? node577 : node564;
									assign node564 = (inp[11]) ? node570 : node565;
										assign node565 = (inp[0]) ? 3'b110 : node566;
											assign node566 = (inp[7]) ? 3'b110 : 3'b110;
										assign node570 = (inp[0]) ? node574 : node571;
											assign node571 = (inp[9]) ? 3'b010 : 3'b010;
											assign node574 = (inp[7]) ? 3'b010 : 3'b011;
									assign node577 = (inp[0]) ? node583 : node578;
										assign node578 = (inp[11]) ? 3'b011 : node579;
											assign node579 = (inp[7]) ? 3'b010 : 3'b010;
										assign node583 = (inp[11]) ? 3'b010 : 3'b011;
						assign node586 = (inp[0]) ? node626 : node587;
							assign node587 = (inp[7]) ? node607 : node588;
								assign node588 = (inp[9]) ? node596 : node589;
									assign node589 = (inp[6]) ? 3'b011 : node590;
										assign node590 = (inp[1]) ? node592 : 3'b111;
											assign node592 = (inp[11]) ? 3'b111 : 3'b011;
									assign node596 = (inp[11]) ? node602 : node597;
										assign node597 = (inp[10]) ? node599 : 3'b010;
											assign node599 = (inp[1]) ? 3'b010 : 3'b110;
										assign node602 = (inp[6]) ? node604 : 3'b010;
											assign node604 = (inp[10]) ? 3'b010 : 3'b110;
								assign node607 = (inp[9]) ? node617 : node608;
									assign node608 = (inp[6]) ? node614 : node609;
										assign node609 = (inp[10]) ? node611 : 3'b010;
											assign node611 = (inp[1]) ? 3'b110 : 3'b010;
										assign node614 = (inp[10]) ? 3'b010 : 3'b110;
									assign node617 = (inp[1]) ? node619 : 3'b111;
										assign node619 = (inp[6]) ? node623 : node620;
											assign node620 = (inp[10]) ? 3'b111 : 3'b011;
											assign node623 = (inp[10]) ? 3'b011 : 3'b111;
							assign node626 = (inp[11]) ? node650 : node627;
								assign node627 = (inp[1]) ? node641 : node628;
									assign node628 = (inp[9]) ? node636 : node629;
										assign node629 = (inp[7]) ? node633 : node630;
											assign node630 = (inp[10]) ? 3'b110 : 3'b010;
											assign node633 = (inp[6]) ? 3'b011 : 3'b011;
										assign node636 = (inp[7]) ? node638 : 3'b111;
											assign node638 = (inp[10]) ? 3'b010 : 3'b110;
									assign node641 = (inp[10]) ? node645 : node642;
										assign node642 = (inp[6]) ? 3'b110 : 3'b010;
										assign node645 = (inp[6]) ? 3'b010 : node646;
											assign node646 = (inp[9]) ? 3'b110 : 3'b110;
								assign node650 = (inp[10]) ? node654 : node651;
									assign node651 = (inp[6]) ? 3'b111 : 3'b011;
									assign node654 = (inp[6]) ? node662 : node655;
										assign node655 = (inp[1]) ? node659 : node656;
											assign node656 = (inp[9]) ? 3'b110 : 3'b110;
											assign node659 = (inp[7]) ? 3'b110 : 3'b111;
										assign node662 = (inp[1]) ? 3'b011 : 3'b010;
			assign node665 = (inp[8]) ? node1019 : node666;
				assign node666 = (inp[3]) ? node862 : node667;
					assign node667 = (inp[5]) ? node757 : node668;
						assign node668 = (inp[0]) ? node712 : node669;
							assign node669 = (inp[10]) ? node697 : node670;
								assign node670 = (inp[6]) ? node682 : node671;
									assign node671 = (inp[1]) ? node677 : node672;
										assign node672 = (inp[7]) ? 3'b100 : node673;
											assign node673 = (inp[9]) ? 3'b100 : 3'b101;
										assign node677 = (inp[11]) ? node679 : 3'b001;
											assign node679 = (inp[7]) ? 3'b000 : 3'b000;
									assign node682 = (inp[11]) ? node690 : node683;
										assign node683 = (inp[1]) ? node687 : node684;
											assign node684 = (inp[9]) ? 3'b000 : 3'b000;
											assign node687 = (inp[9]) ? 3'b101 : 3'b100;
										assign node690 = (inp[1]) ? node694 : node691;
											assign node691 = (inp[9]) ? 3'b101 : 3'b100;
											assign node694 = (inp[9]) ? 3'b100 : 3'b100;
								assign node697 = (inp[1]) ? node705 : node698;
									assign node698 = (inp[6]) ? node702 : node699;
										assign node699 = (inp[11]) ? 3'b100 : 3'b000;
										assign node702 = (inp[7]) ? 3'b100 : 3'b101;
									assign node705 = (inp[6]) ? node707 : 3'b100;
										assign node707 = (inp[11]) ? node709 : 3'b000;
											assign node709 = (inp[9]) ? 3'b000 : 3'b000;
							assign node712 = (inp[10]) ? node738 : node713;
								assign node713 = (inp[6]) ? node725 : node714;
									assign node714 = (inp[1]) ? node720 : node715;
										assign node715 = (inp[11]) ? node717 : 3'b101;
											assign node717 = (inp[7]) ? 3'b000 : 3'b001;
										assign node720 = (inp[9]) ? node722 : 3'b000;
											assign node722 = (inp[7]) ? 3'b001 : 3'b000;
									assign node725 = (inp[1]) ? node733 : node726;
										assign node726 = (inp[11]) ? node730 : node727;
											assign node727 = (inp[9]) ? 3'b001 : 3'b000;
											assign node730 = (inp[7]) ? 3'b100 : 3'b100;
										assign node733 = (inp[11]) ? 3'b101 : node734;
											assign node734 = (inp[9]) ? 3'b100 : 3'b100;
								assign node738 = (inp[6]) ? node746 : node739;
									assign node739 = (inp[7]) ? node743 : node740;
										assign node740 = (inp[11]) ? 3'b101 : 3'b001;
										assign node743 = (inp[9]) ? 3'b101 : 3'b100;
									assign node746 = (inp[11]) ? node752 : node747;
										assign node747 = (inp[1]) ? 3'b001 : node748;
											assign node748 = (inp[9]) ? 3'b101 : 3'b100;
										assign node752 = (inp[9]) ? node754 : 3'b001;
											assign node754 = (inp[7]) ? 3'b001 : 3'b000;
						assign node757 = (inp[10]) ? node809 : node758;
							assign node758 = (inp[6]) ? node784 : node759;
								assign node759 = (inp[11]) ? node773 : node760;
									assign node760 = (inp[1]) ? node768 : node761;
										assign node761 = (inp[7]) ? node765 : node762;
											assign node762 = (inp[9]) ? 3'b100 : 3'b101;
											assign node765 = (inp[9]) ? 3'b101 : 3'b100;
										assign node768 = (inp[7]) ? node770 : 3'b000;
											assign node770 = (inp[0]) ? 3'b001 : 3'b000;
									assign node773 = (inp[1]) ? node779 : node774;
										assign node774 = (inp[7]) ? node776 : 3'b001;
											assign node776 = (inp[9]) ? 3'b001 : 3'b000;
										assign node779 = (inp[9]) ? node781 : 3'b001;
											assign node781 = (inp[7]) ? 3'b001 : 3'b000;
								assign node784 = (inp[11]) ? node798 : node785;
									assign node785 = (inp[1]) ? node793 : node786;
										assign node786 = (inp[9]) ? node790 : node787;
											assign node787 = (inp[7]) ? 3'b000 : 3'b001;
											assign node790 = (inp[7]) ? 3'b001 : 3'b000;
										assign node793 = (inp[7]) ? node795 : 3'b111;
											assign node795 = (inp[9]) ? 3'b110 : 3'b110;
									assign node798 = (inp[9]) ? node804 : node799;
										assign node799 = (inp[7]) ? node801 : 3'b110;
											assign node801 = (inp[1]) ? 3'b110 : 3'b111;
										assign node804 = (inp[1]) ? 3'b111 : node805;
											assign node805 = (inp[0]) ? 3'b110 : 3'b110;
							assign node809 = (inp[6]) ? node835 : node810;
								assign node810 = (inp[11]) ? node822 : node811;
									assign node811 = (inp[1]) ? node817 : node812;
										assign node812 = (inp[7]) ? 3'b001 : node813;
											assign node813 = (inp[9]) ? 3'b000 : 3'b001;
										assign node817 = (inp[7]) ? 3'b111 : node818;
											assign node818 = (inp[0]) ? 3'b110 : 3'b111;
									assign node822 = (inp[0]) ? node828 : node823;
										assign node823 = (inp[1]) ? node825 : 3'b110;
											assign node825 = (inp[7]) ? 3'b110 : 3'b110;
										assign node828 = (inp[9]) ? node832 : node829;
											assign node829 = (inp[7]) ? 3'b111 : 3'b110;
											assign node832 = (inp[7]) ? 3'b110 : 3'b111;
								assign node835 = (inp[1]) ? node847 : node836;
									assign node836 = (inp[11]) ? node842 : node837;
										assign node837 = (inp[7]) ? 3'b110 : node838;
											assign node838 = (inp[9]) ? 3'b111 : 3'b110;
										assign node842 = (inp[7]) ? node844 : 3'b011;
											assign node844 = (inp[9]) ? 3'b010 : 3'b010;
									assign node847 = (inp[0]) ? node855 : node848;
										assign node848 = (inp[11]) ? node852 : node849;
											assign node849 = (inp[9]) ? 3'b010 : 3'b010;
											assign node852 = (inp[7]) ? 3'b010 : 3'b010;
										assign node855 = (inp[9]) ? node859 : node856;
											assign node856 = (inp[7]) ? 3'b011 : 3'b010;
											assign node859 = (inp[7]) ? 3'b010 : 3'b011;
					assign node862 = (inp[5]) ? node936 : node863;
						assign node863 = (inp[6]) ? node899 : node864;
							assign node864 = (inp[10]) ? node882 : node865;
								assign node865 = (inp[11]) ? node875 : node866;
									assign node866 = (inp[1]) ? node872 : node867;
										assign node867 = (inp[0]) ? node869 : 3'b101;
											assign node869 = (inp[9]) ? 3'b100 : 3'b100;
										assign node872 = (inp[0]) ? 3'b001 : 3'b000;
									assign node875 = (inp[7]) ? node879 : node876;
										assign node876 = (inp[9]) ? 3'b000 : 3'b001;
										assign node879 = (inp[9]) ? 3'b001 : 3'b000;
								assign node882 = (inp[11]) ? node892 : node883;
									assign node883 = (inp[1]) ? node889 : node884;
										assign node884 = (inp[7]) ? 3'b000 : node885;
											assign node885 = (inp[9]) ? 3'b000 : 3'b001;
										assign node889 = (inp[9]) ? 3'b110 : 3'b111;
									assign node892 = (inp[7]) ? 3'b111 : node893;
										assign node893 = (inp[9]) ? 3'b110 : node894;
											assign node894 = (inp[0]) ? 3'b110 : 3'b111;
							assign node899 = (inp[10]) ? node919 : node900;
								assign node900 = (inp[11]) ? node908 : node901;
									assign node901 = (inp[1]) ? node903 : 3'b001;
										assign node903 = (inp[7]) ? node905 : 3'b111;
											assign node905 = (inp[9]) ? 3'b111 : 3'b110;
									assign node908 = (inp[0]) ? node914 : node909;
										assign node909 = (inp[7]) ? node911 : 3'b110;
											assign node911 = (inp[1]) ? 3'b110 : 3'b111;
										assign node914 = (inp[7]) ? node916 : 3'b111;
											assign node916 = (inp[9]) ? 3'b110 : 3'b111;
								assign node919 = (inp[11]) ? node929 : node920;
									assign node920 = (inp[1]) ? 3'b010 : node921;
										assign node921 = (inp[9]) ? node925 : node922;
											assign node922 = (inp[7]) ? 3'b110 : 3'b110;
											assign node925 = (inp[0]) ? 3'b110 : 3'b110;
									assign node929 = (inp[9]) ? node931 : 3'b010;
										assign node931 = (inp[0]) ? 3'b011 : node932;
											assign node932 = (inp[1]) ? 3'b010 : 3'b011;
						assign node936 = (inp[9]) ? node978 : node937;
							assign node937 = (inp[11]) ? node961 : node938;
								assign node938 = (inp[10]) ? node948 : node939;
									assign node939 = (inp[0]) ? node943 : node940;
										assign node940 = (inp[1]) ? 3'b011 : 3'b111;
										assign node943 = (inp[6]) ? node945 : 3'b011;
											assign node945 = (inp[1]) ? 3'b111 : 3'b011;
									assign node948 = (inp[6]) ? node954 : node949;
										assign node949 = (inp[1]) ? 3'b111 : node950;
											assign node950 = (inp[0]) ? 3'b010 : 3'b010;
										assign node954 = (inp[1]) ? node958 : node955;
											assign node955 = (inp[0]) ? 3'b110 : 3'b110;
											assign node958 = (inp[7]) ? 3'b010 : 3'b011;
								assign node961 = (inp[10]) ? node967 : node962;
									assign node962 = (inp[6]) ? 3'b110 : node963;
										assign node963 = (inp[1]) ? 3'b011 : 3'b010;
									assign node967 = (inp[6]) ? node973 : node968;
										assign node968 = (inp[7]) ? 3'b111 : node969;
											assign node969 = (inp[0]) ? 3'b110 : 3'b111;
										assign node973 = (inp[0]) ? 3'b011 : node974;
											assign node974 = (inp[7]) ? 3'b010 : 3'b011;
							assign node978 = (inp[1]) ? node994 : node979;
								assign node979 = (inp[0]) ? node985 : node980;
									assign node980 = (inp[11]) ? 3'b110 : node981;
										assign node981 = (inp[10]) ? 3'b010 : 3'b110;
									assign node985 = (inp[7]) ? 3'b110 : node986;
										assign node986 = (inp[6]) ? node990 : node987;
											assign node987 = (inp[11]) ? 3'b011 : 3'b011;
											assign node990 = (inp[11]) ? 3'b111 : 3'b011;
								assign node994 = (inp[7]) ? node1008 : node995;
									assign node995 = (inp[0]) ? node1003 : node996;
										assign node996 = (inp[6]) ? node1000 : node997;
											assign node997 = (inp[10]) ? 3'b110 : 3'b010;
											assign node1000 = (inp[10]) ? 3'b010 : 3'b110;
										assign node1003 = (inp[11]) ? 3'b111 : node1004;
											assign node1004 = (inp[6]) ? 3'b111 : 3'b011;
									assign node1008 = (inp[0]) ? node1014 : node1009;
										assign node1009 = (inp[11]) ? node1011 : 3'b011;
											assign node1011 = (inp[10]) ? 3'b011 : 3'b011;
										assign node1014 = (inp[6]) ? node1016 : 3'b010;
											assign node1016 = (inp[10]) ? 3'b010 : 3'b110;
				assign node1019 = (inp[3]) ? node1187 : node1020;
					assign node1020 = (inp[5]) ? node1102 : node1021;
						assign node1021 = (inp[7]) ? node1061 : node1022;
							assign node1022 = (inp[6]) ? node1046 : node1023;
								assign node1023 = (inp[10]) ? node1035 : node1024;
									assign node1024 = (inp[1]) ? node1028 : node1025;
										assign node1025 = (inp[11]) ? 3'b011 : 3'b110;
										assign node1028 = (inp[9]) ? node1032 : node1029;
											assign node1029 = (inp[0]) ? 3'b010 : 3'b011;
											assign node1032 = (inp[0]) ? 3'b011 : 3'b010;
									assign node1035 = (inp[11]) ? node1041 : node1036;
										assign node1036 = (inp[1]) ? 3'b111 : node1037;
											assign node1037 = (inp[9]) ? 3'b010 : 3'b010;
										assign node1041 = (inp[1]) ? 3'b111 : node1042;
											assign node1042 = (inp[9]) ? 3'b110 : 3'b110;
								assign node1046 = (inp[10]) ? node1054 : node1047;
									assign node1047 = (inp[1]) ? node1049 : 3'b010;
										assign node1049 = (inp[0]) ? node1051 : 3'b110;
											assign node1051 = (inp[9]) ? 3'b111 : 3'b110;
									assign node1054 = (inp[1]) ? node1056 : 3'b010;
										assign node1056 = (inp[0]) ? 3'b011 : node1057;
											assign node1057 = (inp[11]) ? 3'b011 : 3'b010;
							assign node1061 = (inp[10]) ? node1087 : node1062;
								assign node1062 = (inp[6]) ? node1076 : node1063;
									assign node1063 = (inp[1]) ? node1069 : node1064;
										assign node1064 = (inp[11]) ? 3'b011 : node1065;
											assign node1065 = (inp[0]) ? 3'b110 : 3'b110;
										assign node1069 = (inp[9]) ? node1073 : node1070;
											assign node1070 = (inp[0]) ? 3'b011 : 3'b010;
											assign node1073 = (inp[0]) ? 3'b010 : 3'b011;
									assign node1076 = (inp[1]) ? node1080 : node1077;
										assign node1077 = (inp[9]) ? 3'b110 : 3'b011;
										assign node1080 = (inp[9]) ? node1084 : node1081;
											assign node1081 = (inp[0]) ? 3'b111 : 3'b110;
											assign node1084 = (inp[11]) ? 3'b111 : 3'b110;
								assign node1087 = (inp[6]) ? node1095 : node1088;
									assign node1088 = (inp[0]) ? node1092 : node1089;
										assign node1089 = (inp[9]) ? 3'b111 : 3'b110;
										assign node1092 = (inp[9]) ? 3'b110 : 3'b111;
									assign node1095 = (inp[11]) ? node1099 : node1096;
										assign node1096 = (inp[0]) ? 3'b110 : 3'b111;
										assign node1099 = (inp[0]) ? 3'b011 : 3'b010;
						assign node1102 = (inp[6]) ? node1150 : node1103;
							assign node1103 = (inp[10]) ? node1129 : node1104;
								assign node1104 = (inp[11]) ? node1118 : node1105;
									assign node1105 = (inp[1]) ? node1113 : node1106;
										assign node1106 = (inp[0]) ? node1110 : node1107;
											assign node1107 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1110 = (inp[9]) ? 3'b110 : 3'b110;
										assign node1113 = (inp[9]) ? 3'b010 : node1114;
											assign node1114 = (inp[7]) ? 3'b010 : 3'b011;
									assign node1118 = (inp[1]) ? node1124 : node1119;
										assign node1119 = (inp[0]) ? node1121 : 3'b010;
											assign node1121 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1124 = (inp[0]) ? node1126 : 3'b011;
											assign node1126 = (inp[9]) ? 3'b010 : 3'b011;
								assign node1129 = (inp[1]) ? node1139 : node1130;
									assign node1130 = (inp[11]) ? node1136 : node1131;
										assign node1131 = (inp[0]) ? 3'b011 : node1132;
											assign node1132 = (inp[9]) ? 3'b010 : 3'b010;
										assign node1136 = (inp[9]) ? 3'b101 : 3'b100;
									assign node1139 = (inp[7]) ? node1145 : node1140;
										assign node1140 = (inp[11]) ? 3'b100 : node1141;
											assign node1141 = (inp[9]) ? 3'b101 : 3'b100;
										assign node1145 = (inp[0]) ? node1147 : 3'b101;
											assign node1147 = (inp[9]) ? 3'b100 : 3'b101;
							assign node1150 = (inp[10]) ? node1172 : node1151;
								assign node1151 = (inp[11]) ? node1159 : node1152;
									assign node1152 = (inp[1]) ? 3'b100 : node1153;
										assign node1153 = (inp[9]) ? 3'b011 : node1154;
											assign node1154 = (inp[0]) ? 3'b010 : 3'b010;
									assign node1159 = (inp[9]) ? node1165 : node1160;
										assign node1160 = (inp[0]) ? node1162 : 3'b100;
											assign node1162 = (inp[7]) ? 3'b101 : 3'b100;
										assign node1165 = (inp[0]) ? node1169 : node1166;
											assign node1166 = (inp[1]) ? 3'b100 : 3'b101;
											assign node1169 = (inp[1]) ? 3'b101 : 3'b100;
								assign node1172 = (inp[1]) ? node1180 : node1173;
									assign node1173 = (inp[11]) ? node1177 : node1174;
										assign node1174 = (inp[9]) ? 3'b101 : 3'b100;
										assign node1177 = (inp[7]) ? 3'b001 : 3'b000;
									assign node1180 = (inp[9]) ? 3'b001 : node1181;
										assign node1181 = (inp[7]) ? 3'b000 : node1182;
											assign node1182 = (inp[0]) ? 3'b000 : 3'b001;
					assign node1187 = (inp[5]) ? node1287 : node1188;
						assign node1188 = (inp[10]) ? node1232 : node1189;
							assign node1189 = (inp[6]) ? node1209 : node1190;
								assign node1190 = (inp[1]) ? node1200 : node1191;
									assign node1191 = (inp[11]) ? node1197 : node1192;
										assign node1192 = (inp[0]) ? 3'b110 : node1193;
											assign node1193 = (inp[7]) ? 3'b110 : 3'b111;
										assign node1197 = (inp[9]) ? 3'b010 : 3'b011;
									assign node1200 = (inp[7]) ? 3'b010 : node1201;
										assign node1201 = (inp[11]) ? node1205 : node1202;
											assign node1202 = (inp[0]) ? 3'b010 : 3'b010;
											assign node1205 = (inp[0]) ? 3'b010 : 3'b010;
								assign node1209 = (inp[11]) ? node1221 : node1210;
									assign node1210 = (inp[1]) ? node1216 : node1211;
										assign node1211 = (inp[7]) ? 3'b010 : node1212;
											assign node1212 = (inp[9]) ? 3'b010 : 3'b011;
										assign node1216 = (inp[7]) ? node1218 : 3'b100;
											assign node1218 = (inp[9]) ? 3'b101 : 3'b100;
									assign node1221 = (inp[9]) ? node1227 : node1222;
										assign node1222 = (inp[0]) ? 3'b101 : node1223;
											assign node1223 = (inp[7]) ? 3'b100 : 3'b101;
										assign node1227 = (inp[1]) ? 3'b100 : node1228;
											assign node1228 = (inp[0]) ? 3'b101 : 3'b100;
							assign node1232 = (inp[6]) ? node1260 : node1233;
								assign node1233 = (inp[1]) ? node1245 : node1234;
									assign node1234 = (inp[11]) ? node1240 : node1235;
										assign node1235 = (inp[0]) ? node1237 : 3'b011;
											assign node1237 = (inp[9]) ? 3'b010 : 3'b010;
										assign node1240 = (inp[0]) ? 3'b100 : node1241;
											assign node1241 = (inp[9]) ? 3'b101 : 3'b100;
									assign node1245 = (inp[9]) ? node1253 : node1246;
										assign node1246 = (inp[0]) ? node1250 : node1247;
											assign node1247 = (inp[11]) ? 3'b101 : 3'b100;
											assign node1250 = (inp[7]) ? 3'b101 : 3'b100;
										assign node1253 = (inp[0]) ? node1257 : node1254;
											assign node1254 = (inp[7]) ? 3'b101 : 3'b100;
											assign node1257 = (inp[7]) ? 3'b100 : 3'b101;
								assign node1260 = (inp[1]) ? node1272 : node1261;
									assign node1261 = (inp[11]) ? node1267 : node1262;
										assign node1262 = (inp[9]) ? node1264 : 3'b101;
											assign node1264 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1267 = (inp[0]) ? node1269 : 3'b000;
											assign node1269 = (inp[9]) ? 3'b001 : 3'b000;
									assign node1272 = (inp[0]) ? node1280 : node1273;
										assign node1273 = (inp[11]) ? node1277 : node1274;
											assign node1274 = (inp[7]) ? 3'b001 : 3'b000;
											assign node1277 = (inp[7]) ? 3'b000 : 3'b001;
										assign node1280 = (inp[9]) ? node1284 : node1281;
											assign node1281 = (inp[7]) ? 3'b001 : 3'b000;
											assign node1284 = (inp[7]) ? 3'b000 : 3'b001;
						assign node1287 = (inp[0]) ? node1329 : node1288;
							assign node1288 = (inp[11]) ? node1306 : node1289;
								assign node1289 = (inp[9]) ? node1297 : node1290;
									assign node1290 = (inp[7]) ? 3'b100 : node1291;
										assign node1291 = (inp[10]) ? node1293 : 3'b101;
											assign node1293 = (inp[6]) ? 3'b101 : 3'b001;
									assign node1297 = (inp[7]) ? node1301 : node1298;
										assign node1298 = (inp[10]) ? 3'b100 : 3'b000;
										assign node1301 = (inp[6]) ? node1303 : 3'b001;
											assign node1303 = (inp[10]) ? 3'b101 : 3'b001;
								assign node1306 = (inp[10]) ? node1316 : node1307;
									assign node1307 = (inp[6]) ? node1313 : node1308;
										assign node1308 = (inp[1]) ? 3'b000 : node1309;
											assign node1309 = (inp[7]) ? 3'b000 : 3'b001;
										assign node1313 = (inp[9]) ? 3'b101 : 3'b100;
									assign node1316 = (inp[6]) ? node1322 : node1317;
										assign node1317 = (inp[1]) ? 3'b101 : node1318;
											assign node1318 = (inp[9]) ? 3'b100 : 3'b101;
										assign node1322 = (inp[9]) ? node1326 : node1323;
											assign node1323 = (inp[7]) ? 3'b000 : 3'b001;
											assign node1326 = (inp[7]) ? 3'b001 : 3'b000;
							assign node1329 = (inp[1]) ? node1351 : node1330;
								assign node1330 = (inp[11]) ? node1344 : node1331;
									assign node1331 = (inp[9]) ? node1339 : node1332;
										assign node1332 = (inp[7]) ? node1336 : node1333;
											assign node1333 = (inp[10]) ? 3'b100 : 3'b000;
											assign node1336 = (inp[10]) ? 3'b001 : 3'b101;
										assign node1339 = (inp[10]) ? 3'b000 : node1340;
											assign node1340 = (inp[6]) ? 3'b000 : 3'b100;
									assign node1344 = (inp[6]) ? node1348 : node1345;
										assign node1345 = (inp[7]) ? 3'b101 : 3'b100;
										assign node1348 = (inp[7]) ? 3'b100 : 3'b101;
								assign node1351 = (inp[10]) ? node1361 : node1352;
									assign node1352 = (inp[6]) ? node1358 : node1353;
										assign node1353 = (inp[11]) ? node1355 : 3'b000;
											assign node1355 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1358 = (inp[9]) ? 3'b101 : 3'b100;
									assign node1361 = (inp[6]) ? node1369 : node1362;
										assign node1362 = (inp[9]) ? node1366 : node1363;
											assign node1363 = (inp[7]) ? 3'b101 : 3'b100;
											assign node1366 = (inp[7]) ? 3'b100 : 3'b101;
										assign node1369 = (inp[11]) ? 3'b000 : node1370;
											assign node1370 = (inp[7]) ? 3'b000 : 3'b001;
		assign node1374 = (inp[8]) ? node2032 : node1375;
			assign node1375 = (inp[4]) ? node1729 : node1376;
				assign node1376 = (inp[5]) ? node1550 : node1377;
					assign node1377 = (inp[3]) ? node1465 : node1378;
						assign node1378 = (inp[7]) ? node1428 : node1379;
							assign node1379 = (inp[10]) ? node1407 : node1380;
								assign node1380 = (inp[6]) ? node1396 : node1381;
									assign node1381 = (inp[11]) ? node1389 : node1382;
										assign node1382 = (inp[1]) ? node1386 : node1383;
											assign node1383 = (inp[0]) ? 3'b110 : 3'b110;
											assign node1386 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1389 = (inp[0]) ? node1393 : node1390;
											assign node1390 = (inp[9]) ? 3'b010 : 3'b011;
											assign node1393 = (inp[9]) ? 3'b011 : 3'b010;
									assign node1396 = (inp[1]) ? node1402 : node1397;
										assign node1397 = (inp[11]) ? 3'b110 : node1398;
											assign node1398 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1402 = (inp[0]) ? 3'b110 : node1403;
											assign node1403 = (inp[9]) ? 3'b110 : 3'b111;
								assign node1407 = (inp[6]) ? node1419 : node1408;
									assign node1408 = (inp[1]) ? node1414 : node1409;
										assign node1409 = (inp[11]) ? 3'b111 : node1410;
											assign node1410 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1414 = (inp[9]) ? 3'b111 : node1415;
											assign node1415 = (inp[0]) ? 3'b110 : 3'b111;
									assign node1419 = (inp[9]) ? node1423 : node1420;
										assign node1420 = (inp[0]) ? 3'b010 : 3'b011;
										assign node1423 = (inp[11]) ? node1425 : 3'b110;
											assign node1425 = (inp[0]) ? 3'b011 : 3'b010;
							assign node1428 = (inp[6]) ? node1448 : node1429;
								assign node1429 = (inp[10]) ? node1435 : node1430;
									assign node1430 = (inp[9]) ? node1432 : 3'b010;
										assign node1432 = (inp[0]) ? 3'b010 : 3'b111;
									assign node1435 = (inp[11]) ? node1441 : node1436;
										assign node1436 = (inp[1]) ? 3'b111 : node1437;
											assign node1437 = (inp[0]) ? 3'b011 : 3'b010;
										assign node1441 = (inp[1]) ? node1445 : node1442;
											assign node1442 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1445 = (inp[9]) ? 3'b110 : 3'b110;
								assign node1448 = (inp[10]) ? node1458 : node1449;
									assign node1449 = (inp[11]) ? node1453 : node1450;
										assign node1450 = (inp[9]) ? 3'b010 : 3'b111;
										assign node1453 = (inp[0]) ? 3'b111 : node1454;
											assign node1454 = (inp[9]) ? 3'b111 : 3'b110;
									assign node1458 = (inp[11]) ? 3'b011 : node1459;
										assign node1459 = (inp[1]) ? 3'b011 : node1460;
											assign node1460 = (inp[9]) ? 3'b110 : 3'b111;
						assign node1465 = (inp[6]) ? node1501 : node1466;
							assign node1466 = (inp[10]) ? node1486 : node1467;
								assign node1467 = (inp[1]) ? node1479 : node1468;
									assign node1468 = (inp[11]) ? node1474 : node1469;
										assign node1469 = (inp[7]) ? 3'b110 : node1470;
											assign node1470 = (inp[0]) ? 3'b110 : 3'b110;
										assign node1474 = (inp[7]) ? node1476 : 3'b010;
											assign node1476 = (inp[0]) ? 3'b011 : 3'b010;
									assign node1479 = (inp[9]) ? 3'b010 : node1480;
										assign node1480 = (inp[0]) ? node1482 : 3'b011;
											assign node1482 = (inp[11]) ? 3'b010 : 3'b011;
								assign node1486 = (inp[11]) ? node1496 : node1487;
									assign node1487 = (inp[1]) ? node1493 : node1488;
										assign node1488 = (inp[7]) ? 3'b010 : node1489;
											assign node1489 = (inp[9]) ? 3'b010 : 3'b010;
										assign node1493 = (inp[7]) ? 3'b100 : 3'b101;
									assign node1496 = (inp[0]) ? 3'b100 : node1497;
										assign node1497 = (inp[9]) ? 3'b100 : 3'b101;
							assign node1501 = (inp[10]) ? node1527 : node1502;
								assign node1502 = (inp[11]) ? node1514 : node1503;
									assign node1503 = (inp[1]) ? node1509 : node1504;
										assign node1504 = (inp[0]) ? node1506 : 3'b010;
											assign node1506 = (inp[9]) ? 3'b010 : 3'b010;
										assign node1509 = (inp[9]) ? 3'b100 : node1510;
											assign node1510 = (inp[0]) ? 3'b100 : 3'b101;
									assign node1514 = (inp[0]) ? node1522 : node1515;
										assign node1515 = (inp[1]) ? node1519 : node1516;
											assign node1516 = (inp[7]) ? 3'b100 : 3'b100;
											assign node1519 = (inp[9]) ? 3'b101 : 3'b100;
										assign node1522 = (inp[7]) ? node1524 : 3'b100;
											assign node1524 = (inp[1]) ? 3'b100 : 3'b101;
								assign node1527 = (inp[11]) ? node1539 : node1528;
									assign node1528 = (inp[1]) ? node1534 : node1529;
										assign node1529 = (inp[9]) ? node1531 : 3'b100;
											assign node1531 = (inp[0]) ? 3'b100 : 3'b100;
										assign node1534 = (inp[7]) ? 3'b000 : node1535;
											assign node1535 = (inp[9]) ? 3'b000 : 3'b001;
									assign node1539 = (inp[9]) ? node1545 : node1540;
										assign node1540 = (inp[7]) ? node1542 : 3'b001;
											assign node1542 = (inp[0]) ? 3'b001 : 3'b000;
										assign node1545 = (inp[0]) ? 3'b000 : node1546;
											assign node1546 = (inp[7]) ? 3'b001 : 3'b000;
					assign node1550 = (inp[3]) ? node1638 : node1551;
						assign node1551 = (inp[10]) ? node1593 : node1552;
							assign node1552 = (inp[6]) ? node1572 : node1553;
								assign node1553 = (inp[11]) ? node1565 : node1554;
									assign node1554 = (inp[1]) ? node1562 : node1555;
										assign node1555 = (inp[7]) ? node1559 : node1556;
											assign node1556 = (inp[9]) ? 3'b111 : 3'b110;
											assign node1559 = (inp[9]) ? 3'b110 : 3'b111;
										assign node1562 = (inp[0]) ? 3'b010 : 3'b011;
									assign node1565 = (inp[0]) ? 3'b011 : node1566;
										assign node1566 = (inp[7]) ? node1568 : 3'b010;
											assign node1568 = (inp[9]) ? 3'b011 : 3'b010;
								assign node1572 = (inp[1]) ? node1584 : node1573;
									assign node1573 = (inp[11]) ? node1579 : node1574;
										assign node1574 = (inp[7]) ? node1576 : 3'b011;
											assign node1576 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1579 = (inp[0]) ? node1581 : 3'b100;
											assign node1581 = (inp[9]) ? 3'b101 : 3'b100;
									assign node1584 = (inp[0]) ? node1588 : node1585;
										assign node1585 = (inp[7]) ? 3'b100 : 3'b101;
										assign node1588 = (inp[11]) ? node1590 : 3'b100;
											assign node1590 = (inp[9]) ? 3'b100 : 3'b100;
							assign node1593 = (inp[6]) ? node1615 : node1594;
								assign node1594 = (inp[1]) ? node1606 : node1595;
									assign node1595 = (inp[11]) ? node1601 : node1596;
										assign node1596 = (inp[7]) ? 3'b011 : node1597;
											assign node1597 = (inp[0]) ? 3'b010 : 3'b010;
										assign node1601 = (inp[9]) ? 3'b101 : node1602;
											assign node1602 = (inp[0]) ? 3'b100 : 3'b100;
									assign node1606 = (inp[7]) ? 3'b100 : node1607;
										assign node1607 = (inp[9]) ? node1611 : node1608;
											assign node1608 = (inp[0]) ? 3'b100 : 3'b101;
											assign node1611 = (inp[0]) ? 3'b101 : 3'b100;
								assign node1615 = (inp[11]) ? node1625 : node1616;
									assign node1616 = (inp[1]) ? node1620 : node1617;
										assign node1617 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1620 = (inp[0]) ? node1622 : 3'b001;
											assign node1622 = (inp[9]) ? 3'b000 : 3'b000;
									assign node1625 = (inp[9]) ? node1631 : node1626;
										assign node1626 = (inp[7]) ? 3'b000 : node1627;
											assign node1627 = (inp[0]) ? 3'b000 : 3'b001;
										assign node1631 = (inp[7]) ? node1635 : node1632;
											assign node1632 = (inp[0]) ? 3'b001 : 3'b000;
											assign node1635 = (inp[1]) ? 3'b000 : 3'b001;
						assign node1638 = (inp[0]) ? node1682 : node1639;
							assign node1639 = (inp[11]) ? node1661 : node1640;
								assign node1640 = (inp[6]) ? node1648 : node1641;
									assign node1641 = (inp[1]) ? node1645 : node1642;
										assign node1642 = (inp[10]) ? 3'b000 : 3'b100;
										assign node1645 = (inp[10]) ? 3'b100 : 3'b000;
									assign node1648 = (inp[7]) ? node1656 : node1649;
										assign node1649 = (inp[9]) ? node1653 : node1650;
											assign node1650 = (inp[10]) ? 3'b001 : 3'b001;
											assign node1653 = (inp[10]) ? 3'b000 : 3'b100;
										assign node1656 = (inp[9]) ? node1658 : 3'b100;
											assign node1658 = (inp[10]) ? 3'b101 : 3'b001;
								assign node1661 = (inp[6]) ? node1671 : node1662;
									assign node1662 = (inp[10]) ? node1664 : 3'b001;
										assign node1664 = (inp[1]) ? node1668 : node1665;
											assign node1665 = (inp[7]) ? 3'b100 : 3'b101;
											assign node1668 = (inp[9]) ? 3'b100 : 3'b101;
									assign node1671 = (inp[10]) ? node1677 : node1672;
										assign node1672 = (inp[7]) ? node1674 : 3'b101;
											assign node1674 = (inp[1]) ? 3'b100 : 3'b101;
										assign node1677 = (inp[7]) ? 3'b000 : node1678;
											assign node1678 = (inp[9]) ? 3'b000 : 3'b001;
							assign node1682 = (inp[1]) ? node1702 : node1683;
								assign node1683 = (inp[9]) ? node1695 : node1684;
									assign node1684 = (inp[7]) ? node1690 : node1685;
										assign node1685 = (inp[11]) ? node1687 : 3'b000;
											assign node1687 = (inp[10]) ? 3'b000 : 3'b100;
										assign node1690 = (inp[10]) ? node1692 : 3'b001;
											assign node1692 = (inp[11]) ? 3'b101 : 3'b001;
									assign node1695 = (inp[7]) ? 3'b000 : node1696;
										assign node1696 = (inp[11]) ? 3'b001 : node1697;
											assign node1697 = (inp[10]) ? 3'b001 : 3'b101;
								assign node1702 = (inp[7]) ? node1718 : node1703;
									assign node1703 = (inp[9]) ? node1711 : node1704;
										assign node1704 = (inp[6]) ? node1708 : node1705;
											assign node1705 = (inp[10]) ? 3'b100 : 3'b000;
											assign node1708 = (inp[10]) ? 3'b000 : 3'b100;
										assign node1711 = (inp[10]) ? node1715 : node1712;
											assign node1712 = (inp[6]) ? 3'b101 : 3'b001;
											assign node1715 = (inp[6]) ? 3'b001 : 3'b101;
									assign node1718 = (inp[9]) ? node1724 : node1719;
										assign node1719 = (inp[10]) ? node1721 : 3'b101;
											assign node1721 = (inp[6]) ? 3'b001 : 3'b101;
										assign node1724 = (inp[11]) ? 3'b100 : node1725;
											assign node1725 = (inp[6]) ? 3'b000 : 3'b100;
				assign node1729 = (inp[3]) ? node1887 : node1730;
					assign node1730 = (inp[5]) ? node1816 : node1731;
						assign node1731 = (inp[10]) ? node1777 : node1732;
							assign node1732 = (inp[6]) ? node1758 : node1733;
								assign node1733 = (inp[11]) ? node1747 : node1734;
									assign node1734 = (inp[1]) ? node1740 : node1735;
										assign node1735 = (inp[7]) ? 3'b101 : node1736;
											assign node1736 = (inp[9]) ? 3'b100 : 3'b100;
										assign node1740 = (inp[9]) ? node1744 : node1741;
											assign node1741 = (inp[7]) ? 3'b001 : 3'b000;
											assign node1744 = (inp[7]) ? 3'b000 : 3'b001;
									assign node1747 = (inp[9]) ? node1753 : node1748;
										assign node1748 = (inp[7]) ? node1750 : 3'b001;
											assign node1750 = (inp[0]) ? 3'b001 : 3'b000;
										assign node1753 = (inp[7]) ? 3'b000 : node1754;
											assign node1754 = (inp[0]) ? 3'b001 : 3'b000;
								assign node1758 = (inp[1]) ? node1764 : node1759;
									assign node1759 = (inp[11]) ? node1761 : 3'b001;
										assign node1761 = (inp[7]) ? 3'b100 : 3'b101;
									assign node1764 = (inp[11]) ? node1772 : node1765;
										assign node1765 = (inp[7]) ? node1769 : node1766;
											assign node1766 = (inp[0]) ? 3'b100 : 3'b101;
											assign node1769 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1772 = (inp[0]) ? 3'b101 : node1773;
											assign node1773 = (inp[9]) ? 3'b100 : 3'b101;
							assign node1777 = (inp[6]) ? node1795 : node1778;
								assign node1778 = (inp[9]) ? node1788 : node1779;
									assign node1779 = (inp[11]) ? node1781 : 3'b100;
										assign node1781 = (inp[7]) ? node1785 : node1782;
											assign node1782 = (inp[0]) ? 3'b100 : 3'b101;
											assign node1785 = (inp[0]) ? 3'b101 : 3'b100;
									assign node1788 = (inp[1]) ? node1792 : node1789;
										assign node1789 = (inp[11]) ? 3'b100 : 3'b000;
										assign node1792 = (inp[0]) ? 3'b100 : 3'b101;
								assign node1795 = (inp[1]) ? node1805 : node1796;
									assign node1796 = (inp[11]) ? node1802 : node1797;
										assign node1797 = (inp[7]) ? node1799 : 3'b100;
											assign node1799 = (inp[9]) ? 3'b100 : 3'b100;
										assign node1802 = (inp[9]) ? 3'b001 : 3'b000;
									assign node1805 = (inp[0]) ? node1811 : node1806;
										assign node1806 = (inp[7]) ? 3'b000 : node1807;
											assign node1807 = (inp[9]) ? 3'b000 : 3'b001;
										assign node1811 = (inp[11]) ? 3'b001 : node1812;
											assign node1812 = (inp[7]) ? 3'b000 : 3'b000;
						assign node1816 = (inp[10]) ? node1860 : node1817;
							assign node1817 = (inp[6]) ? node1839 : node1818;
								assign node1818 = (inp[1]) ? node1828 : node1819;
									assign node1819 = (inp[11]) ? node1823 : node1820;
										assign node1820 = (inp[7]) ? 3'b101 : 3'b100;
										assign node1823 = (inp[7]) ? 3'b000 : node1824;
											assign node1824 = (inp[9]) ? 3'b001 : 3'b000;
									assign node1828 = (inp[0]) ? node1834 : node1829;
										assign node1829 = (inp[11]) ? 3'b001 : node1830;
											assign node1830 = (inp[7]) ? 3'b000 : 3'b000;
										assign node1834 = (inp[11]) ? 3'b000 : node1835;
											assign node1835 = (inp[7]) ? 3'b000 : 3'b001;
								assign node1839 = (inp[11]) ? node1853 : node1840;
									assign node1840 = (inp[1]) ? node1848 : node1841;
										assign node1841 = (inp[0]) ? node1845 : node1842;
											assign node1842 = (inp[7]) ? 3'b000 : 3'b000;
											assign node1845 = (inp[7]) ? 3'b000 : 3'b001;
										assign node1848 = (inp[9]) ? 3'b111 : node1849;
											assign node1849 = (inp[0]) ? 3'b111 : 3'b110;
									assign node1853 = (inp[7]) ? node1857 : node1854;
										assign node1854 = (inp[9]) ? 3'b111 : 3'b110;
										assign node1857 = (inp[9]) ? 3'b110 : 3'b111;
							assign node1860 = (inp[6]) ? node1872 : node1861;
								assign node1861 = (inp[9]) ? node1869 : node1862;
									assign node1862 = (inp[7]) ? node1864 : 3'b110;
										assign node1864 = (inp[1]) ? 3'b111 : node1865;
											assign node1865 = (inp[11]) ? 3'b111 : 3'b001;
									assign node1869 = (inp[7]) ? 3'b110 : 3'b111;
								assign node1872 = (inp[1]) ? node1880 : node1873;
									assign node1873 = (inp[11]) ? 3'b011 : node1874;
										assign node1874 = (inp[7]) ? 3'b110 : node1875;
											assign node1875 = (inp[9]) ? 3'b111 : 3'b110;
									assign node1880 = (inp[7]) ? node1884 : node1881;
										assign node1881 = (inp[9]) ? 3'b011 : 3'b010;
										assign node1884 = (inp[9]) ? 3'b010 : 3'b011;
					assign node1887 = (inp[5]) ? node1973 : node1888;
						assign node1888 = (inp[10]) ? node1936 : node1889;
							assign node1889 = (inp[6]) ? node1913 : node1890;
								assign node1890 = (inp[11]) ? node1902 : node1891;
									assign node1891 = (inp[1]) ? node1897 : node1892;
										assign node1892 = (inp[7]) ? 3'b100 : node1893;
											assign node1893 = (inp[0]) ? 3'b101 : 3'b100;
										assign node1897 = (inp[0]) ? 3'b000 : node1898;
											assign node1898 = (inp[9]) ? 3'b000 : 3'b000;
									assign node1902 = (inp[0]) ? node1908 : node1903;
										assign node1903 = (inp[7]) ? node1905 : 3'b001;
											assign node1905 = (inp[9]) ? 3'b001 : 3'b000;
										assign node1908 = (inp[1]) ? node1910 : 3'b000;
											assign node1910 = (inp[9]) ? 3'b001 : 3'b000;
								assign node1913 = (inp[11]) ? node1925 : node1914;
									assign node1914 = (inp[1]) ? node1920 : node1915;
										assign node1915 = (inp[7]) ? node1917 : 3'b000;
											assign node1917 = (inp[9]) ? 3'b001 : 3'b000;
										assign node1920 = (inp[0]) ? 3'b110 : node1921;
											assign node1921 = (inp[9]) ? 3'b111 : 3'b110;
									assign node1925 = (inp[0]) ? node1931 : node1926;
										assign node1926 = (inp[1]) ? 3'b111 : node1927;
											assign node1927 = (inp[7]) ? 3'b111 : 3'b110;
										assign node1931 = (inp[1]) ? 3'b110 : node1932;
											assign node1932 = (inp[9]) ? 3'b110 : 3'b110;
							assign node1936 = (inp[6]) ? node1954 : node1937;
								assign node1937 = (inp[1]) ? node1947 : node1938;
									assign node1938 = (inp[11]) ? node1942 : node1939;
										assign node1939 = (inp[7]) ? 3'b001 : 3'b000;
										assign node1942 = (inp[7]) ? 3'b111 : node1943;
											assign node1943 = (inp[9]) ? 3'b111 : 3'b110;
									assign node1947 = (inp[9]) ? node1951 : node1948;
										assign node1948 = (inp[7]) ? 3'b111 : 3'b110;
										assign node1951 = (inp[7]) ? 3'b110 : 3'b111;
								assign node1954 = (inp[1]) ? node1966 : node1955;
									assign node1955 = (inp[11]) ? node1961 : node1956;
										assign node1956 = (inp[7]) ? node1958 : 3'b111;
											assign node1958 = (inp[9]) ? 3'b110 : 3'b111;
										assign node1961 = (inp[0]) ? 3'b010 : node1962;
											assign node1962 = (inp[7]) ? 3'b010 : 3'b011;
									assign node1966 = (inp[9]) ? node1970 : node1967;
										assign node1967 = (inp[7]) ? 3'b011 : 3'b010;
										assign node1970 = (inp[7]) ? 3'b010 : 3'b011;
						assign node1973 = (inp[7]) ? node2011 : node1974;
							assign node1974 = (inp[9]) ? node1994 : node1975;
								assign node1975 = (inp[1]) ? node1987 : node1976;
									assign node1976 = (inp[0]) ? node1982 : node1977;
										assign node1977 = (inp[10]) ? node1979 : 3'b110;
											assign node1979 = (inp[6]) ? 3'b010 : 3'b110;
										assign node1982 = (inp[6]) ? 3'b110 : node1983;
											assign node1983 = (inp[10]) ? 3'b010 : 3'b010;
									assign node1987 = (inp[10]) ? node1991 : node1988;
										assign node1988 = (inp[6]) ? 3'b110 : 3'b010;
										assign node1991 = (inp[6]) ? 3'b010 : 3'b110;
								assign node1994 = (inp[10]) ? node2000 : node1995;
									assign node1995 = (inp[6]) ? 3'b111 : node1996;
										assign node1996 = (inp[11]) ? 3'b011 : 3'b111;
									assign node2000 = (inp[6]) ? node2006 : node2001;
										assign node2001 = (inp[11]) ? 3'b111 : node2002;
											assign node2002 = (inp[1]) ? 3'b111 : 3'b011;
										assign node2006 = (inp[1]) ? 3'b011 : node2007;
											assign node2007 = (inp[11]) ? 3'b011 : 3'b111;
							assign node2011 = (inp[9]) ? node2019 : node2012;
								assign node2012 = (inp[6]) ? 3'b011 : node2013;
									assign node2013 = (inp[10]) ? 3'b111 : node2014;
										assign node2014 = (inp[11]) ? 3'b011 : 3'b111;
								assign node2019 = (inp[6]) ? node2029 : node2020;
									assign node2020 = (inp[10]) ? node2026 : node2021;
										assign node2021 = (inp[11]) ? 3'b010 : node2022;
											assign node2022 = (inp[1]) ? 3'b010 : 3'b110;
										assign node2026 = (inp[1]) ? 3'b110 : 3'b010;
									assign node2029 = (inp[10]) ? 3'b010 : 3'b110;
			assign node2032 = (inp[4]) ? node2372 : node2033;
				assign node2033 = (inp[3]) ? node2205 : node2034;
					assign node2034 = (inp[5]) ? node2120 : node2035;
						assign node2035 = (inp[10]) ? node2077 : node2036;
							assign node2036 = (inp[6]) ? node2050 : node2037;
								assign node2037 = (inp[1]) ? node2043 : node2038;
									assign node2038 = (inp[11]) ? 3'b000 : node2039;
										assign node2039 = (inp[9]) ? 3'b100 : 3'b101;
									assign node2043 = (inp[0]) ? 3'b001 : node2044;
										assign node2044 = (inp[7]) ? node2046 : 3'b000;
											assign node2046 = (inp[9]) ? 3'b001 : 3'b000;
								assign node2050 = (inp[1]) ? node2062 : node2051;
									assign node2051 = (inp[11]) ? node2057 : node2052;
										assign node2052 = (inp[7]) ? 3'b000 : node2053;
											assign node2053 = (inp[9]) ? 3'b000 : 3'b001;
										assign node2057 = (inp[7]) ? 3'b100 : node2058;
											assign node2058 = (inp[9]) ? 3'b100 : 3'b100;
									assign node2062 = (inp[9]) ? node2070 : node2063;
										assign node2063 = (inp[0]) ? node2067 : node2064;
											assign node2064 = (inp[7]) ? 3'b100 : 3'b101;
											assign node2067 = (inp[7]) ? 3'b101 : 3'b100;
										assign node2070 = (inp[11]) ? node2074 : node2071;
											assign node2071 = (inp[0]) ? 3'b100 : 3'b100;
											assign node2074 = (inp[0]) ? 3'b100 : 3'b100;
							assign node2077 = (inp[6]) ? node2103 : node2078;
								assign node2078 = (inp[11]) ? node2092 : node2079;
									assign node2079 = (inp[1]) ? node2085 : node2080;
										assign node2080 = (inp[0]) ? 3'b001 : node2081;
											assign node2081 = (inp[9]) ? 3'b000 : 3'b001;
										assign node2085 = (inp[9]) ? node2089 : node2086;
											assign node2086 = (inp[7]) ? 3'b100 : 3'b101;
											assign node2089 = (inp[7]) ? 3'b101 : 3'b100;
									assign node2092 = (inp[7]) ? node2098 : node2093;
										assign node2093 = (inp[1]) ? node2095 : 3'b100;
											assign node2095 = (inp[0]) ? 3'b100 : 3'b100;
										assign node2098 = (inp[9]) ? 3'b101 : node2099;
											assign node2099 = (inp[0]) ? 3'b101 : 3'b100;
								assign node2103 = (inp[11]) ? node2111 : node2104;
									assign node2104 = (inp[1]) ? 3'b001 : node2105;
										assign node2105 = (inp[9]) ? node2107 : 3'b101;
											assign node2107 = (inp[7]) ? 3'b101 : 3'b100;
									assign node2111 = (inp[1]) ? node2117 : node2112;
										assign node2112 = (inp[9]) ? 3'b000 : node2113;
											assign node2113 = (inp[7]) ? 3'b001 : 3'b000;
										assign node2117 = (inp[9]) ? 3'b001 : 3'b000;
						assign node2120 = (inp[6]) ? node2166 : node2121;
							assign node2121 = (inp[10]) ? node2141 : node2122;
								assign node2122 = (inp[11]) ? node2134 : node2123;
									assign node2123 = (inp[1]) ? node2131 : node2124;
										assign node2124 = (inp[0]) ? node2128 : node2125;
											assign node2125 = (inp[7]) ? 3'b100 : 3'b100;
											assign node2128 = (inp[9]) ? 3'b100 : 3'b100;
										assign node2131 = (inp[0]) ? 3'b000 : 3'b001;
									assign node2134 = (inp[0]) ? node2136 : 3'b001;
										assign node2136 = (inp[7]) ? node2138 : 3'b001;
											assign node2138 = (inp[9]) ? 3'b000 : 3'b001;
								assign node2141 = (inp[1]) ? node2153 : node2142;
									assign node2142 = (inp[11]) ? node2148 : node2143;
										assign node2143 = (inp[9]) ? 3'b001 : node2144;
											assign node2144 = (inp[0]) ? 3'b001 : 3'b000;
										assign node2148 = (inp[0]) ? node2150 : 3'b111;
											assign node2150 = (inp[7]) ? 3'b110 : 3'b110;
									assign node2153 = (inp[11]) ? node2161 : node2154;
										assign node2154 = (inp[0]) ? node2158 : node2155;
											assign node2155 = (inp[9]) ? 3'b110 : 3'b111;
											assign node2158 = (inp[9]) ? 3'b111 : 3'b110;
										assign node2161 = (inp[7]) ? 3'b110 : node2162;
											assign node2162 = (inp[9]) ? 3'b111 : 3'b110;
							assign node2166 = (inp[10]) ? node2186 : node2167;
								assign node2167 = (inp[11]) ? node2179 : node2168;
									assign node2168 = (inp[1]) ? node2174 : node2169;
										assign node2169 = (inp[9]) ? node2171 : 3'b000;
											assign node2171 = (inp[0]) ? 3'b000 : 3'b001;
										assign node2174 = (inp[0]) ? 3'b110 : node2175;
											assign node2175 = (inp[7]) ? 3'b111 : 3'b110;
									assign node2179 = (inp[9]) ? node2183 : node2180;
										assign node2180 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2183 = (inp[7]) ? 3'b110 : 3'b111;
								assign node2186 = (inp[11]) ? node2198 : node2187;
									assign node2187 = (inp[1]) ? node2193 : node2188;
										assign node2188 = (inp[0]) ? node2190 : 3'b110;
											assign node2190 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2193 = (inp[9]) ? node2195 : 3'b010;
											assign node2195 = (inp[7]) ? 3'b010 : 3'b011;
									assign node2198 = (inp[9]) ? node2202 : node2199;
										assign node2199 = (inp[7]) ? 3'b011 : 3'b010;
										assign node2202 = (inp[7]) ? 3'b010 : 3'b011;
					assign node2205 = (inp[5]) ? node2289 : node2206;
						assign node2206 = (inp[10]) ? node2254 : node2207;
							assign node2207 = (inp[6]) ? node2229 : node2208;
								assign node2208 = (inp[11]) ? node2220 : node2209;
									assign node2209 = (inp[1]) ? node2215 : node2210;
										assign node2210 = (inp[7]) ? 3'b101 : node2211;
											assign node2211 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2215 = (inp[0]) ? 3'b001 : node2216;
											assign node2216 = (inp[7]) ? 3'b000 : 3'b000;
									assign node2220 = (inp[7]) ? 3'b001 : node2221;
										assign node2221 = (inp[9]) ? node2225 : node2222;
											assign node2222 = (inp[0]) ? 3'b000 : 3'b001;
											assign node2225 = (inp[1]) ? 3'b000 : 3'b001;
								assign node2229 = (inp[1]) ? node2241 : node2230;
									assign node2230 = (inp[11]) ? node2236 : node2231;
										assign node2231 = (inp[9]) ? node2233 : 3'b001;
											assign node2233 = (inp[0]) ? 3'b001 : 3'b000;
										assign node2236 = (inp[0]) ? 3'b110 : node2237;
											assign node2237 = (inp[9]) ? 3'b111 : 3'b110;
									assign node2241 = (inp[11]) ? node2249 : node2242;
										assign node2242 = (inp[7]) ? node2246 : node2243;
											assign node2243 = (inp[9]) ? 3'b111 : 3'b110;
											assign node2246 = (inp[9]) ? 3'b110 : 3'b111;
										assign node2249 = (inp[9]) ? node2251 : 3'b110;
											assign node2251 = (inp[0]) ? 3'b110 : 3'b111;
							assign node2254 = (inp[6]) ? node2272 : node2255;
								assign node2255 = (inp[11]) ? node2265 : node2256;
									assign node2256 = (inp[1]) ? node2258 : 3'b001;
										assign node2258 = (inp[9]) ? node2262 : node2259;
											assign node2259 = (inp[7]) ? 3'b111 : 3'b110;
											assign node2262 = (inp[7]) ? 3'b110 : 3'b111;
									assign node2265 = (inp[7]) ? node2269 : node2266;
										assign node2266 = (inp[9]) ? 3'b111 : 3'b110;
										assign node2269 = (inp[9]) ? 3'b110 : 3'b111;
								assign node2272 = (inp[11]) ? node2282 : node2273;
									assign node2273 = (inp[1]) ? node2277 : node2274;
										assign node2274 = (inp[0]) ? 3'b110 : 3'b111;
										assign node2277 = (inp[7]) ? node2279 : 3'b010;
											assign node2279 = (inp[9]) ? 3'b010 : 3'b011;
									assign node2282 = (inp[9]) ? node2286 : node2283;
										assign node2283 = (inp[7]) ? 3'b011 : 3'b010;
										assign node2286 = (inp[7]) ? 3'b010 : 3'b011;
						assign node2289 = (inp[10]) ? node2329 : node2290;
							assign node2290 = (inp[6]) ? node2314 : node2291;
								assign node2291 = (inp[1]) ? node2303 : node2292;
									assign node2292 = (inp[11]) ? node2298 : node2293;
										assign node2293 = (inp[9]) ? node2295 : 3'b110;
											assign node2295 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2298 = (inp[7]) ? 3'b011 : node2299;
											assign node2299 = (inp[9]) ? 3'b011 : 3'b010;
									assign node2303 = (inp[0]) ? node2309 : node2304;
										assign node2304 = (inp[9]) ? 3'b010 : node2305;
											assign node2305 = (inp[7]) ? 3'b011 : 3'b010;
										assign node2309 = (inp[7]) ? node2311 : 3'b011;
											assign node2311 = (inp[9]) ? 3'b010 : 3'b011;
								assign node2314 = (inp[11]) ? node2322 : node2315;
									assign node2315 = (inp[1]) ? 3'b111 : node2316;
										assign node2316 = (inp[9]) ? 3'b010 : node2317;
											assign node2317 = (inp[7]) ? 3'b011 : 3'b010;
									assign node2322 = (inp[9]) ? node2326 : node2323;
										assign node2323 = (inp[7]) ? 3'b111 : 3'b110;
										assign node2326 = (inp[7]) ? 3'b110 : 3'b111;
							assign node2329 = (inp[6]) ? node2353 : node2330;
								assign node2330 = (inp[1]) ? node2342 : node2331;
									assign node2331 = (inp[11]) ? node2339 : node2332;
										assign node2332 = (inp[0]) ? node2336 : node2333;
											assign node2333 = (inp[7]) ? 3'b010 : 3'b011;
											assign node2336 = (inp[7]) ? 3'b010 : 3'b010;
										assign node2339 = (inp[9]) ? 3'b111 : 3'b110;
									assign node2342 = (inp[0]) ? node2348 : node2343;
										assign node2343 = (inp[9]) ? node2345 : 3'b111;
											assign node2345 = (inp[11]) ? 3'b111 : 3'b110;
										assign node2348 = (inp[9]) ? 3'b111 : node2349;
											assign node2349 = (inp[7]) ? 3'b111 : 3'b110;
								assign node2353 = (inp[1]) ? node2365 : node2354;
									assign node2354 = (inp[11]) ? node2360 : node2355;
										assign node2355 = (inp[0]) ? node2357 : 3'b110;
											assign node2357 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2360 = (inp[9]) ? node2362 : 3'b011;
											assign node2362 = (inp[7]) ? 3'b010 : 3'b011;
									assign node2365 = (inp[9]) ? node2369 : node2366;
										assign node2366 = (inp[7]) ? 3'b011 : 3'b010;
										assign node2369 = (inp[7]) ? 3'b010 : 3'b011;
				assign node2372 = (inp[3]) ? node2550 : node2373;
					assign node2373 = (inp[5]) ? node2461 : node2374;
						assign node2374 = (inp[11]) ? node2426 : node2375;
							assign node2375 = (inp[0]) ? node2401 : node2376;
								assign node2376 = (inp[6]) ? node2390 : node2377;
									assign node2377 = (inp[10]) ? node2383 : node2378;
										assign node2378 = (inp[7]) ? node2380 : 3'b110;
											assign node2380 = (inp[9]) ? 3'b110 : 3'b111;
										assign node2383 = (inp[7]) ? node2387 : node2384;
											assign node2384 = (inp[9]) ? 3'b111 : 3'b110;
											assign node2387 = (inp[9]) ? 3'b110 : 3'b111;
									assign node2390 = (inp[1]) ? node2398 : node2391;
										assign node2391 = (inp[10]) ? node2395 : node2392;
											assign node2392 = (inp[9]) ? 3'b010 : 3'b010;
											assign node2395 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2398 = (inp[10]) ? 3'b010 : 3'b110;
								assign node2401 = (inp[6]) ? node2415 : node2402;
									assign node2402 = (inp[7]) ? node2408 : node2403;
										assign node2403 = (inp[10]) ? 3'b011 : node2404;
											assign node2404 = (inp[1]) ? 3'b011 : 3'b111;
										assign node2408 = (inp[9]) ? node2412 : node2409;
											assign node2409 = (inp[10]) ? 3'b111 : 3'b011;
											assign node2412 = (inp[1]) ? 3'b010 : 3'b110;
									assign node2415 = (inp[1]) ? node2421 : node2416;
										assign node2416 = (inp[9]) ? node2418 : 3'b110;
											assign node2418 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2421 = (inp[10]) ? 3'b011 : node2422;
											assign node2422 = (inp[7]) ? 3'b111 : 3'b110;
							assign node2426 = (inp[6]) ? node2442 : node2427;
								assign node2427 = (inp[10]) ? node2435 : node2428;
									assign node2428 = (inp[7]) ? node2432 : node2429;
										assign node2429 = (inp[9]) ? 3'b011 : 3'b010;
										assign node2432 = (inp[9]) ? 3'b010 : 3'b011;
									assign node2435 = (inp[1]) ? 3'b111 : node2436;
										assign node2436 = (inp[9]) ? 3'b110 : node2437;
											assign node2437 = (inp[7]) ? 3'b111 : 3'b110;
								assign node2442 = (inp[10]) ? node2452 : node2443;
									assign node2443 = (inp[0]) ? 3'b110 : node2444;
										assign node2444 = (inp[9]) ? node2448 : node2445;
											assign node2445 = (inp[7]) ? 3'b111 : 3'b110;
											assign node2448 = (inp[7]) ? 3'b110 : 3'b111;
									assign node2452 = (inp[0]) ? 3'b010 : node2453;
										assign node2453 = (inp[1]) ? node2457 : node2454;
											assign node2454 = (inp[7]) ? 3'b011 : 3'b010;
											assign node2457 = (inp[9]) ? 3'b010 : 3'b011;
						assign node2461 = (inp[10]) ? node2505 : node2462;
							assign node2462 = (inp[6]) ? node2486 : node2463;
								assign node2463 = (inp[11]) ? node2475 : node2464;
									assign node2464 = (inp[1]) ? node2472 : node2465;
										assign node2465 = (inp[9]) ? node2469 : node2466;
											assign node2466 = (inp[7]) ? 3'b111 : 3'b110;
											assign node2469 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2472 = (inp[0]) ? 3'b010 : 3'b011;
									assign node2475 = (inp[1]) ? node2481 : node2476;
										assign node2476 = (inp[9]) ? 3'b010 : node2477;
											assign node2477 = (inp[7]) ? 3'b011 : 3'b010;
										assign node2481 = (inp[0]) ? node2483 : 3'b011;
											assign node2483 = (inp[9]) ? 3'b010 : 3'b010;
								assign node2486 = (inp[11]) ? node2498 : node2487;
									assign node2487 = (inp[1]) ? node2493 : node2488;
										assign node2488 = (inp[9]) ? node2490 : 3'b010;
											assign node2490 = (inp[7]) ? 3'b010 : 3'b011;
										assign node2493 = (inp[0]) ? 3'b101 : node2494;
											assign node2494 = (inp[9]) ? 3'b100 : 3'b100;
									assign node2498 = (inp[9]) ? node2502 : node2499;
										assign node2499 = (inp[7]) ? 3'b101 : 3'b100;
										assign node2502 = (inp[7]) ? 3'b100 : 3'b101;
							assign node2505 = (inp[6]) ? node2523 : node2506;
								assign node2506 = (inp[11]) ? node2516 : node2507;
									assign node2507 = (inp[1]) ? node2511 : node2508;
										assign node2508 = (inp[0]) ? 3'b010 : 3'b011;
										assign node2511 = (inp[9]) ? 3'b101 : node2512;
											assign node2512 = (inp[7]) ? 3'b101 : 3'b100;
									assign node2516 = (inp[7]) ? node2520 : node2517;
										assign node2517 = (inp[0]) ? 3'b100 : 3'b101;
										assign node2520 = (inp[9]) ? 3'b100 : 3'b101;
								assign node2523 = (inp[1]) ? node2537 : node2524;
									assign node2524 = (inp[11]) ? node2530 : node2525;
										assign node2525 = (inp[7]) ? 3'b101 : node2526;
											assign node2526 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2530 = (inp[9]) ? node2534 : node2531;
											assign node2531 = (inp[7]) ? 3'b001 : 3'b000;
											assign node2534 = (inp[7]) ? 3'b000 : 3'b001;
									assign node2537 = (inp[0]) ? node2545 : node2538;
										assign node2538 = (inp[11]) ? node2542 : node2539;
											assign node2539 = (inp[9]) ? 3'b001 : 3'b000;
											assign node2542 = (inp[9]) ? 3'b000 : 3'b001;
										assign node2545 = (inp[7]) ? node2547 : 3'b000;
											assign node2547 = (inp[9]) ? 3'b000 : 3'b001;
					assign node2550 = (inp[5]) ? node2630 : node2551;
						assign node2551 = (inp[6]) ? node2593 : node2552;
							assign node2552 = (inp[10]) ? node2572 : node2553;
								assign node2553 = (inp[1]) ? node2565 : node2554;
									assign node2554 = (inp[11]) ? node2562 : node2555;
										assign node2555 = (inp[0]) ? node2559 : node2556;
											assign node2556 = (inp[7]) ? 3'b111 : 3'b110;
											assign node2559 = (inp[7]) ? 3'b110 : 3'b111;
										assign node2562 = (inp[9]) ? 3'b010 : 3'b011;
									assign node2565 = (inp[9]) ? node2569 : node2566;
										assign node2566 = (inp[7]) ? 3'b011 : 3'b010;
										assign node2569 = (inp[7]) ? 3'b010 : 3'b011;
								assign node2572 = (inp[1]) ? node2582 : node2573;
									assign node2573 = (inp[11]) ? node2579 : node2574;
										assign node2574 = (inp[7]) ? node2576 : 3'b011;
											assign node2576 = (inp[9]) ? 3'b010 : 3'b011;
										assign node2579 = (inp[9]) ? 3'b100 : 3'b101;
									assign node2582 = (inp[0]) ? node2588 : node2583;
										assign node2583 = (inp[11]) ? 3'b100 : node2584;
											assign node2584 = (inp[9]) ? 3'b100 : 3'b101;
										assign node2588 = (inp[11]) ? node2590 : 3'b101;
											assign node2590 = (inp[7]) ? 3'b100 : 3'b100;
							assign node2593 = (inp[10]) ? node2617 : node2594;
								assign node2594 = (inp[1]) ? node2604 : node2595;
									assign node2595 = (inp[11]) ? node2597 : 3'b011;
										assign node2597 = (inp[0]) ? node2601 : node2598;
											assign node2598 = (inp[7]) ? 3'b101 : 3'b100;
											assign node2601 = (inp[7]) ? 3'b100 : 3'b101;
									assign node2604 = (inp[11]) ? node2612 : node2605;
										assign node2605 = (inp[0]) ? node2609 : node2606;
											assign node2606 = (inp[7]) ? 3'b100 : 3'b100;
											assign node2609 = (inp[9]) ? 3'b100 : 3'b100;
										assign node2612 = (inp[9]) ? 3'b100 : node2613;
											assign node2613 = (inp[7]) ? 3'b101 : 3'b100;
								assign node2617 = (inp[11]) ? node2623 : node2618;
									assign node2618 = (inp[1]) ? 3'b001 : node2619;
										assign node2619 = (inp[9]) ? 3'b100 : 3'b101;
									assign node2623 = (inp[1]) ? node2625 : 3'b001;
										assign node2625 = (inp[9]) ? 3'b000 : node2626;
											assign node2626 = (inp[7]) ? 3'b001 : 3'b000;
						assign node2630 = (inp[10]) ? node2674 : node2631;
							assign node2631 = (inp[6]) ? node2655 : node2632;
								assign node2632 = (inp[1]) ? node2644 : node2633;
									assign node2633 = (inp[11]) ? node2639 : node2634;
										assign node2634 = (inp[7]) ? node2636 : 3'b100;
											assign node2636 = (inp[9]) ? 3'b100 : 3'b101;
										assign node2639 = (inp[9]) ? node2641 : 3'b001;
											assign node2641 = (inp[7]) ? 3'b000 : 3'b001;
									assign node2644 = (inp[0]) ? node2650 : node2645;
										assign node2645 = (inp[7]) ? 3'b000 : node2646;
											assign node2646 = (inp[9]) ? 3'b001 : 3'b000;
										assign node2650 = (inp[11]) ? node2652 : 3'b001;
											assign node2652 = (inp[7]) ? 3'b000 : 3'b001;
								assign node2655 = (inp[11]) ? node2667 : node2656;
									assign node2656 = (inp[1]) ? node2662 : node2657;
										assign node2657 = (inp[0]) ? 3'b000 : node2658;
											assign node2658 = (inp[7]) ? 3'b000 : 3'b001;
										assign node2662 = (inp[7]) ? node2664 : 3'b100;
											assign node2664 = (inp[9]) ? 3'b100 : 3'b101;
									assign node2667 = (inp[7]) ? node2671 : node2668;
										assign node2668 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2671 = (inp[9]) ? 3'b100 : 3'b101;
							assign node2674 = (inp[6]) ? node2694 : node2675;
								assign node2675 = (inp[11]) ? node2687 : node2676;
									assign node2676 = (inp[1]) ? node2682 : node2677;
										assign node2677 = (inp[7]) ? node2679 : 3'b000;
											assign node2679 = (inp[9]) ? 3'b000 : 3'b001;
										assign node2682 = (inp[0]) ? node2684 : 3'b100;
											assign node2684 = (inp[7]) ? 3'b101 : 3'b100;
									assign node2687 = (inp[7]) ? node2691 : node2688;
										assign node2688 = (inp[9]) ? 3'b101 : 3'b100;
										assign node2691 = (inp[9]) ? 3'b100 : 3'b101;
								assign node2694 = (inp[11]) ? node2708 : node2695;
									assign node2695 = (inp[1]) ? node2703 : node2696;
										assign node2696 = (inp[9]) ? node2700 : node2697;
											assign node2697 = (inp[7]) ? 3'b101 : 3'b100;
											assign node2700 = (inp[7]) ? 3'b100 : 3'b101;
										assign node2703 = (inp[9]) ? 3'b001 : node2704;
											assign node2704 = (inp[7]) ? 3'b001 : 3'b000;
									assign node2708 = (inp[9]) ? node2710 : 3'b001;
										assign node2710 = (inp[7]) ? 3'b000 : 3'b001;

endmodule