module dtc_split25_bm30 (
	input  wire [14-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node7;
	wire [8-1:0] node9;
	wire [8-1:0] node11;
	wire [8-1:0] node14;
	wire [8-1:0] node15;
	wire [8-1:0] node16;
	wire [8-1:0] node18;
	wire [8-1:0] node22;
	wire [8-1:0] node24;
	wire [8-1:0] node25;
	wire [8-1:0] node28;
	wire [8-1:0] node31;
	wire [8-1:0] node32;
	wire [8-1:0] node33;
	wire [8-1:0] node35;
	wire [8-1:0] node38;
	wire [8-1:0] node39;
	wire [8-1:0] node41;
	wire [8-1:0] node44;
	wire [8-1:0] node46;
	wire [8-1:0] node49;
	wire [8-1:0] node50;
	wire [8-1:0] node53;
	wire [8-1:0] node54;
	wire [8-1:0] node55;
	wire [8-1:0] node56;
	wire [8-1:0] node60;
	wire [8-1:0] node61;
	wire [8-1:0] node65;
	wire [8-1:0] node68;
	wire [8-1:0] node69;
	wire [8-1:0] node70;
	wire [8-1:0] node71;
	wire [8-1:0] node73;
	wire [8-1:0] node76;
	wire [8-1:0] node77;
	wire [8-1:0] node79;
	wire [8-1:0] node82;
	wire [8-1:0] node84;
	wire [8-1:0] node87;
	wire [8-1:0] node88;
	wire [8-1:0] node90;
	wire [8-1:0] node91;
	wire [8-1:0] node94;
	wire [8-1:0] node97;
	wire [8-1:0] node98;
	wire [8-1:0] node100;
	wire [8-1:0] node103;
	wire [8-1:0] node104;
	wire [8-1:0] node109;
	wire [8-1:0] node110;
	wire [8-1:0] node111;
	wire [8-1:0] node112;
	wire [8-1:0] node115;
	wire [8-1:0] node116;
	wire [8-1:0] node118;
	wire [8-1:0] node121;
	wire [8-1:0] node122;
	wire [8-1:0] node125;
	wire [8-1:0] node128;
	wire [8-1:0] node129;
	wire [8-1:0] node130;
	wire [8-1:0] node131;
	wire [8-1:0] node133;
	wire [8-1:0] node136;
	wire [8-1:0] node139;
	wire [8-1:0] node140;
	wire [8-1:0] node142;
	wire [8-1:0] node144;
	wire [8-1:0] node147;
	wire [8-1:0] node148;
	wire [8-1:0] node149;
	wire [8-1:0] node154;
	wire [8-1:0] node155;
	wire [8-1:0] node156;
	wire [8-1:0] node158;
	wire [8-1:0] node161;
	wire [8-1:0] node163;
	wire [8-1:0] node166;
	wire [8-1:0] node167;
	wire [8-1:0] node169;
	wire [8-1:0] node172;
	wire [8-1:0] node173;
	wire [8-1:0] node177;
	wire [8-1:0] node178;
	wire [8-1:0] node179;
	wire [8-1:0] node180;
	wire [8-1:0] node182;
	wire [8-1:0] node183;
	wire [8-1:0] node185;
	wire [8-1:0] node189;
	wire [8-1:0] node190;
	wire [8-1:0] node191;
	wire [8-1:0] node196;
	wire [8-1:0] node197;
	wire [8-1:0] node198;
	wire [8-1:0] node199;
	wire [8-1:0] node202;
	wire [8-1:0] node204;
	wire [8-1:0] node207;
	wire [8-1:0] node209;
	wire [8-1:0] node212;
	wire [8-1:0] node213;
	wire [8-1:0] node216;
	wire [8-1:0] node217;
	wire [8-1:0] node218;
	wire [8-1:0] node219;
	wire [8-1:0] node224;
	wire [8-1:0] node226;
	wire [8-1:0] node227;
	wire [8-1:0] node231;
	wire [8-1:0] node232;
	wire [8-1:0] node233;
	wire [8-1:0] node234;
	wire [8-1:0] node235;
	wire [8-1:0] node239;
	wire [8-1:0] node241;
	wire [8-1:0] node244;
	wire [8-1:0] node245;
	wire [8-1:0] node246;
	wire [8-1:0] node247;
	wire [8-1:0] node251;
	wire [8-1:0] node253;
	wire [8-1:0] node256;
	wire [8-1:0] node259;
	wire [8-1:0] node260;
	wire [8-1:0] node261;
	wire [8-1:0] node262;
	wire [8-1:0] node266;
	wire [8-1:0] node269;
	wire [8-1:0] node270;
	wire [8-1:0] node271;
	wire [8-1:0] node272;
	wire [8-1:0] node274;
	wire [8-1:0] node277;
	wire [8-1:0] node279;
	wire [8-1:0] node282;
	wire [8-1:0] node285;
	wire [8-1:0] node288;
	wire [8-1:0] node289;
	wire [8-1:0] node290;
	wire [8-1:0] node291;
	wire [8-1:0] node292;
	wire [8-1:0] node293;
	wire [8-1:0] node294;
	wire [8-1:0] node295;
	wire [8-1:0] node299;
	wire [8-1:0] node301;
	wire [8-1:0] node303;
	wire [8-1:0] node304;
	wire [8-1:0] node308;
	wire [8-1:0] node309;
	wire [8-1:0] node311;
	wire [8-1:0] node312;
	wire [8-1:0] node315;
	wire [8-1:0] node317;
	wire [8-1:0] node320;
	wire [8-1:0] node321;
	wire [8-1:0] node324;
	wire [8-1:0] node326;
	wire [8-1:0] node329;
	wire [8-1:0] node330;
	wire [8-1:0] node331;
	wire [8-1:0] node332;
	wire [8-1:0] node335;
	wire [8-1:0] node338;
	wire [8-1:0] node339;
	wire [8-1:0] node341;
	wire [8-1:0] node344;
	wire [8-1:0] node347;
	wire [8-1:0] node348;
	wire [8-1:0] node349;
	wire [8-1:0] node350;
	wire [8-1:0] node355;
	wire [8-1:0] node356;
	wire [8-1:0] node357;
	wire [8-1:0] node361;
	wire [8-1:0] node364;
	wire [8-1:0] node365;
	wire [8-1:0] node366;
	wire [8-1:0] node367;
	wire [8-1:0] node368;
	wire [8-1:0] node371;
	wire [8-1:0] node372;
	wire [8-1:0] node376;
	wire [8-1:0] node377;
	wire [8-1:0] node380;
	wire [8-1:0] node381;
	wire [8-1:0] node385;
	wire [8-1:0] node386;
	wire [8-1:0] node390;
	wire [8-1:0] node391;
	wire [8-1:0] node392;
	wire [8-1:0] node393;
	wire [8-1:0] node395;
	wire [8-1:0] node399;
	wire [8-1:0] node401;
	wire [8-1:0] node403;
	wire [8-1:0] node406;
	wire [8-1:0] node407;
	wire [8-1:0] node408;
	wire [8-1:0] node411;
	wire [8-1:0] node412;
	wire [8-1:0] node414;
	wire [8-1:0] node417;
	wire [8-1:0] node419;
	wire [8-1:0] node422;
	wire [8-1:0] node423;
	wire [8-1:0] node426;
	wire [8-1:0] node427;
	wire [8-1:0] node430;
	wire [8-1:0] node431;
	wire [8-1:0] node435;
	wire [8-1:0] node436;
	wire [8-1:0] node437;
	wire [8-1:0] node438;
	wire [8-1:0] node439;
	wire [8-1:0] node440;
	wire [8-1:0] node441;
	wire [8-1:0] node445;
	wire [8-1:0] node448;
	wire [8-1:0] node449;
	wire [8-1:0] node453;
	wire [8-1:0] node454;
	wire [8-1:0] node456;
	wire [8-1:0] node459;
	wire [8-1:0] node460;
	wire [8-1:0] node464;
	wire [8-1:0] node465;
	wire [8-1:0] node466;
	wire [8-1:0] node467;
	wire [8-1:0] node469;
	wire [8-1:0] node472;
	wire [8-1:0] node474;
	wire [8-1:0] node475;
	wire [8-1:0] node479;
	wire [8-1:0] node480;
	wire [8-1:0] node483;
	wire [8-1:0] node486;
	wire [8-1:0] node487;
	wire [8-1:0] node488;
	wire [8-1:0] node489;
	wire [8-1:0] node493;
	wire [8-1:0] node494;
	wire [8-1:0] node498;
	wire [8-1:0] node499;
	wire [8-1:0] node501;
	wire [8-1:0] node505;
	wire [8-1:0] node506;
	wire [8-1:0] node507;
	wire [8-1:0] node508;
	wire [8-1:0] node511;
	wire [8-1:0] node512;
	wire [8-1:0] node513;
	wire [8-1:0] node516;
	wire [8-1:0] node519;
	wire [8-1:0] node522;
	wire [8-1:0] node523;
	wire [8-1:0] node524;
	wire [8-1:0] node527;
	wire [8-1:0] node529;
	wire [8-1:0] node532;
	wire [8-1:0] node533;
	wire [8-1:0] node534;
	wire [8-1:0] node538;
	wire [8-1:0] node541;
	wire [8-1:0] node542;
	wire [8-1:0] node543;
	wire [8-1:0] node544;
	wire [8-1:0] node547;
	wire [8-1:0] node550;
	wire [8-1:0] node551;
	wire [8-1:0] node552;
	wire [8-1:0] node556;
	wire [8-1:0] node557;
	wire [8-1:0] node559;
	wire [8-1:0] node562;
	wire [8-1:0] node565;
	wire [8-1:0] node566;
	wire [8-1:0] node567;
	wire [8-1:0] node568;
	wire [8-1:0] node570;
	wire [8-1:0] node573;
	wire [8-1:0] node576;
	wire [8-1:0] node577;
	wire [8-1:0] node579;
	wire [8-1:0] node583;
	wire [8-1:0] node585;
	wire [8-1:0] node586;
	wire [8-1:0] node589;
	wire [8-1:0] node592;
	wire [8-1:0] node593;
	wire [8-1:0] node594;
	wire [8-1:0] node595;
	wire [8-1:0] node596;
	wire [8-1:0] node598;
	wire [8-1:0] node599;
	wire [8-1:0] node603;
	wire [8-1:0] node604;
	wire [8-1:0] node607;
	wire [8-1:0] node610;
	wire [8-1:0] node611;
	wire [8-1:0] node612;
	wire [8-1:0] node613;
	wire [8-1:0] node615;
	wire [8-1:0] node616;
	wire [8-1:0] node619;
	wire [8-1:0] node623;
	wire [8-1:0] node624;
	wire [8-1:0] node625;
	wire [8-1:0] node627;
	wire [8-1:0] node630;
	wire [8-1:0] node631;
	wire [8-1:0] node635;
	wire [8-1:0] node636;
	wire [8-1:0] node640;
	wire [8-1:0] node641;
	wire [8-1:0] node642;
	wire [8-1:0] node646;
	wire [8-1:0] node647;
	wire [8-1:0] node648;
	wire [8-1:0] node649;
	wire [8-1:0] node654;
	wire [8-1:0] node655;
	wire [8-1:0] node656;
	wire [8-1:0] node661;
	wire [8-1:0] node662;
	wire [8-1:0] node663;
	wire [8-1:0] node664;
	wire [8-1:0] node666;
	wire [8-1:0] node667;
	wire [8-1:0] node671;
	wire [8-1:0] node672;
	wire [8-1:0] node676;
	wire [8-1:0] node677;
	wire [8-1:0] node678;
	wire [8-1:0] node680;
	wire [8-1:0] node682;
	wire [8-1:0] node685;
	wire [8-1:0] node688;
	wire [8-1:0] node690;
	wire [8-1:0] node693;
	wire [8-1:0] node694;
	wire [8-1:0] node695;
	wire [8-1:0] node697;
	wire [8-1:0] node700;
	wire [8-1:0] node701;
	wire [8-1:0] node703;
	wire [8-1:0] node704;
	wire [8-1:0] node709;
	wire [8-1:0] node710;
	wire [8-1:0] node711;
	wire [8-1:0] node712;
	wire [8-1:0] node715;
	wire [8-1:0] node719;
	wire [8-1:0] node720;
	wire [8-1:0] node724;
	wire [8-1:0] node725;
	wire [8-1:0] node726;
	wire [8-1:0] node727;
	wire [8-1:0] node728;
	wire [8-1:0] node730;
	wire [8-1:0] node732;
	wire [8-1:0] node734;
	wire [8-1:0] node737;
	wire [8-1:0] node738;
	wire [8-1:0] node740;
	wire [8-1:0] node743;
	wire [8-1:0] node746;
	wire [8-1:0] node747;
	wire [8-1:0] node748;
	wire [8-1:0] node750;
	wire [8-1:0] node751;
	wire [8-1:0] node755;
	wire [8-1:0] node756;
	wire [8-1:0] node757;
	wire [8-1:0] node762;
	wire [8-1:0] node763;
	wire [8-1:0] node764;
	wire [8-1:0] node768;
	wire [8-1:0] node769;
	wire [8-1:0] node773;
	wire [8-1:0] node774;
	wire [8-1:0] node775;
	wire [8-1:0] node776;
	wire [8-1:0] node778;
	wire [8-1:0] node781;
	wire [8-1:0] node783;
	wire [8-1:0] node786;
	wire [8-1:0] node787;
	wire [8-1:0] node788;
	wire [8-1:0] node790;
	wire [8-1:0] node793;
	wire [8-1:0] node794;
	wire [8-1:0] node798;
	wire [8-1:0] node801;
	wire [8-1:0] node802;
	wire [8-1:0] node803;
	wire [8-1:0] node806;
	wire [8-1:0] node808;
	wire [8-1:0] node811;
	wire [8-1:0] node812;
	wire [8-1:0] node814;
	wire [8-1:0] node815;
	wire [8-1:0] node819;
	wire [8-1:0] node821;
	wire [8-1:0] node824;
	wire [8-1:0] node825;
	wire [8-1:0] node826;
	wire [8-1:0] node827;
	wire [8-1:0] node829;
	wire [8-1:0] node831;
	wire [8-1:0] node834;
	wire [8-1:0] node835;
	wire [8-1:0] node836;
	wire [8-1:0] node838;
	wire [8-1:0] node842;
	wire [8-1:0] node845;
	wire [8-1:0] node846;
	wire [8-1:0] node847;
	wire [8-1:0] node848;
	wire [8-1:0] node849;
	wire [8-1:0] node854;
	wire [8-1:0] node855;
	wire [8-1:0] node856;
	wire [8-1:0] node859;
	wire [8-1:0] node862;
	wire [8-1:0] node864;
	wire [8-1:0] node867;
	wire [8-1:0] node869;
	wire [8-1:0] node870;
	wire [8-1:0] node872;
	wire [8-1:0] node876;
	wire [8-1:0] node877;
	wire [8-1:0] node878;
	wire [8-1:0] node880;
	wire [8-1:0] node881;
	wire [8-1:0] node882;
	wire [8-1:0] node886;
	wire [8-1:0] node889;
	wire [8-1:0] node890;
	wire [8-1:0] node891;
	wire [8-1:0] node893;
	wire [8-1:0] node896;
	wire [8-1:0] node900;
	wire [8-1:0] node901;
	wire [8-1:0] node902;
	wire [8-1:0] node903;
	wire [8-1:0] node904;
	wire [8-1:0] node908;
	wire [8-1:0] node911;
	wire [8-1:0] node912;
	wire [8-1:0] node915;
	wire [8-1:0] node918;
	wire [8-1:0] node919;
	wire [8-1:0] node921;
	wire [8-1:0] node922;
	wire [8-1:0] node925;
	wire [8-1:0] node928;
	wire [8-1:0] node929;
	wire [8-1:0] node933;
	wire [8-1:0] node934;
	wire [8-1:0] node935;
	wire [8-1:0] node936;
	wire [8-1:0] node937;
	wire [8-1:0] node938;
	wire [8-1:0] node940;
	wire [8-1:0] node941;
	wire [8-1:0] node945;
	wire [8-1:0] node946;
	wire [8-1:0] node947;
	wire [8-1:0] node951;
	wire [8-1:0] node952;
	wire [8-1:0] node956;
	wire [8-1:0] node957;
	wire [8-1:0] node958;
	wire [8-1:0] node959;
	wire [8-1:0] node960;
	wire [8-1:0] node963;
	wire [8-1:0] node964;
	wire [8-1:0] node967;
	wire [8-1:0] node970;
	wire [8-1:0] node973;
	wire [8-1:0] node974;
	wire [8-1:0] node975;
	wire [8-1:0] node979;
	wire [8-1:0] node980;
	wire [8-1:0] node983;
	wire [8-1:0] node986;
	wire [8-1:0] node987;
	wire [8-1:0] node988;
	wire [8-1:0] node989;
	wire [8-1:0] node993;
	wire [8-1:0] node994;
	wire [8-1:0] node996;
	wire [8-1:0] node999;
	wire [8-1:0] node1001;
	wire [8-1:0] node1004;
	wire [8-1:0] node1005;
	wire [8-1:0] node1007;
	wire [8-1:0] node1010;
	wire [8-1:0] node1011;
	wire [8-1:0] node1013;
	wire [8-1:0] node1017;
	wire [8-1:0] node1018;
	wire [8-1:0] node1019;
	wire [8-1:0] node1020;
	wire [8-1:0] node1021;
	wire [8-1:0] node1025;
	wire [8-1:0] node1026;
	wire [8-1:0] node1030;
	wire [8-1:0] node1031;
	wire [8-1:0] node1032;
	wire [8-1:0] node1034;
	wire [8-1:0] node1035;
	wire [8-1:0] node1039;
	wire [8-1:0] node1040;
	wire [8-1:0] node1044;
	wire [8-1:0] node1045;
	wire [8-1:0] node1046;
	wire [8-1:0] node1049;
	wire [8-1:0] node1053;
	wire [8-1:0] node1054;
	wire [8-1:0] node1055;
	wire [8-1:0] node1056;
	wire [8-1:0] node1057;
	wire [8-1:0] node1061;
	wire [8-1:0] node1064;
	wire [8-1:0] node1065;
	wire [8-1:0] node1069;
	wire [8-1:0] node1070;
	wire [8-1:0] node1074;
	wire [8-1:0] node1075;
	wire [8-1:0] node1076;
	wire [8-1:0] node1077;
	wire [8-1:0] node1078;
	wire [8-1:0] node1079;
	wire [8-1:0] node1080;
	wire [8-1:0] node1084;
	wire [8-1:0] node1086;
	wire [8-1:0] node1089;
	wire [8-1:0] node1090;
	wire [8-1:0] node1091;
	wire [8-1:0] node1094;
	wire [8-1:0] node1095;
	wire [8-1:0] node1099;
	wire [8-1:0] node1100;
	wire [8-1:0] node1101;
	wire [8-1:0] node1105;
	wire [8-1:0] node1107;
	wire [8-1:0] node1109;
	wire [8-1:0] node1112;
	wire [8-1:0] node1113;
	wire [8-1:0] node1114;
	wire [8-1:0] node1115;
	wire [8-1:0] node1116;
	wire [8-1:0] node1119;
	wire [8-1:0] node1122;
	wire [8-1:0] node1123;
	wire [8-1:0] node1126;
	wire [8-1:0] node1129;
	wire [8-1:0] node1130;
	wire [8-1:0] node1132;
	wire [8-1:0] node1133;
	wire [8-1:0] node1137;
	wire [8-1:0] node1138;
	wire [8-1:0] node1141;
	wire [8-1:0] node1144;
	wire [8-1:0] node1145;
	wire [8-1:0] node1146;
	wire [8-1:0] node1148;
	wire [8-1:0] node1152;
	wire [8-1:0] node1155;
	wire [8-1:0] node1156;
	wire [8-1:0] node1157;
	wire [8-1:0] node1158;
	wire [8-1:0] node1159;
	wire [8-1:0] node1160;
	wire [8-1:0] node1164;
	wire [8-1:0] node1167;
	wire [8-1:0] node1169;
	wire [8-1:0] node1172;
	wire [8-1:0] node1173;
	wire [8-1:0] node1174;
	wire [8-1:0] node1175;
	wire [8-1:0] node1180;
	wire [8-1:0] node1181;
	wire [8-1:0] node1182;
	wire [8-1:0] node1185;
	wire [8-1:0] node1188;
	wire [8-1:0] node1189;
	wire [8-1:0] node1192;
	wire [8-1:0] node1195;
	wire [8-1:0] node1196;
	wire [8-1:0] node1197;
	wire [8-1:0] node1198;
	wire [8-1:0] node1199;
	wire [8-1:0] node1203;
	wire [8-1:0] node1206;
	wire [8-1:0] node1207;
	wire [8-1:0] node1211;
	wire [8-1:0] node1212;
	wire [8-1:0] node1213;
	wire [8-1:0] node1214;
	wire [8-1:0] node1217;
	wire [8-1:0] node1218;
	wire [8-1:0] node1222;
	wire [8-1:0] node1225;
	wire [8-1:0] node1226;
	wire [8-1:0] node1228;
	wire [8-1:0] node1231;
	wire [8-1:0] node1232;
	wire [8-1:0] node1236;
	wire [8-1:0] node1237;
	wire [8-1:0] node1238;
	wire [8-1:0] node1239;
	wire [8-1:0] node1240;
	wire [8-1:0] node1243;
	wire [8-1:0] node1244;
	wire [8-1:0] node1248;
	wire [8-1:0] node1249;
	wire [8-1:0] node1251;
	wire [8-1:0] node1252;
	wire [8-1:0] node1255;
	wire [8-1:0] node1258;
	wire [8-1:0] node1260;
	wire [8-1:0] node1263;
	wire [8-1:0] node1264;
	wire [8-1:0] node1265;
	wire [8-1:0] node1267;
	wire [8-1:0] node1270;
	wire [8-1:0] node1271;
	wire [8-1:0] node1274;
	wire [8-1:0] node1276;
	wire [8-1:0] node1279;
	wire [8-1:0] node1280;
	wire [8-1:0] node1282;
	wire [8-1:0] node1285;
	wire [8-1:0] node1288;
	wire [8-1:0] node1289;
	wire [8-1:0] node1290;
	wire [8-1:0] node1291;
	wire [8-1:0] node1294;
	wire [8-1:0] node1295;
	wire [8-1:0] node1296;
	wire [8-1:0] node1299;
	wire [8-1:0] node1301;
	wire [8-1:0] node1304;
	wire [8-1:0] node1305;
	wire [8-1:0] node1306;
	wire [8-1:0] node1309;
	wire [8-1:0] node1312;
	wire [8-1:0] node1315;
	wire [8-1:0] node1316;
	wire [8-1:0] node1318;
	wire [8-1:0] node1319;
	wire [8-1:0] node1322;
	wire [8-1:0] node1323;
	wire [8-1:0] node1326;
	wire [8-1:0] node1329;
	wire [8-1:0] node1330;
	wire [8-1:0] node1331;
	wire [8-1:0] node1335;
	wire [8-1:0] node1336;
	wire [8-1:0] node1339;
	wire [8-1:0] node1341;
	wire [8-1:0] node1344;
	wire [8-1:0] node1345;
	wire [8-1:0] node1346;
	wire [8-1:0] node1347;
	wire [8-1:0] node1348;
	wire [8-1:0] node1351;
	wire [8-1:0] node1353;
	wire [8-1:0] node1356;
	wire [8-1:0] node1358;
	wire [8-1:0] node1360;
	wire [8-1:0] node1363;
	wire [8-1:0] node1364;
	wire [8-1:0] node1365;
	wire [8-1:0] node1366;
	wire [8-1:0] node1369;
	wire [8-1:0] node1373;
	wire [8-1:0] node1375;
	wire [8-1:0] node1378;
	wire [8-1:0] node1379;
	wire [8-1:0] node1380;
	wire [8-1:0] node1383;
	wire [8-1:0] node1384;
	wire [8-1:0] node1387;
	wire [8-1:0] node1388;
	wire [8-1:0] node1392;
	wire [8-1:0] node1393;
	wire [8-1:0] node1395;
	wire [8-1:0] node1398;
	wire [8-1:0] node1399;
	wire [8-1:0] node1400;
	wire [8-1:0] node1404;
	wire [8-1:0] node1405;
	wire [8-1:0] node1408;
	wire [8-1:0] node1411;
	wire [8-1:0] node1412;
	wire [8-1:0] node1413;
	wire [8-1:0] node1414;
	wire [8-1:0] node1415;
	wire [8-1:0] node1416;
	wire [8-1:0] node1417;
	wire [8-1:0] node1419;
	wire [8-1:0] node1422;
	wire [8-1:0] node1423;
	wire [8-1:0] node1425;
	wire [8-1:0] node1428;
	wire [8-1:0] node1430;
	wire [8-1:0] node1433;
	wire [8-1:0] node1434;
	wire [8-1:0] node1435;
	wire [8-1:0] node1437;
	wire [8-1:0] node1440;
	wire [8-1:0] node1442;
	wire [8-1:0] node1446;
	wire [8-1:0] node1447;
	wire [8-1:0] node1448;
	wire [8-1:0] node1449;
	wire [8-1:0] node1451;
	wire [8-1:0] node1452;
	wire [8-1:0] node1456;
	wire [8-1:0] node1457;
	wire [8-1:0] node1458;
	wire [8-1:0] node1463;
	wire [8-1:0] node1464;
	wire [8-1:0] node1465;
	wire [8-1:0] node1468;
	wire [8-1:0] node1469;
	wire [8-1:0] node1473;
	wire [8-1:0] node1475;
	wire [8-1:0] node1478;
	wire [8-1:0] node1479;
	wire [8-1:0] node1480;
	wire [8-1:0] node1483;
	wire [8-1:0] node1485;
	wire [8-1:0] node1486;
	wire [8-1:0] node1489;
	wire [8-1:0] node1492;
	wire [8-1:0] node1494;
	wire [8-1:0] node1495;
	wire [8-1:0] node1499;
	wire [8-1:0] node1500;
	wire [8-1:0] node1501;
	wire [8-1:0] node1502;
	wire [8-1:0] node1503;
	wire [8-1:0] node1504;
	wire [8-1:0] node1509;
	wire [8-1:0] node1510;
	wire [8-1:0] node1511;
	wire [8-1:0] node1514;
	wire [8-1:0] node1516;
	wire [8-1:0] node1519;
	wire [8-1:0] node1520;
	wire [8-1:0] node1523;
	wire [8-1:0] node1526;
	wire [8-1:0] node1527;
	wire [8-1:0] node1528;
	wire [8-1:0] node1530;
	wire [8-1:0] node1532;
	wire [8-1:0] node1535;
	wire [8-1:0] node1536;
	wire [8-1:0] node1537;
	wire [8-1:0] node1542;
	wire [8-1:0] node1543;
	wire [8-1:0] node1545;
	wire [8-1:0] node1548;
	wire [8-1:0] node1551;
	wire [8-1:0] node1552;
	wire [8-1:0] node1553;
	wire [8-1:0] node1554;
	wire [8-1:0] node1556;
	wire [8-1:0] node1559;
	wire [8-1:0] node1561;
	wire [8-1:0] node1564;
	wire [8-1:0] node1565;
	wire [8-1:0] node1566;
	wire [8-1:0] node1570;
	wire [8-1:0] node1572;
	wire [8-1:0] node1573;
	wire [8-1:0] node1577;
	wire [8-1:0] node1578;
	wire [8-1:0] node1579;
	wire [8-1:0] node1583;
	wire [8-1:0] node1585;
	wire [8-1:0] node1588;
	wire [8-1:0] node1589;
	wire [8-1:0] node1591;
	wire [8-1:0] node1593;
	wire [8-1:0] node1596;
	wire [8-1:0] node1597;
	wire [8-1:0] node1598;
	wire [8-1:0] node1599;
	wire [8-1:0] node1601;
	wire [8-1:0] node1602;
	wire [8-1:0] node1606;
	wire [8-1:0] node1607;
	wire [8-1:0] node1610;
	wire [8-1:0] node1613;
	wire [8-1:0] node1614;
	wire [8-1:0] node1615;
	wire [8-1:0] node1618;
	wire [8-1:0] node1621;
	wire [8-1:0] node1623;
	wire [8-1:0] node1625;
	wire [8-1:0] node1627;
	wire [8-1:0] node1630;
	wire [8-1:0] node1631;
	wire [8-1:0] node1632;
	wire [8-1:0] node1633;
	wire [8-1:0] node1634;
	wire [8-1:0] node1638;
	wire [8-1:0] node1640;
	wire [8-1:0] node1643;
	wire [8-1:0] node1646;
	wire [8-1:0] node1647;
	wire [8-1:0] node1648;
	wire [8-1:0] node1652;
	wire [8-1:0] node1653;
	wire [8-1:0] node1657;
	wire [8-1:0] node1658;
	wire [8-1:0] node1659;
	wire [8-1:0] node1660;
	wire [8-1:0] node1661;
	wire [8-1:0] node1662;
	wire [8-1:0] node1663;
	wire [8-1:0] node1665;
	wire [8-1:0] node1668;
	wire [8-1:0] node1671;
	wire [8-1:0] node1672;
	wire [8-1:0] node1673;
	wire [8-1:0] node1676;
	wire [8-1:0] node1679;
	wire [8-1:0] node1680;
	wire [8-1:0] node1682;
	wire [8-1:0] node1686;
	wire [8-1:0] node1687;
	wire [8-1:0] node1688;
	wire [8-1:0] node1691;
	wire [8-1:0] node1694;
	wire [8-1:0] node1695;
	wire [8-1:0] node1696;
	wire [8-1:0] node1698;
	wire [8-1:0] node1701;
	wire [8-1:0] node1703;
	wire [8-1:0] node1706;
	wire [8-1:0] node1708;
	wire [8-1:0] node1711;
	wire [8-1:0] node1712;
	wire [8-1:0] node1713;
	wire [8-1:0] node1715;
	wire [8-1:0] node1718;
	wire [8-1:0] node1720;
	wire [8-1:0] node1723;
	wire [8-1:0] node1724;
	wire [8-1:0] node1725;
	wire [8-1:0] node1728;
	wire [8-1:0] node1731;
	wire [8-1:0] node1732;
	wire [8-1:0] node1734;
	wire [8-1:0] node1738;
	wire [8-1:0] node1739;
	wire [8-1:0] node1740;
	wire [8-1:0] node1741;
	wire [8-1:0] node1742;
	wire [8-1:0] node1744;
	wire [8-1:0] node1747;
	wire [8-1:0] node1748;
	wire [8-1:0] node1749;
	wire [8-1:0] node1753;
	wire [8-1:0] node1756;
	wire [8-1:0] node1758;
	wire [8-1:0] node1759;
	wire [8-1:0] node1763;
	wire [8-1:0] node1764;
	wire [8-1:0] node1767;
	wire [8-1:0] node1768;
	wire [8-1:0] node1771;
	wire [8-1:0] node1774;
	wire [8-1:0] node1775;
	wire [8-1:0] node1776;
	wire [8-1:0] node1777;
	wire [8-1:0] node1780;
	wire [8-1:0] node1783;
	wire [8-1:0] node1784;
	wire [8-1:0] node1785;
	wire [8-1:0] node1788;
	wire [8-1:0] node1792;
	wire [8-1:0] node1793;
	wire [8-1:0] node1796;
	wire [8-1:0] node1799;
	wire [8-1:0] node1800;
	wire [8-1:0] node1801;
	wire [8-1:0] node1802;
	wire [8-1:0] node1803;
	wire [8-1:0] node1804;
	wire [8-1:0] node1806;
	wire [8-1:0] node1809;
	wire [8-1:0] node1810;
	wire [8-1:0] node1813;
	wire [8-1:0] node1816;
	wire [8-1:0] node1817;
	wire [8-1:0] node1820;
	wire [8-1:0] node1821;
	wire [8-1:0] node1822;
	wire [8-1:0] node1826;
	wire [8-1:0] node1829;
	wire [8-1:0] node1830;
	wire [8-1:0] node1832;
	wire [8-1:0] node1834;
	wire [8-1:0] node1837;
	wire [8-1:0] node1838;
	wire [8-1:0] node1841;
	wire [8-1:0] node1844;
	wire [8-1:0] node1845;
	wire [8-1:0] node1846;
	wire [8-1:0] node1847;
	wire [8-1:0] node1849;
	wire [8-1:0] node1852;
	wire [8-1:0] node1853;
	wire [8-1:0] node1854;
	wire [8-1:0] node1859;
	wire [8-1:0] node1861;
	wire [8-1:0] node1862;
	wire [8-1:0] node1863;
	wire [8-1:0] node1867;
	wire [8-1:0] node1868;
	wire [8-1:0] node1872;
	wire [8-1:0] node1873;
	wire [8-1:0] node1874;
	wire [8-1:0] node1877;
	wire [8-1:0] node1880;
	wire [8-1:0] node1883;
	wire [8-1:0] node1884;
	wire [8-1:0] node1885;
	wire [8-1:0] node1886;
	wire [8-1:0] node1887;
	wire [8-1:0] node1888;
	wire [8-1:0] node1891;
	wire [8-1:0] node1892;
	wire [8-1:0] node1895;
	wire [8-1:0] node1898;
	wire [8-1:0] node1901;
	wire [8-1:0] node1902;
	wire [8-1:0] node1905;
	wire [8-1:0] node1906;
	wire [8-1:0] node1909;
	wire [8-1:0] node1912;
	wire [8-1:0] node1913;
	wire [8-1:0] node1914;
	wire [8-1:0] node1915;
	wire [8-1:0] node1918;
	wire [8-1:0] node1921;
	wire [8-1:0] node1922;
	wire [8-1:0] node1924;
	wire [8-1:0] node1928;
	wire [8-1:0] node1929;
	wire [8-1:0] node1932;
	wire [8-1:0] node1935;
	wire [8-1:0] node1936;
	wire [8-1:0] node1937;
	wire [8-1:0] node1939;
	wire [8-1:0] node1942;
	wire [8-1:0] node1943;
	wire [8-1:0] node1944;
	wire [8-1:0] node1949;
	wire [8-1:0] node1952;
	wire [8-1:0] node1953;
	wire [8-1:0] node1954;
	wire [8-1:0] node1955;
	wire [8-1:0] node1956;
	wire [8-1:0] node1957;
	wire [8-1:0] node1958;
	wire [8-1:0] node1959;
	wire [8-1:0] node1960;
	wire [8-1:0] node1961;
	wire [8-1:0] node1965;
	wire [8-1:0] node1966;
	wire [8-1:0] node1969;
	wire [8-1:0] node1970;
	wire [8-1:0] node1974;
	wire [8-1:0] node1975;
	wire [8-1:0] node1978;
	wire [8-1:0] node1981;
	wire [8-1:0] node1982;
	wire [8-1:0] node1983;
	wire [8-1:0] node1985;
	wire [8-1:0] node1988;
	wire [8-1:0] node1990;
	wire [8-1:0] node1993;
	wire [8-1:0] node1995;
	wire [8-1:0] node1997;
	wire [8-1:0] node2000;
	wire [8-1:0] node2001;
	wire [8-1:0] node2002;
	wire [8-1:0] node2003;
	wire [8-1:0] node2004;
	wire [8-1:0] node2005;
	wire [8-1:0] node2007;
	wire [8-1:0] node2010;
	wire [8-1:0] node2012;
	wire [8-1:0] node2015;
	wire [8-1:0] node2016;
	wire [8-1:0] node2017;
	wire [8-1:0] node2022;
	wire [8-1:0] node2023;
	wire [8-1:0] node2025;
	wire [8-1:0] node2028;
	wire [8-1:0] node2030;
	wire [8-1:0] node2033;
	wire [8-1:0] node2034;
	wire [8-1:0] node2035;
	wire [8-1:0] node2037;
	wire [8-1:0] node2039;
	wire [8-1:0] node2042;
	wire [8-1:0] node2045;
	wire [8-1:0] node2046;
	wire [8-1:0] node2047;
	wire [8-1:0] node2048;
	wire [8-1:0] node2052;
	wire [8-1:0] node2054;
	wire [8-1:0] node2057;
	wire [8-1:0] node2058;
	wire [8-1:0] node2062;
	wire [8-1:0] node2063;
	wire [8-1:0] node2064;
	wire [8-1:0] node2066;
	wire [8-1:0] node2069;
	wire [8-1:0] node2070;
	wire [8-1:0] node2073;
	wire [8-1:0] node2076;
	wire [8-1:0] node2077;
	wire [8-1:0] node2079;
	wire [8-1:0] node2082;
	wire [8-1:0] node2083;
	wire [8-1:0] node2085;
	wire [8-1:0] node2089;
	wire [8-1:0] node2090;
	wire [8-1:0] node2091;
	wire [8-1:0] node2092;
	wire [8-1:0] node2093;
	wire [8-1:0] node2094;
	wire [8-1:0] node2095;
	wire [8-1:0] node2099;
	wire [8-1:0] node2101;
	wire [8-1:0] node2104;
	wire [8-1:0] node2105;
	wire [8-1:0] node2107;
	wire [8-1:0] node2110;
	wire [8-1:0] node2111;
	wire [8-1:0] node2114;
	wire [8-1:0] node2117;
	wire [8-1:0] node2118;
	wire [8-1:0] node2119;
	wire [8-1:0] node2121;
	wire [8-1:0] node2124;
	wire [8-1:0] node2127;
	wire [8-1:0] node2128;
	wire [8-1:0] node2129;
	wire [8-1:0] node2133;
	wire [8-1:0] node2134;
	wire [8-1:0] node2138;
	wire [8-1:0] node2139;
	wire [8-1:0] node2140;
	wire [8-1:0] node2141;
	wire [8-1:0] node2144;
	wire [8-1:0] node2145;
	wire [8-1:0] node2146;
	wire [8-1:0] node2151;
	wire [8-1:0] node2152;
	wire [8-1:0] node2155;
	wire [8-1:0] node2157;
	wire [8-1:0] node2160;
	wire [8-1:0] node2161;
	wire [8-1:0] node2162;
	wire [8-1:0] node2164;
	wire [8-1:0] node2166;
	wire [8-1:0] node2169;
	wire [8-1:0] node2170;
	wire [8-1:0] node2174;
	wire [8-1:0] node2176;
	wire [8-1:0] node2177;
	wire [8-1:0] node2180;
	wire [8-1:0] node2183;
	wire [8-1:0] node2184;
	wire [8-1:0] node2185;
	wire [8-1:0] node2186;
	wire [8-1:0] node2187;
	wire [8-1:0] node2188;
	wire [8-1:0] node2191;
	wire [8-1:0] node2194;
	wire [8-1:0] node2197;
	wire [8-1:0] node2198;
	wire [8-1:0] node2202;
	wire [8-1:0] node2203;
	wire [8-1:0] node2204;
	wire [8-1:0] node2205;
	wire [8-1:0] node2209;
	wire [8-1:0] node2210;
	wire [8-1:0] node2211;
	wire [8-1:0] node2215;
	wire [8-1:0] node2216;
	wire [8-1:0] node2220;
	wire [8-1:0] node2221;
	wire [8-1:0] node2222;
	wire [8-1:0] node2224;
	wire [8-1:0] node2227;
	wire [8-1:0] node2228;
	wire [8-1:0] node2231;
	wire [8-1:0] node2235;
	wire [8-1:0] node2236;
	wire [8-1:0] node2237;
	wire [8-1:0] node2238;
	wire [8-1:0] node2240;
	wire [8-1:0] node2241;
	wire [8-1:0] node2245;
	wire [8-1:0] node2246;
	wire [8-1:0] node2250;
	wire [8-1:0] node2251;
	wire [8-1:0] node2253;
	wire [8-1:0] node2255;
	wire [8-1:0] node2258;
	wire [8-1:0] node2259;
	wire [8-1:0] node2261;
	wire [8-1:0] node2264;
	wire [8-1:0] node2266;
	wire [8-1:0] node2269;
	wire [8-1:0] node2270;
	wire [8-1:0] node2271;
	wire [8-1:0] node2272;
	wire [8-1:0] node2276;
	wire [8-1:0] node2279;
	wire [8-1:0] node2280;
	wire [8-1:0] node2282;
	wire [8-1:0] node2285;
	wire [8-1:0] node2287;
	wire [8-1:0] node2290;
	wire [8-1:0] node2291;
	wire [8-1:0] node2292;
	wire [8-1:0] node2293;
	wire [8-1:0] node2294;
	wire [8-1:0] node2295;
	wire [8-1:0] node2296;
	wire [8-1:0] node2298;
	wire [8-1:0] node2300;
	wire [8-1:0] node2304;
	wire [8-1:0] node2306;
	wire [8-1:0] node2309;
	wire [8-1:0] node2310;
	wire [8-1:0] node2311;
	wire [8-1:0] node2312;
	wire [8-1:0] node2316;
	wire [8-1:0] node2318;
	wire [8-1:0] node2322;
	wire [8-1:0] node2323;
	wire [8-1:0] node2324;
	wire [8-1:0] node2325;
	wire [8-1:0] node2326;
	wire [8-1:0] node2329;
	wire [8-1:0] node2332;
	wire [8-1:0] node2333;
	wire [8-1:0] node2336;
	wire [8-1:0] node2338;
	wire [8-1:0] node2341;
	wire [8-1:0] node2342;
	wire [8-1:0] node2345;
	wire [8-1:0] node2346;
	wire [8-1:0] node2350;
	wire [8-1:0] node2351;
	wire [8-1:0] node2354;
	wire [8-1:0] node2355;
	wire [8-1:0] node2358;
	wire [8-1:0] node2359;
	wire [8-1:0] node2363;
	wire [8-1:0] node2364;
	wire [8-1:0] node2365;
	wire [8-1:0] node2367;
	wire [8-1:0] node2368;
	wire [8-1:0] node2370;
	wire [8-1:0] node2373;
	wire [8-1:0] node2376;
	wire [8-1:0] node2377;
	wire [8-1:0] node2378;
	wire [8-1:0] node2381;
	wire [8-1:0] node2384;
	wire [8-1:0] node2385;
	wire [8-1:0] node2387;
	wire [8-1:0] node2390;
	wire [8-1:0] node2391;
	wire [8-1:0] node2395;
	wire [8-1:0] node2396;
	wire [8-1:0] node2397;
	wire [8-1:0] node2398;
	wire [8-1:0] node2400;
	wire [8-1:0] node2401;
	wire [8-1:0] node2405;
	wire [8-1:0] node2407;
	wire [8-1:0] node2410;
	wire [8-1:0] node2411;
	wire [8-1:0] node2412;
	wire [8-1:0] node2413;
	wire [8-1:0] node2419;
	wire [8-1:0] node2420;
	wire [8-1:0] node2421;
	wire [8-1:0] node2424;
	wire [8-1:0] node2426;
	wire [8-1:0] node2427;
	wire [8-1:0] node2431;
	wire [8-1:0] node2433;
	wire [8-1:0] node2435;
	wire [8-1:0] node2438;
	wire [8-1:0] node2439;
	wire [8-1:0] node2440;
	wire [8-1:0] node2441;
	wire [8-1:0] node2442;
	wire [8-1:0] node2443;
	wire [8-1:0] node2444;
	wire [8-1:0] node2449;
	wire [8-1:0] node2452;
	wire [8-1:0] node2453;
	wire [8-1:0] node2455;
	wire [8-1:0] node2456;
	wire [8-1:0] node2461;
	wire [8-1:0] node2462;
	wire [8-1:0] node2463;
	wire [8-1:0] node2464;
	wire [8-1:0] node2467;
	wire [8-1:0] node2469;
	wire [8-1:0] node2472;
	wire [8-1:0] node2473;
	wire [8-1:0] node2475;
	wire [8-1:0] node2476;
	wire [8-1:0] node2480;
	wire [8-1:0] node2481;
	wire [8-1:0] node2485;
	wire [8-1:0] node2486;
	wire [8-1:0] node2487;
	wire [8-1:0] node2488;
	wire [8-1:0] node2491;
	wire [8-1:0] node2494;
	wire [8-1:0] node2496;
	wire [8-1:0] node2499;
	wire [8-1:0] node2500;
	wire [8-1:0] node2501;
	wire [8-1:0] node2502;
	wire [8-1:0] node2506;
	wire [8-1:0] node2508;
	wire [8-1:0] node2511;
	wire [8-1:0] node2514;
	wire [8-1:0] node2515;
	wire [8-1:0] node2516;
	wire [8-1:0] node2517;
	wire [8-1:0] node2518;
	wire [8-1:0] node2521;
	wire [8-1:0] node2524;
	wire [8-1:0] node2525;
	wire [8-1:0] node2528;
	wire [8-1:0] node2529;
	wire [8-1:0] node2530;
	wire [8-1:0] node2535;
	wire [8-1:0] node2536;
	wire [8-1:0] node2537;
	wire [8-1:0] node2538;
	wire [8-1:0] node2541;
	wire [8-1:0] node2543;
	wire [8-1:0] node2546;
	wire [8-1:0] node2549;
	wire [8-1:0] node2552;
	wire [8-1:0] node2553;
	wire [8-1:0] node2554;
	wire [8-1:0] node2555;
	wire [8-1:0] node2558;
	wire [8-1:0] node2559;
	wire [8-1:0] node2562;
	wire [8-1:0] node2563;
	wire [8-1:0] node2567;
	wire [8-1:0] node2568;
	wire [8-1:0] node2569;
	wire [8-1:0] node2571;
	wire [8-1:0] node2575;
	wire [8-1:0] node2576;
	wire [8-1:0] node2579;
	wire [8-1:0] node2582;
	wire [8-1:0] node2583;
	wire [8-1:0] node2584;
	wire [8-1:0] node2585;
	wire [8-1:0] node2586;
	wire [8-1:0] node2591;
	wire [8-1:0] node2592;
	wire [8-1:0] node2595;
	wire [8-1:0] node2598;
	wire [8-1:0] node2599;
	wire [8-1:0] node2602;
	wire [8-1:0] node2605;
	wire [8-1:0] node2606;
	wire [8-1:0] node2607;
	wire [8-1:0] node2608;
	wire [8-1:0] node2609;
	wire [8-1:0] node2610;
	wire [8-1:0] node2611;
	wire [8-1:0] node2612;
	wire [8-1:0] node2615;
	wire [8-1:0] node2616;
	wire [8-1:0] node2620;
	wire [8-1:0] node2621;
	wire [8-1:0] node2625;
	wire [8-1:0] node2626;
	wire [8-1:0] node2627;
	wire [8-1:0] node2628;
	wire [8-1:0] node2632;
	wire [8-1:0] node2633;
	wire [8-1:0] node2637;
	wire [8-1:0] node2638;
	wire [8-1:0] node2642;
	wire [8-1:0] node2643;
	wire [8-1:0] node2644;
	wire [8-1:0] node2645;
	wire [8-1:0] node2648;
	wire [8-1:0] node2649;
	wire [8-1:0] node2653;
	wire [8-1:0] node2654;
	wire [8-1:0] node2657;
	wire [8-1:0] node2660;
	wire [8-1:0] node2661;
	wire [8-1:0] node2662;
	wire [8-1:0] node2663;
	wire [8-1:0] node2667;
	wire [8-1:0] node2668;
	wire [8-1:0] node2673;
	wire [8-1:0] node2674;
	wire [8-1:0] node2675;
	wire [8-1:0] node2676;
	wire [8-1:0] node2677;
	wire [8-1:0] node2678;
	wire [8-1:0] node2683;
	wire [8-1:0] node2684;
	wire [8-1:0] node2688;
	wire [8-1:0] node2689;
	wire [8-1:0] node2690;
	wire [8-1:0] node2691;
	wire [8-1:0] node2696;
	wire [8-1:0] node2697;
	wire [8-1:0] node2701;
	wire [8-1:0] node2702;
	wire [8-1:0] node2704;
	wire [8-1:0] node2705;
	wire [8-1:0] node2709;
	wire [8-1:0] node2710;
	wire [8-1:0] node2714;
	wire [8-1:0] node2715;
	wire [8-1:0] node2716;
	wire [8-1:0] node2717;
	wire [8-1:0] node2718;
	wire [8-1:0] node2720;
	wire [8-1:0] node2721;
	wire [8-1:0] node2725;
	wire [8-1:0] node2726;
	wire [8-1:0] node2727;
	wire [8-1:0] node2729;
	wire [8-1:0] node2732;
	wire [8-1:0] node2735;
	wire [8-1:0] node2736;
	wire [8-1:0] node2738;
	wire [8-1:0] node2741;
	wire [8-1:0] node2742;
	wire [8-1:0] node2746;
	wire [8-1:0] node2747;
	wire [8-1:0] node2748;
	wire [8-1:0] node2751;
	wire [8-1:0] node2752;
	wire [8-1:0] node2756;
	wire [8-1:0] node2758;
	wire [8-1:0] node2759;
	wire [8-1:0] node2760;
	wire [8-1:0] node2765;
	wire [8-1:0] node2766;
	wire [8-1:0] node2767;
	wire [8-1:0] node2768;
	wire [8-1:0] node2770;
	wire [8-1:0] node2773;
	wire [8-1:0] node2776;
	wire [8-1:0] node2777;
	wire [8-1:0] node2781;
	wire [8-1:0] node2782;
	wire [8-1:0] node2783;
	wire [8-1:0] node2784;
	wire [8-1:0] node2787;
	wire [8-1:0] node2790;
	wire [8-1:0] node2793;
	wire [8-1:0] node2794;
	wire [8-1:0] node2796;
	wire [8-1:0] node2799;
	wire [8-1:0] node2800;
	wire [8-1:0] node2804;
	wire [8-1:0] node2805;
	wire [8-1:0] node2806;
	wire [8-1:0] node2807;
	wire [8-1:0] node2808;
	wire [8-1:0] node2811;
	wire [8-1:0] node2813;
	wire [8-1:0] node2816;
	wire [8-1:0] node2817;
	wire [8-1:0] node2818;
	wire [8-1:0] node2822;
	wire [8-1:0] node2823;
	wire [8-1:0] node2827;
	wire [8-1:0] node2828;
	wire [8-1:0] node2829;
	wire [8-1:0] node2832;
	wire [8-1:0] node2834;
	wire [8-1:0] node2837;
	wire [8-1:0] node2838;
	wire [8-1:0] node2839;
	wire [8-1:0] node2842;
	wire [8-1:0] node2845;
	wire [8-1:0] node2848;
	wire [8-1:0] node2849;
	wire [8-1:0] node2850;
	wire [8-1:0] node2853;
	wire [8-1:0] node2854;
	wire [8-1:0] node2855;
	wire [8-1:0] node2858;
	wire [8-1:0] node2861;
	wire [8-1:0] node2862;
	wire [8-1:0] node2866;
	wire [8-1:0] node2867;
	wire [8-1:0] node2868;
	wire [8-1:0] node2871;
	wire [8-1:0] node2872;
	wire [8-1:0] node2873;
	wire [8-1:0] node2877;
	wire [8-1:0] node2880;
	wire [8-1:0] node2881;
	wire [8-1:0] node2882;
	wire [8-1:0] node2883;
	wire [8-1:0] node2887;
	wire [8-1:0] node2888;
	wire [8-1:0] node2892;
	wire [8-1:0] node2893;
	wire [8-1:0] node2895;
	wire [8-1:0] node2899;
	wire [8-1:0] node2900;
	wire [8-1:0] node2901;
	wire [8-1:0] node2902;
	wire [8-1:0] node2903;
	wire [8-1:0] node2904;
	wire [8-1:0] node2905;
	wire [8-1:0] node2908;
	wire [8-1:0] node2911;
	wire [8-1:0] node2912;
	wire [8-1:0] node2913;
	wire [8-1:0] node2917;
	wire [8-1:0] node2919;
	wire [8-1:0] node2922;
	wire [8-1:0] node2923;
	wire [8-1:0] node2924;
	wire [8-1:0] node2925;
	wire [8-1:0] node2928;
	wire [8-1:0] node2931;
	wire [8-1:0] node2932;
	wire [8-1:0] node2935;
	wire [8-1:0] node2937;
	wire [8-1:0] node2940;
	wire [8-1:0] node2941;
	wire [8-1:0] node2942;
	wire [8-1:0] node2944;
	wire [8-1:0] node2947;
	wire [8-1:0] node2950;
	wire [8-1:0] node2951;
	wire [8-1:0] node2953;
	wire [8-1:0] node2956;
	wire [8-1:0] node2959;
	wire [8-1:0] node2960;
	wire [8-1:0] node2961;
	wire [8-1:0] node2962;
	wire [8-1:0] node2963;
	wire [8-1:0] node2964;
	wire [8-1:0] node2969;
	wire [8-1:0] node2972;
	wire [8-1:0] node2973;
	wire [8-1:0] node2976;
	wire [8-1:0] node2978;
	wire [8-1:0] node2981;
	wire [8-1:0] node2982;
	wire [8-1:0] node2983;
	wire [8-1:0] node2984;
	wire [8-1:0] node2987;
	wire [8-1:0] node2990;
	wire [8-1:0] node2993;
	wire [8-1:0] node2994;
	wire [8-1:0] node2995;
	wire [8-1:0] node2998;
	wire [8-1:0] node3001;
	wire [8-1:0] node3002;
	wire [8-1:0] node3005;
	wire [8-1:0] node3007;
	wire [8-1:0] node3010;
	wire [8-1:0] node3011;
	wire [8-1:0] node3012;
	wire [8-1:0] node3014;
	wire [8-1:0] node3016;
	wire [8-1:0] node3018;
	wire [8-1:0] node3021;
	wire [8-1:0] node3022;
	wire [8-1:0] node3024;
	wire [8-1:0] node3027;
	wire [8-1:0] node3028;
	wire [8-1:0] node3032;
	wire [8-1:0] node3033;
	wire [8-1:0] node3034;
	wire [8-1:0] node3035;
	wire [8-1:0] node3036;
	wire [8-1:0] node3040;
	wire [8-1:0] node3043;
	wire [8-1:0] node3046;
	wire [8-1:0] node3047;
	wire [8-1:0] node3048;
	wire [8-1:0] node3051;
	wire [8-1:0] node3053;
	wire [8-1:0] node3056;
	wire [8-1:0] node3057;
	wire [8-1:0] node3060;
	wire [8-1:0] node3063;
	wire [8-1:0] node3064;
	wire [8-1:0] node3065;
	wire [8-1:0] node3066;
	wire [8-1:0] node3067;
	wire [8-1:0] node3068;
	wire [8-1:0] node3070;
	wire [8-1:0] node3073;
	wire [8-1:0] node3075;
	wire [8-1:0] node3076;
	wire [8-1:0] node3080;
	wire [8-1:0] node3081;
	wire [8-1:0] node3082;
	wire [8-1:0] node3087;
	wire [8-1:0] node3088;
	wire [8-1:0] node3090;
	wire [8-1:0] node3093;
	wire [8-1:0] node3094;
	wire [8-1:0] node3095;
	wire [8-1:0] node3099;
	wire [8-1:0] node3102;
	wire [8-1:0] node3103;
	wire [8-1:0] node3104;
	wire [8-1:0] node3105;
	wire [8-1:0] node3106;
	wire [8-1:0] node3108;
	wire [8-1:0] node3112;
	wire [8-1:0] node3115;
	wire [8-1:0] node3116;
	wire [8-1:0] node3119;
	wire [8-1:0] node3122;
	wire [8-1:0] node3123;
	wire [8-1:0] node3124;
	wire [8-1:0] node3126;
	wire [8-1:0] node3129;
	wire [8-1:0] node3130;
	wire [8-1:0] node3134;
	wire [8-1:0] node3135;
	wire [8-1:0] node3136;
	wire [8-1:0] node3140;
	wire [8-1:0] node3142;
	wire [8-1:0] node3145;
	wire [8-1:0] node3146;
	wire [8-1:0] node3147;
	wire [8-1:0] node3148;
	wire [8-1:0] node3149;
	wire [8-1:0] node3150;
	wire [8-1:0] node3152;
	wire [8-1:0] node3156;
	wire [8-1:0] node3158;
	wire [8-1:0] node3160;
	wire [8-1:0] node3163;
	wire [8-1:0] node3164;
	wire [8-1:0] node3166;
	wire [8-1:0] node3169;
	wire [8-1:0] node3171;
	wire [8-1:0] node3174;
	wire [8-1:0] node3175;
	wire [8-1:0] node3176;
	wire [8-1:0] node3177;
	wire [8-1:0] node3178;
	wire [8-1:0] node3182;
	wire [8-1:0] node3185;
	wire [8-1:0] node3186;
	wire [8-1:0] node3189;
	wire [8-1:0] node3192;
	wire [8-1:0] node3193;
	wire [8-1:0] node3195;
	wire [8-1:0] node3196;
	wire [8-1:0] node3200;
	wire [8-1:0] node3202;
	wire [8-1:0] node3205;
	wire [8-1:0] node3206;
	wire [8-1:0] node3207;
	wire [8-1:0] node3208;
	wire [8-1:0] node3211;
	wire [8-1:0] node3214;
	wire [8-1:0] node3215;
	wire [8-1:0] node3216;
	wire [8-1:0] node3220;
	wire [8-1:0] node3223;
	wire [8-1:0] node3224;
	wire [8-1:0] node3225;
	wire [8-1:0] node3229;
	wire [8-1:0] node3232;
	wire [8-1:0] node3233;
	wire [8-1:0] node3234;
	wire [8-1:0] node3235;
	wire [8-1:0] node3238;
	wire [8-1:0] node3239;
	wire [8-1:0] node3240;
	wire [8-1:0] node3241;
	wire [8-1:0] node3242;
	wire [8-1:0] node3243;
	wire [8-1:0] node3245;
	wire [8-1:0] node3249;
	wire [8-1:0] node3251;
	wire [8-1:0] node3254;
	wire [8-1:0] node3255;
	wire [8-1:0] node3256;
	wire [8-1:0] node3260;
	wire [8-1:0] node3263;
	wire [8-1:0] node3264;
	wire [8-1:0] node3265;
	wire [8-1:0] node3266;
	wire [8-1:0] node3269;
	wire [8-1:0] node3272;
	wire [8-1:0] node3274;
	wire [8-1:0] node3276;
	wire [8-1:0] node3279;
	wire [8-1:0] node3280;
	wire [8-1:0] node3282;
	wire [8-1:0] node3285;
	wire [8-1:0] node3286;
	wire [8-1:0] node3290;
	wire [8-1:0] node3291;
	wire [8-1:0] node3292;
	wire [8-1:0] node3293;
	wire [8-1:0] node3295;
	wire [8-1:0] node3297;
	wire [8-1:0] node3300;
	wire [8-1:0] node3301;
	wire [8-1:0] node3305;
	wire [8-1:0] node3306;
	wire [8-1:0] node3307;
	wire [8-1:0] node3308;
	wire [8-1:0] node3313;
	wire [8-1:0] node3314;
	wire [8-1:0] node3318;
	wire [8-1:0] node3319;
	wire [8-1:0] node3320;
	wire [8-1:0] node3322;
	wire [8-1:0] node3325;
	wire [8-1:0] node3326;
	wire [8-1:0] node3329;
	wire [8-1:0] node3332;
	wire [8-1:0] node3333;
	wire [8-1:0] node3334;
	wire [8-1:0] node3335;
	wire [8-1:0] node3338;
	wire [8-1:0] node3342;
	wire [8-1:0] node3344;
	wire [8-1:0] node3346;
	wire [8-1:0] node3349;
	wire [8-1:0] node3350;
	wire [8-1:0] node3351;
	wire [8-1:0] node3352;
	wire [8-1:0] node3353;
	wire [8-1:0] node3356;
	wire [8-1:0] node3357;
	wire [8-1:0] node3358;
	wire [8-1:0] node3363;
	wire [8-1:0] node3364;
	wire [8-1:0] node3365;
	wire [8-1:0] node3368;
	wire [8-1:0] node3370;
	wire [8-1:0] node3373;
	wire [8-1:0] node3376;
	wire [8-1:0] node3377;
	wire [8-1:0] node3378;
	wire [8-1:0] node3379;
	wire [8-1:0] node3380;
	wire [8-1:0] node3383;
	wire [8-1:0] node3386;
	wire [8-1:0] node3389;
	wire [8-1:0] node3391;
	wire [8-1:0] node3392;
	wire [8-1:0] node3396;
	wire [8-1:0] node3397;
	wire [8-1:0] node3398;
	wire [8-1:0] node3399;
	wire [8-1:0] node3402;
	wire [8-1:0] node3406;
	wire [8-1:0] node3407;
	wire [8-1:0] node3408;
	wire [8-1:0] node3410;
	wire [8-1:0] node3413;
	wire [8-1:0] node3414;
	wire [8-1:0] node3417;
	wire [8-1:0] node3421;
	wire [8-1:0] node3422;
	wire [8-1:0] node3423;
	wire [8-1:0] node3424;
	wire [8-1:0] node3425;
	wire [8-1:0] node3428;
	wire [8-1:0] node3430;
	wire [8-1:0] node3433;
	wire [8-1:0] node3436;
	wire [8-1:0] node3437;
	wire [8-1:0] node3438;
	wire [8-1:0] node3440;
	wire [8-1:0] node3443;
	wire [8-1:0] node3444;
	wire [8-1:0] node3448;
	wire [8-1:0] node3449;
	wire [8-1:0] node3450;
	wire [8-1:0] node3453;
	wire [8-1:0] node3454;
	wire [8-1:0] node3459;
	wire [8-1:0] node3460;
	wire [8-1:0] node3461;
	wire [8-1:0] node3462;
	wire [8-1:0] node3465;
	wire [8-1:0] node3466;
	wire [8-1:0] node3469;
	wire [8-1:0] node3471;
	wire [8-1:0] node3474;
	wire [8-1:0] node3477;
	wire [8-1:0] node3478;
	wire [8-1:0] node3479;
	wire [8-1:0] node3480;
	wire [8-1:0] node3481;
	wire [8-1:0] node3484;
	wire [8-1:0] node3487;
	wire [8-1:0] node3488;
	wire [8-1:0] node3493;
	wire [8-1:0] node3494;
	wire [8-1:0] node3495;
	wire [8-1:0] node3497;
	wire [8-1:0] node3499;
	wire [8-1:0] node3503;
	wire [8-1:0] node3504;
	wire [8-1:0] node3507;
	wire [8-1:0] node3508;
	wire [8-1:0] node3512;
	wire [8-1:0] node3513;
	wire [8-1:0] node3514;
	wire [8-1:0] node3516;
	wire [8-1:0] node3517;
	wire [8-1:0] node3518;
	wire [8-1:0] node3519;
	wire [8-1:0] node3521;
	wire [8-1:0] node3522;
	wire [8-1:0] node3524;
	wire [8-1:0] node3527;
	wire [8-1:0] node3530;
	wire [8-1:0] node3532;
	wire [8-1:0] node3535;
	wire [8-1:0] node3537;
	wire [8-1:0] node3540;
	wire [8-1:0] node3541;
	wire [8-1:0] node3542;
	wire [8-1:0] node3543;
	wire [8-1:0] node3545;
	wire [8-1:0] node3547;
	wire [8-1:0] node3550;
	wire [8-1:0] node3553;
	wire [8-1:0] node3554;
	wire [8-1:0] node3558;
	wire [8-1:0] node3559;
	wire [8-1:0] node3561;
	wire [8-1:0] node3564;
	wire [8-1:0] node3566;
	wire [8-1:0] node3568;
	wire [8-1:0] node3571;
	wire [8-1:0] node3572;
	wire [8-1:0] node3573;
	wire [8-1:0] node3574;
	wire [8-1:0] node3575;
	wire [8-1:0] node3577;
	wire [8-1:0] node3580;
	wire [8-1:0] node3583;
	wire [8-1:0] node3584;
	wire [8-1:0] node3587;
	wire [8-1:0] node3589;
	wire [8-1:0] node3590;
	wire [8-1:0] node3593;
	wire [8-1:0] node3596;
	wire [8-1:0] node3597;
	wire [8-1:0] node3598;
	wire [8-1:0] node3601;
	wire [8-1:0] node3604;
	wire [8-1:0] node3605;
	wire [8-1:0] node3608;
	wire [8-1:0] node3611;
	wire [8-1:0] node3612;
	wire [8-1:0] node3613;
	wire [8-1:0] node3614;
	wire [8-1:0] node3615;
	wire [8-1:0] node3619;
	wire [8-1:0] node3620;
	wire [8-1:0] node3622;
	wire [8-1:0] node3626;
	wire [8-1:0] node3627;
	wire [8-1:0] node3629;
	wire [8-1:0] node3631;
	wire [8-1:0] node3634;
	wire [8-1:0] node3635;
	wire [8-1:0] node3639;
	wire [8-1:0] node3640;
	wire [8-1:0] node3641;
	wire [8-1:0] node3644;
	wire [8-1:0] node3645;
	wire [8-1:0] node3647;
	wire [8-1:0] node3651;
	wire [8-1:0] node3652;
	wire [8-1:0] node3653;
	wire [8-1:0] node3655;
	wire [8-1:0] node3658;
	wire [8-1:0] node3659;
	wire [8-1:0] node3662;
	wire [8-1:0] node3664;
	wire [8-1:0] node3667;
	wire [8-1:0] node3670;
	wire [8-1:0] node3671;
	wire [8-1:0] node3673;
	wire [8-1:0] node3674;
	wire [8-1:0] node3675;
	wire [8-1:0] node3677;
	wire [8-1:0] node3679;
	wire [8-1:0] node3682;
	wire [8-1:0] node3683;
	wire [8-1:0] node3685;
	wire [8-1:0] node3687;
	wire [8-1:0] node3690;
	wire [8-1:0] node3692;
	wire [8-1:0] node3695;
	wire [8-1:0] node3696;
	wire [8-1:0] node3697;
	wire [8-1:0] node3698;
	wire [8-1:0] node3700;
	wire [8-1:0] node3702;
	wire [8-1:0] node3705;
	wire [8-1:0] node3708;
	wire [8-1:0] node3709;
	wire [8-1:0] node3711;
	wire [8-1:0] node3712;
	wire [8-1:0] node3716;
	wire [8-1:0] node3718;
	wire [8-1:0] node3721;
	wire [8-1:0] node3722;
	wire [8-1:0] node3724;
	wire [8-1:0] node3726;
	wire [8-1:0] node3729;
	wire [8-1:0] node3732;
	wire [8-1:0] node3733;
	wire [8-1:0] node3734;
	wire [8-1:0] node3735;
	wire [8-1:0] node3736;
	wire [8-1:0] node3739;
	wire [8-1:0] node3740;
	wire [8-1:0] node3743;
	wire [8-1:0] node3745;
	wire [8-1:0] node3748;
	wire [8-1:0] node3750;
	wire [8-1:0] node3751;
	wire [8-1:0] node3755;
	wire [8-1:0] node3756;
	wire [8-1:0] node3757;
	wire [8-1:0] node3758;
	wire [8-1:0] node3759;
	wire [8-1:0] node3763;
	wire [8-1:0] node3764;
	wire [8-1:0] node3768;
	wire [8-1:0] node3769;
	wire [8-1:0] node3770;
	wire [8-1:0] node3773;
	wire [8-1:0] node3776;
	wire [8-1:0] node3777;
	wire [8-1:0] node3781;
	wire [8-1:0] node3782;
	wire [8-1:0] node3785;
	wire [8-1:0] node3788;
	wire [8-1:0] node3789;
	wire [8-1:0] node3790;
	wire [8-1:0] node3791;
	wire [8-1:0] node3792;
	wire [8-1:0] node3796;
	wire [8-1:0] node3797;
	wire [8-1:0] node3800;
	wire [8-1:0] node3803;
	wire [8-1:0] node3804;
	wire [8-1:0] node3807;
	wire [8-1:0] node3810;
	wire [8-1:0] node3811;
	wire [8-1:0] node3812;
	wire [8-1:0] node3813;
	wire [8-1:0] node3814;
	wire [8-1:0] node3816;
	wire [8-1:0] node3820;
	wire [8-1:0] node3821;
	wire [8-1:0] node3824;
	wire [8-1:0] node3827;
	wire [8-1:0] node3828;
	wire [8-1:0] node3830;
	wire [8-1:0] node3831;
	wire [8-1:0] node3835;
	wire [8-1:0] node3836;
	wire [8-1:0] node3839;
	wire [8-1:0] node3841;
	wire [8-1:0] node3844;
	wire [8-1:0] node3845;
	wire [8-1:0] node3848;

	assign outp = (inp[7]) ? node1952 : node1;
		assign node1 = (inp[13]) ? node933 : node2;
			assign node2 = (inp[4]) ? node288 : node3;
				assign node3 = (inp[11]) ? node109 : node4;
					assign node4 = (inp[0]) ? node68 : node5;
						assign node5 = (inp[2]) ? node31 : node6;
							assign node6 = (inp[8]) ? node14 : node7;
								assign node7 = (inp[1]) ? node9 : 8'b01111111;
									assign node9 = (inp[3]) ? node11 : 8'b00111110;
										assign node11 = (inp[10]) ? 8'b01111111 : 8'b00111110;
								assign node14 = (inp[1]) ? node22 : node15;
									assign node15 = (inp[12]) ? 8'b00111011 : node16;
										assign node16 = (inp[9]) ? node18 : 8'b00111011;
											assign node18 = (inp[10]) ? 8'b01111111 : 8'b00111011;
									assign node22 = (inp[5]) ? node24 : 8'b00111010;
										assign node24 = (inp[10]) ? node28 : node25;
											assign node25 = (inp[3]) ? 8'b00111011 : 8'b00111010;
											assign node28 = (inp[3]) ? 8'b01111111 : 8'b00111110;
							assign node31 = (inp[1]) ? node49 : node32;
								assign node32 = (inp[8]) ? node38 : node33;
									assign node33 = (inp[5]) ? node35 : 8'b00101111;
										assign node35 = (inp[6]) ? 8'b01111111 : 8'b00101111;
									assign node38 = (inp[6]) ? node44 : node39;
										assign node39 = (inp[10]) ? node41 : 8'b00101011;
											assign node41 = (inp[5]) ? 8'b00101111 : 8'b00101011;
										assign node44 = (inp[5]) ? node46 : 8'b00101011;
											assign node46 = (inp[10]) ? 8'b01111111 : 8'b00111011;
								assign node49 = (inp[5]) ? node53 : node50;
									assign node50 = (inp[8]) ? 8'b00101010 : 8'b00101110;
									assign node53 = (inp[6]) ? node65 : node54;
										assign node54 = (inp[3]) ? node60 : node55;
											assign node55 = (inp[9]) ? 8'b00101110 : node56;
												assign node56 = (inp[10]) ? 8'b00101110 : 8'b00101010;
											assign node60 = (inp[10]) ? 8'b00101111 : node61;
												assign node61 = (inp[12]) ? 8'b00101011 : 8'b00101111;
										assign node65 = (inp[3]) ? 8'b01111111 : 8'b00111110;
						assign node68 = (inp[5]) ? 8'b01111111 : node69;
							assign node69 = (inp[6]) ? node87 : node70;
								assign node70 = (inp[8]) ? node76 : node71;
									assign node71 = (inp[1]) ? node73 : 8'b01111111;
										assign node73 = (inp[3]) ? 8'b00111110 : 8'b01111111;
									assign node76 = (inp[10]) ? node82 : node77;
										assign node77 = (inp[3]) ? node79 : 8'b01111111;
											assign node79 = (inp[1]) ? 8'b00111110 : 8'b01111111;
										assign node82 = (inp[1]) ? node84 : 8'b00111011;
											assign node84 = (inp[9]) ? 8'b00111011 : 8'b00111010;
								assign node87 = (inp[2]) ? node97 : node88;
									assign node88 = (inp[3]) ? node90 : 8'b01111111;
										assign node90 = (inp[1]) ? node94 : node91;
											assign node91 = (inp[9]) ? 8'b01111111 : 8'b00111011;
											assign node94 = (inp[9]) ? 8'b00111110 : 8'b00111010;
									assign node97 = (inp[1]) ? node103 : node98;
										assign node98 = (inp[8]) ? node100 : 8'b00101111;
											assign node100 = (inp[10]) ? 8'b00101011 : 8'b00101111;
										assign node103 = (inp[3]) ? 8'b00101110 : node104;
											assign node104 = (inp[8]) ? 8'b00101011 : 8'b00101111;
					assign node109 = (inp[8]) ? node177 : node110;
						assign node110 = (inp[1]) ? node128 : node111;
							assign node111 = (inp[2]) ? node115 : node112;
								assign node112 = (inp[12]) ? 8'b01111111 : 8'b00101111;
								assign node115 = (inp[12]) ? node121 : node116;
									assign node116 = (inp[0]) ? node118 : 8'b00111110;
										assign node118 = (inp[5]) ? 8'b00101110 : 8'b00111110;
									assign node121 = (inp[6]) ? node125 : node122;
										assign node122 = (inp[0]) ? 8'b00111110 : 8'b00101111;
										assign node125 = (inp[5]) ? 8'b00111110 : 8'b00101111;
							assign node128 = (inp[0]) ? node154 : node129;
								assign node129 = (inp[2]) ? node139 : node130;
									assign node130 = (inp[12]) ? node136 : node131;
										assign node131 = (inp[5]) ? node133 : 8'b00101110;
											assign node133 = (inp[3]) ? 8'b00101011 : 8'b00101110;
										assign node136 = (inp[9]) ? 8'b00111011 : 8'b00111110;
									assign node139 = (inp[12]) ? node147 : node140;
										assign node140 = (inp[5]) ? node142 : 8'b00111011;
											assign node142 = (inp[6]) ? node144 : 8'b00111010;
												assign node144 = (inp[3]) ? 8'b00101010 : 8'b00101011;
										assign node147 = (inp[9]) ? 8'b00101110 : node148;
											assign node148 = (inp[6]) ? 8'b00111011 : node149;
												assign node149 = (inp[3]) ? 8'b00101011 : 8'b00101110;
								assign node154 = (inp[12]) ? node166 : node155;
									assign node155 = (inp[2]) ? node161 : node156;
										assign node156 = (inp[3]) ? node158 : 8'b00101011;
											assign node158 = (inp[5]) ? 8'b00101011 : 8'b00101110;
										assign node161 = (inp[6]) ? node163 : 8'b00101010;
											assign node163 = (inp[3]) ? 8'b00111011 : 8'b00101010;
									assign node166 = (inp[2]) ? node172 : node167;
										assign node167 = (inp[3]) ? node169 : 8'b00111011;
											assign node169 = (inp[5]) ? 8'b00111011 : 8'b00111110;
										assign node172 = (inp[5]) ? 8'b00111010 : node173;
											assign node173 = (inp[6]) ? 8'b00101011 : 8'b00111010;
						assign node177 = (inp[5]) ? node231 : node178;
							assign node178 = (inp[2]) ? node196 : node179;
								assign node179 = (inp[12]) ? node189 : node180;
									assign node180 = (inp[1]) ? node182 : 8'b00101011;
										assign node182 = (inp[3]) ? 8'b00101010 : node183;
											assign node183 = (inp[0]) ? node185 : 8'b00101010;
												assign node185 = (inp[10]) ? 8'b00001111 : 8'b00001011;
									assign node189 = (inp[1]) ? 8'b00111010 : node190;
										assign node190 = (inp[3]) ? 8'b00111011 : node191;
											assign node191 = (inp[10]) ? 8'b00111011 : 8'b00011111;
								assign node196 = (inp[12]) ? node212 : node197;
									assign node197 = (inp[1]) ? node207 : node198;
										assign node198 = (inp[10]) ? node202 : node199;
											assign node199 = (inp[9]) ? 8'b00001110 : 8'b00011110;
											assign node202 = (inp[3]) ? node204 : 8'b00111010;
												assign node204 = (inp[6]) ? 8'b00111010 : 8'b00101010;
										assign node207 = (inp[0]) ? node209 : 8'b00011111;
											assign node209 = (inp[3]) ? 8'b00001111 : 8'b00011010;
									assign node212 = (inp[0]) ? node216 : node213;
										assign node213 = (inp[1]) ? 8'b00101010 : 8'b00101011;
										assign node216 = (inp[6]) ? node224 : node217;
											assign node217 = (inp[3]) ? 8'b00011111 : node218;
												assign node218 = (inp[10]) ? 8'b00111010 : node219;
													assign node219 = (inp[1]) ? 8'b00011010 : 8'b00011110;
											assign node224 = (inp[10]) ? node226 : 8'b00001111;
												assign node226 = (inp[3]) ? 8'b00101010 : node227;
													assign node227 = (inp[1]) ? 8'b00001111 : 8'b00101011;
							assign node231 = (inp[2]) ? node259 : node232;
								assign node232 = (inp[12]) ? node244 : node233;
									assign node233 = (inp[1]) ? node239 : node234;
										assign node234 = (inp[0]) ? 8'b00001111 : node235;
											assign node235 = (inp[6]) ? 8'b00101011 : 8'b00001111;
										assign node239 = (inp[3]) ? node241 : 8'b00001110;
											assign node241 = (inp[10]) ? 8'b00001011 : 8'b00001111;
									assign node244 = (inp[10]) ? node256 : node245;
										assign node245 = (inp[3]) ? node251 : node246;
											assign node246 = (inp[0]) ? 8'b00011011 : node247;
												assign node247 = (inp[1]) ? 8'b00111010 : 8'b00111011;
											assign node251 = (inp[9]) ? node253 : 8'b00011111;
												assign node253 = (inp[0]) ? 8'b00011011 : 8'b00011111;
										assign node256 = (inp[1]) ? 8'b00011110 : 8'b00011111;
								assign node259 = (inp[1]) ? node269 : node260;
									assign node260 = (inp[0]) ? node266 : node261;
										assign node261 = (inp[10]) ? 8'b00011110 : node262;
											assign node262 = (inp[6]) ? 8'b00101010 : 8'b00111010;
										assign node266 = (inp[12]) ? 8'b00011110 : 8'b00001110;
									assign node269 = (inp[0]) ? node285 : node270;
										assign node270 = (inp[10]) ? node282 : node271;
											assign node271 = (inp[9]) ? node277 : node272;
												assign node272 = (inp[3]) ? node274 : 8'b00101010;
													assign node274 = (inp[6]) ? 8'b00011110 : 8'b00001111;
												assign node277 = (inp[6]) ? node279 : 8'b00011111;
													assign node279 = (inp[3]) ? 8'b00001110 : 8'b00001111;
											assign node282 = (inp[6]) ? 8'b00001011 : 8'b00011010;
										assign node285 = (inp[12]) ? 8'b00011010 : 8'b00001010;
				assign node288 = (inp[9]) ? node592 : node289;
					assign node289 = (inp[8]) ? node435 : node290;
						assign node290 = (inp[10]) ? node364 : node291;
							assign node291 = (inp[11]) ? node329 : node292;
								assign node292 = (inp[2]) ? node308 : node293;
									assign node293 = (inp[6]) ? node299 : node294;
										assign node294 = (inp[3]) ? 8'b00001011 : node295;
											assign node295 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node299 = (inp[12]) ? node301 : 8'b00011010;
											assign node301 = (inp[1]) ? node303 : 8'b00011011;
												assign node303 = (inp[5]) ? 8'b10011001 : node304;
													assign node304 = (inp[0]) ? 8'b00011000 : 8'b00011010;
									assign node308 = (inp[0]) ? node320 : node309;
										assign node309 = (inp[5]) ? node311 : 8'b00000010;
											assign node311 = (inp[12]) ? node315 : node312;
												assign node312 = (inp[3]) ? 8'b10000001 : 8'b10000010;
												assign node315 = (inp[3]) ? node317 : 8'b10010000;
													assign node317 = (inp[1]) ? 8'b10010001 : 8'b00011011;
										assign node320 = (inp[3]) ? node324 : node321;
											assign node321 = (inp[1]) ? 8'b10010001 : 8'b10010000;
											assign node324 = (inp[1]) ? node326 : 8'b00011011;
												assign node326 = (inp[6]) ? 8'b10000010 : 8'b10010000;
								assign node329 = (inp[3]) ? node347 : node330;
									assign node330 = (inp[0]) ? node338 : node331;
										assign node331 = (inp[1]) ? node335 : node332;
											assign node332 = (inp[6]) ? 8'b00000010 : 8'b11110111;
											assign node335 = (inp[2]) ? 8'b00000010 : 8'b00001010;
										assign node338 = (inp[1]) ? node344 : node339;
											assign node339 = (inp[5]) ? node341 : 8'b00000010;
												assign node341 = (inp[2]) ? 8'b10100101 : 8'b11110111;
											assign node344 = (inp[2]) ? 8'b10100100 : 8'b10100101;
									assign node347 = (inp[1]) ? node355 : node348;
										assign node348 = (inp[12]) ? 8'b00001011 : node349;
											assign node349 = (inp[6]) ? 8'b00001011 : node350;
												assign node350 = (inp[2]) ? 8'b00001010 : 8'b00011010;
										assign node355 = (inp[6]) ? node361 : node356;
											assign node356 = (inp[12]) ? 8'b00000010 : node357;
												assign node357 = (inp[5]) ? 8'b10110100 : 8'b11110111;
											assign node361 = (inp[0]) ? 8'b00000010 : 8'b00001010;
							assign node364 = (inp[11]) ? node390 : node365;
								assign node365 = (inp[5]) ? node385 : node366;
									assign node366 = (inp[2]) ? node376 : node367;
										assign node367 = (inp[6]) ? node371 : node368;
											assign node368 = (inp[3]) ? 8'b00001111 : 8'b00001110;
											assign node371 = (inp[1]) ? 8'b00011110 : node372;
												assign node372 = (inp[0]) ? 8'b00011110 : 8'b00011111;
										assign node376 = (inp[0]) ? node380 : node377;
											assign node377 = (inp[1]) ? 8'b00001110 : 8'b00001111;
											assign node380 = (inp[6]) ? 8'b00001111 : node381;
												assign node381 = (inp[1]) ? 8'b00011111 : 8'b00011110;
									assign node385 = (inp[3]) ? 8'b00011111 : node386;
										assign node386 = (inp[1]) ? 8'b00011111 : 8'b00011110;
								assign node390 = (inp[1]) ? node406 : node391;
									assign node391 = (inp[3]) ? node399 : node392;
										assign node392 = (inp[12]) ? 8'b00001110 : node393;
											assign node393 = (inp[2]) ? node395 : 8'b00001110;
												assign node395 = (inp[0]) ? 8'b00001011 : 8'b00011011;
										assign node399 = (inp[5]) ? node401 : 8'b00001111;
											assign node401 = (inp[6]) ? node403 : 8'b00011110;
												assign node403 = (inp[12]) ? 8'b00011110 : 8'b00001110;
									assign node406 = (inp[0]) ? node422 : node407;
										assign node407 = (inp[12]) ? node411 : node408;
											assign node408 = (inp[6]) ? 8'b00001011 : 8'b00011011;
											assign node411 = (inp[6]) ? node417 : node412;
												assign node412 = (inp[5]) ? node414 : 8'b00001110;
													assign node414 = (inp[3]) ? 8'b00001011 : 8'b00001110;
												assign node417 = (inp[3]) ? node419 : 8'b00011110;
													assign node419 = (inp[2]) ? 8'b00011010 : 8'b00011011;
										assign node422 = (inp[12]) ? node426 : node423;
											assign node423 = (inp[2]) ? 8'b00001010 : 8'b00001011;
											assign node426 = (inp[3]) ? node430 : node427;
												assign node427 = (inp[5]) ? 8'b00011011 : 8'b00001011;
												assign node430 = (inp[2]) ? 8'b00011011 : node431;
													assign node431 = (inp[6]) ? 8'b00011011 : 8'b00001011;
						assign node435 = (inp[5]) ? node505 : node436;
							assign node436 = (inp[0]) ? node464 : node437;
								assign node437 = (inp[1]) ? node453 : node438;
									assign node438 = (inp[3]) ? node448 : node439;
										assign node439 = (inp[6]) ? node445 : node440;
											assign node440 = (inp[12]) ? 8'b00000010 : node441;
												assign node441 = (inp[10]) ? 8'b10000010 : 8'b11110111;
											assign node445 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node448 = (inp[11]) ? 8'b00011010 : node449;
											assign node449 = (inp[6]) ? 8'b00011011 : 8'b00001011;
									assign node453 = (inp[12]) ? node459 : node454;
										assign node454 = (inp[11]) ? node456 : 8'b10000010;
											assign node456 = (inp[2]) ? 8'b11110111 : 8'b00001010;
										assign node459 = (inp[2]) ? 8'b00000010 : node460;
											assign node460 = (inp[6]) ? 8'b00011010 : 8'b00000010;
								assign node464 = (inp[10]) ? node486 : node465;
									assign node465 = (inp[11]) ? node479 : node466;
										assign node466 = (inp[2]) ? node472 : node467;
											assign node467 = (inp[6]) ? node469 : 8'b10000100;
												assign node469 = (inp[12]) ? 8'b10011101 : 8'b10011100;
											assign node472 = (inp[6]) ? node474 : 8'b10010100;
												assign node474 = (inp[12]) ? 8'b10000100 : node475;
													assign node475 = (inp[1]) ? 8'b10000101 : 8'b10000100;
										assign node479 = (inp[1]) ? node483 : node480;
											assign node480 = (inp[6]) ? 8'b10101100 : 8'b10101101;
											assign node483 = (inp[2]) ? 8'b10100000 : 8'b10110000;
									assign node486 = (inp[11]) ? node498 : node487;
										assign node487 = (inp[3]) ? node493 : node488;
											assign node488 = (inp[2]) ? 8'b10010000 : node489;
												assign node489 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node493 = (inp[1]) ? 8'b00000010 : node494;
												assign node494 = (inp[12]) ? 8'b00011011 : 8'b00001011;
										assign node498 = (inp[12]) ? 8'b00001011 : node499;
											assign node499 = (inp[2]) ? node501 : 8'b10101101;
												assign node501 = (inp[6]) ? 8'b11110111 : 8'b10100101;
							assign node505 = (inp[11]) ? node541 : node506;
								assign node506 = (inp[3]) ? node522 : node507;
									assign node507 = (inp[6]) ? node511 : node508;
										assign node508 = (inp[2]) ? 8'b10010100 : 8'b10000100;
										assign node511 = (inp[2]) ? node519 : node512;
											assign node512 = (inp[12]) ? node516 : node513;
												assign node513 = (inp[0]) ? 8'b10011101 : 8'b10011100;
												assign node516 = (inp[0]) ? 8'b10011100 : 8'b00011010;
											assign node519 = (inp[0]) ? 8'b10010100 : 8'b10010000;
									assign node522 = (inp[6]) ? node532 : node523;
										assign node523 = (inp[0]) ? node527 : node524;
											assign node524 = (inp[10]) ? 8'b10000101 : 8'b10000001;
											assign node527 = (inp[1]) ? node529 : 8'b10011101;
												assign node529 = (inp[2]) ? 8'b10010101 : 8'b10000101;
										assign node532 = (inp[10]) ? node538 : node533;
											assign node533 = (inp[2]) ? 8'b00011011 : node534;
												assign node534 = (inp[12]) ? 8'b10011001 : 8'b10011101;
											assign node538 = (inp[2]) ? 8'b10010101 : 8'b10011101;
								assign node541 = (inp[3]) ? node565 : node542;
									assign node542 = (inp[12]) ? node550 : node543;
										assign node543 = (inp[2]) ? node547 : node544;
											assign node544 = (inp[6]) ? 8'b10101001 : 8'b10110001;
											assign node547 = (inp[1]) ? 8'b10100000 : 8'b10100001;
										assign node550 = (inp[6]) ? node556 : node551;
											assign node551 = (inp[10]) ? 8'b10100100 : node552;
												assign node552 = (inp[2]) ? 8'b10110001 : 8'b10100001;
											assign node556 = (inp[2]) ? node562 : node557;
												assign node557 = (inp[0]) ? node559 : 8'b00011010;
													assign node559 = (inp[1]) ? 8'b10111001 : 8'b10111100;
												assign node562 = (inp[0]) ? 8'b10110000 : 8'b11110101;
									assign node565 = (inp[1]) ? node583 : node566;
										assign node566 = (inp[10]) ? node576 : node567;
											assign node567 = (inp[0]) ? node573 : node568;
												assign node568 = (inp[12]) ? node570 : 8'b00011010;
													assign node570 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node573 = (inp[12]) ? 8'b10101101 : 8'b10101100;
											assign node576 = (inp[0]) ? 8'b10111100 : node577;
												assign node577 = (inp[6]) ? node579 : 8'b10101101;
													assign node579 = (inp[2]) ? 8'b10111100 : 8'b11111101;
										assign node583 = (inp[12]) ? node585 : 8'b10110100;
											assign node585 = (inp[0]) ? node589 : node586;
												assign node586 = (inp[10]) ? 8'b10100001 : 8'b10100101;
												assign node589 = (inp[2]) ? 8'b10110000 : 8'b10111001;
					assign node592 = (inp[11]) ? node724 : node593;
						assign node593 = (inp[3]) ? node661 : node594;
							assign node594 = (inp[0]) ? node610 : node595;
								assign node595 = (inp[6]) ? node603 : node596;
									assign node596 = (inp[10]) ? node598 : 8'b00101010;
										assign node598 = (inp[5]) ? 8'b00101110 : node599;
											assign node599 = (inp[8]) ? 8'b00101010 : 8'b00101110;
									assign node603 = (inp[2]) ? node607 : node604;
										assign node604 = (inp[5]) ? 8'b00111110 : 8'b00111010;
										assign node607 = (inp[5]) ? 8'b00111010 : 8'b00101010;
								assign node610 = (inp[1]) ? node640 : node611;
									assign node611 = (inp[6]) ? node623 : node612;
										assign node612 = (inp[2]) ? 8'b00111010 : node613;
											assign node613 = (inp[12]) ? node615 : 8'b00101110;
												assign node615 = (inp[10]) ? node619 : node616;
													assign node616 = (inp[8]) ? 8'b00101110 : 8'b00101010;
													assign node619 = (inp[8]) ? 8'b00101010 : 8'b00101110;
										assign node623 = (inp[2]) ? node635 : node624;
											assign node624 = (inp[5]) ? node630 : node625;
												assign node625 = (inp[8]) ? node627 : 8'b00111110;
													assign node627 = (inp[10]) ? 8'b00111010 : 8'b00111110;
												assign node630 = (inp[10]) ? 8'b00111110 : node631;
													assign node631 = (inp[8]) ? 8'b00111110 : 8'b00111010;
											assign node635 = (inp[12]) ? 8'b00111110 : node636;
												assign node636 = (inp[8]) ? 8'b00101010 : 8'b00101110;
									assign node640 = (inp[12]) ? node646 : node641;
										assign node641 = (inp[5]) ? 8'b01111111 : node642;
											assign node642 = (inp[10]) ? 8'b00101111 : 8'b01111111;
										assign node646 = (inp[6]) ? node654 : node647;
											assign node647 = (inp[2]) ? 8'b00111011 : node648;
												assign node648 = (inp[10]) ? 8'b00101111 : node649;
													assign node649 = (inp[8]) ? 8'b00101111 : 8'b00101011;
											assign node654 = (inp[10]) ? 8'b01111111 : node655;
												assign node655 = (inp[5]) ? 8'b00111011 : node656;
													assign node656 = (inp[2]) ? 8'b00101011 : 8'b00111011;
							assign node661 = (inp[1]) ? node693 : node662;
								assign node662 = (inp[10]) ? node676 : node663;
									assign node663 = (inp[8]) ? node671 : node664;
										assign node664 = (inp[5]) ? node666 : 8'b00101011;
											assign node666 = (inp[6]) ? 8'b00111011 : node667;
												assign node667 = (inp[2]) ? 8'b00111011 : 8'b00101011;
										assign node671 = (inp[0]) ? 8'b01111111 : node672;
											assign node672 = (inp[6]) ? 8'b00111011 : 8'b00101011;
									assign node676 = (inp[5]) ? node688 : node677;
										assign node677 = (inp[8]) ? node685 : node678;
											assign node678 = (inp[0]) ? node680 : 8'b01111111;
												assign node680 = (inp[12]) ? node682 : 8'b00101111;
													assign node682 = (inp[6]) ? 8'b00101111 : 8'b00101111;
											assign node685 = (inp[6]) ? 8'b00101011 : 8'b00111011;
										assign node688 = (inp[12]) ? node690 : 8'b01111111;
											assign node690 = (inp[0]) ? 8'b01111111 : 8'b00101111;
								assign node693 = (inp[5]) ? node709 : node694;
									assign node694 = (inp[12]) ? node700 : node695;
										assign node695 = (inp[2]) ? node697 : 8'b00111110;
											assign node697 = (inp[10]) ? 8'b00101010 : 8'b00111010;
										assign node700 = (inp[0]) ? 8'b00101110 : node701;
											assign node701 = (inp[10]) ? node703 : 8'b00101010;
												assign node703 = (inp[8]) ? 8'b00101010 : node704;
													assign node704 = (inp[6]) ? 8'b00111110 : 8'b00101110;
									assign node709 = (inp[6]) ? node719 : node710;
										assign node710 = (inp[10]) ? 8'b00101111 : node711;
											assign node711 = (inp[8]) ? node715 : node712;
												assign node712 = (inp[2]) ? 8'b00111011 : 8'b00101011;
												assign node715 = (inp[2]) ? 8'b00101011 : 8'b00101111;
										assign node719 = (inp[10]) ? 8'b01111111 : node720;
											assign node720 = (inp[8]) ? 8'b01111111 : 8'b00111011;
						assign node724 = (inp[8]) ? node824 : node725;
							assign node725 = (inp[10]) ? node773 : node726;
								assign node726 = (inp[1]) ? node746 : node727;
									assign node727 = (inp[3]) ? node737 : node728;
										assign node728 = (inp[2]) ? node730 : 8'b00101010;
											assign node730 = (inp[0]) ? node732 : 8'b00101010;
												assign node732 = (inp[6]) ? node734 : 8'b00011111;
													assign node734 = (inp[5]) ? 8'b00001111 : 8'b00011111;
										assign node737 = (inp[2]) ? node743 : node738;
											assign node738 = (inp[12]) ? node740 : 8'b00101011;
												assign node740 = (inp[6]) ? 8'b00111011 : 8'b00101011;
											assign node743 = (inp[6]) ? 8'b00101010 : 8'b00101011;
									assign node746 = (inp[5]) ? node762 : node747;
										assign node747 = (inp[0]) ? node755 : node748;
											assign node748 = (inp[3]) ? node750 : 8'b00101010;
												assign node750 = (inp[2]) ? 8'b00101010 : node751;
													assign node751 = (inp[6]) ? 8'b00111010 : 8'b00101010;
											assign node755 = (inp[12]) ? 8'b00111010 : node756;
												assign node756 = (inp[2]) ? 8'b00001110 : node757;
													assign node757 = (inp[3]) ? 8'b00011111 : 8'b00011110;
										assign node762 = (inp[2]) ? node768 : node763;
											assign node763 = (inp[3]) ? 8'b00001111 : node764;
												assign node764 = (inp[0]) ? 8'b00001111 : 8'b00101010;
											assign node768 = (inp[6]) ? 8'b00011110 : node769;
												assign node769 = (inp[0]) ? 8'b00001110 : 8'b00001111;
								assign node773 = (inp[2]) ? node801 : node774;
									assign node774 = (inp[0]) ? node786 : node775;
										assign node775 = (inp[1]) ? node781 : node776;
											assign node776 = (inp[6]) ? node778 : 8'b00111110;
												assign node778 = (inp[12]) ? 8'b01111111 : 8'b00101111;
											assign node781 = (inp[6]) ? node783 : 8'b00101110;
												assign node783 = (inp[12]) ? 8'b00111110 : 8'b00101110;
										assign node786 = (inp[1]) ? node798 : node787;
											assign node787 = (inp[3]) ? node793 : node788;
												assign node788 = (inp[12]) ? node790 : 8'b00101110;
													assign node790 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node793 = (inp[6]) ? 8'b00101111 : node794;
													assign node794 = (inp[12]) ? 8'b00101111 : 8'b00111110;
											assign node798 = (inp[12]) ? 8'b00111011 : 8'b00101011;
									assign node801 = (inp[5]) ? node811 : node802;
										assign node802 = (inp[0]) ? node806 : node803;
											assign node803 = (inp[12]) ? 8'b00101110 : 8'b00111110;
											assign node806 = (inp[6]) ? node808 : 8'b00111011;
												assign node808 = (inp[3]) ? 8'b00101111 : 8'b00101110;
										assign node811 = (inp[3]) ? node819 : node812;
											assign node812 = (inp[0]) ? node814 : 8'b00111011;
												assign node814 = (inp[1]) ? 8'b00101010 : node815;
													assign node815 = (inp[12]) ? 8'b00111011 : 8'b00101011;
											assign node819 = (inp[6]) ? node821 : 8'b00111110;
												assign node821 = (inp[12]) ? 8'b00111010 : 8'b00101010;
							assign node824 = (inp[5]) ? node876 : node825;
								assign node825 = (inp[0]) ? node845 : node826;
									assign node826 = (inp[6]) ? node834 : node827;
										assign node827 = (inp[3]) ? node829 : 8'b00011111;
											assign node829 = (inp[12]) ? node831 : 8'b00111010;
												assign node831 = (inp[1]) ? 8'b00101010 : 8'b00101011;
										assign node834 = (inp[2]) ? node842 : node835;
											assign node835 = (inp[12]) ? 8'b00111010 : node836;
												assign node836 = (inp[10]) ? node838 : 8'b00101010;
													assign node838 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node842 = (inp[3]) ? 8'b00101011 : 8'b00101010;
									assign node845 = (inp[12]) ? node867 : node846;
										assign node846 = (inp[10]) ? node854 : node847;
											assign node847 = (inp[2]) ? 8'b00011011 : node848;
												assign node848 = (inp[6]) ? 8'b00001110 : node849;
													assign node849 = (inp[3]) ? 8'b00011110 : 8'b00011010;
											assign node854 = (inp[3]) ? node862 : node855;
												assign node855 = (inp[6]) ? node859 : node856;
													assign node856 = (inp[1]) ? 8'b00001110 : 8'b00001111;
													assign node859 = (inp[2]) ? 8'b00011111 : 8'b00001111;
												assign node862 = (inp[6]) ? node864 : 8'b00011111;
													assign node864 = (inp[2]) ? 8'b00011010 : 8'b00101010;
										assign node867 = (inp[10]) ? node869 : 8'b00001111;
											assign node869 = (inp[1]) ? 8'b00001111 : node870;
												assign node870 = (inp[3]) ? node872 : 8'b00101010;
													assign node872 = (inp[2]) ? 8'b00101011 : 8'b00111011;
								assign node876 = (inp[2]) ? node900 : node877;
									assign node877 = (inp[1]) ? node889 : node878;
										assign node878 = (inp[10]) ? node880 : 8'b00101010;
											assign node880 = (inp[3]) ? node886 : node881;
												assign node881 = (inp[6]) ? 8'b00001110 : node882;
													assign node882 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node886 = (inp[6]) ? 8'b00011111 : 8'b00001111;
										assign node889 = (inp[12]) ? 8'b00001011 : node890;
											assign node890 = (inp[6]) ? node896 : node891;
												assign node891 = (inp[3]) ? node893 : 8'b00011111;
													assign node893 = (inp[0]) ? 8'b00011010 : 8'b00011110;
												assign node896 = (inp[10]) ? 8'b00001011 : 8'b00001111;
									assign node900 = (inp[3]) ? node918 : node901;
										assign node901 = (inp[0]) ? node911 : node902;
											assign node902 = (inp[12]) ? node908 : node903;
												assign node903 = (inp[6]) ? 8'b00001111 : node904;
													assign node904 = (inp[1]) ? 8'b00011111 : 8'b00011011;
												assign node908 = (inp[6]) ? 8'b00011011 : 8'b00001110;
											assign node911 = (inp[10]) ? node915 : node912;
												assign node912 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node915 = (inp[12]) ? 8'b00011011 : 8'b00001011;
										assign node918 = (inp[12]) ? node928 : node919;
											assign node919 = (inp[6]) ? node921 : 8'b00011010;
												assign node921 = (inp[1]) ? node925 : node922;
													assign node922 = (inp[0]) ? 8'b00001110 : 8'b00101010;
													assign node925 = (inp[0]) ? 8'b00001010 : 8'b00001010;
											assign node928 = (inp[0]) ? 8'b00011110 : node929;
												assign node929 = (inp[1]) ? 8'b00011110 : 8'b00111010;
			assign node933 = (inp[0]) ? node1411 : node934;
				assign node934 = (inp[5]) ? node1074 : node935;
					assign node935 = (inp[8]) ? node1017 : node936;
						assign node936 = (inp[4]) ? node956 : node937;
							assign node937 = (inp[1]) ? node945 : node938;
								assign node938 = (inp[2]) ? node940 : 8'b00011111;
									assign node940 = (inp[12]) ? 8'b00001111 : node941;
										assign node941 = (inp[11]) ? 8'b00011110 : 8'b00001111;
								assign node945 = (inp[2]) ? node951 : node946;
									assign node946 = (inp[12]) ? 8'b00011110 : node947;
										assign node947 = (inp[6]) ? 8'b00001110 : 8'b00011110;
									assign node951 = (inp[12]) ? 8'b00001110 : node952;
										assign node952 = (inp[11]) ? 8'b00011011 : 8'b00001110;
							assign node956 = (inp[10]) ? node986 : node957;
								assign node957 = (inp[12]) ? node973 : node958;
									assign node958 = (inp[2]) ? node970 : node959;
										assign node959 = (inp[3]) ? node963 : node960;
											assign node960 = (inp[6]) ? 8'b00001010 : 8'b11110111;
											assign node963 = (inp[6]) ? node967 : node964;
												assign node964 = (inp[11]) ? 8'b00011010 : 8'b00001011;
												assign node967 = (inp[11]) ? 8'b00001011 : 8'b00011011;
										assign node970 = (inp[11]) ? 8'b11110111 : 8'b10000010;
									assign node973 = (inp[3]) ? node979 : node974;
										assign node974 = (inp[2]) ? 8'b00000010 : node975;
											assign node975 = (inp[6]) ? 8'b00011010 : 8'b00000010;
										assign node979 = (inp[1]) ? node983 : node980;
											assign node980 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node983 = (inp[6]) ? 8'b00011010 : 8'b00000010;
								assign node986 = (inp[12]) ? node1004 : node987;
									assign node987 = (inp[11]) ? node993 : node988;
										assign node988 = (inp[3]) ? 8'b00001111 : node989;
											assign node989 = (inp[1]) ? 8'b00011110 : 8'b00001110;
										assign node993 = (inp[3]) ? node999 : node994;
											assign node994 = (inp[6]) ? node996 : 8'b00011011;
												assign node996 = (inp[2]) ? 8'b00011011 : 8'b00001110;
											assign node999 = (inp[1]) ? node1001 : 8'b00011110;
												assign node1001 = (inp[2]) ? 8'b00011011 : 8'b00001110;
									assign node1004 = (inp[3]) ? node1010 : node1005;
										assign node1005 = (inp[6]) ? node1007 : 8'b00001110;
											assign node1007 = (inp[9]) ? 8'b00001110 : 8'b00011110;
										assign node1010 = (inp[1]) ? 8'b00001110 : node1011;
											assign node1011 = (inp[6]) ? node1013 : 8'b00001111;
												assign node1013 = (inp[2]) ? 8'b00001111 : 8'b00011111;
						assign node1017 = (inp[1]) ? node1053 : node1018;
							assign node1018 = (inp[4]) ? node1030 : node1019;
								assign node1019 = (inp[2]) ? node1025 : node1020;
									assign node1020 = (inp[12]) ? 8'b00011011 : node1021;
										assign node1021 = (inp[11]) ? 8'b00001011 : 8'b00011011;
									assign node1025 = (inp[12]) ? 8'b00001011 : node1026;
										assign node1026 = (inp[11]) ? 8'b00011010 : 8'b00001011;
								assign node1030 = (inp[3]) ? node1044 : node1031;
									assign node1031 = (inp[2]) ? node1039 : node1032;
										assign node1032 = (inp[6]) ? node1034 : 8'b10000010;
											assign node1034 = (inp[12]) ? 8'b00011010 : node1035;
												assign node1035 = (inp[11]) ? 8'b00001010 : 8'b00011010;
										assign node1039 = (inp[12]) ? 8'b00000010 : node1040;
											assign node1040 = (inp[11]) ? 8'b11110111 : 8'b10000010;
									assign node1044 = (inp[2]) ? 8'b00001011 : node1045;
										assign node1045 = (inp[11]) ? node1049 : node1046;
											assign node1046 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node1049 = (inp[6]) ? 8'b00001011 : 8'b00011010;
							assign node1053 = (inp[2]) ? node1069 : node1054;
								assign node1054 = (inp[6]) ? node1064 : node1055;
									assign node1055 = (inp[4]) ? node1061 : node1056;
										assign node1056 = (inp[12]) ? 8'b00011010 : node1057;
											assign node1057 = (inp[11]) ? 8'b00001010 : 8'b00011010;
										assign node1061 = (inp[12]) ? 8'b00000010 : 8'b11110111;
									assign node1064 = (inp[12]) ? 8'b00011010 : node1065;
										assign node1065 = (inp[11]) ? 8'b00001010 : 8'b00011010;
								assign node1069 = (inp[12]) ? 8'b00000010 : node1070;
									assign node1070 = (inp[11]) ? 8'b11110111 : 8'b10000010;
					assign node1074 = (inp[9]) ? node1236 : node1075;
						assign node1075 = (inp[8]) ? node1155 : node1076;
							assign node1076 = (inp[4]) ? node1112 : node1077;
								assign node1077 = (inp[2]) ? node1089 : node1078;
									assign node1078 = (inp[1]) ? node1084 : node1079;
										assign node1079 = (inp[10]) ? 8'b00011111 : node1080;
											assign node1080 = (inp[11]) ? 8'b00001111 : 8'b00011111;
										assign node1084 = (inp[3]) ? node1086 : 8'b00011110;
											assign node1086 = (inp[11]) ? 8'b00011011 : 8'b00011111;
									assign node1089 = (inp[6]) ? node1099 : node1090;
										assign node1090 = (inp[11]) ? node1094 : node1091;
											assign node1091 = (inp[3]) ? 8'b00001111 : 8'b00001110;
											assign node1094 = (inp[12]) ? 8'b00001110 : node1095;
												assign node1095 = (inp[1]) ? 8'b00011010 : 8'b00011110;
										assign node1099 = (inp[11]) ? node1105 : node1100;
											assign node1100 = (inp[3]) ? 8'b00011111 : node1101;
												assign node1101 = (inp[1]) ? 8'b00011110 : 8'b00011111;
											assign node1105 = (inp[1]) ? node1107 : 8'b00001110;
												assign node1107 = (inp[12]) ? node1109 : 8'b00001011;
													assign node1109 = (inp[3]) ? 8'b00011010 : 8'b00011011;
								assign node1112 = (inp[10]) ? node1144 : node1113;
									assign node1113 = (inp[3]) ? node1129 : node1114;
										assign node1114 = (inp[2]) ? node1122 : node1115;
											assign node1115 = (inp[6]) ? node1119 : node1116;
												assign node1116 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node1119 = (inp[1]) ? 8'b00001010 : 8'b00011010;
											assign node1122 = (inp[12]) ? node1126 : node1123;
												assign node1123 = (inp[6]) ? 8'b10100101 : 8'b11110111;
												assign node1126 = (inp[6]) ? 8'b10010000 : 8'b00000010;
										assign node1129 = (inp[1]) ? node1137 : node1130;
											assign node1130 = (inp[6]) ? node1132 : 8'b00001011;
												assign node1132 = (inp[12]) ? 8'b00011011 : node1133;
													assign node1133 = (inp[11]) ? 8'b00001011 : 8'b00011011;
											assign node1137 = (inp[11]) ? node1141 : node1138;
												assign node1138 = (inp[6]) ? 8'b10011001 : 8'b10000001;
												assign node1141 = (inp[6]) ? 8'b10100100 : 8'b10110100;
									assign node1144 = (inp[3]) ? node1152 : node1145;
										assign node1145 = (inp[12]) ? 8'b00001110 : node1146;
											assign node1146 = (inp[2]) ? node1148 : 8'b00001110;
												assign node1148 = (inp[6]) ? 8'b00001011 : 8'b00011011;
										assign node1152 = (inp[6]) ? 8'b00011110 : 8'b00001111;
							assign node1155 = (inp[10]) ? node1195 : node1156;
								assign node1156 = (inp[1]) ? node1172 : node1157;
									assign node1157 = (inp[4]) ? node1167 : node1158;
										assign node1158 = (inp[12]) ? node1164 : node1159;
											assign node1159 = (inp[11]) ? 8'b00001011 : node1160;
												assign node1160 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node1164 = (inp[2]) ? 8'b00011010 : 8'b00011011;
										assign node1167 = (inp[11]) ? node1169 : 8'b10000010;
											assign node1169 = (inp[6]) ? 8'b00001010 : 8'b00011010;
									assign node1172 = (inp[11]) ? node1180 : node1173;
										assign node1173 = (inp[3]) ? 8'b10000001 : node1174;
											assign node1174 = (inp[6]) ? 8'b10010000 : node1175;
												assign node1175 = (inp[4]) ? 8'b00000010 : 8'b00011010;
										assign node1180 = (inp[6]) ? node1188 : node1181;
											assign node1181 = (inp[12]) ? node1185 : node1182;
												assign node1182 = (inp[4]) ? 8'b11110111 : 8'b10110100;
												assign node1185 = (inp[2]) ? 8'b00000010 : 8'b10100101;
											assign node1188 = (inp[12]) ? node1192 : node1189;
												assign node1189 = (inp[3]) ? 8'b10100100 : 8'b10100101;
												assign node1192 = (inp[3]) ? 8'b10110100 : 8'b11110101;
								assign node1195 = (inp[11]) ? node1211 : node1196;
									assign node1196 = (inp[6]) ? node1206 : node1197;
										assign node1197 = (inp[1]) ? node1203 : node1198;
											assign node1198 = (inp[4]) ? 8'b10001101 : node1199;
												assign node1199 = (inp[2]) ? 8'b10001101 : 8'b10011101;
											assign node1203 = (inp[3]) ? 8'b10000101 : 8'b10000100;
										assign node1206 = (inp[4]) ? 8'b10010100 : node1207;
											assign node1207 = (inp[1]) ? 8'b10011100 : 8'b10011101;
									assign node1211 = (inp[1]) ? node1225 : node1212;
										assign node1212 = (inp[3]) ? node1222 : node1213;
											assign node1213 = (inp[4]) ? node1217 : node1214;
												assign node1214 = (inp[2]) ? 8'b10111100 : 8'b11111101;
												assign node1217 = (inp[2]) ? 8'b10110001 : node1218;
													assign node1218 = (inp[6]) ? 8'b10111100 : 8'b10100100;
											assign node1222 = (inp[2]) ? 8'b10101100 : 8'b10101101;
										assign node1225 = (inp[6]) ? node1231 : node1226;
											assign node1226 = (inp[12]) ? node1228 : 8'b10110000;
												assign node1228 = (inp[3]) ? 8'b10100001 : 8'b10100100;
											assign node1231 = (inp[12]) ? 8'b10111001 : node1232;
												assign node1232 = (inp[2]) ? 8'b10100001 : 8'b10101001;
						assign node1236 = (inp[11]) ? node1288 : node1237;
							assign node1237 = (inp[4]) ? node1263 : node1238;
								assign node1238 = (inp[8]) ? node1248 : node1239;
									assign node1239 = (inp[3]) ? node1243 : node1240;
										assign node1240 = (inp[1]) ? 8'b10111100 : 8'b11111101;
										assign node1243 = (inp[6]) ? 8'b11111101 : node1244;
											assign node1244 = (inp[2]) ? 8'b10101101 : 8'b11111101;
									assign node1248 = (inp[10]) ? node1258 : node1249;
										assign node1249 = (inp[2]) ? node1251 : 8'b10111001;
											assign node1251 = (inp[1]) ? node1255 : node1252;
												assign node1252 = (inp[6]) ? 8'b10111001 : 8'b10101001;
												assign node1255 = (inp[3]) ? 8'b10110001 : 8'b10110000;
										assign node1258 = (inp[2]) ? node1260 : 8'b11111101;
											assign node1260 = (inp[1]) ? 8'b10100100 : 8'b10101101;
								assign node1263 = (inp[10]) ? node1279 : node1264;
									assign node1264 = (inp[6]) ? node1270 : node1265;
										assign node1265 = (inp[3]) ? node1267 : 8'b10100000;
											assign node1267 = (inp[1]) ? 8'b10100001 : 8'b10101001;
										assign node1270 = (inp[3]) ? node1274 : node1271;
											assign node1271 = (inp[2]) ? 8'b10110000 : 8'b10111000;
											assign node1274 = (inp[1]) ? node1276 : 8'b10111001;
												assign node1276 = (inp[12]) ? 8'b10110001 : 8'b10111001;
									assign node1279 = (inp[3]) ? node1285 : node1280;
										assign node1280 = (inp[8]) ? node1282 : 8'b10101100;
											assign node1282 = (inp[6]) ? 8'b10111100 : 8'b10100100;
										assign node1285 = (inp[6]) ? 8'b11111101 : 8'b10101101;
							assign node1288 = (inp[8]) ? node1344 : node1289;
								assign node1289 = (inp[1]) ? node1315 : node1290;
									assign node1290 = (inp[10]) ? node1294 : node1291;
										assign node1291 = (inp[4]) ? 8'b10101001 : 8'b10101101;
										assign node1294 = (inp[4]) ? node1304 : node1295;
											assign node1295 = (inp[2]) ? node1299 : node1296;
												assign node1296 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node1299 = (inp[12]) ? node1301 : 8'b10111100;
													assign node1301 = (inp[3]) ? 8'b10111100 : 8'b10101101;
											assign node1304 = (inp[2]) ? node1312 : node1305;
												assign node1305 = (inp[6]) ? node1309 : node1306;
													assign node1306 = (inp[3]) ? 8'b10111100 : 8'b10101100;
													assign node1309 = (inp[3]) ? 8'b10101101 : 8'b10101100;
												assign node1312 = (inp[6]) ? 8'b10101001 : 8'b10101101;
									assign node1315 = (inp[12]) ? node1329 : node1316;
										assign node1316 = (inp[4]) ? node1318 : 8'b10101001;
											assign node1318 = (inp[6]) ? node1322 : node1319;
												assign node1319 = (inp[3]) ? 8'b10111000 : 8'b10111001;
												assign node1322 = (inp[2]) ? node1326 : node1323;
													assign node1323 = (inp[10]) ? 8'b10101100 : 8'b10101000;
													assign node1326 = (inp[3]) ? 8'b10101000 : 8'b10101001;
										assign node1329 = (inp[6]) ? node1335 : node1330;
											assign node1330 = (inp[2]) ? 8'b10101100 : node1331;
												assign node1331 = (inp[4]) ? 8'b10101001 : 8'b10111001;
											assign node1335 = (inp[3]) ? node1339 : node1336;
												assign node1336 = (inp[2]) ? 8'b10111001 : 8'b10111000;
												assign node1339 = (inp[2]) ? node1341 : 8'b10011101;
													assign node1341 = (inp[10]) ? 8'b10111000 : 8'b10010000;
								assign node1344 = (inp[2]) ? node1378 : node1345;
									assign node1345 = (inp[10]) ? node1363 : node1346;
										assign node1346 = (inp[1]) ? node1356 : node1347;
											assign node1347 = (inp[3]) ? node1351 : node1348;
												assign node1348 = (inp[12]) ? 8'b10100000 : 8'b10010101;
												assign node1351 = (inp[12]) ? node1353 : 8'b10111000;
													assign node1353 = (inp[4]) ? 8'b10101001 : 8'b10111001;
											assign node1356 = (inp[3]) ? node1358 : 8'b10101000;
												assign node1358 = (inp[4]) ? node1360 : 8'b10001101;
													assign node1360 = (inp[12]) ? 8'b10000101 : 8'b10010100;
										assign node1363 = (inp[3]) ? node1373 : node1364;
											assign node1364 = (inp[6]) ? 8'b10011100 : node1365;
												assign node1365 = (inp[1]) ? node1369 : node1366;
													assign node1366 = (inp[12]) ? 8'b10011101 : 8'b10001101;
													assign node1369 = (inp[4]) ? 8'b10000100 : 8'b10001100;
											assign node1373 = (inp[1]) ? node1375 : 8'b10001101;
												assign node1375 = (inp[4]) ? 8'b10011001 : 8'b10001001;
									assign node1378 = (inp[1]) ? node1392 : node1379;
										assign node1379 = (inp[4]) ? node1383 : node1380;
											assign node1380 = (inp[10]) ? 8'b10001100 : 8'b10101000;
											assign node1383 = (inp[3]) ? node1387 : node1384;
												assign node1384 = (inp[10]) ? 8'b10010001 : 8'b10000101;
												assign node1387 = (inp[12]) ? 8'b10001101 : node1388;
													assign node1388 = (inp[10]) ? 8'b10011100 : 8'b10111000;
										assign node1392 = (inp[10]) ? node1398 : node1393;
											assign node1393 = (inp[3]) ? node1395 : 8'b10100000;
												assign node1395 = (inp[6]) ? 8'b10000100 : 8'b10010100;
											assign node1398 = (inp[3]) ? node1404 : node1399;
												assign node1399 = (inp[4]) ? 8'b10010001 : node1400;
													assign node1400 = (inp[12]) ? 8'b10010001 : 8'b10000001;
												assign node1404 = (inp[6]) ? node1408 : node1405;
													assign node1405 = (inp[12]) ? 8'b10000001 : 8'b10010000;
													assign node1408 = (inp[12]) ? 8'b10010000 : 8'b10000000;
				assign node1411 = (inp[11]) ? node1657 : node1412;
					assign node1412 = (inp[5]) ? node1588 : node1413;
						assign node1413 = (inp[9]) ? node1499 : node1414;
							assign node1414 = (inp[4]) ? node1446 : node1415;
								assign node1415 = (inp[2]) ? node1433 : node1416;
									assign node1416 = (inp[1]) ? node1422 : node1417;
										assign node1417 = (inp[8]) ? node1419 : 8'b11111101;
											assign node1419 = (inp[10]) ? 8'b10111001 : 8'b11111101;
										assign node1422 = (inp[3]) ? node1428 : node1423;
											assign node1423 = (inp[8]) ? node1425 : 8'b11111101;
												assign node1425 = (inp[10]) ? 8'b10111001 : 8'b11111101;
											assign node1428 = (inp[8]) ? node1430 : 8'b10111100;
												assign node1430 = (inp[12]) ? 8'b10111100 : 8'b10111000;
									assign node1433 = (inp[6]) ? 8'b10101101 : node1434;
										assign node1434 = (inp[1]) ? node1440 : node1435;
											assign node1435 = (inp[12]) ? node1437 : 8'b11111101;
												assign node1437 = (inp[3]) ? 8'b11111101 : 8'b10111001;
											assign node1440 = (inp[3]) ? node1442 : 8'b11110101;
												assign node1442 = (inp[8]) ? 8'b10110100 : 8'b10111100;
								assign node1446 = (inp[2]) ? node1478 : node1447;
									assign node1447 = (inp[6]) ? node1463 : node1448;
										assign node1448 = (inp[10]) ? node1456 : node1449;
											assign node1449 = (inp[8]) ? node1451 : 8'b10100001;
												assign node1451 = (inp[3]) ? 8'b10101101 : node1452;
													assign node1452 = (inp[1]) ? 8'b10100101 : 8'b10100100;
											assign node1456 = (inp[8]) ? 8'b10101001 : node1457;
												assign node1457 = (inp[3]) ? 8'b10101100 : node1458;
													assign node1458 = (inp[1]) ? 8'b10101101 : 8'b10101100;
										assign node1463 = (inp[8]) ? node1473 : node1464;
											assign node1464 = (inp[10]) ? node1468 : node1465;
												assign node1465 = (inp[1]) ? 8'b10111000 : 8'b10111001;
												assign node1468 = (inp[3]) ? 8'b11111101 : node1469;
													assign node1469 = (inp[1]) ? 8'b11111101 : 8'b10111100;
											assign node1473 = (inp[10]) ? node1475 : 8'b10111100;
												assign node1475 = (inp[12]) ? 8'b10111001 : 8'b10111000;
									assign node1478 = (inp[6]) ? node1492 : node1479;
										assign node1479 = (inp[1]) ? node1483 : node1480;
											assign node1480 = (inp[3]) ? 8'b10111001 : 8'b10110000;
											assign node1483 = (inp[3]) ? node1485 : 8'b11110101;
												assign node1485 = (inp[12]) ? node1489 : node1486;
													assign node1486 = (inp[10]) ? 8'b10111100 : 8'b10110100;
													assign node1489 = (inp[10]) ? 8'b10110000 : 8'b10110000;
										assign node1492 = (inp[1]) ? node1494 : 8'b10100000;
											assign node1494 = (inp[10]) ? 8'b10100001 : node1495;
												assign node1495 = (inp[8]) ? 8'b10100101 : 8'b10100001;
							assign node1499 = (inp[8]) ? node1551 : node1500;
								assign node1500 = (inp[10]) ? node1526 : node1501;
									assign node1501 = (inp[4]) ? node1509 : node1502;
										assign node1502 = (inp[2]) ? 8'b00001111 : node1503;
											assign node1503 = (inp[6]) ? 8'b00011111 : node1504;
												assign node1504 = (inp[1]) ? 8'b00011110 : 8'b00011111;
										assign node1509 = (inp[2]) ? node1519 : node1510;
											assign node1510 = (inp[6]) ? node1514 : node1511;
												assign node1511 = (inp[3]) ? 8'b00001011 : 8'b10000010;
												assign node1514 = (inp[3]) ? node1516 : 8'b00011010;
													assign node1516 = (inp[1]) ? 8'b00011010 : 8'b00011011;
											assign node1519 = (inp[6]) ? node1523 : node1520;
												assign node1520 = (inp[1]) ? 8'b10010000 : 8'b00011011;
												assign node1523 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node1526 = (inp[6]) ? node1542 : node1527;
										assign node1527 = (inp[2]) ? node1535 : node1528;
											assign node1528 = (inp[4]) ? node1530 : 8'b00011111;
												assign node1530 = (inp[12]) ? node1532 : 8'b00001111;
													assign node1532 = (inp[3]) ? 8'b00001110 : 8'b00001111;
											assign node1535 = (inp[12]) ? 8'b00011111 : node1536;
												assign node1536 = (inp[1]) ? 8'b00011111 : node1537;
													assign node1537 = (inp[4]) ? 8'b00011110 : 8'b00011111;
										assign node1542 = (inp[2]) ? node1548 : node1543;
											assign node1543 = (inp[12]) ? node1545 : 8'b00011110;
												assign node1545 = (inp[4]) ? 8'b00011111 : 8'b00011110;
											assign node1548 = (inp[3]) ? 8'b00001110 : 8'b00001111;
								assign node1551 = (inp[10]) ? node1577 : node1552;
									assign node1552 = (inp[2]) ? node1564 : node1553;
										assign node1553 = (inp[4]) ? node1559 : node1554;
											assign node1554 = (inp[3]) ? node1556 : 8'b10011101;
												assign node1556 = (inp[1]) ? 8'b10011100 : 8'b10011101;
											assign node1559 = (inp[6]) ? node1561 : 8'b10000100;
												assign node1561 = (inp[12]) ? 8'b10011100 : 8'b10011101;
										assign node1564 = (inp[6]) ? node1570 : node1565;
											assign node1565 = (inp[3]) ? 8'b10010100 : node1566;
												assign node1566 = (inp[1]) ? 8'b10010101 : 8'b10010100;
											assign node1570 = (inp[4]) ? node1572 : 8'b10001101;
												assign node1572 = (inp[1]) ? 8'b10000100 : node1573;
													assign node1573 = (inp[3]) ? 8'b10001101 : 8'b10000100;
									assign node1577 = (inp[2]) ? node1583 : node1578;
										assign node1578 = (inp[3]) ? 8'b00001011 : node1579;
											assign node1579 = (inp[4]) ? 8'b10000010 : 8'b00011011;
										assign node1583 = (inp[3]) ? node1585 : 8'b10010000;
											assign node1585 = (inp[1]) ? 8'b10010000 : 8'b00011011;
						assign node1588 = (inp[4]) ? node1596 : node1589;
							assign node1589 = (inp[8]) ? node1591 : 8'b11111101;
								assign node1591 = (inp[2]) ? node1593 : 8'b11111101;
									assign node1593 = (inp[1]) ? 8'b11110101 : 8'b11111101;
							assign node1596 = (inp[6]) ? node1630 : node1597;
								assign node1597 = (inp[2]) ? node1613 : node1598;
									assign node1598 = (inp[8]) ? node1606 : node1599;
										assign node1599 = (inp[10]) ? node1601 : 8'b10100001;
											assign node1601 = (inp[1]) ? 8'b10101101 : node1602;
												assign node1602 = (inp[3]) ? 8'b10101101 : 8'b10101100;
										assign node1606 = (inp[3]) ? node1610 : node1607;
											assign node1607 = (inp[1]) ? 8'b10100101 : 8'b10100100;
											assign node1610 = (inp[1]) ? 8'b10100101 : 8'b10101101;
									assign node1613 = (inp[10]) ? node1621 : node1614;
										assign node1614 = (inp[8]) ? node1618 : node1615;
											assign node1615 = (inp[1]) ? 8'b10110001 : 8'b10110000;
											assign node1618 = (inp[1]) ? 8'b11110101 : 8'b10110100;
										assign node1621 = (inp[3]) ? node1623 : 8'b10111100;
											assign node1623 = (inp[12]) ? node1625 : 8'b11111101;
												assign node1625 = (inp[1]) ? node1627 : 8'b11111101;
													assign node1627 = (inp[8]) ? 8'b11110101 : 8'b11111101;
								assign node1630 = (inp[8]) ? node1646 : node1631;
									assign node1631 = (inp[10]) ? node1643 : node1632;
										assign node1632 = (inp[2]) ? node1638 : node1633;
											assign node1633 = (inp[1]) ? 8'b10111001 : node1634;
												assign node1634 = (inp[3]) ? 8'b10111001 : 8'b10111000;
											assign node1638 = (inp[9]) ? node1640 : 8'b10111001;
												assign node1640 = (inp[1]) ? 8'b10110001 : 8'b10110000;
										assign node1643 = (inp[3]) ? 8'b11111101 : 8'b10111100;
									assign node1646 = (inp[2]) ? node1652 : node1647;
										assign node1647 = (inp[1]) ? 8'b11111101 : node1648;
											assign node1648 = (inp[10]) ? 8'b10111100 : 8'b11111101;
										assign node1652 = (inp[1]) ? 8'b11110101 : node1653;
											assign node1653 = (inp[3]) ? 8'b11111101 : 8'b10110100;
					assign node1657 = (inp[12]) ? node1799 : node1658;
						assign node1658 = (inp[8]) ? node1738 : node1659;
							assign node1659 = (inp[5]) ? node1711 : node1660;
								assign node1660 = (inp[9]) ? node1686 : node1661;
									assign node1661 = (inp[1]) ? node1671 : node1662;
										assign node1662 = (inp[2]) ? node1668 : node1663;
											assign node1663 = (inp[4]) ? node1665 : 8'b10101101;
												assign node1665 = (inp[3]) ? 8'b10101001 : 8'b10101000;
											assign node1668 = (inp[6]) ? 8'b10111100 : 8'b10101100;
										assign node1671 = (inp[4]) ? node1679 : node1672;
											assign node1672 = (inp[6]) ? node1676 : node1673;
												assign node1673 = (inp[3]) ? 8'b10101001 : 8'b10101000;
												assign node1676 = (inp[3]) ? 8'b10111001 : 8'b10111000;
											assign node1679 = (inp[2]) ? 8'b10010101 : node1680;
												assign node1680 = (inp[3]) ? node1682 : 8'b10001101;
													assign node1682 = (inp[6]) ? 8'b10101000 : 8'b10111001;
									assign node1686 = (inp[4]) ? node1694 : node1687;
										assign node1687 = (inp[1]) ? node1691 : node1688;
											assign node1688 = (inp[10]) ? 8'b00001111 : 8'b00011110;
											assign node1691 = (inp[3]) ? 8'b00001011 : 8'b00001010;
										assign node1694 = (inp[10]) ? node1706 : node1695;
											assign node1695 = (inp[2]) ? node1701 : node1696;
												assign node1696 = (inp[6]) ? node1698 : 8'b10110100;
													assign node1698 = (inp[1]) ? 8'b00001010 : 8'b00001010;
												assign node1701 = (inp[1]) ? node1703 : 8'b11110111;
													assign node1703 = (inp[6]) ? 8'b10110100 : 8'b10100100;
											assign node1706 = (inp[6]) ? node1708 : 8'b00001011;
												assign node1708 = (inp[1]) ? 8'b00011010 : 8'b00011110;
								assign node1711 = (inp[2]) ? node1723 : node1712;
									assign node1712 = (inp[1]) ? node1718 : node1713;
										assign node1713 = (inp[4]) ? node1715 : 8'b10101101;
											assign node1715 = (inp[10]) ? 8'b10111001 : 8'b10010101;
										assign node1718 = (inp[4]) ? node1720 : 8'b10101001;
											assign node1720 = (inp[6]) ? 8'b10101001 : 8'b10111000;
									assign node1723 = (inp[3]) ? node1731 : node1724;
										assign node1724 = (inp[10]) ? node1728 : node1725;
											assign node1725 = (inp[9]) ? 8'b10000101 : 8'b10000100;
											assign node1728 = (inp[4]) ? 8'b10101001 : 8'b10101100;
										assign node1731 = (inp[1]) ? 8'b10101000 : node1732;
											assign node1732 = (inp[6]) ? node1734 : 8'b10101100;
												assign node1734 = (inp[10]) ? 8'b10101100 : 8'b10101000;
							assign node1738 = (inp[1]) ? node1774 : node1739;
								assign node1739 = (inp[5]) ? node1763 : node1740;
									assign node1740 = (inp[9]) ? node1756 : node1741;
										assign node1741 = (inp[10]) ? node1747 : node1742;
											assign node1742 = (inp[3]) ? node1744 : 8'b10010001;
												assign node1744 = (inp[6]) ? 8'b10001101 : 8'b10011100;
											assign node1747 = (inp[3]) ? node1753 : node1748;
												assign node1748 = (inp[2]) ? 8'b10000101 : node1749;
													assign node1749 = (inp[4]) ? 8'b10101000 : 8'b10101001;
												assign node1753 = (inp[6]) ? 8'b10111000 : 8'b10101000;
										assign node1756 = (inp[10]) ? node1758 : 8'b10101100;
											assign node1758 = (inp[6]) ? 8'b00011010 : node1759;
												assign node1759 = (inp[4]) ? 8'b00001010 : 8'b00001011;
									assign node1763 = (inp[4]) ? node1767 : node1764;
										assign node1764 = (inp[2]) ? 8'b10001100 : 8'b10001101;
										assign node1767 = (inp[3]) ? node1771 : node1768;
											assign node1768 = (inp[2]) ? 8'b10000001 : 8'b10010001;
											assign node1771 = (inp[2]) ? 8'b10001100 : 8'b10001101;
								assign node1774 = (inp[5]) ? node1792 : node1775;
									assign node1775 = (inp[9]) ? node1783 : node1776;
										assign node1776 = (inp[3]) ? node1780 : node1777;
											assign node1777 = (inp[10]) ? 8'b10010100 : 8'b10000000;
											assign node1780 = (inp[10]) ? 8'b10101000 : 8'b10001100;
										assign node1783 = (inp[10]) ? 8'b11110111 : node1784;
											assign node1784 = (inp[2]) ? node1788 : node1785;
												assign node1785 = (inp[4]) ? 8'b10101001 : 8'b10101100;
												assign node1788 = (inp[6]) ? 8'b10110001 : 8'b10100000;
									assign node1792 = (inp[6]) ? node1796 : node1793;
										assign node1793 = (inp[2]) ? 8'b10000000 : 8'b10010000;
										assign node1796 = (inp[2]) ? 8'b10000000 : 8'b10001001;
						assign node1799 = (inp[8]) ? node1883 : node1800;
							assign node1800 = (inp[9]) ? node1844 : node1801;
								assign node1801 = (inp[2]) ? node1829 : node1802;
									assign node1802 = (inp[6]) ? node1816 : node1803;
										assign node1803 = (inp[10]) ? node1809 : node1804;
											assign node1804 = (inp[5]) ? node1806 : 8'b10100000;
												assign node1806 = (inp[1]) ? 8'b10000101 : 8'b10100000;
											assign node1809 = (inp[1]) ? node1813 : node1810;
												assign node1810 = (inp[3]) ? 8'b10101101 : 8'b10101100;
												assign node1813 = (inp[3]) ? 8'b10101100 : 8'b10101001;
										assign node1816 = (inp[4]) ? node1820 : node1817;
											assign node1817 = (inp[1]) ? 8'b10111001 : 8'b11111101;
											assign node1820 = (inp[1]) ? node1826 : node1821;
												assign node1821 = (inp[3]) ? 8'b10111001 : node1822;
													assign node1822 = (inp[5]) ? 8'b10111000 : 8'b10111100;
												assign node1826 = (inp[10]) ? 8'b10111001 : 8'b10011101;
									assign node1829 = (inp[1]) ? node1837 : node1830;
										assign node1830 = (inp[6]) ? node1832 : 8'b10111100;
											assign node1832 = (inp[4]) ? node1834 : 8'b10111100;
												assign node1834 = (inp[10]) ? 8'b10111100 : 8'b10111000;
										assign node1837 = (inp[4]) ? node1841 : node1838;
											assign node1838 = (inp[5]) ? 8'b10111000 : 8'b10111001;
											assign node1841 = (inp[3]) ? 8'b10010100 : 8'b10111000;
								assign node1844 = (inp[5]) ? node1872 : node1845;
									assign node1845 = (inp[1]) ? node1859 : node1846;
										assign node1846 = (inp[10]) ? node1852 : node1847;
											assign node1847 = (inp[4]) ? node1849 : 8'b00011111;
												assign node1849 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node1852 = (inp[6]) ? 8'b00011111 : node1853;
												assign node1853 = (inp[4]) ? 8'b00001110 : node1854;
													assign node1854 = (inp[2]) ? 8'b00011110 : 8'b00011111;
										assign node1859 = (inp[10]) ? node1861 : 8'b00000010;
											assign node1861 = (inp[4]) ? node1867 : node1862;
												assign node1862 = (inp[3]) ? 8'b00011011 : node1863;
													assign node1863 = (inp[6]) ? 8'b00011011 : 8'b00011010;
												assign node1867 = (inp[6]) ? 8'b00011011 : node1868;
													assign node1868 = (inp[3]) ? 8'b00011011 : 8'b00001011;
									assign node1872 = (inp[1]) ? node1880 : node1873;
										assign node1873 = (inp[4]) ? node1877 : node1874;
											assign node1874 = (inp[2]) ? 8'b10111100 : 8'b11111101;
											assign node1877 = (inp[10]) ? 8'b10111001 : 8'b10111000;
										assign node1880 = (inp[2]) ? 8'b10111000 : 8'b10111001;
							assign node1883 = (inp[5]) ? node1935 : node1884;
								assign node1884 = (inp[10]) ? node1912 : node1885;
									assign node1885 = (inp[9]) ? node1901 : node1886;
										assign node1886 = (inp[1]) ? node1898 : node1887;
											assign node1887 = (inp[3]) ? node1891 : node1888;
												assign node1888 = (inp[4]) ? 8'b10010001 : 8'b10011100;
												assign node1891 = (inp[2]) ? node1895 : node1892;
													assign node1892 = (inp[6]) ? 8'b10011101 : 8'b10001101;
													assign node1895 = (inp[6]) ? 8'b10001101 : 8'b10011100;
											assign node1898 = (inp[3]) ? 8'b10010001 : 8'b10011001;
										assign node1901 = (inp[1]) ? node1905 : node1902;
											assign node1902 = (inp[4]) ? 8'b10101101 : 8'b10111100;
											assign node1905 = (inp[6]) ? node1909 : node1906;
												assign node1906 = (inp[3]) ? 8'b10110001 : 8'b10110000;
												assign node1909 = (inp[4]) ? 8'b10100100 : 8'b10111100;
									assign node1912 = (inp[9]) ? node1928 : node1913;
										assign node1913 = (inp[1]) ? node1921 : node1914;
											assign node1914 = (inp[6]) ? node1918 : node1915;
												assign node1915 = (inp[2]) ? 8'b10111000 : 8'b10111001;
												assign node1918 = (inp[2]) ? 8'b10101001 : 8'b10111001;
											assign node1921 = (inp[2]) ? 8'b10010101 : node1922;
												assign node1922 = (inp[3]) ? node1924 : 8'b10011101;
													assign node1924 = (inp[4]) ? 8'b10100000 : 8'b10111000;
										assign node1928 = (inp[2]) ? node1932 : node1929;
											assign node1929 = (inp[1]) ? 8'b11111101 : 8'b00011011;
											assign node1932 = (inp[4]) ? 8'b11110101 : 8'b10100101;
								assign node1935 = (inp[1]) ? node1949 : node1936;
									assign node1936 = (inp[3]) ? node1942 : node1937;
										assign node1937 = (inp[2]) ? node1939 : 8'b10000100;
											assign node1939 = (inp[4]) ? 8'b10010001 : 8'b10011100;
										assign node1942 = (inp[2]) ? 8'b10011100 : node1943;
											assign node1943 = (inp[6]) ? 8'b10011101 : node1944;
												assign node1944 = (inp[4]) ? 8'b10001101 : 8'b10011101;
									assign node1949 = (inp[2]) ? 8'b10010000 : 8'b10011001;
		assign node1952 = (inp[4]) ? node3232 : node1953;
			assign node1953 = (inp[13]) ? node2605 : node1954;
				assign node1954 = (inp[9]) ? node2290 : node1955;
					assign node1955 = (inp[11]) ? node2089 : node1956;
						assign node1956 = (inp[5]) ? node2000 : node1957;
							assign node1957 = (inp[3]) ? node1981 : node1958;
								assign node1958 = (inp[0]) ? node1974 : node1959;
									assign node1959 = (inp[1]) ? node1965 : node1960;
										assign node1960 = (inp[6]) ? 8'b00101011 : node1961;
											assign node1961 = (inp[2]) ? 8'b00101011 : 8'b00111011;
										assign node1965 = (inp[8]) ? node1969 : node1966;
											assign node1966 = (inp[10]) ? 8'b00101010 : 8'b00101110;
											assign node1969 = (inp[2]) ? 8'b00101010 : node1970;
												assign node1970 = (inp[6]) ? 8'b00101010 : 8'b00111010;
									assign node1974 = (inp[10]) ? node1978 : node1975;
										assign node1975 = (inp[6]) ? 8'b00101111 : 8'b01111111;
										assign node1978 = (inp[6]) ? 8'b00101011 : 8'b00111011;
								assign node1981 = (inp[6]) ? node1993 : node1982;
									assign node1982 = (inp[10]) ? node1988 : node1983;
										assign node1983 = (inp[8]) ? node1985 : 8'b00111110;
											assign node1985 = (inp[2]) ? 8'b00101010 : 8'b00111010;
										assign node1988 = (inp[2]) ? node1990 : 8'b00111010;
											assign node1990 = (inp[0]) ? 8'b00111010 : 8'b00101010;
									assign node1993 = (inp[8]) ? node1995 : 8'b00101110;
										assign node1995 = (inp[0]) ? node1997 : 8'b00101010;
											assign node1997 = (inp[12]) ? 8'b00101010 : 8'b00101110;
							assign node2000 = (inp[0]) ? node2062 : node2001;
								assign node2001 = (inp[12]) ? node2033 : node2002;
									assign node2002 = (inp[10]) ? node2022 : node2003;
										assign node2003 = (inp[8]) ? node2015 : node2004;
											assign node2004 = (inp[3]) ? node2010 : node2005;
												assign node2005 = (inp[1]) ? node2007 : 8'b00101111;
													assign node2007 = (inp[6]) ? 8'b00101110 : 8'b00101110;
												assign node2010 = (inp[1]) ? node2012 : 8'b00111110;
													assign node2012 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node2015 = (inp[1]) ? 8'b00111010 : node2016;
												assign node2016 = (inp[3]) ? 8'b00101010 : node2017;
													assign node2017 = (inp[2]) ? 8'b00111011 : 8'b00101011;
										assign node2022 = (inp[8]) ? node2028 : node2023;
											assign node2023 = (inp[1]) ? node2025 : 8'b00111011;
												assign node2025 = (inp[3]) ? 8'b00111011 : 8'b00111010;
											assign node2028 = (inp[2]) ? node2030 : 8'b01111111;
												assign node2030 = (inp[6]) ? 8'b01111111 : 8'b00101111;
									assign node2033 = (inp[3]) ? node2045 : node2034;
										assign node2034 = (inp[1]) ? node2042 : node2035;
											assign node2035 = (inp[10]) ? node2037 : 8'b00111011;
												assign node2037 = (inp[8]) ? node2039 : 8'b00101011;
													assign node2039 = (inp[2]) ? 8'b00101111 : 8'b00101111;
											assign node2042 = (inp[6]) ? 8'b00111010 : 8'b00101010;
										assign node2045 = (inp[1]) ? node2057 : node2046;
											assign node2046 = (inp[6]) ? node2052 : node2047;
												assign node2047 = (inp[2]) ? 8'b00101110 : node2048;
													assign node2048 = (inp[8]) ? 8'b00111110 : 8'b00111010;
												assign node2052 = (inp[10]) ? node2054 : 8'b00111010;
													assign node2054 = (inp[8]) ? 8'b00111110 : 8'b00111010;
											assign node2057 = (inp[10]) ? 8'b00111011 : node2058;
												assign node2058 = (inp[8]) ? 8'b00111011 : 8'b00101111;
								assign node2062 = (inp[1]) ? node2076 : node2063;
									assign node2063 = (inp[3]) ? node2069 : node2064;
										assign node2064 = (inp[10]) ? node2066 : 8'b00101111;
											assign node2066 = (inp[8]) ? 8'b01111111 : 8'b00111011;
										assign node2069 = (inp[6]) ? node2073 : node2070;
											assign node2070 = (inp[10]) ? 8'b00111010 : 8'b00111110;
											assign node2073 = (inp[2]) ? 8'b00111110 : 8'b00101110;
									assign node2076 = (inp[10]) ? node2082 : node2077;
										assign node2077 = (inp[6]) ? node2079 : 8'b01111111;
											assign node2079 = (inp[2]) ? 8'b01111111 : 8'b00101111;
										assign node2082 = (inp[8]) ? 8'b01111111 : node2083;
											assign node2083 = (inp[6]) ? node2085 : 8'b00111011;
												assign node2085 = (inp[2]) ? 8'b00111011 : 8'b00101011;
						assign node2089 = (inp[10]) ? node2183 : node2090;
							assign node2090 = (inp[8]) ? node2138 : node2091;
								assign node2091 = (inp[12]) ? node2117 : node2092;
									assign node2092 = (inp[3]) ? node2104 : node2093;
										assign node2093 = (inp[1]) ? node2099 : node2094;
											assign node2094 = (inp[6]) ? 8'b00111110 : node2095;
												assign node2095 = (inp[2]) ? 8'b00111110 : 8'b00101111;
											assign node2099 = (inp[0]) ? node2101 : 8'b00101110;
												assign node2101 = (inp[5]) ? 8'b00101010 : 8'b00101011;
										assign node2104 = (inp[2]) ? node2110 : node2105;
											assign node2105 = (inp[1]) ? node2107 : 8'b00111011;
												assign node2107 = (inp[0]) ? 8'b00111010 : 8'b00111011;
											assign node2110 = (inp[5]) ? node2114 : node2111;
												assign node2111 = (inp[0]) ? 8'b00101011 : 8'b00111011;
												assign node2114 = (inp[0]) ? 8'b00101010 : 8'b00101011;
									assign node2117 = (inp[3]) ? node2127 : node2118;
										assign node2118 = (inp[5]) ? node2124 : node2119;
											assign node2119 = (inp[1]) ? node2121 : 8'b00101111;
												assign node2121 = (inp[2]) ? 8'b00101110 : 8'b00111110;
											assign node2124 = (inp[6]) ? 8'b00111011 : 8'b01111111;
										assign node2127 = (inp[6]) ? node2133 : node2128;
											assign node2128 = (inp[5]) ? 8'b00101110 : node2129;
												assign node2129 = (inp[2]) ? 8'b00111011 : 8'b00111110;
											assign node2133 = (inp[0]) ? 8'b00101110 : node2134;
												assign node2134 = (inp[5]) ? 8'b00101011 : 8'b00101110;
								assign node2138 = (inp[12]) ? node2160 : node2139;
									assign node2139 = (inp[5]) ? node2151 : node2140;
										assign node2140 = (inp[6]) ? node2144 : node2141;
											assign node2141 = (inp[0]) ? 8'b00001111 : 8'b00101011;
											assign node2144 = (inp[3]) ? 8'b00011011 : node2145;
												assign node2145 = (inp[1]) ? 8'b00011111 : node2146;
													assign node2146 = (inp[0]) ? 8'b00011110 : 8'b00111010;
										assign node2151 = (inp[0]) ? node2155 : node2152;
											assign node2152 = (inp[1]) ? 8'b00011110 : 8'b00001111;
											assign node2155 = (inp[1]) ? node2157 : 8'b00001110;
												assign node2157 = (inp[2]) ? 8'b00001010 : 8'b00001011;
									assign node2160 = (inp[6]) ? node2174 : node2161;
										assign node2161 = (inp[2]) ? node2169 : node2162;
											assign node2162 = (inp[1]) ? node2164 : 8'b00111010;
												assign node2164 = (inp[3]) ? node2166 : 8'b00111010;
													assign node2166 = (inp[5]) ? 8'b00011111 : 8'b00111010;
											assign node2169 = (inp[0]) ? 8'b00011010 : node2170;
												assign node2170 = (inp[1]) ? 8'b00101010 : 8'b00101011;
										assign node2174 = (inp[5]) ? node2176 : 8'b00101010;
											assign node2176 = (inp[3]) ? node2180 : node2177;
												assign node2177 = (inp[1]) ? 8'b00101010 : 8'b00101011;
												assign node2180 = (inp[1]) ? 8'b00001111 : 8'b00001110;
							assign node2183 = (inp[5]) ? node2235 : node2184;
								assign node2184 = (inp[8]) ? node2202 : node2185;
									assign node2185 = (inp[0]) ? node2197 : node2186;
										assign node2186 = (inp[12]) ? node2194 : node2187;
											assign node2187 = (inp[3]) ? node2191 : node2188;
												assign node2188 = (inp[1]) ? 8'b00011111 : 8'b00111010;
												assign node2191 = (inp[1]) ? 8'b00101010 : 8'b00011111;
											assign node2194 = (inp[6]) ? 8'b00101010 : 8'b00101011;
										assign node2197 = (inp[3]) ? 8'b00011111 : node2198;
											assign node2198 = (inp[12]) ? 8'b00001111 : 8'b00111010;
									assign node2202 = (inp[1]) ? node2220 : node2203;
										assign node2203 = (inp[3]) ? node2209 : node2204;
											assign node2204 = (inp[2]) ? 8'b00111010 : node2205;
												assign node2205 = (inp[0]) ? 8'b00101011 : 8'b00111011;
											assign node2209 = (inp[12]) ? node2215 : node2210;
												assign node2210 = (inp[6]) ? 8'b00011111 : node2211;
													assign node2211 = (inp[2]) ? 8'b00011111 : 8'b00101010;
												assign node2215 = (inp[6]) ? 8'b00101010 : node2216;
													assign node2216 = (inp[2]) ? 8'b00011111 : 8'b00111010;
										assign node2220 = (inp[2]) ? 8'b00101010 : node2221;
											assign node2221 = (inp[3]) ? node2227 : node2222;
												assign node2222 = (inp[0]) ? node2224 : 8'b00101010;
													assign node2224 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node2227 = (inp[0]) ? node2231 : node2228;
													assign node2228 = (inp[6]) ? 8'b00011111 : 8'b00101010;
													assign node2231 = (inp[12]) ? 8'b00101010 : 8'b00101010;
								assign node2235 = (inp[1]) ? node2269 : node2236;
									assign node2236 = (inp[8]) ? node2250 : node2237;
										assign node2237 = (inp[0]) ? node2245 : node2238;
											assign node2238 = (inp[12]) ? node2240 : 8'b00111010;
												assign node2240 = (inp[2]) ? 8'b00101011 : node2241;
													assign node2241 = (inp[3]) ? 8'b00111010 : 8'b00111011;
											assign node2245 = (inp[2]) ? 8'b00011111 : node2246;
												assign node2246 = (inp[12]) ? 8'b00111010 : 8'b00011111;
										assign node2250 = (inp[3]) ? node2258 : node2251;
											assign node2251 = (inp[12]) ? node2253 : 8'b00011110;
												assign node2253 = (inp[2]) ? node2255 : 8'b00001111;
													assign node2255 = (inp[0]) ? 8'b00011110 : 8'b00001110;
											assign node2258 = (inp[2]) ? node2264 : node2259;
												assign node2259 = (inp[12]) ? node2261 : 8'b00011011;
													assign node2261 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node2264 = (inp[6]) ? node2266 : 8'b00011011;
													assign node2266 = (inp[12]) ? 8'b00011011 : 8'b00001011;
									assign node2269 = (inp[8]) ? node2279 : node2270;
										assign node2270 = (inp[12]) ? node2276 : node2271;
											assign node2271 = (inp[2]) ? 8'b00001110 : node2272;
												assign node2272 = (inp[6]) ? 8'b00011110 : 8'b00001111;
											assign node2276 = (inp[0]) ? 8'b00011110 : 8'b00011111;
										assign node2279 = (inp[12]) ? node2285 : node2280;
											assign node2280 = (inp[0]) ? node2282 : 8'b00011010;
												assign node2282 = (inp[2]) ? 8'b00001010 : 8'b00001011;
											assign node2285 = (inp[2]) ? node2287 : 8'b00011110;
												assign node2287 = (inp[0]) ? 8'b00011010 : 8'b00011011;
					assign node2290 = (inp[8]) ? node2438 : node2291;
						assign node2291 = (inp[10]) ? node2363 : node2292;
							assign node2292 = (inp[11]) ? node2322 : node2293;
								assign node2293 = (inp[6]) ? node2309 : node2294;
									assign node2294 = (inp[0]) ? node2304 : node2295;
										assign node2295 = (inp[2]) ? 8'b00001110 : node2296;
											assign node2296 = (inp[12]) ? node2298 : 8'b00011110;
												assign node2298 = (inp[3]) ? node2300 : 8'b00011111;
													assign node2300 = (inp[1]) ? 8'b00011111 : 8'b00011110;
										assign node2304 = (inp[3]) ? node2306 : 8'b00011111;
											assign node2306 = (inp[5]) ? 8'b00011111 : 8'b00011110;
									assign node2309 = (inp[3]) ? 8'b00001110 : node2310;
										assign node2310 = (inp[5]) ? node2316 : node2311;
											assign node2311 = (inp[0]) ? 8'b00001111 : node2312;
												assign node2312 = (inp[1]) ? 8'b00001110 : 8'b00001111;
											assign node2316 = (inp[2]) ? node2318 : 8'b00001111;
												assign node2318 = (inp[0]) ? 8'b00011111 : 8'b00011110;
								assign node2322 = (inp[6]) ? node2350 : node2323;
									assign node2323 = (inp[12]) ? node2341 : node2324;
										assign node2324 = (inp[1]) ? node2332 : node2325;
											assign node2325 = (inp[5]) ? node2329 : node2326;
												assign node2326 = (inp[0]) ? 8'b00001110 : 8'b00011110;
												assign node2329 = (inp[3]) ? 8'b00001110 : 8'b00001111;
											assign node2332 = (inp[0]) ? node2336 : node2333;
												assign node2333 = (inp[2]) ? 8'b00011011 : 8'b00001110;
												assign node2336 = (inp[2]) ? node2338 : 8'b00001011;
													assign node2338 = (inp[3]) ? 8'b00001011 : 8'b00001010;
										assign node2341 = (inp[0]) ? node2345 : node2342;
											assign node2342 = (inp[1]) ? 8'b00011110 : 8'b00001111;
											assign node2345 = (inp[1]) ? 8'b00011010 : node2346;
												assign node2346 = (inp[3]) ? 8'b00011011 : 8'b00011110;
									assign node2350 = (inp[5]) ? node2354 : node2351;
										assign node2351 = (inp[12]) ? 8'b00001011 : 8'b00011011;
										assign node2354 = (inp[1]) ? node2358 : node2355;
											assign node2355 = (inp[2]) ? 8'b00011110 : 8'b00001110;
											assign node2358 = (inp[0]) ? 8'b00011010 : node2359;
												assign node2359 = (inp[3]) ? 8'b00011010 : 8'b00011011;
							assign node2363 = (inp[1]) ? node2395 : node2364;
								assign node2364 = (inp[3]) ? node2376 : node2365;
									assign node2365 = (inp[11]) ? node2367 : 8'b00001011;
										assign node2367 = (inp[2]) ? node2373 : node2368;
											assign node2368 = (inp[12]) ? node2370 : 8'b00011010;
												assign node2370 = (inp[6]) ? 8'b00001011 : 8'b00011011;
											assign node2373 = (inp[12]) ? 8'b00011010 : 8'b00001010;
									assign node2376 = (inp[11]) ? node2384 : node2377;
										assign node2377 = (inp[2]) ? node2381 : node2378;
											assign node2378 = (inp[6]) ? 8'b00000010 : 8'b00011010;
											assign node2381 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node2384 = (inp[2]) ? node2390 : node2385;
											assign node2385 = (inp[12]) ? node2387 : 8'b11110111;
												assign node2387 = (inp[6]) ? 8'b00000010 : 8'b00011010;
											assign node2390 = (inp[6]) ? 8'b11110111 : node2391;
												assign node2391 = (inp[12]) ? 8'b11110101 : 8'b10100101;
								assign node2395 = (inp[11]) ? node2419 : node2396;
									assign node2396 = (inp[0]) ? node2410 : node2397;
										assign node2397 = (inp[12]) ? node2405 : node2398;
											assign node2398 = (inp[5]) ? node2400 : 8'b10000010;
												assign node2400 = (inp[6]) ? 8'b10010001 : node2401;
													assign node2401 = (inp[2]) ? 8'b10000010 : 8'b00011010;
											assign node2405 = (inp[3]) ? node2407 : 8'b00000010;
												assign node2407 = (inp[2]) ? 8'b00000010 : 8'b00011010;
										assign node2410 = (inp[6]) ? 8'b10000001 : node2411;
											assign node2411 = (inp[2]) ? 8'b10010001 : node2412;
												assign node2412 = (inp[5]) ? 8'b10011001 : node2413;
													assign node2413 = (inp[3]) ? 8'b00011010 : 8'b10011001;
									assign node2419 = (inp[12]) ? node2431 : node2420;
										assign node2420 = (inp[6]) ? node2424 : node2421;
											assign node2421 = (inp[3]) ? 8'b11110111 : 8'b10101101;
											assign node2424 = (inp[5]) ? node2426 : 8'b10110100;
												assign node2426 = (inp[3]) ? 8'b10100100 : node2427;
													assign node2427 = (inp[0]) ? 8'b10100100 : 8'b10100101;
										assign node2431 = (inp[5]) ? node2433 : 8'b00000010;
											assign node2433 = (inp[3]) ? node2435 : 8'b00011010;
												assign node2435 = (inp[2]) ? 8'b10110100 : 8'b11111101;
						assign node2438 = (inp[5]) ? node2514 : node2439;
							assign node2439 = (inp[0]) ? node2461 : node2440;
								assign node2440 = (inp[6]) ? node2452 : node2441;
									assign node2441 = (inp[2]) ? node2449 : node2442;
										assign node2442 = (inp[1]) ? 8'b00011010 : node2443;
											assign node2443 = (inp[3]) ? 8'b00011010 : node2444;
												assign node2444 = (inp[11]) ? 8'b00001011 : 8'b00011011;
										assign node2449 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node2452 = (inp[12]) ? 8'b00000010 : node2453;
										assign node2453 = (inp[11]) ? node2455 : 8'b10000010;
											assign node2455 = (inp[3]) ? 8'b11110111 : node2456;
												assign node2456 = (inp[1]) ? 8'b11110111 : 8'b00011010;
								assign node2461 = (inp[10]) ? node2485 : node2462;
									assign node2462 = (inp[11]) ? node2472 : node2463;
										assign node2463 = (inp[1]) ? node2467 : node2464;
											assign node2464 = (inp[6]) ? 8'b10001101 : 8'b10011101;
											assign node2467 = (inp[6]) ? node2469 : 8'b10010100;
												assign node2469 = (inp[3]) ? 8'b10000100 : 8'b10000101;
										assign node2472 = (inp[2]) ? node2480 : node2473;
											assign node2473 = (inp[3]) ? node2475 : 8'b10111001;
												assign node2475 = (inp[6]) ? 8'b10100100 : node2476;
													assign node2476 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node2480 = (inp[6]) ? 8'b10100100 : node2481;
												assign node2481 = (inp[12]) ? 8'b10110001 : 8'b10100001;
									assign node2485 = (inp[1]) ? node2499 : node2486;
										assign node2486 = (inp[3]) ? node2494 : node2487;
											assign node2487 = (inp[11]) ? node2491 : node2488;
												assign node2488 = (inp[6]) ? 8'b00001011 : 8'b00011011;
												assign node2491 = (inp[12]) ? 8'b00011011 : 8'b00011010;
											assign node2494 = (inp[2]) ? node2496 : 8'b00011010;
												assign node2496 = (inp[11]) ? 8'b00000010 : 8'b10000010;
										assign node2499 = (inp[11]) ? node2511 : node2500;
											assign node2500 = (inp[3]) ? node2506 : node2501;
												assign node2501 = (inp[6]) ? 8'b10000001 : node2502;
													assign node2502 = (inp[2]) ? 8'b10010001 : 8'b10011001;
												assign node2506 = (inp[6]) ? node2508 : 8'b10010000;
													assign node2508 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node2511 = (inp[6]) ? 8'b10110100 : 8'b10100101;
							assign node2514 = (inp[11]) ? node2552 : node2515;
								assign node2515 = (inp[2]) ? node2535 : node2516;
									assign node2516 = (inp[6]) ? node2524 : node2517;
										assign node2517 = (inp[10]) ? node2521 : node2518;
											assign node2518 = (inp[0]) ? 8'b10011101 : 8'b00011010;
											assign node2521 = (inp[1]) ? 8'b10011101 : 8'b10011100;
										assign node2524 = (inp[3]) ? node2528 : node2525;
											assign node2525 = (inp[1]) ? 8'b10000100 : 8'b10001101;
											assign node2528 = (inp[1]) ? 8'b10000101 : node2529;
												assign node2529 = (inp[0]) ? 8'b10000100 : node2530;
													assign node2530 = (inp[10]) ? 8'b10000100 : 8'b10000010;
									assign node2535 = (inp[10]) ? node2549 : node2536;
										assign node2536 = (inp[0]) ? node2546 : node2537;
											assign node2537 = (inp[6]) ? node2541 : node2538;
												assign node2538 = (inp[1]) ? 8'b10000001 : 8'b10000010;
												assign node2541 = (inp[1]) ? node2543 : 8'b10010000;
													assign node2543 = (inp[3]) ? 8'b10010001 : 8'b10010000;
											assign node2546 = (inp[1]) ? 8'b10010101 : 8'b10010100;
										assign node2549 = (inp[6]) ? 8'b10010100 : 8'b10000100;
								assign node2552 = (inp[1]) ? node2582 : node2553;
									assign node2553 = (inp[3]) ? node2567 : node2554;
										assign node2554 = (inp[2]) ? node2558 : node2555;
											assign node2555 = (inp[6]) ? 8'b10101101 : 8'b11111101;
											assign node2558 = (inp[10]) ? node2562 : node2559;
												assign node2559 = (inp[6]) ? 8'b00011010 : 8'b10101100;
												assign node2562 = (inp[6]) ? 8'b10101100 : node2563;
													assign node2563 = (inp[0]) ? 8'b10111100 : 8'b10101100;
										assign node2567 = (inp[0]) ? node2575 : node2568;
											assign node2568 = (inp[10]) ? 8'b10101100 : node2569;
												assign node2569 = (inp[2]) ? node2571 : 8'b11110111;
													assign node2571 = (inp[6]) ? 8'b10100101 : 8'b11110111;
											assign node2575 = (inp[2]) ? node2579 : node2576;
												assign node2576 = (inp[10]) ? 8'b10111100 : 8'b10110001;
												assign node2579 = (inp[12]) ? 8'b10110001 : 8'b10100001;
									assign node2582 = (inp[0]) ? node2598 : node2583;
										assign node2583 = (inp[10]) ? node2591 : node2584;
											assign node2584 = (inp[6]) ? 8'b10110100 : node2585;
												assign node2585 = (inp[2]) ? 8'b10100101 : node2586;
													assign node2586 = (inp[12]) ? 8'b11111101 : 8'b10101101;
											assign node2591 = (inp[12]) ? node2595 : node2592;
												assign node2592 = (inp[3]) ? 8'b10110000 : 8'b10110001;
												assign node2595 = (inp[3]) ? 8'b10100001 : 8'b10110001;
										assign node2598 = (inp[2]) ? node2602 : node2599;
											assign node2599 = (inp[12]) ? 8'b10100001 : 8'b10110000;
											assign node2602 = (inp[12]) ? 8'b10110000 : 8'b10100000;
				assign node2605 = (inp[5]) ? node2899 : node2606;
					assign node2606 = (inp[0]) ? node2714 : node2607;
						assign node2607 = (inp[12]) ? node2673 : node2608;
							assign node2608 = (inp[11]) ? node2642 : node2609;
								assign node2609 = (inp[10]) ? node2625 : node2610;
									assign node2610 = (inp[8]) ? node2620 : node2611;
										assign node2611 = (inp[6]) ? node2615 : node2612;
											assign node2612 = (inp[2]) ? 8'b00001110 : 8'b00011110;
											assign node2615 = (inp[9]) ? 8'b00001110 : node2616;
												assign node2616 = (inp[3]) ? 8'b00001110 : 8'b00001111;
										assign node2620 = (inp[3]) ? 8'b10000010 : node2621;
											assign node2621 = (inp[9]) ? 8'b10000010 : 8'b00001011;
									assign node2625 = (inp[2]) ? node2637 : node2626;
										assign node2626 = (inp[6]) ? node2632 : node2627;
											assign node2627 = (inp[3]) ? 8'b00011010 : node2628;
												assign node2628 = (inp[1]) ? 8'b00011010 : 8'b00011011;
											assign node2632 = (inp[1]) ? 8'b10000010 : node2633;
												assign node2633 = (inp[3]) ? 8'b10000010 : 8'b00001011;
										assign node2637 = (inp[1]) ? 8'b10000010 : node2638;
											assign node2638 = (inp[3]) ? 8'b10000010 : 8'b00001011;
								assign node2642 = (inp[10]) ? node2660 : node2643;
									assign node2643 = (inp[3]) ? node2653 : node2644;
										assign node2644 = (inp[1]) ? node2648 : node2645;
											assign node2645 = (inp[8]) ? 8'b00011010 : 8'b00011110;
											assign node2648 = (inp[6]) ? 8'b00011011 : node2649;
												assign node2649 = (inp[2]) ? 8'b00011011 : 8'b00001110;
										assign node2653 = (inp[6]) ? node2657 : node2654;
											assign node2654 = (inp[8]) ? 8'b00001010 : 8'b00011011;
											assign node2657 = (inp[8]) ? 8'b11110111 : 8'b00011011;
									assign node2660 = (inp[1]) ? 8'b11110111 : node2661;
										assign node2661 = (inp[3]) ? node2667 : node2662;
											assign node2662 = (inp[6]) ? 8'b00011010 : node2663;
												assign node2663 = (inp[2]) ? 8'b00011010 : 8'b00001011;
											assign node2667 = (inp[6]) ? 8'b11110111 : node2668;
												assign node2668 = (inp[9]) ? 8'b11110111 : 8'b00001010;
							assign node2673 = (inp[2]) ? node2701 : node2674;
								assign node2674 = (inp[6]) ? node2688 : node2675;
									assign node2675 = (inp[3]) ? node2683 : node2676;
										assign node2676 = (inp[1]) ? 8'b00011110 : node2677;
											assign node2677 = (inp[8]) ? 8'b00011011 : node2678;
												assign node2678 = (inp[10]) ? 8'b00011011 : 8'b00011111;
										assign node2683 = (inp[8]) ? 8'b00011010 : node2684;
											assign node2684 = (inp[9]) ? 8'b00011110 : 8'b00011010;
									assign node2688 = (inp[8]) ? node2696 : node2689;
										assign node2689 = (inp[10]) ? 8'b00001011 : node2690;
											assign node2690 = (inp[1]) ? 8'b00001110 : node2691;
												assign node2691 = (inp[9]) ? 8'b00001111 : 8'b00001110;
										assign node2696 = (inp[1]) ? 8'b00000010 : node2697;
											assign node2697 = (inp[3]) ? 8'b00000010 : 8'b00001011;
								assign node2701 = (inp[8]) ? node2709 : node2702;
									assign node2702 = (inp[10]) ? node2704 : 8'b00001110;
										assign node2704 = (inp[1]) ? 8'b00000010 : node2705;
											assign node2705 = (inp[3]) ? 8'b00000010 : 8'b00001011;
									assign node2709 = (inp[1]) ? 8'b00000010 : node2710;
										assign node2710 = (inp[3]) ? 8'b00000010 : 8'b00001011;
						assign node2714 = (inp[9]) ? node2804 : node2715;
							assign node2715 = (inp[6]) ? node2765 : node2716;
								assign node2716 = (inp[10]) ? node2746 : node2717;
									assign node2717 = (inp[12]) ? node2725 : node2718;
										assign node2718 = (inp[11]) ? node2720 : 8'b10111100;
											assign node2720 = (inp[2]) ? 8'b10101001 : node2721;
												assign node2721 = (inp[8]) ? 8'b10001100 : 8'b10101100;
										assign node2725 = (inp[3]) ? node2735 : node2726;
											assign node2726 = (inp[2]) ? node2732 : node2727;
												assign node2727 = (inp[8]) ? node2729 : 8'b11111101;
													assign node2729 = (inp[11]) ? 8'b10011101 : 8'b11111101;
												assign node2732 = (inp[8]) ? 8'b10011100 : 8'b10111100;
											assign node2735 = (inp[11]) ? node2741 : node2736;
												assign node2736 = (inp[8]) ? node2738 : 8'b10111100;
													assign node2738 = (inp[2]) ? 8'b10110100 : 8'b10111100;
												assign node2741 = (inp[2]) ? 8'b10111001 : node2742;
													assign node2742 = (inp[8]) ? 8'b10011100 : 8'b10111100;
									assign node2746 = (inp[2]) ? node2756 : node2747;
										assign node2747 = (inp[3]) ? node2751 : node2748;
											assign node2748 = (inp[11]) ? 8'b10101001 : 8'b10111001;
											assign node2751 = (inp[12]) ? 8'b10111000 : node2752;
												assign node2752 = (inp[11]) ? 8'b10101000 : 8'b10111000;
										assign node2756 = (inp[11]) ? node2758 : 8'b10110001;
											assign node2758 = (inp[3]) ? 8'b10000101 : node2759;
												assign node2759 = (inp[1]) ? 8'b10000100 : node2760;
													assign node2760 = (inp[12]) ? 8'b10111000 : 8'b10101000;
								assign node2765 = (inp[11]) ? node2781 : node2766;
									assign node2766 = (inp[3]) ? node2776 : node2767;
										assign node2767 = (inp[10]) ? node2773 : node2768;
											assign node2768 = (inp[8]) ? node2770 : 8'b10101101;
												assign node2770 = (inp[1]) ? 8'b10100101 : 8'b10101101;
											assign node2773 = (inp[1]) ? 8'b10100001 : 8'b10101001;
										assign node2776 = (inp[10]) ? 8'b10100000 : node2777;
											assign node2777 = (inp[8]) ? 8'b10100100 : 8'b10101100;
									assign node2781 = (inp[12]) ? node2793 : node2782;
										assign node2782 = (inp[3]) ? node2790 : node2783;
											assign node2783 = (inp[8]) ? node2787 : node2784;
												assign node2784 = (inp[10]) ? 8'b10111000 : 8'b10111100;
												assign node2787 = (inp[2]) ? 8'b10010000 : 8'b10010100;
											assign node2790 = (inp[10]) ? 8'b10010101 : 8'b10010001;
										assign node2793 = (inp[3]) ? node2799 : node2794;
											assign node2794 = (inp[1]) ? node2796 : 8'b10001101;
												assign node2796 = (inp[2]) ? 8'b10000101 : 8'b10000001;
											assign node2799 = (inp[10]) ? 8'b10100000 : node2800;
												assign node2800 = (inp[8]) ? 8'b10000100 : 8'b10101100;
							assign node2804 = (inp[8]) ? node2848 : node2805;
								assign node2805 = (inp[10]) ? node2827 : node2806;
									assign node2806 = (inp[6]) ? node2816 : node2807;
										assign node2807 = (inp[3]) ? node2811 : node2808;
											assign node2808 = (inp[2]) ? 8'b00011010 : 8'b00011111;
											assign node2811 = (inp[11]) ? node2813 : 8'b00011110;
												assign node2813 = (inp[12]) ? 8'b00011110 : 8'b00001110;
										assign node2816 = (inp[12]) ? node2822 : node2817;
											assign node2817 = (inp[3]) ? 8'b00011011 : node2818;
												assign node2818 = (inp[11]) ? 8'b00011110 : 8'b00001111;
											assign node2822 = (inp[3]) ? 8'b00001110 : node2823;
												assign node2823 = (inp[11]) ? 8'b00001011 : 8'b00001111;
									assign node2827 = (inp[6]) ? node2837 : node2828;
										assign node2828 = (inp[3]) ? node2832 : node2829;
											assign node2829 = (inp[1]) ? 8'b10011001 : 8'b00011011;
											assign node2832 = (inp[1]) ? node2834 : 8'b00011010;
												assign node2834 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node2837 = (inp[12]) ? node2845 : node2838;
											assign node2838 = (inp[11]) ? node2842 : node2839;
												assign node2839 = (inp[3]) ? 8'b10000010 : 8'b10000001;
												assign node2842 = (inp[1]) ? 8'b11110111 : 8'b00011010;
											assign node2845 = (inp[3]) ? 8'b00000010 : 8'b10000001;
								assign node2848 = (inp[11]) ? node2866 : node2849;
									assign node2849 = (inp[10]) ? node2853 : node2850;
										assign node2850 = (inp[6]) ? 8'b10001101 : 8'b10011101;
										assign node2853 = (inp[1]) ? node2861 : node2854;
											assign node2854 = (inp[3]) ? node2858 : node2855;
												assign node2855 = (inp[12]) ? 8'b00001011 : 8'b00011011;
												assign node2858 = (inp[2]) ? 8'b10010000 : 8'b00011010;
											assign node2861 = (inp[6]) ? 8'b10000001 : node2862;
												assign node2862 = (inp[2]) ? 8'b10010001 : 8'b10011001;
									assign node2866 = (inp[2]) ? node2880 : node2867;
										assign node2867 = (inp[1]) ? node2871 : node2868;
											assign node2868 = (inp[6]) ? 8'b00001011 : 8'b00011011;
											assign node2871 = (inp[3]) ? node2877 : node2872;
												assign node2872 = (inp[6]) ? 8'b10100001 : node2873;
													assign node2873 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node2877 = (inp[10]) ? 8'b00011010 : 8'b10111100;
										assign node2880 = (inp[3]) ? node2892 : node2881;
											assign node2881 = (inp[1]) ? node2887 : node2882;
												assign node2882 = (inp[10]) ? 8'b00011010 : node2883;
													assign node2883 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node2887 = (inp[6]) ? 8'b10100101 : node2888;
													assign node2888 = (inp[10]) ? 8'b10110100 : 8'b10100000;
											assign node2892 = (inp[6]) ? 8'b10100100 : node2893;
												assign node2893 = (inp[12]) ? node2895 : 8'b10100101;
													assign node2895 = (inp[1]) ? 8'b10110001 : 8'b11110101;
					assign node2899 = (inp[11]) ? node3063 : node2900;
						assign node2900 = (inp[0]) ? node3010 : node2901;
							assign node2901 = (inp[9]) ? node2959 : node2902;
								assign node2902 = (inp[8]) ? node2922 : node2903;
									assign node2903 = (inp[10]) ? node2911 : node2904;
										assign node2904 = (inp[6]) ? node2908 : node2905;
											assign node2905 = (inp[2]) ? 8'b00001111 : 8'b00011110;
											assign node2908 = (inp[2]) ? 8'b00011110 : 8'b00001110;
										assign node2911 = (inp[3]) ? node2917 : node2912;
											assign node2912 = (inp[2]) ? 8'b00011011 : node2913;
												assign node2913 = (inp[6]) ? 8'b00000010 : 8'b00011010;
											assign node2917 = (inp[6]) ? node2919 : 8'b00000010;
												assign node2919 = (inp[1]) ? 8'b10010001 : 8'b10010000;
									assign node2922 = (inp[10]) ? node2940 : node2923;
										assign node2923 = (inp[3]) ? node2931 : node2924;
											assign node2924 = (inp[1]) ? node2928 : node2925;
												assign node2925 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node2928 = (inp[6]) ? 8'b10000010 : 8'b00011010;
											assign node2931 = (inp[1]) ? node2935 : node2932;
												assign node2932 = (inp[12]) ? 8'b00011010 : 8'b10000010;
												assign node2935 = (inp[2]) ? node2937 : 8'b10011001;
													assign node2937 = (inp[6]) ? 8'b10010001 : 8'b10000001;
										assign node2940 = (inp[1]) ? node2950 : node2941;
											assign node2941 = (inp[3]) ? node2947 : node2942;
												assign node2942 = (inp[12]) ? node2944 : 8'b10001101;
													assign node2944 = (inp[6]) ? 8'b10001101 : 8'b10011101;
												assign node2947 = (inp[12]) ? 8'b10000100 : 8'b10011100;
											assign node2950 = (inp[3]) ? node2956 : node2951;
												assign node2951 = (inp[12]) ? node2953 : 8'b10000100;
													assign node2953 = (inp[6]) ? 8'b10000100 : 8'b10011100;
												assign node2956 = (inp[12]) ? 8'b10010101 : 8'b10000101;
								assign node2959 = (inp[6]) ? node2981 : node2960;
									assign node2960 = (inp[2]) ? node2972 : node2961;
										assign node2961 = (inp[8]) ? node2969 : node2962;
											assign node2962 = (inp[10]) ? 8'b10111001 : node2963;
												assign node2963 = (inp[1]) ? 8'b11111101 : node2964;
													assign node2964 = (inp[3]) ? 8'b10111100 : 8'b11111101;
											assign node2969 = (inp[1]) ? 8'b10111000 : 8'b10111001;
										assign node2972 = (inp[3]) ? node2976 : node2973;
											assign node2973 = (inp[10]) ? 8'b10101101 : 8'b10101001;
											assign node2976 = (inp[10]) ? node2978 : 8'b10100001;
												assign node2978 = (inp[8]) ? 8'b10100100 : 8'b10100000;
									assign node2981 = (inp[2]) ? node2993 : node2982;
										assign node2982 = (inp[10]) ? node2990 : node2983;
											assign node2983 = (inp[8]) ? node2987 : node2984;
												assign node2984 = (inp[1]) ? 8'b10101100 : 8'b10101101;
												assign node2987 = (inp[3]) ? 8'b10100000 : 8'b10101001;
											assign node2990 = (inp[8]) ? 8'b10100100 : 8'b10100000;
										assign node2993 = (inp[3]) ? node3001 : node2994;
											assign node2994 = (inp[10]) ? node2998 : node2995;
												assign node2995 = (inp[8]) ? 8'b10110000 : 8'b10111100;
												assign node2998 = (inp[8]) ? 8'b10110100 : 8'b10110000;
											assign node3001 = (inp[1]) ? node3005 : node3002;
												assign node3002 = (inp[10]) ? 8'b10110100 : 8'b10110000;
												assign node3005 = (inp[10]) ? node3007 : 8'b11111101;
													assign node3007 = (inp[8]) ? 8'b11110101 : 8'b10110001;
							assign node3010 = (inp[3]) ? node3032 : node3011;
								assign node3011 = (inp[2]) ? node3021 : node3012;
									assign node3012 = (inp[6]) ? node3014 : 8'b11111101;
										assign node3014 = (inp[1]) ? node3016 : 8'b10101101;
											assign node3016 = (inp[10]) ? node3018 : 8'b10101101;
												assign node3018 = (inp[8]) ? 8'b10100101 : 8'b10100001;
									assign node3021 = (inp[1]) ? node3027 : node3022;
										assign node3022 = (inp[10]) ? node3024 : 8'b11111101;
											assign node3024 = (inp[8]) ? 8'b11111101 : 8'b10111001;
										assign node3027 = (inp[8]) ? 8'b11110101 : node3028;
											assign node3028 = (inp[10]) ? 8'b10110001 : 8'b11111101;
								assign node3032 = (inp[1]) ? node3046 : node3033;
									assign node3033 = (inp[8]) ? node3043 : node3034;
										assign node3034 = (inp[10]) ? node3040 : node3035;
											assign node3035 = (inp[2]) ? 8'b10111100 : node3036;
												assign node3036 = (inp[6]) ? 8'b10101100 : 8'b10111100;
											assign node3040 = (inp[12]) ? 8'b10110000 : 8'b10111000;
										assign node3043 = (inp[2]) ? 8'b10110100 : 8'b10100100;
									assign node3046 = (inp[8]) ? node3056 : node3047;
										assign node3047 = (inp[10]) ? node3051 : node3048;
											assign node3048 = (inp[6]) ? 8'b10101101 : 8'b11111101;
											assign node3051 = (inp[12]) ? node3053 : 8'b10100001;
												assign node3053 = (inp[2]) ? 8'b10110001 : 8'b10111001;
										assign node3056 = (inp[6]) ? node3060 : node3057;
											assign node3057 = (inp[2]) ? 8'b11110101 : 8'b11111101;
											assign node3060 = (inp[2]) ? 8'b11110101 : 8'b10100101;
						assign node3063 = (inp[8]) ? node3145 : node3064;
							assign node3064 = (inp[10]) ? node3102 : node3065;
								assign node3065 = (inp[0]) ? node3087 : node3066;
									assign node3066 = (inp[9]) ? node3080 : node3067;
										assign node3067 = (inp[3]) ? node3073 : node3068;
											assign node3068 = (inp[12]) ? node3070 : 8'b00011011;
												assign node3070 = (inp[1]) ? 8'b00001110 : 8'b00001111;
											assign node3073 = (inp[2]) ? node3075 : 8'b00001110;
												assign node3075 = (inp[12]) ? 8'b00011011 : node3076;
													assign node3076 = (inp[6]) ? 8'b00001011 : 8'b00011011;
										assign node3080 = (inp[12]) ? 8'b10111100 : node3081;
											assign node3081 = (inp[1]) ? 8'b10101001 : node3082;
												assign node3082 = (inp[6]) ? 8'b10111100 : 8'b10111001;
									assign node3087 = (inp[2]) ? node3093 : node3088;
										assign node3088 = (inp[6]) ? node3090 : 8'b10111001;
											assign node3090 = (inp[1]) ? 8'b10111000 : 8'b10111001;
										assign node3093 = (inp[12]) ? node3099 : node3094;
											assign node3094 = (inp[1]) ? 8'b10101000 : node3095;
												assign node3095 = (inp[3]) ? 8'b10101001 : 8'b10101100;
											assign node3099 = (inp[1]) ? 8'b10111000 : 8'b10111100;
								assign node3102 = (inp[3]) ? node3122 : node3103;
									assign node3103 = (inp[1]) ? node3115 : node3104;
										assign node3104 = (inp[12]) ? node3112 : node3105;
											assign node3105 = (inp[6]) ? 8'b10111000 : node3106;
												assign node3106 = (inp[0]) ? node3108 : 8'b10111000;
													assign node3108 = (inp[2]) ? 8'b10101000 : 8'b10101001;
											assign node3112 = (inp[2]) ? 8'b10101001 : 8'b10111001;
										assign node3115 = (inp[6]) ? node3119 : node3116;
											assign node3116 = (inp[9]) ? 8'b10100000 : 8'b00000010;
											assign node3119 = (inp[0]) ? 8'b10010100 : 8'b11110101;
									assign node3122 = (inp[12]) ? node3134 : node3123;
										assign node3123 = (inp[2]) ? node3129 : node3124;
											assign node3124 = (inp[6]) ? node3126 : 8'b00001010;
												assign node3126 = (inp[1]) ? 8'b10010100 : 8'b10010101;
											assign node3129 = (inp[0]) ? 8'b10000101 : node3130;
												assign node3130 = (inp[6]) ? 8'b10000101 : 8'b10010101;
										assign node3134 = (inp[0]) ? node3140 : node3135;
											assign node3135 = (inp[9]) ? 8'b10011101 : node3136;
												assign node3136 = (inp[2]) ? 8'b11110101 : 8'b11111101;
											assign node3140 = (inp[2]) ? node3142 : 8'b10111000;
												assign node3142 = (inp[1]) ? 8'b10010100 : 8'b10010101;
							assign node3145 = (inp[0]) ? node3205 : node3146;
								assign node3146 = (inp[9]) ? node3174 : node3147;
									assign node3147 = (inp[6]) ? node3163 : node3148;
										assign node3148 = (inp[2]) ? node3156 : node3149;
											assign node3149 = (inp[12]) ? 8'b10111100 : node3150;
												assign node3150 = (inp[10]) ? node3152 : 8'b10101101;
													assign node3152 = (inp[1]) ? 8'b10101001 : 8'b10101101;
											assign node3156 = (inp[10]) ? node3158 : 8'b00011010;
												assign node3158 = (inp[3]) ? node3160 : 8'b10101101;
													assign node3160 = (inp[12]) ? 8'b10100001 : 8'b10110001;
										assign node3163 = (inp[2]) ? node3169 : node3164;
											assign node3164 = (inp[12]) ? node3166 : 8'b11110111;
												assign node3166 = (inp[10]) ? 8'b10100100 : 8'b00000010;
											assign node3169 = (inp[1]) ? node3171 : 8'b11110101;
												assign node3171 = (inp[3]) ? 8'b10110100 : 8'b10110001;
									assign node3174 = (inp[2]) ? node3192 : node3175;
										assign node3175 = (inp[6]) ? node3185 : node3176;
											assign node3176 = (inp[10]) ? node3182 : node3177;
												assign node3177 = (inp[3]) ? 8'b10111000 : node3178;
													assign node3178 = (inp[1]) ? 8'b10111000 : 8'b10111001;
												assign node3182 = (inp[1]) ? 8'b10001100 : 8'b10011100;
											assign node3185 = (inp[1]) ? node3189 : node3186;
												assign node3186 = (inp[3]) ? 8'b10100000 : 8'b10101001;
												assign node3189 = (inp[12]) ? 8'b10000101 : 8'b10010001;
										assign node3192 = (inp[1]) ? node3200 : node3193;
											assign node3193 = (inp[3]) ? node3195 : 8'b10101000;
												assign node3195 = (inp[6]) ? 8'b10010101 : node3196;
													assign node3196 = (inp[12]) ? 8'b10100000 : 8'b10010101;
											assign node3200 = (inp[10]) ? node3202 : 8'b10010101;
												assign node3202 = (inp[12]) ? 8'b10000001 : 8'b10010001;
								assign node3205 = (inp[1]) ? node3223 : node3206;
									assign node3206 = (inp[3]) ? node3214 : node3207;
										assign node3207 = (inp[2]) ? node3211 : node3208;
											assign node3208 = (inp[6]) ? 8'b10001101 : 8'b10011101;
											assign node3211 = (inp[12]) ? 8'b10011100 : 8'b10001100;
										assign node3214 = (inp[2]) ? node3220 : node3215;
											assign node3215 = (inp[6]) ? 8'b10000100 : node3216;
												assign node3216 = (inp[12]) ? 8'b10011100 : 8'b10001100;
											assign node3220 = (inp[12]) ? 8'b10010001 : 8'b10000001;
									assign node3223 = (inp[2]) ? node3229 : node3224;
										assign node3224 = (inp[6]) ? 8'b10000001 : node3225;
											assign node3225 = (inp[12]) ? 8'b10011001 : 8'b10001001;
										assign node3229 = (inp[12]) ? 8'b10010000 : 8'b10000000;
			assign node3232 = (inp[11]) ? node3512 : node3233;
				assign node3233 = (inp[5]) ? node3349 : node3234;
					assign node3234 = (inp[0]) ? node3238 : node3235;
						assign node3235 = (inp[12]) ? 8'b00000010 : 8'b10000010;
						assign node3238 = (inp[13]) ? node3290 : node3239;
							assign node3239 = (inp[3]) ? node3263 : node3240;
								assign node3240 = (inp[1]) ? node3254 : node3241;
									assign node3241 = (inp[2]) ? node3249 : node3242;
										assign node3242 = (inp[12]) ? 8'b00000010 : node3243;
											assign node3243 = (inp[6]) ? node3245 : 8'b10000010;
												assign node3245 = (inp[9]) ? 8'b10000100 : 8'b10000010;
										assign node3249 = (inp[6]) ? node3251 : 8'b10010000;
											assign node3251 = (inp[10]) ? 8'b10000010 : 8'b10000100;
									assign node3254 = (inp[2]) ? node3260 : node3255;
										assign node3255 = (inp[10]) ? 8'b10000001 : node3256;
											assign node3256 = (inp[8]) ? 8'b10000101 : 8'b10000001;
										assign node3260 = (inp[6]) ? 8'b10000001 : 8'b10010001;
								assign node3263 = (inp[6]) ? node3279 : node3264;
									assign node3264 = (inp[2]) ? node3272 : node3265;
										assign node3265 = (inp[8]) ? node3269 : node3266;
											assign node3266 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node3269 = (inp[10]) ? 8'b10000010 : 8'b10000100;
										assign node3272 = (inp[1]) ? node3274 : 8'b10010000;
											assign node3274 = (inp[12]) ? node3276 : 8'b10010000;
												assign node3276 = (inp[10]) ? 8'b10010000 : 8'b10010100;
									assign node3279 = (inp[12]) ? node3285 : node3280;
										assign node3280 = (inp[8]) ? node3282 : 8'b10000010;
											assign node3282 = (inp[10]) ? 8'b10000010 : 8'b10000100;
										assign node3285 = (inp[10]) ? 8'b00000010 : node3286;
											assign node3286 = (inp[8]) ? 8'b10000100 : 8'b00000010;
							assign node3290 = (inp[9]) ? node3318 : node3291;
								assign node3291 = (inp[8]) ? node3305 : node3292;
									assign node3292 = (inp[6]) ? node3300 : node3293;
										assign node3293 = (inp[2]) ? node3295 : 8'b10100000;
											assign node3295 = (inp[1]) ? node3297 : 8'b10110000;
												assign node3297 = (inp[3]) ? 8'b10110000 : 8'b10110001;
										assign node3300 = (inp[3]) ? 8'b10100000 : node3301;
											assign node3301 = (inp[1]) ? 8'b10100001 : 8'b10100000;
									assign node3305 = (inp[10]) ? node3313 : node3306;
										assign node3306 = (inp[3]) ? 8'b10100100 : node3307;
											assign node3307 = (inp[2]) ? 8'b11110101 : node3308;
												assign node3308 = (inp[1]) ? 8'b10100101 : 8'b10100100;
										assign node3313 = (inp[6]) ? 8'b10100000 : node3314;
											assign node3314 = (inp[2]) ? 8'b10110000 : 8'b10100001;
								assign node3318 = (inp[10]) ? node3332 : node3319;
									assign node3319 = (inp[8]) ? node3325 : node3320;
										assign node3320 = (inp[1]) ? node3322 : 8'b10000010;
											assign node3322 = (inp[12]) ? 8'b10000001 : 8'b10010000;
										assign node3325 = (inp[3]) ? node3329 : node3326;
											assign node3326 = (inp[1]) ? 8'b10000101 : 8'b10000100;
											assign node3329 = (inp[12]) ? 8'b10000100 : 8'b10010100;
									assign node3332 = (inp[3]) ? node3342 : node3333;
										assign node3333 = (inp[1]) ? 8'b10000001 : node3334;
											assign node3334 = (inp[6]) ? node3338 : node3335;
												assign node3335 = (inp[2]) ? 8'b10010000 : 8'b10000010;
												assign node3338 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node3342 = (inp[12]) ? node3344 : 8'b10000010;
											assign node3344 = (inp[2]) ? node3346 : 8'b00000010;
												assign node3346 = (inp[6]) ? 8'b00000010 : 8'b10010000;
					assign node3349 = (inp[8]) ? node3421 : node3350;
						assign node3350 = (inp[13]) ? node3376 : node3351;
							assign node3351 = (inp[1]) ? node3363 : node3352;
								assign node3352 = (inp[2]) ? node3356 : node3353;
									assign node3353 = (inp[12]) ? 8'b00000010 : 8'b10000010;
									assign node3356 = (inp[6]) ? 8'b10010000 : node3357;
										assign node3357 = (inp[0]) ? 8'b10010000 : node3358;
											assign node3358 = (inp[9]) ? 8'b10000010 : 8'b00000010;
								assign node3363 = (inp[0]) ? node3373 : node3364;
									assign node3364 = (inp[3]) ? node3368 : node3365;
										assign node3365 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node3368 = (inp[6]) ? node3370 : 8'b10000001;
											assign node3370 = (inp[2]) ? 8'b10010001 : 8'b10000001;
									assign node3373 = (inp[2]) ? 8'b10010001 : 8'b10000001;
							assign node3376 = (inp[2]) ? node3396 : node3377;
								assign node3377 = (inp[9]) ? node3389 : node3378;
									assign node3378 = (inp[0]) ? node3386 : node3379;
										assign node3379 = (inp[1]) ? node3383 : node3380;
											assign node3380 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node3383 = (inp[3]) ? 8'b10000001 : 8'b10000010;
										assign node3386 = (inp[1]) ? 8'b10100001 : 8'b10100000;
									assign node3389 = (inp[1]) ? node3391 : 8'b10100000;
										assign node3391 = (inp[3]) ? 8'b10100001 : node3392;
											assign node3392 = (inp[0]) ? 8'b10100001 : 8'b10100000;
								assign node3396 = (inp[1]) ? node3406 : node3397;
									assign node3397 = (inp[0]) ? 8'b10110000 : node3398;
										assign node3398 = (inp[6]) ? node3402 : node3399;
											assign node3399 = (inp[9]) ? 8'b10100000 : 8'b00000010;
											assign node3402 = (inp[9]) ? 8'b10110000 : 8'b10010000;
									assign node3406 = (inp[0]) ? 8'b10110001 : node3407;
										assign node3407 = (inp[9]) ? node3413 : node3408;
											assign node3408 = (inp[3]) ? node3410 : 8'b10010000;
												assign node3410 = (inp[6]) ? 8'b10010001 : 8'b10000001;
											assign node3413 = (inp[3]) ? node3417 : node3414;
												assign node3414 = (inp[12]) ? 8'b10110000 : 8'b10100000;
												assign node3417 = (inp[6]) ? 8'b10110001 : 8'b10100001;
						assign node3421 = (inp[2]) ? node3459 : node3422;
							assign node3422 = (inp[13]) ? node3436 : node3423;
								assign node3423 = (inp[0]) ? node3433 : node3424;
									assign node3424 = (inp[10]) ? node3428 : node3425;
										assign node3425 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node3428 = (inp[3]) ? node3430 : 8'b10000100;
											assign node3430 = (inp[1]) ? 8'b10000101 : 8'b10000100;
									assign node3433 = (inp[1]) ? 8'b10000101 : 8'b10000100;
								assign node3436 = (inp[1]) ? node3448 : node3437;
									assign node3437 = (inp[9]) ? node3443 : node3438;
										assign node3438 = (inp[10]) ? node3440 : 8'b10000010;
											assign node3440 = (inp[0]) ? 8'b10100100 : 8'b10000100;
										assign node3443 = (inp[10]) ? 8'b10100100 : node3444;
											assign node3444 = (inp[0]) ? 8'b10100100 : 8'b10100000;
									assign node3448 = (inp[0]) ? 8'b10100101 : node3449;
										assign node3449 = (inp[12]) ? node3453 : node3450;
											assign node3450 = (inp[9]) ? 8'b10100100 : 8'b10000100;
											assign node3453 = (inp[6]) ? 8'b10100001 : node3454;
												assign node3454 = (inp[10]) ? 8'b10000101 : 8'b10000001;
							assign node3459 = (inp[1]) ? node3477 : node3460;
								assign node3460 = (inp[0]) ? node3474 : node3461;
									assign node3461 = (inp[10]) ? node3465 : node3462;
										assign node3462 = (inp[6]) ? 8'b10010000 : 8'b10000010;
										assign node3465 = (inp[6]) ? node3469 : node3466;
											assign node3466 = (inp[3]) ? 8'b10000100 : 8'b10100100;
											assign node3469 = (inp[3]) ? node3471 : 8'b10010100;
												assign node3471 = (inp[9]) ? 8'b10110100 : 8'b10010100;
									assign node3474 = (inp[13]) ? 8'b10110100 : 8'b10010100;
								assign node3477 = (inp[13]) ? node3493 : node3478;
									assign node3478 = (inp[0]) ? 8'b10010101 : node3479;
										assign node3479 = (inp[3]) ? node3487 : node3480;
											assign node3480 = (inp[10]) ? node3484 : node3481;
												assign node3481 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node3484 = (inp[6]) ? 8'b10010100 : 8'b10000100;
											assign node3487 = (inp[6]) ? 8'b10010001 : node3488;
												assign node3488 = (inp[10]) ? 8'b10000101 : 8'b10000001;
									assign node3493 = (inp[10]) ? node3503 : node3494;
										assign node3494 = (inp[0]) ? 8'b11110101 : node3495;
											assign node3495 = (inp[9]) ? node3497 : 8'b10000010;
												assign node3497 = (inp[6]) ? node3499 : 8'b10100001;
													assign node3499 = (inp[3]) ? 8'b10110001 : 8'b10110000;
										assign node3503 = (inp[9]) ? node3507 : node3504;
											assign node3504 = (inp[12]) ? 8'b10010100 : 8'b11110101;
											assign node3507 = (inp[6]) ? 8'b11110101 : node3508;
												assign node3508 = (inp[0]) ? 8'b11110101 : 8'b10100101;
				assign node3512 = (inp[12]) ? node3670 : node3513;
					assign node3513 = (inp[5]) ? node3571 : node3514;
						assign node3514 = (inp[0]) ? node3516 : 8'b11110111;
							assign node3516 = (inp[1]) ? node3540 : node3517;
								assign node3517 = (inp[6]) ? node3535 : node3518;
									assign node3518 = (inp[2]) ? node3530 : node3519;
										assign node3519 = (inp[8]) ? node3521 : 8'b11110111;
											assign node3521 = (inp[10]) ? node3527 : node3522;
												assign node3522 = (inp[13]) ? node3524 : 8'b10110001;
													assign node3524 = (inp[9]) ? 8'b10110001 : 8'b10010001;
												assign node3527 = (inp[13]) ? 8'b10010101 : 8'b11110111;
										assign node3530 = (inp[8]) ? node3532 : 8'b10100101;
											assign node3532 = (inp[10]) ? 8'b10100101 : 8'b10100001;
									assign node3535 = (inp[13]) ? node3537 : 8'b11110111;
										assign node3537 = (inp[9]) ? 8'b11110111 : 8'b10010101;
								assign node3540 = (inp[3]) ? node3558 : node3541;
									assign node3541 = (inp[10]) ? node3553 : node3542;
										assign node3542 = (inp[2]) ? node3550 : node3543;
											assign node3543 = (inp[8]) ? node3545 : 8'b10010100;
												assign node3545 = (inp[6]) ? node3547 : 8'b10110000;
													assign node3547 = (inp[13]) ? 8'b10010000 : 8'b10110000;
											assign node3550 = (inp[9]) ? 8'b10100000 : 8'b10100100;
										assign node3553 = (inp[6]) ? 8'b10110100 : node3554;
											assign node3554 = (inp[2]) ? 8'b10100100 : 8'b10110100;
									assign node3558 = (inp[8]) ? node3564 : node3559;
										assign node3559 = (inp[2]) ? node3561 : 8'b11110111;
											assign node3561 = (inp[6]) ? 8'b11110111 : 8'b10100101;
										assign node3564 = (inp[10]) ? node3566 : 8'b10110001;
											assign node3566 = (inp[13]) ? node3568 : 8'b10100101;
												assign node3568 = (inp[9]) ? 8'b11110111 : 8'b10010101;
						assign node3571 = (inp[1]) ? node3611 : node3572;
							assign node3572 = (inp[0]) ? node3596 : node3573;
								assign node3573 = (inp[6]) ? node3583 : node3574;
									assign node3574 = (inp[10]) ? node3580 : node3575;
										assign node3575 = (inp[13]) ? node3577 : 8'b11110111;
											assign node3577 = (inp[2]) ? 8'b11110111 : 8'b10010101;
										assign node3580 = (inp[8]) ? 8'b10110001 : 8'b11110111;
									assign node3583 = (inp[2]) ? node3587 : node3584;
										assign node3584 = (inp[9]) ? 8'b10010101 : 8'b11110111;
										assign node3587 = (inp[10]) ? node3589 : 8'b10100101;
											assign node3589 = (inp[8]) ? node3593 : node3590;
												assign node3590 = (inp[13]) ? 8'b10000101 : 8'b10100101;
												assign node3593 = (inp[9]) ? 8'b10000001 : 8'b10100001;
								assign node3596 = (inp[13]) ? node3604 : node3597;
									assign node3597 = (inp[8]) ? node3601 : node3598;
										assign node3598 = (inp[2]) ? 8'b10100101 : 8'b11110111;
										assign node3601 = (inp[2]) ? 8'b10100001 : 8'b10110001;
									assign node3604 = (inp[8]) ? node3608 : node3605;
										assign node3605 = (inp[2]) ? 8'b10000101 : 8'b10010101;
										assign node3608 = (inp[2]) ? 8'b10000001 : 8'b10010001;
							assign node3611 = (inp[2]) ? node3639 : node3612;
								assign node3612 = (inp[8]) ? node3626 : node3613;
									assign node3613 = (inp[13]) ? node3619 : node3614;
										assign node3614 = (inp[0]) ? 8'b10110100 : node3615;
											assign node3615 = (inp[3]) ? 8'b10110100 : 8'b11110111;
										assign node3619 = (inp[0]) ? 8'b10010100 : node3620;
											assign node3620 = (inp[3]) ? node3622 : 8'b11110111;
												assign node3622 = (inp[9]) ? 8'b10010100 : 8'b10110100;
									assign node3626 = (inp[9]) ? node3634 : node3627;
										assign node3627 = (inp[13]) ? node3629 : 8'b10110000;
											assign node3629 = (inp[10]) ? node3631 : 8'b11110111;
												assign node3631 = (inp[3]) ? 8'b10110000 : 8'b10110001;
										assign node3634 = (inp[0]) ? 8'b10010000 : node3635;
											assign node3635 = (inp[3]) ? 8'b10110100 : 8'b10010101;
								assign node3639 = (inp[13]) ? node3651 : node3640;
									assign node3640 = (inp[8]) ? node3644 : node3641;
										assign node3641 = (inp[0]) ? 8'b10100100 : 8'b10110100;
										assign node3644 = (inp[0]) ? 8'b10100000 : node3645;
											assign node3645 = (inp[3]) ? node3647 : 8'b11110111;
												assign node3647 = (inp[10]) ? 8'b10100000 : 8'b10100100;
									assign node3651 = (inp[0]) ? node3667 : node3652;
										assign node3652 = (inp[9]) ? node3658 : node3653;
											assign node3653 = (inp[6]) ? node3655 : 8'b11110111;
												assign node3655 = (inp[3]) ? 8'b10100100 : 8'b10100101;
											assign node3658 = (inp[6]) ? node3662 : node3659;
												assign node3659 = (inp[3]) ? 8'b10010100 : 8'b10010101;
												assign node3662 = (inp[3]) ? node3664 : 8'b10000101;
													assign node3664 = (inp[8]) ? 8'b10000000 : 8'b10000100;
										assign node3667 = (inp[8]) ? 8'b10000000 : 8'b10000100;
					assign node3670 = (inp[0]) ? node3732 : node3671;
						assign node3671 = (inp[5]) ? node3673 : 8'b00000010;
							assign node3673 = (inp[2]) ? node3695 : node3674;
								assign node3674 = (inp[9]) ? node3682 : node3675;
									assign node3675 = (inp[3]) ? node3677 : 8'b00000010;
										assign node3677 = (inp[1]) ? node3679 : 8'b00000010;
											assign node3679 = (inp[8]) ? 8'b10100001 : 8'b10100101;
									assign node3682 = (inp[13]) ? node3690 : node3683;
										assign node3683 = (inp[8]) ? node3685 : 8'b00000010;
											assign node3685 = (inp[10]) ? node3687 : 8'b00000010;
												assign node3687 = (inp[3]) ? 8'b10100001 : 8'b10100100;
										assign node3690 = (inp[10]) ? node3692 : 8'b10100000;
											assign node3692 = (inp[8]) ? 8'b10000100 : 8'b10100000;
								assign node3695 = (inp[6]) ? node3721 : node3696;
									assign node3696 = (inp[3]) ? node3708 : node3697;
										assign node3697 = (inp[9]) ? node3705 : node3698;
											assign node3698 = (inp[13]) ? node3700 : 8'b00000010;
												assign node3700 = (inp[10]) ? node3702 : 8'b00000010;
													assign node3702 = (inp[8]) ? 8'b10100100 : 8'b00000010;
											assign node3705 = (inp[8]) ? 8'b10000100 : 8'b10100000;
										assign node3708 = (inp[1]) ? node3716 : node3709;
											assign node3709 = (inp[13]) ? node3711 : 8'b00000010;
												assign node3711 = (inp[9]) ? 8'b10100000 : node3712;
													assign node3712 = (inp[8]) ? 8'b10100100 : 8'b00000010;
											assign node3716 = (inp[13]) ? node3718 : 8'b10100101;
												assign node3718 = (inp[9]) ? 8'b10000101 : 8'b10100101;
									assign node3721 = (inp[1]) ? node3729 : node3722;
										assign node3722 = (inp[9]) ? node3724 : 8'b11110101;
											assign node3724 = (inp[8]) ? node3726 : 8'b10010101;
												assign node3726 = (inp[13]) ? 8'b10010001 : 8'b10110001;
										assign node3729 = (inp[3]) ? 8'b10110100 : 8'b11110101;
						assign node3732 = (inp[2]) ? node3788 : node3733;
							assign node3733 = (inp[1]) ? node3755 : node3734;
								assign node3734 = (inp[9]) ? node3748 : node3735;
									assign node3735 = (inp[8]) ? node3739 : node3736;
										assign node3736 = (inp[13]) ? 8'b10100000 : 8'b00000010;
										assign node3739 = (inp[10]) ? node3743 : node3740;
											assign node3740 = (inp[13]) ? 8'b10000100 : 8'b10100100;
											assign node3743 = (inp[6]) ? node3745 : 8'b00000010;
												assign node3745 = (inp[13]) ? 8'b10100000 : 8'b10100100;
									assign node3748 = (inp[5]) ? node3750 : 8'b00000010;
										assign node3750 = (inp[8]) ? 8'b10100100 : node3751;
											assign node3751 = (inp[10]) ? 8'b00000010 : 8'b10100000;
								assign node3755 = (inp[5]) ? node3781 : node3756;
									assign node3756 = (inp[3]) ? node3768 : node3757;
										assign node3757 = (inp[13]) ? node3763 : node3758;
											assign node3758 = (inp[10]) ? 8'b10100101 : node3759;
												assign node3759 = (inp[8]) ? 8'b10100001 : 8'b10100101;
											assign node3763 = (inp[9]) ? 8'b10100101 : node3764;
												assign node3764 = (inp[10]) ? 8'b10000101 : 8'b10000001;
										assign node3768 = (inp[9]) ? node3776 : node3769;
											assign node3769 = (inp[10]) ? node3773 : node3770;
												assign node3770 = (inp[13]) ? 8'b10100000 : 8'b10100100;
												assign node3773 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node3776 = (inp[6]) ? 8'b00000010 : node3777;
												assign node3777 = (inp[8]) ? 8'b10100100 : 8'b00000010;
									assign node3781 = (inp[8]) ? node3785 : node3782;
										assign node3782 = (inp[13]) ? 8'b10000101 : 8'b10100101;
										assign node3785 = (inp[13]) ? 8'b10000001 : 8'b10100001;
							assign node3788 = (inp[13]) ? node3810 : node3789;
								assign node3789 = (inp[5]) ? node3803 : node3790;
									assign node3790 = (inp[6]) ? node3796 : node3791;
										assign node3791 = (inp[10]) ? 8'b11110101 : node3792;
											assign node3792 = (inp[9]) ? 8'b11110101 : 8'b10110001;
										assign node3796 = (inp[1]) ? node3800 : node3797;
											assign node3797 = (inp[8]) ? 8'b10100100 : 8'b00000010;
											assign node3800 = (inp[8]) ? 8'b10100001 : 8'b10100101;
									assign node3803 = (inp[1]) ? node3807 : node3804;
										assign node3804 = (inp[8]) ? 8'b10110001 : 8'b11110101;
										assign node3807 = (inp[8]) ? 8'b10110000 : 8'b10110100;
								assign node3810 = (inp[5]) ? node3844 : node3811;
									assign node3811 = (inp[6]) ? node3827 : node3812;
										assign node3812 = (inp[9]) ? node3820 : node3813;
											assign node3813 = (inp[3]) ? 8'b10010001 : node3814;
												assign node3814 = (inp[8]) ? node3816 : 8'b10010100;
													assign node3816 = (inp[10]) ? 8'b10010100 : 8'b10010000;
											assign node3820 = (inp[8]) ? node3824 : node3821;
												assign node3821 = (inp[10]) ? 8'b11110101 : 8'b10110100;
												assign node3824 = (inp[3]) ? 8'b10110001 : 8'b10110000;
										assign node3827 = (inp[3]) ? node3835 : node3828;
											assign node3828 = (inp[1]) ? node3830 : 8'b10100100;
												assign node3830 = (inp[10]) ? 8'b10100101 : node3831;
													assign node3831 = (inp[8]) ? 8'b10100001 : 8'b10100101;
											assign node3835 = (inp[8]) ? node3839 : node3836;
												assign node3836 = (inp[9]) ? 8'b00000010 : 8'b10100000;
												assign node3839 = (inp[1]) ? node3841 : 8'b10000100;
													assign node3841 = (inp[9]) ? 8'b10100100 : 8'b10100000;
									assign node3844 = (inp[1]) ? node3848 : node3845;
										assign node3845 = (inp[8]) ? 8'b10010001 : 8'b10010101;
										assign node3848 = (inp[8]) ? 8'b10010000 : 8'b10010100;

endmodule