module dtc_split25_bm85 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node8;
	wire [3-1:0] node10;
	wire [3-1:0] node12;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node25;
	wire [3-1:0] node26;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node38;
	wire [3-1:0] node39;
	wire [3-1:0] node42;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node60;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node76;
	wire [3-1:0] node79;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node85;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node96;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node126;
	wire [3-1:0] node128;
	wire [3-1:0] node129;
	wire [3-1:0] node130;
	wire [3-1:0] node134;
	wire [3-1:0] node137;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node145;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node155;
	wire [3-1:0] node156;
	wire [3-1:0] node158;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node178;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node203;

	assign outp = (inp[0]) ? node46 : node1;
		assign node1 = (inp[9]) ? node3 : 3'b000;
			assign node3 = (inp[6]) ? 3'b000 : node4;
				assign node4 = (inp[4]) ? node16 : node5;
					assign node5 = (inp[7]) ? 3'b000 : node6;
						assign node6 = (inp[1]) ? node8 : 3'b000;
							assign node8 = (inp[3]) ? node10 : 3'b000;
								assign node10 = (inp[2]) ? node12 : 3'b000;
									assign node12 = (inp[8]) ? 3'b000 : 3'b000;
					assign node16 = (inp[3]) ? node18 : 3'b000;
						assign node18 = (inp[1]) ? node30 : node19;
							assign node19 = (inp[10]) ? node25 : node20;
								assign node20 = (inp[2]) ? node22 : 3'b000;
									assign node22 = (inp[5]) ? 3'b011 : 3'b010;
								assign node25 = (inp[7]) ? 3'b000 : node26;
									assign node26 = (inp[5]) ? 3'b001 : 3'b000;
							assign node30 = (inp[2]) ? node38 : node31;
								assign node31 = (inp[10]) ? node35 : node32;
									assign node32 = (inp[7]) ? 3'b000 : 3'b010;
									assign node35 = (inp[7]) ? 3'b000 : 3'b001;
								assign node38 = (inp[5]) ? node42 : node39;
									assign node39 = (inp[8]) ? 3'b110 : 3'b010;
									assign node42 = (inp[7]) ? 3'b000 : 3'b101;
		assign node46 = (inp[6]) ? node166 : node47;
			assign node47 = (inp[3]) ? node103 : node48;
				assign node48 = (inp[4]) ? node60 : node49;
					assign node49 = (inp[10]) ? node51 : 3'b000;
						assign node51 = (inp[5]) ? node53 : 3'b000;
							assign node53 = (inp[8]) ? 3'b000 : node54;
								assign node54 = (inp[9]) ? node56 : 3'b000;
									assign node56 = (inp[2]) ? 3'b100 : 3'b000;
					assign node60 = (inp[5]) ? node82 : node61;
						assign node61 = (inp[9]) ? node67 : node62;
							assign node62 = (inp[7]) ? 3'b100 : node63;
								assign node63 = (inp[1]) ? 3'b100 : 3'b000;
							assign node67 = (inp[2]) ? node75 : node68;
								assign node68 = (inp[7]) ? node72 : node69;
									assign node69 = (inp[11]) ? 3'b000 : 3'b000;
									assign node72 = (inp[11]) ? 3'b100 : 3'b100;
								assign node75 = (inp[7]) ? node79 : node76;
									assign node76 = (inp[10]) ? 3'b100 : 3'b100;
									assign node79 = (inp[11]) ? 3'b000 : 3'b100;
						assign node82 = (inp[7]) ? node96 : node83;
							assign node83 = (inp[2]) ? node89 : node84;
								assign node84 = (inp[9]) ? 3'b000 : node85;
									assign node85 = (inp[1]) ? 3'b000 : 3'b000;
								assign node89 = (inp[10]) ? node93 : node90;
									assign node90 = (inp[1]) ? 3'b110 : 3'b100;
									assign node93 = (inp[9]) ? 3'b100 : 3'b000;
							assign node96 = (inp[9]) ? node98 : 3'b100;
								assign node98 = (inp[11]) ? 3'b000 : node99;
									assign node99 = (inp[10]) ? 3'b100 : 3'b000;
				assign node103 = (inp[7]) ? node137 : node104;
					assign node104 = (inp[4]) ? node126 : node105;
						assign node105 = (inp[9]) ? node117 : node106;
							assign node106 = (inp[10]) ? node112 : node107;
								assign node107 = (inp[1]) ? node109 : 3'b001;
									assign node109 = (inp[2]) ? 3'b101 : 3'b001;
								assign node112 = (inp[5]) ? 3'b101 : node113;
									assign node113 = (inp[8]) ? 3'b101 : 3'b001;
							assign node117 = (inp[1]) ? node123 : node118;
								assign node118 = (inp[2]) ? 3'b010 : node119;
									assign node119 = (inp[11]) ? 3'b110 : 3'b010;
								assign node123 = (inp[5]) ? 3'b011 : 3'b001;
						assign node126 = (inp[9]) ? node128 : 3'b111;
							assign node128 = (inp[10]) ? node134 : node129;
								assign node129 = (inp[1]) ? 3'b111 : node130;
									assign node130 = (inp[8]) ? 3'b011 : 3'b111;
								assign node134 = (inp[5]) ? 3'b111 : 3'b101;
					assign node137 = (inp[9]) ? node139 : 3'b001;
						assign node139 = (inp[8]) ? node155 : node140;
							assign node140 = (inp[5]) ? node148 : node141;
								assign node141 = (inp[2]) ? node145 : node142;
									assign node142 = (inp[1]) ? 3'b001 : 3'b000;
									assign node145 = (inp[10]) ? 3'b110 : 3'b100;
								assign node148 = (inp[4]) ? node152 : node149;
									assign node149 = (inp[2]) ? 3'b001 : 3'b010;
									assign node152 = (inp[2]) ? 3'b111 : 3'b011;
							assign node155 = (inp[10]) ? node161 : node156;
								assign node156 = (inp[4]) ? node158 : 3'b101;
									assign node158 = (inp[5]) ? 3'b001 : 3'b001;
								assign node161 = (inp[4]) ? node163 : 3'b001;
									assign node163 = (inp[5]) ? 3'b111 : 3'b110;
			assign node166 = (inp[3]) ? node168 : 3'b000;
				assign node168 = (inp[9]) ? node170 : 3'b000;
					assign node170 = (inp[7]) ? node198 : node171;
						assign node171 = (inp[4]) ? node183 : node172;
							assign node172 = (inp[5]) ? node178 : node173;
								assign node173 = (inp[1]) ? node175 : 3'b000;
									assign node175 = (inp[2]) ? 3'b000 : 3'b000;
								assign node178 = (inp[11]) ? node180 : 3'b000;
									assign node180 = (inp[2]) ? 3'b110 : 3'b010;
							assign node183 = (inp[8]) ? node191 : node184;
								assign node184 = (inp[1]) ? node188 : node185;
									assign node185 = (inp[10]) ? 3'b110 : 3'b100;
									assign node188 = (inp[2]) ? 3'b101 : 3'b110;
								assign node191 = (inp[1]) ? node195 : node192;
									assign node192 = (inp[10]) ? 3'b010 : 3'b000;
									assign node195 = (inp[10]) ? 3'b101 : 3'b010;
						assign node198 = (inp[2]) ? node200 : 3'b000;
							assign node200 = (inp[4]) ? node202 : 3'b000;
								assign node202 = (inp[8]) ? 3'b000 : node203;
									assign node203 = (inp[5]) ? 3'b100 : 3'b000;

endmodule