module dtc_split25_bm40 (
	input  wire [16-1:0] inp,
	output wire [40-1:0] outp
);

	wire [40-1:0] node1;
	wire [40-1:0] node2;
	wire [40-1:0] node3;
	wire [40-1:0] node5;
	wire [40-1:0] node6;
	wire [40-1:0] node8;
	wire [40-1:0] node10;
	wire [40-1:0] node15;
	wire [40-1:0] node17;
	wire [40-1:0] node18;
	wire [40-1:0] node19;
	wire [40-1:0] node20;
	wire [40-1:0] node21;
	wire [40-1:0] node24;
	wire [40-1:0] node27;
	wire [40-1:0] node28;
	wire [40-1:0] node31;
	wire [40-1:0] node33;
	wire [40-1:0] node34;
	wire [40-1:0] node36;
	wire [40-1:0] node39;
	wire [40-1:0] node40;
	wire [40-1:0] node43;
	wire [40-1:0] node46;
	wire [40-1:0] node47;
	wire [40-1:0] node49;
	wire [40-1:0] node50;
	wire [40-1:0] node51;
	wire [40-1:0] node53;
	wire [40-1:0] node54;
	wire [40-1:0] node56;
	wire [40-1:0] node61;
	wire [40-1:0] node62;
	wire [40-1:0] node64;
	wire [40-1:0] node65;
	wire [40-1:0] node67;
	wire [40-1:0] node70;
	wire [40-1:0] node71;
	wire [40-1:0] node74;
	wire [40-1:0] node77;
	wire [40-1:0] node79;
	wire [40-1:0] node82;
	wire [40-1:0] node83;
	wire [40-1:0] node86;
	wire [40-1:0] node87;
	wire [40-1:0] node89;
	wire [40-1:0] node91;
	wire [40-1:0] node93;
	wire [40-1:0] node96;
	wire [40-1:0] node97;
	wire [40-1:0] node99;
	wire [40-1:0] node101;
	wire [40-1:0] node102;
	wire [40-1:0] node105;
	wire [40-1:0] node108;
	wire [40-1:0] node110;
	wire [40-1:0] node113;
	wire [40-1:0] node114;
	wire [40-1:0] node116;
	wire [40-1:0] node118;
	wire [40-1:0] node119;
	wire [40-1:0] node120;
	wire [40-1:0] node122;
	wire [40-1:0] node124;
	wire [40-1:0] node125;
	wire [40-1:0] node129;
	wire [40-1:0] node130;
	wire [40-1:0] node132;
	wire [40-1:0] node134;
	wire [40-1:0] node137;
	wire [40-1:0] node138;
	wire [40-1:0] node139;
	wire [40-1:0] node145;
	wire [40-1:0] node146;
	wire [40-1:0] node148;
	wire [40-1:0] node150;
	wire [40-1:0] node151;
	wire [40-1:0] node153;
	wire [40-1:0] node156;
	wire [40-1:0] node157;
	wire [40-1:0] node160;
	wire [40-1:0] node163;
	wire [40-1:0] node164;
	wire [40-1:0] node167;
	wire [40-1:0] node168;
	wire [40-1:0] node170;
	wire [40-1:0] node172;
	wire [40-1:0] node174;
	wire [40-1:0] node175;
	wire [40-1:0] node179;
	wire [40-1:0] node180;
	wire [40-1:0] node182;
	wire [40-1:0] node184;
	wire [40-1:0] node186;
	wire [40-1:0] node189;
	wire [40-1:0] node191;
	wire [40-1:0] node194;
	wire [40-1:0] node195;
	wire [40-1:0] node196;
	wire [40-1:0] node199;
	wire [40-1:0] node200;
	wire [40-1:0] node201;
	wire [40-1:0] node202;
	wire [40-1:0] node203;
	wire [40-1:0] node206;
	wire [40-1:0] node209;
	wire [40-1:0] node210;
	wire [40-1:0] node213;
	wire [40-1:0] node216;
	wire [40-1:0] node217;
	wire [40-1:0] node218;
	wire [40-1:0] node221;
	wire [40-1:0] node224;
	wire [40-1:0] node225;
	wire [40-1:0] node228;
	wire [40-1:0] node231;
	wire [40-1:0] node232;
	wire [40-1:0] node233;
	wire [40-1:0] node234;
	wire [40-1:0] node237;
	wire [40-1:0] node240;
	wire [40-1:0] node241;
	wire [40-1:0] node244;
	wire [40-1:0] node247;
	wire [40-1:0] node248;
	wire [40-1:0] node249;
	wire [40-1:0] node252;
	wire [40-1:0] node255;
	wire [40-1:0] node256;
	wire [40-1:0] node259;
	wire [40-1:0] node262;
	wire [40-1:0] node263;
	wire [40-1:0] node266;
	wire [40-1:0] node268;
	wire [40-1:0] node269;
	wire [40-1:0] node270;
	wire [40-1:0] node271;
	wire [40-1:0] node272;
	wire [40-1:0] node273;
	wire [40-1:0] node274;
	wire [40-1:0] node275;
	wire [40-1:0] node276;
	wire [40-1:0] node279;
	wire [40-1:0] node282;
	wire [40-1:0] node283;
	wire [40-1:0] node286;
	wire [40-1:0] node289;
	wire [40-1:0] node290;
	wire [40-1:0] node291;
	wire [40-1:0] node294;
	wire [40-1:0] node297;
	wire [40-1:0] node298;
	wire [40-1:0] node301;
	wire [40-1:0] node304;
	wire [40-1:0] node305;
	wire [40-1:0] node306;
	wire [40-1:0] node307;
	wire [40-1:0] node310;
	wire [40-1:0] node313;
	wire [40-1:0] node314;
	wire [40-1:0] node317;
	wire [40-1:0] node320;
	wire [40-1:0] node321;
	wire [40-1:0] node322;
	wire [40-1:0] node325;
	wire [40-1:0] node328;
	wire [40-1:0] node329;
	wire [40-1:0] node333;
	wire [40-1:0] node334;
	wire [40-1:0] node335;
	wire [40-1:0] node336;
	wire [40-1:0] node337;
	wire [40-1:0] node340;
	wire [40-1:0] node343;
	wire [40-1:0] node344;
	wire [40-1:0] node347;
	wire [40-1:0] node350;
	wire [40-1:0] node351;
	wire [40-1:0] node352;
	wire [40-1:0] node355;
	wire [40-1:0] node358;
	wire [40-1:0] node359;
	wire [40-1:0] node362;
	wire [40-1:0] node365;
	wire [40-1:0] node366;
	wire [40-1:0] node367;
	wire [40-1:0] node368;
	wire [40-1:0] node371;
	wire [40-1:0] node374;
	wire [40-1:0] node375;
	wire [40-1:0] node378;
	wire [40-1:0] node381;
	wire [40-1:0] node382;
	wire [40-1:0] node383;
	wire [40-1:0] node386;
	wire [40-1:0] node389;
	wire [40-1:0] node390;
	wire [40-1:0] node394;
	wire [40-1:0] node395;
	wire [40-1:0] node397;
	wire [40-1:0] node398;
	wire [40-1:0] node399;
	wire [40-1:0] node400;
	wire [40-1:0] node404;
	wire [40-1:0] node405;
	wire [40-1:0] node410;
	wire [40-1:0] node411;
	wire [40-1:0] node412;
	wire [40-1:0] node413;
	wire [40-1:0] node414;
	wire [40-1:0] node417;
	wire [40-1:0] node420;
	wire [40-1:0] node421;
	wire [40-1:0] node424;
	wire [40-1:0] node427;
	wire [40-1:0] node428;
	wire [40-1:0] node429;
	wire [40-1:0] node432;
	wire [40-1:0] node435;
	wire [40-1:0] node436;
	wire [40-1:0] node439;
	wire [40-1:0] node442;
	wire [40-1:0] node443;
	wire [40-1:0] node444;
	wire [40-1:0] node445;
	wire [40-1:0] node448;
	wire [40-1:0] node451;
	wire [40-1:0] node452;
	wire [40-1:0] node455;
	wire [40-1:0] node458;
	wire [40-1:0] node459;
	wire [40-1:0] node460;
	wire [40-1:0] node463;
	wire [40-1:0] node466;
	wire [40-1:0] node467;
	wire [40-1:0] node470;
	wire [40-1:0] node473;
	wire [40-1:0] node474;
	wire [40-1:0] node475;
	wire [40-1:0] node476;
	wire [40-1:0] node478;
	wire [40-1:0] node479;
	wire [40-1:0] node481;
	wire [40-1:0] node484;
	wire [40-1:0] node486;
	wire [40-1:0] node489;
	wire [40-1:0] node490;
	wire [40-1:0] node491;
	wire [40-1:0] node493;
	wire [40-1:0] node499;
	wire [40-1:0] node500;
	wire [40-1:0] node502;
	wire [40-1:0] node504;
	wire [40-1:0] node506;
	wire [40-1:0] node507;
	wire [40-1:0] node511;
	wire [40-1:0] node512;
	wire [40-1:0] node513;
	wire [40-1:0] node514;
	wire [40-1:0] node515;
	wire [40-1:0] node518;
	wire [40-1:0] node521;
	wire [40-1:0] node522;
	wire [40-1:0] node525;
	wire [40-1:0] node528;
	wire [40-1:0] node529;
	wire [40-1:0] node530;
	wire [40-1:0] node533;
	wire [40-1:0] node536;
	wire [40-1:0] node537;
	wire [40-1:0] node540;
	wire [40-1:0] node543;
	wire [40-1:0] node544;
	wire [40-1:0] node545;
	wire [40-1:0] node546;
	wire [40-1:0] node549;
	wire [40-1:0] node552;
	wire [40-1:0] node553;
	wire [40-1:0] node557;
	wire [40-1:0] node558;
	wire [40-1:0] node559;
	wire [40-1:0] node563;
	wire [40-1:0] node564;
	wire [40-1:0] node567;
	wire [40-1:0] node570;
	wire [40-1:0] node571;
	wire [40-1:0] node572;
	wire [40-1:0] node574;
	wire [40-1:0] node575;
	wire [40-1:0] node577;
	wire [40-1:0] node579;
	wire [40-1:0] node582;
	wire [40-1:0] node583;
	wire [40-1:0] node585;
	wire [40-1:0] node587;
	wire [40-1:0] node590;
	wire [40-1:0] node591;
	wire [40-1:0] node592;
	wire [40-1:0] node595;
	wire [40-1:0] node598;
	wire [40-1:0] node599;
	wire [40-1:0] node603;
	wire [40-1:0] node604;
	wire [40-1:0] node605;
	wire [40-1:0] node606;
	wire [40-1:0] node608;
	wire [40-1:0] node611;
	wire [40-1:0] node612;
	wire [40-1:0] node616;
	wire [40-1:0] node617;
	wire [40-1:0] node619;
	wire [40-1:0] node622;
	wire [40-1:0] node623;
	wire [40-1:0] node628;
	wire [40-1:0] node629;
	wire [40-1:0] node630;
	wire [40-1:0] node632;
	wire [40-1:0] node633;
	wire [40-1:0] node634;
	wire [40-1:0] node635;
	wire [40-1:0] node638;
	wire [40-1:0] node641;
	wire [40-1:0] node642;
	wire [40-1:0] node645;
	wire [40-1:0] node648;
	wire [40-1:0] node649;
	wire [40-1:0] node650;
	wire [40-1:0] node653;
	wire [40-1:0] node656;
	wire [40-1:0] node657;
	wire [40-1:0] node660;
	wire [40-1:0] node663;
	wire [40-1:0] node664;
	wire [40-1:0] node665;
	wire [40-1:0] node666;
	wire [40-1:0] node667;
	wire [40-1:0] node670;
	wire [40-1:0] node673;
	wire [40-1:0] node674;
	wire [40-1:0] node677;
	wire [40-1:0] node680;
	wire [40-1:0] node681;
	wire [40-1:0] node682;
	wire [40-1:0] node685;
	wire [40-1:0] node688;
	wire [40-1:0] node689;
	wire [40-1:0] node692;
	wire [40-1:0] node696;
	wire [40-1:0] node697;
	wire [40-1:0] node699;
	wire [40-1:0] node700;
	wire [40-1:0] node701;
	wire [40-1:0] node703;
	wire [40-1:0] node706;
	wire [40-1:0] node707;
	wire [40-1:0] node710;
	wire [40-1:0] node713;
	wire [40-1:0] node714;
	wire [40-1:0] node715;
	wire [40-1:0] node718;
	wire [40-1:0] node721;
	wire [40-1:0] node722;
	wire [40-1:0] node725;
	wire [40-1:0] node728;
	wire [40-1:0] node729;
	wire [40-1:0] node730;
	wire [40-1:0] node731;
	wire [40-1:0] node732;
	wire [40-1:0] node735;
	wire [40-1:0] node738;
	wire [40-1:0] node739;
	wire [40-1:0] node742;
	wire [40-1:0] node745;
	wire [40-1:0] node746;
	wire [40-1:0] node747;
	wire [40-1:0] node750;
	wire [40-1:0] node753;
	wire [40-1:0] node754;
	wire [40-1:0] node757;

	assign outp = (inp[9]) ? node194 : node1;
		assign node1 = (inp[1]) ? node15 : node2;
			assign node2 = (inp[3]) ? 40'b0000000000000000000000000000000000000000 : node3;
				assign node3 = (inp[8]) ? node5 : 40'b0000000000000000000000000000000000000000;
					assign node5 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node6;
						assign node6 = (inp[4]) ? node8 : 40'b0000000000000000000000000000000000000000;
							assign node8 = (inp[7]) ? node10 : 40'b0000000000000000000000000000000000000000;
								assign node10 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000100000000000000000000000;
			assign node15 = (inp[4]) ? node17 : 40'b0000000001000000000000000000000000000000;
				assign node17 = (inp[7]) ? node113 : node18;
					assign node18 = (inp[8]) ? node46 : node19;
						assign node19 = (inp[14]) ? node27 : node20;
							assign node20 = (inp[3]) ? node24 : node21;
								assign node21 = (inp[11]) ? 40'b0000000000000010000001000000000000000000 : 40'b0000000000000010000000000100000000000000;
								assign node24 = (inp[11]) ? 40'b0000000000000001010000000100000000000000 : 40'b0000000000100010000000000000000000000000;
							assign node27 = (inp[3]) ? node31 : node28;
								assign node28 = (inp[11]) ? 40'b0000000000000000000001000000000010000000 : 40'b0000000000000000000000000100000010000000;
								assign node31 = (inp[11]) ? node33 : 40'b0000000000100000000000000000000010000000;
									assign node33 = (inp[13]) ? node39 : node34;
										assign node34 = (inp[10]) ? node36 : 40'b0000000000000000000000000000000000000000;
											assign node36 = (inp[0]) ? 40'b0000000000000000010000010000000010000000 : 40'b0000000000000000000000000000000000000000;
										assign node39 = (inp[0]) ? node43 : node40;
											assign node40 = (inp[10]) ? 40'b0000000000000010010000010000000010000000 : 40'b0000000000000000000000000000000000000000;
											assign node43 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000010010000010000000000000000;
						assign node46 = (inp[14]) ? node82 : node47;
							assign node47 = (inp[0]) ? node49 : 40'b0000000000000000000000000000000000000000;
								assign node49 = (inp[3]) ? node61 : node50;
									assign node50 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node51;
										assign node51 = (inp[6]) ? node53 : 40'b0000000000000000000000000000000000000000;
											assign node53 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node54;
												assign node54 = (inp[2]) ? node56 : 40'b0000000000000000000000000000000000000000;
													assign node56 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node61 = (inp[10]) ? node77 : node62;
										assign node62 = (inp[15]) ? node64 : 40'b0000000000000000000000000000000000000000;
											assign node64 = (inp[2]) ? node70 : node65;
												assign node65 = (inp[5]) ? node67 : 40'b0000000000000000000000000000000000000000;
													assign node67 = (inp[6]) ? 40'b0000000010000010010000100000000000000000 : 40'b0000000000000000000000000000000000000000;
												assign node70 = (inp[5]) ? node74 : node71;
													assign node71 = (inp[11]) ? 40'b0000000000000001010000000000010000000010 : 40'b0000000000000010010000100000000000000010;
													assign node74 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000001010000000000001000000000;
										assign node77 = (inp[13]) ? node79 : 40'b0000000000000000000000000000000000000000;
											assign node79 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000001000000000;
							assign node82 = (inp[3]) ? node86 : node83;
								assign node83 = (inp[11]) ? 40'b0000000000001000010000100100000001000000 : 40'b0000000000000000010100100100000001000000;
								assign node86 = (inp[0]) ? node96 : node87;
									assign node87 = (inp[12]) ? node89 : 40'b0000000000000000000000000000000000000000;
										assign node89 = (inp[2]) ? node91 : 40'b0000000000000000000000000000000000000000;
											assign node91 = (inp[5]) ? node93 : 40'b0000000000000000000000000000000000000000;
												assign node93 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000100000000000001000000;
									assign node96 = (inp[10]) ? node108 : node97;
										assign node97 = (inp[15]) ? node99 : 40'b0000000000000000000000000000000000000000;
											assign node99 = (inp[12]) ? node101 : 40'b0000000000000000000000000000000000000000;
												assign node101 = (inp[5]) ? node105 : node102;
													assign node102 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node105 = (inp[11]) ? 40'b0000000010001000010000000000000001000000 : 40'b0000000000000001010100000000001001000000;
										assign node108 = (inp[13]) ? node110 : 40'b0000000000000000000000000000000000000000;
											assign node110 = (inp[11]) ? 40'b0000000010001000000000000000000001000010 : 40'b0000000000000000000100000000001001000010;
					assign node113 = (inp[14]) ? node145 : node114;
						assign node114 = (inp[0]) ? node116 : 40'b0000000000000000000000000000000000000000;
							assign node116 = (inp[8]) ? node118 : 40'b0000000000000000000000000000000000000000;
								assign node118 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node119;
									assign node119 = (inp[3]) ? node129 : node120;
										assign node120 = (inp[15]) ? node122 : 40'b0000000000000000000000000000000000000000;
											assign node122 = (inp[2]) ? node124 : 40'b0000000000000000000000000000000000000000;
												assign node124 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : node125;
													assign node125 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node129 = (inp[10]) ? node137 : node130;
											assign node130 = (inp[12]) ? node132 : 40'b0000000000000000000000000000000000000000;
												assign node132 = (inp[2]) ? node134 : 40'b0000000000000000000000000000000000000000;
													assign node134 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
											assign node137 = (inp[13]) ? 40'b0000000000000000000000010000000100000000 : node138;
												assign node138 = (inp[2]) ? 40'b0000000000000000000000000000000000000000 : node139;
													assign node139 = (inp[15]) ? 40'b0000000010000000000000100000000110000000 : 40'b0000000000000000000000000000000000000000;
						assign node145 = (inp[8]) ? node163 : node146;
							assign node146 = (inp[3]) ? node148 : 40'b0000000000000000000000000000000000000000;
								assign node148 = (inp[11]) ? node150 : 40'b0000000000000000000000000000000000000000;
									assign node150 = (inp[10]) ? node156 : node151;
										assign node151 = (inp[0]) ? node153 : 40'b0000000000000000000000000000000000000000;
											assign node153 = (inp[13]) ? 40'b0000000000000010000000010000000100000000 : 40'b0000000000000000000000000000000000000000;
										assign node156 = (inp[0]) ? node160 : node157;
											assign node157 = (inp[13]) ? 40'b0000000000000010000000010000000110000000 : 40'b0000000000000000000000000000000000000000;
											assign node160 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000010000000110000000;
							assign node163 = (inp[3]) ? node167 : node164;
								assign node164 = (inp[11]) ? 40'b0100000000000000000000100100000100000001 : 40'b0100000000000000000000101100000100000000;
								assign node167 = (inp[13]) ? node179 : node168;
									assign node168 = (inp[15]) ? node170 : 40'b0000000000000000000000000000000000000000;
										assign node170 = (inp[12]) ? node172 : 40'b0000000000000000000000000000000000000000;
											assign node172 = (inp[2]) ? node174 : 40'b0000000000000000000000000000000000000000;
												assign node174 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node175;
													assign node175 = (inp[0]) ? 40'b0100000000000000000000100000000110000011 : 40'b0000000000000000000000000000000000000000;
									assign node179 = (inp[10]) ? node189 : node180;
										assign node180 = (inp[11]) ? node182 : 40'b0000000000000000000000000000000000000000;
											assign node182 = (inp[12]) ? node184 : 40'b0000000000000000000000000000000000000000;
												assign node184 = (inp[5]) ? node186 : 40'b0000000000000000000000000000000000000000;
													assign node186 = (inp[15]) ? 40'b0100000000000000000000000000000000000001 : 40'b0000000000000000000000000000000000000000;
										assign node189 = (inp[0]) ? node191 : 40'b0000000000000000000000000000000000000000;
											assign node191 = (inp[11]) ? 40'b0100000000000000000000010000000100000001 : 40'b0100000000000000000000011000000100000000;
		assign node194 = (inp[1]) ? node262 : node195;
			assign node195 = (inp[8]) ? node199 : node196;
				assign node196 = (inp[4]) ? 40'b0000000001000000000000000000000000000100 : 40'b0000000000000000000000000000000000000100;
				assign node199 = (inp[7]) ? node231 : node200;
					assign node200 = (inp[14]) ? node216 : node201;
						assign node201 = (inp[11]) ? node209 : node202;
							assign node202 = (inp[3]) ? node206 : node203;
								assign node203 = (inp[4]) ? 40'b0000000001000010010100100000001001000100 : 40'b0000000000000010010100100000001001000100;
								assign node206 = (inp[4]) ? 40'b0000000001000000010100100000001011000100 : 40'b0000000000000000010100100000001011000100;
							assign node209 = (inp[3]) ? node213 : node210;
								assign node210 = (inp[4]) ? 40'b0000000001000010010100100000000001000110 : 40'b0000000000000010010100100000000001000110;
								assign node213 = (inp[4]) ? 40'b0000000001000000010100100000000011000110 : 40'b0000000000000000010100100000000011000110;
						assign node216 = (inp[11]) ? node224 : node217;
							assign node217 = (inp[3]) ? node221 : node218;
								assign node218 = (inp[4]) ? 40'b0000000001001010010000100000001001000100 : 40'b0000000000001010010000100000001001000100;
								assign node221 = (inp[4]) ? 40'b0000000001001000010000100000001011000100 : 40'b0000000000001000010000100000001011000100;
							assign node224 = (inp[3]) ? node228 : node225;
								assign node225 = (inp[4]) ? 40'b0000000001001010010000100000000001000110 : 40'b0000000000001010010000100000000001000110;
								assign node228 = (inp[4]) ? 40'b0000000001001000010000100000000011000110 : 40'b0000000000001000010000100000000011000110;
					assign node231 = (inp[14]) ? node247 : node232;
						assign node232 = (inp[3]) ? node240 : node233;
							assign node233 = (inp[11]) ? node237 : node234;
								assign node234 = (inp[4]) ? 40'b0100000001000010000000101000001100000100 : 40'b0100000000000010000000101000001100000100;
								assign node237 = (inp[4]) ? 40'b0100000001000010000000101000000100000110 : 40'b0100000000000010000000101000000100000110;
							assign node240 = (inp[11]) ? node244 : node241;
								assign node241 = (inp[4]) ? 40'b0100000001000000000000101000001110000100 : 40'b0100000000000000000000101000001110000100;
								assign node244 = (inp[4]) ? 40'b0100000001000000000000101000000110000110 : 40'b0100000000000000000000101000000110000110;
						assign node247 = (inp[3]) ? node255 : node248;
							assign node248 = (inp[11]) ? node252 : node249;
								assign node249 = (inp[4]) ? 40'b0100000001000010000000100000001100000101 : 40'b0100000000000010000000100000001100000101;
								assign node252 = (inp[4]) ? 40'b0100000001000010000000100000000100000111 : 40'b0100000000000010000000100000000100000111;
							assign node255 = (inp[11]) ? node259 : node256;
								assign node256 = (inp[4]) ? 40'b0100000001000000000000100000001110000101 : 40'b0100000000000000000000100000001110000101;
								assign node259 = (inp[4]) ? 40'b0100000001000000000000100000000110000111 : 40'b0100000000000000000000100000000110000111;
			assign node262 = (inp[4]) ? node266 : node263;
				assign node263 = (inp[8]) ? 40'b0000000001000000000000000000000000000000 : 40'b0000100001000000000000000000000000000000;
				assign node266 = (inp[8]) ? node268 : 40'b0000100000000000000000000000000000000000;
					assign node268 = (inp[7]) ? node570 : node269;
						assign node269 = (inp[3]) ? node473 : node270;
							assign node270 = (inp[14]) ? node394 : node271;
								assign node271 = (inp[13]) ? node333 : node272;
									assign node272 = (inp[10]) ? node304 : node273;
										assign node273 = (inp[0]) ? node289 : node274;
											assign node274 = (inp[15]) ? node282 : node275;
												assign node275 = (inp[5]) ? node279 : node276;
													assign node276 = (inp[12]) ? 40'b0001000000011101010010000010101000000000 : 40'b1001000000011101010010000010101000000000;
													assign node279 = (inp[11]) ? 40'b1001000000010101010010000001101000000000 : 40'b1001000000010101010010000001101000010000;
												assign node282 = (inp[11]) ? node286 : node283;
													assign node283 = (inp[12]) ? 40'b0001000000000101010010000011101000010000 : 40'b1001000000001101010110000010101000010000;
													assign node286 = (inp[6]) ? 40'b0001000000000101010010000001101000000000 : 40'b1001000000001101010010000010101000000000;
											assign node289 = (inp[5]) ? node297 : node290;
												assign node290 = (inp[11]) ? node294 : node291;
													assign node291 = (inp[15]) ? 40'b0000000000001101010010000010101000010000 : 40'b1000000000011101010010000010101000010000;
													assign node294 = (inp[6]) ? 40'b0000000000001101010010000010101000000000 : 40'b1000000000001101010010000010101000000000;
												assign node297 = (inp[2]) ? node301 : node298;
													assign node298 = (inp[11]) ? 40'b1000000000000101010110000010101000000000 : 40'b1000000000010101010110000010101000010000;
													assign node301 = (inp[15]) ? 40'b0000000000000101010110000011101000010000 : 40'b0000000000010101010110000011101000000000;
										assign node304 = (inp[0]) ? node320 : node305;
											assign node305 = (inp[5]) ? node313 : node306;
												assign node306 = (inp[6]) ? node310 : node307;
													assign node307 = (inp[15]) ? 40'b1001000000000001010010000000101000000000 : 40'b1001000000010001010010000000101000000000;
													assign node310 = (inp[12]) ? 40'b0001000000001001010010000010101000000000 : 40'b1001000000001001010010000010101000000000;
												assign node313 = (inp[2]) ? node317 : node314;
													assign node314 = (inp[11]) ? 40'b0001000000001001010010000011101000000000 : 40'b0001000000011001010010000010101000010000;
													assign node317 = (inp[6]) ? 40'b0001000000000001010110000011101000010000 : 40'b0001000000010001010110000010101000000000;
											assign node320 = (inp[11]) ? node328 : node321;
												assign node321 = (inp[5]) ? node325 : node322;
													assign node322 = (inp[15]) ? 40'b1000000000001001010010000010101000010000 : 40'b1000000000011001010010000010101000010000;
													assign node325 = (inp[2]) ? 40'b0000000000010001010110000011101000010000 : 40'b0000000000010001010010000001101000010000;
												assign node328 = (inp[2]) ? 40'b1000000000010001010010000001101000000000 : node329;
													assign node329 = (inp[12]) ? 40'b0000000000011001010010000010101000000000 : 40'b1000000000000001010010000000101000000000;
									assign node333 = (inp[15]) ? node365 : node334;
										assign node334 = (inp[0]) ? node350 : node335;
											assign node335 = (inp[10]) ? node343 : node336;
												assign node336 = (inp[5]) ? node340 : node337;
													assign node337 = (inp[11]) ? 40'b1001000000011101010010000010001000000000 : 40'b1001000000010101010010000000001000010000;
													assign node340 = (inp[2]) ? 40'b0001000000010101010110000011001000010000 : 40'b1001000000010101010110000010001000000000;
												assign node343 = (inp[2]) ? node347 : node344;
													assign node344 = (inp[6]) ? 40'b0001000000011001010010000010001000000000 : 40'b0001000000011001010110000010001000000000;
													assign node347 = (inp[11]) ? 40'b0001000000010001010010000001001000000000 : 40'b0001000000010001010010000001001000010000;
											assign node350 = (inp[11]) ? node358 : node351;
												assign node351 = (inp[6]) ? node355 : node352;
													assign node352 = (inp[10]) ? 40'b1000000000010001010110000010001000010000 : 40'b0000000000010101010010000010001000010000;
													assign node355 = (inp[2]) ? 40'b0000000000010001010010000001001000010000 : 40'b1000000000010001010010000001001000010000;
												assign node358 = (inp[2]) ? node362 : node359;
													assign node359 = (inp[10]) ? 40'b1000000000010001010010000000001000000000 : 40'b1000000000010101010010000000001000000000;
													assign node362 = (inp[5]) ? 40'b0000000000010101010010000001001000000000 : 40'b0000000000011101010010000011001000000000;
										assign node365 = (inp[0]) ? node381 : node366;
											assign node366 = (inp[5]) ? node374 : node367;
												assign node367 = (inp[11]) ? node371 : node368;
													assign node368 = (inp[12]) ? 40'b0001000000001001010010000010001000010000 : 40'b1001000000000101010010000000001000010000;
													assign node371 = (inp[2]) ? 40'b1001000000000101010010000001001000000000 : 40'b1001000000000001010010000000001000000000;
												assign node374 = (inp[12]) ? node378 : node375;
													assign node375 = (inp[6]) ? 40'b0001000000000101010110000011001000000000 : 40'b0001000000000101010110000010001000000000;
													assign node378 = (inp[10]) ? 40'b0001000000001001010110000010001000000000 : 40'b0001000000001101010110000010001000000000;
											assign node381 = (inp[10]) ? node389 : node382;
												assign node382 = (inp[11]) ? node386 : node383;
													assign node383 = (inp[5]) ? 40'b0000000000001101010110000010001000010000 : 40'b1000000000000101010010000010001000010000;
													assign node386 = (inp[12]) ? 40'b0000000000000101010010000001001000000000 : 40'b1000000000000101010010000010001000000000;
												assign node389 = (inp[12]) ? 40'b0000000000001001010110000010001000010000 : node390;
													assign node390 = (inp[11]) ? 40'b0000000000000001010110000010001000000000 : 40'b1000000000000001010110000010001000010000;
								assign node394 = (inp[11]) ? node410 : node395;
									assign node395 = (inp[2]) ? node397 : 40'b0000000000000000000000000000000000000000;
										assign node397 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node398;
											assign node398 = (inp[15]) ? node404 : node399;
												assign node399 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node400;
													assign node400 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000010100001000000000000000000000;
												assign node404 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : node405;
													assign node405 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
									assign node410 = (inp[10]) ? node442 : node411;
										assign node411 = (inp[15]) ? node427 : node412;
											assign node412 = (inp[6]) ? node420 : node413;
												assign node413 = (inp[0]) ? node417 : node414;
													assign node414 = (inp[13]) ? 40'b1001010000010100000100000010000000000000 : 40'b1001010000010100000100000010100000000000;
													assign node417 = (inp[5]) ? 40'b1000010000010100000100000010000000000000 : 40'b1000010000010100000000000000000000000000;
												assign node420 = (inp[0]) ? node424 : node421;
													assign node421 = (inp[12]) ? 40'b0001010000011100000000000011100000000000 : 40'b1001010000010100000000000001000000000000;
													assign node424 = (inp[12]) ? 40'b0000010000011100000000000010100000000000 : 40'b0000010000010100000100000011000000000000;
											assign node427 = (inp[13]) ? node435 : node428;
												assign node428 = (inp[0]) ? node432 : node429;
													assign node429 = (inp[5]) ? 40'b0001010000000100000100000011100000000000 : 40'b1001010000001100000100000010100000000000;
													assign node432 = (inp[12]) ? 40'b0000010000001100000000000010100000000000 : 40'b0000010000000100000100000010100000000000;
												assign node435 = (inp[0]) ? node439 : node436;
													assign node436 = (inp[6]) ? 40'b0001010000001100000000000011000000000000 : 40'b1001010000000100000000000001000000000000;
													assign node439 = (inp[5]) ? 40'b0000010000001100000100000010000000000000 : 40'b1000010000000100000000000000000000000000;
										assign node442 = (inp[13]) ? node458 : node443;
											assign node443 = (inp[15]) ? node451 : node444;
												assign node444 = (inp[2]) ? node448 : node445;
													assign node445 = (inp[5]) ? 40'b1000010000010000000000000001100000000000 : 40'b1001010000011000000000000010100000000000;
													assign node448 = (inp[12]) ? 40'b1001010000010000000000000001100000000000 : 40'b0001010000010000000100000010100000000000;
												assign node451 = (inp[0]) ? node455 : node452;
													assign node452 = (inp[12]) ? 40'b0001010000000000000100000011100000000000 : 40'b1001010000000000000000000000100000000000;
													assign node455 = (inp[6]) ? 40'b0000010000001000000000000010100000000000 : 40'b1000010000000000000000000000100000000000;
											assign node458 = (inp[15]) ? node466 : node459;
												assign node459 = (inp[6]) ? node463 : node460;
													assign node460 = (inp[5]) ? 40'b0001010000010000000100000010000000000000 : 40'b1001010000010000000000000000000000000000;
													assign node463 = (inp[0]) ? 40'b0000010000010000000000000001000000000000 : 40'b0001010000011000000000000010000000000000;
												assign node466 = (inp[0]) ? node470 : node467;
													assign node467 = (inp[12]) ? 40'b0001010000001000000000000010000000000000 : 40'b0001010000000000000100000010000000000000;
													assign node470 = (inp[2]) ? 40'b1000010000000000000000000001000000000000 : 40'b0000010000001000000000000010000000000000;
							assign node473 = (inp[11]) ? node499 : node474;
								assign node474 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node475;
									assign node475 = (inp[0]) ? node489 : node476;
										assign node476 = (inp[10]) ? node478 : 40'b0000000000000000000000000000000000000000;
											assign node478 = (inp[15]) ? node484 : node479;
												assign node479 = (inp[13]) ? node481 : 40'b0000000000000000000000000000000000000000;
													assign node481 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : 40'b1001000000010000000000000000000000100000;
												assign node484 = (inp[5]) ? node486 : 40'b0000000000000000000000000000000000000000;
													assign node486 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b0001000000000000000100000010100000100000;
										assign node489 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node490;
											assign node490 = (inp[6]) ? 40'b0000000000000000000000000000000000000000 : node491;
												assign node491 = (inp[15]) ? node493 : 40'b0000000000000000000000000000000000000000;
													assign node493 = (inp[12]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000000000000100000100000010100000100000;
								assign node499 = (inp[14]) ? node511 : node500;
									assign node500 = (inp[12]) ? node502 : 40'b0000000000000000000000000000000000000000;
										assign node502 = (inp[5]) ? node504 : 40'b0000000000000000000000000000000000000000;
											assign node504 = (inp[2]) ? node506 : 40'b0000000000000000000000000000000000000000;
												assign node506 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : node507;
													assign node507 = (inp[0]) ? 40'b1000000000010100001000000000100000010000 : 40'b1001000000010000001000000000100000010000;
									assign node511 = (inp[0]) ? node543 : node512;
										assign node512 = (inp[10]) ? node528 : node513;
											assign node513 = (inp[13]) ? node521 : node514;
												assign node514 = (inp[15]) ? node518 : node515;
													assign node515 = (inp[12]) ? 40'b0011000000011100000000000010100000000000 : 40'b0011000000010100000100000010100000000000;
													assign node518 = (inp[12]) ? 40'b0011000000001100000000000010100000000000 : 40'b0011000000001100000000000010100000000000;
												assign node521 = (inp[2]) ? node525 : node522;
													assign node522 = (inp[12]) ? 40'b0011000000011100000000000011000000000000 : 40'b1011000000001100000000000010000000000000;
													assign node525 = (inp[12]) ? 40'b0011000000000100000000000001000000000000 : 40'b0011000000010100000100000011000000000000;
											assign node528 = (inp[13]) ? node536 : node529;
												assign node529 = (inp[5]) ? node533 : node530;
													assign node530 = (inp[2]) ? 40'b1011000000000000000100000010100000000000 : 40'b1011000000011000000000000010100000000000;
													assign node533 = (inp[2]) ? 40'b0011000000000000000100000011100000000000 : 40'b1011000000000000000100000010100000000000;
												assign node536 = (inp[15]) ? node540 : node537;
													assign node537 = (inp[6]) ? 40'b0011000000010000000100000010000000000000 : 40'b1011000000010000000000000000000000000000;
													assign node540 = (inp[5]) ? 40'b0011000000001000000100000010000000000000 : 40'b0011000000001000000000000010000000000000;
										assign node543 = (inp[15]) ? node557 : node544;
											assign node544 = (inp[13]) ? node552 : node545;
												assign node545 = (inp[10]) ? node549 : node546;
													assign node546 = (inp[2]) ? 40'b0010000000011100000100000010100000000000 : 40'b1010000000011100000000000010100000000000;
													assign node549 = (inp[5]) ? 40'b0010000000010000000100000011100000000000 : 40'b1010000000010000000000000000100000000000;
												assign node552 = (inp[6]) ? 40'b1010000000010100000000000001000000000000 : node553;
													assign node553 = (inp[5]) ? 40'b1010000000010100000100000010000000000000 : 40'b1010000000010100000000000000000000000000;
											assign node557 = (inp[12]) ? node563 : node558;
												assign node558 = (inp[13]) ? 40'b1010000000000000000000000000000000000000 : node559;
													assign node559 = (inp[6]) ? 40'b0010000000001000000000000010100000000000 : 40'b1010000000000100000100000010100000000000;
												assign node563 = (inp[2]) ? node567 : node564;
													assign node564 = (inp[10]) ? 40'b0010000000001000000000000010000000000000 : 40'b0010000000001100000000000010000000000000;
													assign node567 = (inp[13]) ? 40'b1010000000000000000000000001000000000000 : 40'b0010000000001100000000000011100000000000;
						assign node570 = (inp[3]) ? node628 : node571;
							assign node571 = (inp[11]) ? node603 : node572;
								assign node572 = (inp[14]) ? node574 : 40'b0000000000000000000000000000000000000000;
									assign node574 = (inp[10]) ? node582 : node575;
										assign node575 = (inp[15]) ? node577 : 40'b0000000000000000000000000000000000000000;
											assign node577 = (inp[13]) ? node579 : 40'b0000000000000000000000000000000000000000;
												assign node579 = (inp[0]) ? 40'b0000001100001100000000000011000000000000 : 40'b0000000000000000000000000000000000000000;
										assign node582 = (inp[0]) ? node590 : node583;
											assign node583 = (inp[13]) ? node585 : 40'b0000000000000000000000000000000000000000;
												assign node585 = (inp[15]) ? node587 : 40'b0000000000000000000000000000000000000000;
													assign node587 = (inp[5]) ? 40'b0001001100000000000100000011000000000000 : 40'b1001001100000000000000000010000000000000;
											assign node590 = (inp[6]) ? node598 : node591;
												assign node591 = (inp[15]) ? node595 : node592;
													assign node592 = (inp[13]) ? 40'b1000001100010000000000000000000000000000 : 40'b0000000000000000000000000000000000000000;
													assign node595 = (inp[13]) ? 40'b0000000000000000000000000000000000000000 : 40'b1000001100000000000000000001100000000000;
												assign node598 = (inp[5]) ? 40'b0000000000000000000000000000000000000000 : node599;
													assign node599 = (inp[13]) ? 40'b0000001100011000000000000010000000000000 : 40'b0000001100001000000000000010100000000000;
								assign node603 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node604;
									assign node604 = (inp[15]) ? node616 : node605;
										assign node605 = (inp[10]) ? node611 : node606;
											assign node606 = (inp[0]) ? node608 : 40'b0000000000000000000000000000000000000000;
												assign node608 = (inp[13]) ? 40'b1000001000010100000000000000000000001000 : 40'b1000001000010100000000000000100000001000;
											assign node611 = (inp[0]) ? 40'b0000000000000000000000000000000000000000 : node612;
												assign node612 = (inp[13]) ? 40'b1001001000010000000000000000000000001000 : 40'b1001001000010000000000000000100000001000;
										assign node616 = (inp[0]) ? node622 : node617;
											assign node617 = (inp[10]) ? node619 : 40'b0000000000000000000000000000000000000000;
												assign node619 = (inp[13]) ? 40'b0001001000000000000100000010000000001000 : 40'b0001001000000000000100000010100000001000;
											assign node622 = (inp[10]) ? 40'b0000000000000000000000000000000000000000 : node623;
												assign node623 = (inp[13]) ? 40'b0000001000000100000100000010000000001000 : 40'b0000001000000100000100000010100000001000;
							assign node628 = (inp[13]) ? node696 : node629;
								assign node629 = (inp[11]) ? node663 : node630;
									assign node630 = (inp[14]) ? node632 : 40'b0000000000000000000000000000000000000000;
										assign node632 = (inp[0]) ? node648 : node633;
											assign node633 = (inp[15]) ? node641 : node634;
												assign node634 = (inp[10]) ? node638 : node635;
													assign node635 = (inp[5]) ? 40'b0001001000010100000100000010100000000000 : 40'b0001001000010100000000000001100000000000;
													assign node638 = (inp[5]) ? 40'b1001001000010000000000000001100000000000 : 40'b1001001000010000000000000010100000000000;
												assign node641 = (inp[2]) ? node645 : node642;
													assign node642 = (inp[5]) ? 40'b1001001000000100000000000001100000000000 : 40'b1001001000001100000000000010100000000000;
													assign node645 = (inp[6]) ? 40'b0001001000000000000100000011100000000000 : 40'b1001001000000000000000000001100000000000;
											assign node648 = (inp[15]) ? node656 : node649;
												assign node649 = (inp[6]) ? node653 : node650;
													assign node650 = (inp[12]) ? 40'b0000001000011000000100000010100000000000 : 40'b0000001000010000000100000010100000000000;
													assign node653 = (inp[5]) ? 40'b0000001000010000000000000001100000000000 : 40'b0000001000011000000000000010100000000000;
												assign node656 = (inp[5]) ? node660 : node657;
													assign node657 = (inp[6]) ? 40'b0000001000001000000000000010100000000000 : 40'b1000001000000000000000000001100000000000;
													assign node660 = (inp[6]) ? 40'b0000001000000100000000000001100000000000 : 40'b0000001000000100000100000010100000000000;
									assign node663 = (inp[14]) ? 40'b0000000000000000000000000000000000000000 : node664;
										assign node664 = (inp[0]) ? node680 : node665;
											assign node665 = (inp[15]) ? node673 : node666;
												assign node666 = (inp[10]) ? node670 : node667;
													assign node667 = (inp[2]) ? 40'b1001001000010100000100000010100000001000 : 40'b0001001000011100000000000010100000001000;
													assign node670 = (inp[2]) ? 40'b1001001000010000000000000001100000001000 : 40'b1001001000010000000000000010100000001000;
												assign node673 = (inp[6]) ? node677 : node674;
													assign node674 = (inp[12]) ? 40'b0001001000001000000100000010100000001000 : 40'b1001001000000000000100000010100000001000;
													assign node677 = (inp[2]) ? 40'b0001001000000000000000000011100000001000 : 40'b0001001000001000000000000010100000001000;
											assign node680 = (inp[10]) ? node688 : node681;
												assign node681 = (inp[15]) ? node685 : node682;
													assign node682 = (inp[12]) ? 40'b0000001000011100000000000010100000001000 : 40'b1000001000010100000100000010100000001000;
													assign node685 = (inp[6]) ? 40'b0000001000001100000000000010100000001000 : 40'b1000001000000100000000000000100000001000;
												assign node688 = (inp[5]) ? node692 : node689;
													assign node689 = (inp[2]) ? 40'b0000001000011000000100000010100000001000 : 40'b0000001000011000000000000010100000001000;
													assign node692 = (inp[15]) ? 40'b0000001000000000000100000010100000001000 : 40'b0000001000010000000000000001100000001000;
								assign node696 = (inp[14]) ? node728 : node697;
									assign node697 = (inp[11]) ? node699 : 40'b0000000000000000000000000000000000000000;
										assign node699 = (inp[10]) ? node713 : node700;
											assign node700 = (inp[0]) ? node706 : node701;
												assign node701 = (inp[12]) ? node703 : 40'b1001001000010100000000000000000000001000;
													assign node703 = (inp[5]) ? 40'b0001001000010100000100000011000000001000 : 40'b0001001000011100000000000011000000001000;
												assign node706 = (inp[15]) ? node710 : node707;
													assign node707 = (inp[5]) ? 40'b0000001000010100000100000010000000001000 : 40'b1000001000011100000000000010000000001000;
													assign node710 = (inp[12]) ? 40'b0000001000001100000000000010000000001000 : 40'b1000001000000100000100000010000000001000;
											assign node713 = (inp[15]) ? node721 : node714;
												assign node714 = (inp[12]) ? node718 : node715;
													assign node715 = (inp[2]) ? 40'b0000001000010000000100000010000000001000 : 40'b1001001000010000000000000000000000001000;
													assign node718 = (inp[0]) ? 40'b0000001000011000000000000011000000001000 : 40'b0001001000011000000000000010000000001000;
												assign node721 = (inp[6]) ? node725 : node722;
													assign node722 = (inp[5]) ? 40'b0001001000000000000100000010000000001000 : 40'b1000001000000000000000000000000000001000;
													assign node725 = (inp[5]) ? 40'b0001001000000000000000000011000000001000 : 40'b0000001000001000000000000010000000001000;
									assign node728 = (inp[11]) ? 40'b0000000000000000000000000000000000000000 : node729;
										assign node729 = (inp[10]) ? node745 : node730;
											assign node730 = (inp[0]) ? node738 : node731;
												assign node731 = (inp[15]) ? node735 : node732;
													assign node732 = (inp[5]) ? 40'b1001001000010100000000000000000000000000 : 40'b0001001000011100000000000010000000000000;
													assign node735 = (inp[2]) ? 40'b0001001000000100000100000010000000000000 : 40'b1001001000001100000000000010000000000000;
												assign node738 = (inp[15]) ? node742 : node739;
													assign node739 = (inp[2]) ? 40'b0000001000010100000000000001000000000000 : 40'b0000001000011100000000000010000000000000;
													assign node742 = (inp[6]) ? 40'b0000001000000100000000000001000000000000 : 40'b1000001000000100000000000000000000000000;
											assign node745 = (inp[15]) ? node753 : node746;
												assign node746 = (inp[6]) ? node750 : node747;
													assign node747 = (inp[12]) ? 40'b0000001000011000000100000010000000000000 : 40'b0000001000010000000100000010000000000000;
													assign node750 = (inp[12]) ? 40'b0001001000011000000000000011000000000000 : 40'b1000001000010000000000000000000000000000;
												assign node753 = (inp[2]) ? node757 : node754;
													assign node754 = (inp[5]) ? 40'b0000001000001000000100000010000000000000 : 40'b0000001000001000000000000010000000000000;
													assign node757 = (inp[12]) ? 40'b0001001000000000000000000001000000000000 : 40'b0001001000000000000100000010000000000000;

endmodule