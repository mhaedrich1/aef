module dtc_split125_bm91 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node18;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node30;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node39;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node44;
	wire [3-1:0] node48;
	wire [3-1:0] node49;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node60;
	wire [3-1:0] node63;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node81;
	wire [3-1:0] node82;
	wire [3-1:0] node83;
	wire [3-1:0] node84;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node102;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node114;
	wire [3-1:0] node115;
	wire [3-1:0] node116;
	wire [3-1:0] node119;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node149;
	wire [3-1:0] node150;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node165;
	wire [3-1:0] node168;
	wire [3-1:0] node170;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node176;
	wire [3-1:0] node179;
	wire [3-1:0] node181;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node186;
	wire [3-1:0] node189;
	wire [3-1:0] node192;
	wire [3-1:0] node194;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node211;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node217;
	wire [3-1:0] node220;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node224;
	wire [3-1:0] node229;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node239;
	wire [3-1:0] node243;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node250;
	wire [3-1:0] node252;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node261;
	wire [3-1:0] node264;
	wire [3-1:0] node265;
	wire [3-1:0] node267;
	wire [3-1:0] node268;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node282;
	wire [3-1:0] node283;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node287;
	wire [3-1:0] node289;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node296;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node302;
	wire [3-1:0] node303;
	wire [3-1:0] node306;
	wire [3-1:0] node307;
	wire [3-1:0] node311;
	wire [3-1:0] node312;
	wire [3-1:0] node314;
	wire [3-1:0] node315;
	wire [3-1:0] node316;
	wire [3-1:0] node320;
	wire [3-1:0] node323;
	wire [3-1:0] node325;
	wire [3-1:0] node327;
	wire [3-1:0] node330;
	wire [3-1:0] node331;
	wire [3-1:0] node332;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node339;
	wire [3-1:0] node340;
	wire [3-1:0] node342;
	wire [3-1:0] node345;

	assign outp = (inp[3]) ? node264 : node1;
		assign node1 = (inp[9]) ? node123 : node2;
			assign node2 = (inp[1]) ? node70 : node3;
				assign node3 = (inp[5]) ? node33 : node4;
					assign node4 = (inp[0]) ? node22 : node5;
						assign node5 = (inp[11]) ? node11 : node6;
							assign node6 = (inp[10]) ? 3'b000 : node7;
								assign node7 = (inp[8]) ? 3'b001 : 3'b000;
							assign node11 = (inp[10]) ? 3'b001 : node12;
								assign node12 = (inp[8]) ? node18 : node13;
									assign node13 = (inp[6]) ? 3'b000 : node14;
										assign node14 = (inp[2]) ? 3'b000 : 3'b001;
									assign node18 = (inp[7]) ? 3'b000 : 3'b001;
						assign node22 = (inp[7]) ? node24 : 3'b000;
							assign node24 = (inp[6]) ? node28 : node25;
								assign node25 = (inp[4]) ? 3'b001 : 3'b000;
								assign node28 = (inp[10]) ? node30 : 3'b000;
									assign node30 = (inp[4]) ? 3'b000 : 3'b001;
					assign node33 = (inp[11]) ? node53 : node34;
						assign node34 = (inp[8]) ? node48 : node35;
							assign node35 = (inp[10]) ? node39 : node36;
								assign node36 = (inp[4]) ? 3'b000 : 3'b001;
								assign node39 = (inp[7]) ? node41 : 3'b001;
									assign node41 = (inp[2]) ? 3'b000 : node42;
										assign node42 = (inp[6]) ? node44 : 3'b001;
											assign node44 = (inp[4]) ? 3'b001 : 3'b000;
							assign node48 = (inp[2]) ? 3'b001 : node49;
								assign node49 = (inp[4]) ? 3'b001 : 3'b000;
						assign node53 = (inp[2]) ? node63 : node54;
							assign node54 = (inp[6]) ? node56 : 3'b000;
								assign node56 = (inp[0]) ? node60 : node57;
									assign node57 = (inp[4]) ? 3'b000 : 3'b001;
									assign node60 = (inp[4]) ? 3'b001 : 3'b000;
							assign node63 = (inp[4]) ? 3'b000 : node64;
								assign node64 = (inp[6]) ? 3'b000 : node65;
									assign node65 = (inp[7]) ? 3'b001 : 3'b000;
				assign node70 = (inp[8]) ? node90 : node71;
					assign node71 = (inp[6]) ? node81 : node72;
						assign node72 = (inp[7]) ? node74 : 3'b001;
							assign node74 = (inp[4]) ? node76 : 3'b000;
								assign node76 = (inp[5]) ? 3'b001 : node77;
									assign node77 = (inp[10]) ? 3'b000 : 3'b001;
						assign node81 = (inp[11]) ? 3'b000 : node82;
							assign node82 = (inp[2]) ? 3'b001 : node83;
								assign node83 = (inp[5]) ? 3'b000 : node84;
									assign node84 = (inp[4]) ? 3'b000 : 3'b001;
					assign node90 = (inp[6]) ? node114 : node91;
						assign node91 = (inp[4]) ? node105 : node92;
							assign node92 = (inp[2]) ? node100 : node93;
								assign node93 = (inp[10]) ? 3'b001 : node94;
									assign node94 = (inp[11]) ? node96 : 3'b001;
										assign node96 = (inp[7]) ? 3'b000 : 3'b001;
								assign node100 = (inp[5]) ? node102 : 3'b000;
									assign node102 = (inp[7]) ? 3'b000 : 3'b001;
							assign node105 = (inp[5]) ? 3'b000 : node106;
								assign node106 = (inp[7]) ? 3'b001 : node107;
									assign node107 = (inp[10]) ? 3'b000 : node108;
										assign node108 = (inp[11]) ? 3'b001 : 3'b000;
						assign node114 = (inp[7]) ? 3'b001 : node115;
							assign node115 = (inp[5]) ? node119 : node116;
								assign node116 = (inp[0]) ? 3'b000 : 3'b001;
								assign node119 = (inp[0]) ? 3'b001 : 3'b000;
			assign node123 = (inp[4]) ? node197 : node124;
				assign node124 = (inp[6]) ? node158 : node125;
					assign node125 = (inp[0]) ? node141 : node126;
						assign node126 = (inp[1]) ? node132 : node127;
							assign node127 = (inp[5]) ? node129 : 3'b010;
								assign node129 = (inp[7]) ? 3'b010 : 3'b100;
							assign node132 = (inp[2]) ? node138 : node133;
								assign node133 = (inp[11]) ? node135 : 3'b101;
									assign node135 = (inp[10]) ? 3'b110 : 3'b010;
								assign node138 = (inp[10]) ? 3'b001 : 3'b101;
						assign node141 = (inp[5]) ? node149 : node142;
							assign node142 = (inp[8]) ? node146 : node143;
								assign node143 = (inp[1]) ? 3'b101 : 3'b001;
								assign node146 = (inp[11]) ? 3'b000 : 3'b001;
							assign node149 = (inp[11]) ? 3'b110 : node150;
								assign node150 = (inp[10]) ? 3'b111 : node151;
									assign node151 = (inp[2]) ? 3'b101 : node152;
										assign node152 = (inp[8]) ? 3'b101 : 3'b110;
					assign node158 = (inp[1]) ? node184 : node159;
						assign node159 = (inp[5]) ? node173 : node160;
							assign node160 = (inp[2]) ? node168 : node161;
								assign node161 = (inp[0]) ? node165 : node162;
									assign node162 = (inp[8]) ? 3'b101 : 3'b001;
									assign node165 = (inp[11]) ? 3'b001 : 3'b011;
								assign node168 = (inp[7]) ? node170 : 3'b101;
									assign node170 = (inp[10]) ? 3'b111 : 3'b001;
							assign node173 = (inp[0]) ? node179 : node174;
								assign node174 = (inp[7]) ? node176 : 3'b110;
									assign node176 = (inp[11]) ? 3'b110 : 3'b010;
								assign node179 = (inp[2]) ? node181 : 3'b101;
									assign node181 = (inp[7]) ? 3'b001 : 3'b101;
						assign node184 = (inp[5]) ? node192 : node185;
							assign node185 = (inp[10]) ? node189 : node186;
								assign node186 = (inp[7]) ? 3'b001 : 3'b011;
								assign node189 = (inp[8]) ? 3'b111 : 3'b011;
							assign node192 = (inp[8]) ? node194 : 3'b001;
								assign node194 = (inp[0]) ? 3'b011 : 3'b001;
				assign node197 = (inp[0]) ? node235 : node198;
					assign node198 = (inp[6]) ? node220 : node199;
						assign node199 = (inp[5]) ? node211 : node200;
							assign node200 = (inp[11]) ? 3'b100 : node201;
								assign node201 = (inp[10]) ? node203 : 3'b100;
									assign node203 = (inp[8]) ? node207 : node204;
										assign node204 = (inp[1]) ? 3'b000 : 3'b100;
										assign node207 = (inp[1]) ? 3'b100 : 3'b000;
							assign node211 = (inp[1]) ? node213 : 3'b000;
								assign node213 = (inp[2]) ? node217 : node214;
									assign node214 = (inp[7]) ? 3'b010 : 3'b000;
									assign node217 = (inp[11]) ? 3'b110 : 3'b100;
						assign node220 = (inp[11]) ? node232 : node221;
							assign node221 = (inp[8]) ? node229 : node222;
								assign node222 = (inp[7]) ? 3'b110 : node223;
									assign node223 = (inp[5]) ? 3'b100 : node224;
										assign node224 = (inp[1]) ? 3'b110 : 3'b100;
								assign node229 = (inp[1]) ? 3'b110 : 3'b010;
							assign node232 = (inp[7]) ? 3'b001 : 3'b100;
					assign node235 = (inp[6]) ? node255 : node236;
						assign node236 = (inp[7]) ? node250 : node237;
							assign node237 = (inp[8]) ? node243 : node238;
								assign node238 = (inp[1]) ? 3'b100 : node239;
									assign node239 = (inp[5]) ? 3'b000 : 3'b010;
								assign node243 = (inp[5]) ? node245 : 3'b100;
									assign node245 = (inp[11]) ? 3'b010 : node246;
										assign node246 = (inp[10]) ? 3'b100 : 3'b110;
							assign node250 = (inp[1]) ? node252 : 3'b010;
								assign node252 = (inp[5]) ? 3'b010 : 3'b110;
						assign node255 = (inp[5]) ? node259 : node256;
							assign node256 = (inp[7]) ? 3'b101 : 3'b001;
							assign node259 = (inp[1]) ? node261 : 3'b010;
								assign node261 = (inp[8]) ? 3'b001 : 3'b110;
		assign node264 = (inp[6]) ? node282 : node265;
			assign node265 = (inp[0]) ? node267 : 3'b000;
				assign node267 = (inp[4]) ? 3'b000 : node268;
					assign node268 = (inp[9]) ? node270 : 3'b000;
						assign node270 = (inp[1]) ? node272 : 3'b000;
							assign node272 = (inp[8]) ? node276 : node273;
								assign node273 = (inp[7]) ? 3'b100 : 3'b000;
								assign node276 = (inp[5]) ? node278 : 3'b100;
									assign node278 = (inp[2]) ? 3'b100 : 3'b000;
			assign node282 = (inp[9]) ? node330 : node283;
				assign node283 = (inp[4]) ? node299 : node284;
					assign node284 = (inp[0]) ? node292 : node285;
						assign node285 = (inp[2]) ? node287 : 3'b010;
							assign node287 = (inp[1]) ? node289 : 3'b010;
								assign node289 = (inp[11]) ? 3'b011 : 3'b010;
						assign node292 = (inp[5]) ? node294 : 3'b011;
							assign node294 = (inp[1]) ? node296 : 3'b010;
								assign node296 = (inp[7]) ? 3'b011 : 3'b010;
					assign node299 = (inp[0]) ? node311 : node300;
						assign node300 = (inp[11]) ? node302 : 3'b000;
							assign node302 = (inp[7]) ? node306 : node303;
								assign node303 = (inp[5]) ? 3'b100 : 3'b000;
								assign node306 = (inp[10]) ? 3'b000 : node307;
									assign node307 = (inp[2]) ? 3'b100 : 3'b110;
						assign node311 = (inp[10]) ? node323 : node312;
							assign node312 = (inp[7]) ? node314 : 3'b010;
								assign node314 = (inp[1]) ? node320 : node315;
									assign node315 = (inp[5]) ? 3'b010 : node316;
										assign node316 = (inp[2]) ? 3'b010 : 3'b110;
									assign node320 = (inp[5]) ? 3'b110 : 3'b101;
							assign node323 = (inp[7]) ? node325 : 3'b100;
								assign node325 = (inp[1]) ? node327 : 3'b100;
									assign node327 = (inp[8]) ? 3'b110 : 3'b010;
				assign node330 = (inp[4]) ? 3'b000 : node331;
					assign node331 = (inp[5]) ? node339 : node332;
						assign node332 = (inp[0]) ? node334 : 3'b000;
							assign node334 = (inp[7]) ? node336 : 3'b010;
								assign node336 = (inp[1]) ? 3'b110 : 3'b010;
						assign node339 = (inp[0]) ? node345 : node340;
							assign node340 = (inp[10]) ? node342 : 3'b000;
								assign node342 = (inp[2]) ? 3'b100 : 3'b000;
							assign node345 = (inp[8]) ? 3'b100 : 3'b010;

endmodule