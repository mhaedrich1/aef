module dtc_split33_bm39 (
	input  wire [14-1:0] inp,
	output wire [14-1:0] outp
);

	wire [14-1:0] node1;
	wire [14-1:0] node3;
	wire [14-1:0] node4;
	wire [14-1:0] node5;
	wire [14-1:0] node6;
	wire [14-1:0] node7;
	wire [14-1:0] node8;
	wire [14-1:0] node9;
	wire [14-1:0] node10;
	wire [14-1:0] node12;
	wire [14-1:0] node14;
	wire [14-1:0] node16;
	wire [14-1:0] node19;
	wire [14-1:0] node20;
	wire [14-1:0] node21;
	wire [14-1:0] node22;
	wire [14-1:0] node24;
	wire [14-1:0] node28;
	wire [14-1:0] node29;
	wire [14-1:0] node32;
	wire [14-1:0] node33;
	wire [14-1:0] node37;
	wire [14-1:0] node38;
	wire [14-1:0] node40;
	wire [14-1:0] node43;
	wire [14-1:0] node46;
	wire [14-1:0] node47;
	wire [14-1:0] node48;
	wire [14-1:0] node50;
	wire [14-1:0] node53;
	wire [14-1:0] node54;
	wire [14-1:0] node56;
	wire [14-1:0] node59;
	wire [14-1:0] node60;
	wire [14-1:0] node61;
	wire [14-1:0] node65;
	wire [14-1:0] node66;
	wire [14-1:0] node70;
	wire [14-1:0] node71;
	wire [14-1:0] node72;
	wire [14-1:0] node74;
	wire [14-1:0] node77;
	wire [14-1:0] node78;
	wire [14-1:0] node82;
	wire [14-1:0] node83;
	wire [14-1:0] node85;
	wire [14-1:0] node87;
	wire [14-1:0] node90;
	wire [14-1:0] node93;
	wire [14-1:0] node94;
	wire [14-1:0] node95;
	wire [14-1:0] node96;
	wire [14-1:0] node97;
	wire [14-1:0] node100;
	wire [14-1:0] node103;
	wire [14-1:0] node104;
	wire [14-1:0] node107;
	wire [14-1:0] node110;
	wire [14-1:0] node111;
	wire [14-1:0] node112;
	wire [14-1:0] node115;
	wire [14-1:0] node116;
	wire [14-1:0] node119;
	wire [14-1:0] node122;
	wire [14-1:0] node123;
	wire [14-1:0] node125;
	wire [14-1:0] node126;
	wire [14-1:0] node130;
	wire [14-1:0] node131;
	wire [14-1:0] node134;
	wire [14-1:0] node137;
	wire [14-1:0] node138;
	wire [14-1:0] node139;
	wire [14-1:0] node140;
	wire [14-1:0] node142;
	wire [14-1:0] node145;
	wire [14-1:0] node149;
	wire [14-1:0] node151;
	wire [14-1:0] node152;
	wire [14-1:0] node153;
	wire [14-1:0] node156;
	wire [14-1:0] node159;
	wire [14-1:0] node161;
	wire [14-1:0] node164;
	wire [14-1:0] node165;
	wire [14-1:0] node166;
	wire [14-1:0] node167;
	wire [14-1:0] node168;
	wire [14-1:0] node169;
	wire [14-1:0] node173;
	wire [14-1:0] node174;
	wire [14-1:0] node177;
	wire [14-1:0] node179;
	wire [14-1:0] node182;
	wire [14-1:0] node183;
	wire [14-1:0] node184;
	wire [14-1:0] node186;
	wire [14-1:0] node188;
	wire [14-1:0] node192;
	wire [14-1:0] node193;
	wire [14-1:0] node195;
	wire [14-1:0] node198;
	wire [14-1:0] node200;
	wire [14-1:0] node203;
	wire [14-1:0] node204;
	wire [14-1:0] node205;
	wire [14-1:0] node206;
	wire [14-1:0] node207;
	wire [14-1:0] node212;
	wire [14-1:0] node213;
	wire [14-1:0] node214;
	wire [14-1:0] node217;
	wire [14-1:0] node220;
	wire [14-1:0] node222;
	wire [14-1:0] node224;
	wire [14-1:0] node227;
	wire [14-1:0] node229;
	wire [14-1:0] node231;
	wire [14-1:0] node232;
	wire [14-1:0] node234;
	wire [14-1:0] node237;
	wire [14-1:0] node238;
	wire [14-1:0] node242;
	wire [14-1:0] node243;
	wire [14-1:0] node244;
	wire [14-1:0] node246;
	wire [14-1:0] node247;
	wire [14-1:0] node249;
	wire [14-1:0] node252;
	wire [14-1:0] node253;
	wire [14-1:0] node256;
	wire [14-1:0] node259;
	wire [14-1:0] node260;
	wire [14-1:0] node262;
	wire [14-1:0] node267;
	wire [14-1:0] node268;
	wire [14-1:0] node269;
	wire [14-1:0] node270;
	wire [14-1:0] node271;
	wire [14-1:0] node272;
	wire [14-1:0] node273;
	wire [14-1:0] node275;
	wire [14-1:0] node279;
	wire [14-1:0] node281;
	wire [14-1:0] node282;
	wire [14-1:0] node285;
	wire [14-1:0] node288;
	wire [14-1:0] node289;
	wire [14-1:0] node290;
	wire [14-1:0] node291;
	wire [14-1:0] node295;
	wire [14-1:0] node296;
	wire [14-1:0] node300;
	wire [14-1:0] node301;
	wire [14-1:0] node302;
	wire [14-1:0] node305;
	wire [14-1:0] node308;
	wire [14-1:0] node311;
	wire [14-1:0] node312;
	wire [14-1:0] node313;
	wire [14-1:0] node315;
	wire [14-1:0] node318;
	wire [14-1:0] node320;
	wire [14-1:0] node323;
	wire [14-1:0] node324;
	wire [14-1:0] node325;
	wire [14-1:0] node328;
	wire [14-1:0] node329;
	wire [14-1:0] node334;
	wire [14-1:0] node336;
	wire [14-1:0] node337;
	wire [14-1:0] node338;
	wire [14-1:0] node339;
	wire [14-1:0] node340;
	wire [14-1:0] node343;
	wire [14-1:0] node346;
	wire [14-1:0] node349;
	wire [14-1:0] node350;
	wire [14-1:0] node353;
	wire [14-1:0] node354;
	wire [14-1:0] node355;
	wire [14-1:0] node361;
	wire [14-1:0] node362;
	wire [14-1:0] node364;
	wire [14-1:0] node365;
	wire [14-1:0] node366;
	wire [14-1:0] node367;
	wire [14-1:0] node370;
	wire [14-1:0] node373;
	wire [14-1:0] node374;
	wire [14-1:0] node378;
	wire [14-1:0] node379;
	wire [14-1:0] node380;
	wire [14-1:0] node381;
	wire [14-1:0] node385;
	wire [14-1:0] node388;
	wire [14-1:0] node390;
	wire [14-1:0] node394;
	wire [14-1:0] node395;
	wire [14-1:0] node396;
	wire [14-1:0] node397;
	wire [14-1:0] node398;
	wire [14-1:0] node399;
	wire [14-1:0] node400;
	wire [14-1:0] node402;
	wire [14-1:0] node404;
	wire [14-1:0] node405;
	wire [14-1:0] node409;
	wire [14-1:0] node410;
	wire [14-1:0] node412;
	wire [14-1:0] node416;
	wire [14-1:0] node417;
	wire [14-1:0] node418;
	wire [14-1:0] node420;
	wire [14-1:0] node421;
	wire [14-1:0] node424;
	wire [14-1:0] node427;
	wire [14-1:0] node428;
	wire [14-1:0] node432;
	wire [14-1:0] node433;
	wire [14-1:0] node437;
	wire [14-1:0] node438;
	wire [14-1:0] node439;
	wire [14-1:0] node440;
	wire [14-1:0] node444;
	wire [14-1:0] node445;
	wire [14-1:0] node448;
	wire [14-1:0] node450;
	wire [14-1:0] node453;
	wire [14-1:0] node454;
	wire [14-1:0] node455;
	wire [14-1:0] node456;
	wire [14-1:0] node460;
	wire [14-1:0] node464;
	wire [14-1:0] node465;
	wire [14-1:0] node466;
	wire [14-1:0] node467;
	wire [14-1:0] node468;
	wire [14-1:0] node469;
	wire [14-1:0] node472;
	wire [14-1:0] node473;
	wire [14-1:0] node477;
	wire [14-1:0] node480;
	wire [14-1:0] node483;
	wire [14-1:0] node484;
	wire [14-1:0] node487;
	wire [14-1:0] node489;
	wire [14-1:0] node493;
	wire [14-1:0] node494;
	wire [14-1:0] node495;
	wire [14-1:0] node496;
	wire [14-1:0] node497;
	wire [14-1:0] node498;
	wire [14-1:0] node501;
	wire [14-1:0] node502;
	wire [14-1:0] node506;
	wire [14-1:0] node507;
	wire [14-1:0] node508;
	wire [14-1:0] node511;
	wire [14-1:0] node515;
	wire [14-1:0] node516;
	wire [14-1:0] node517;
	wire [14-1:0] node520;
	wire [14-1:0] node521;
	wire [14-1:0] node524;
	wire [14-1:0] node527;
	wire [14-1:0] node528;
	wire [14-1:0] node532;
	wire [14-1:0] node534;
	wire [14-1:0] node535;
	wire [14-1:0] node536;
	wire [14-1:0] node537;
	wire [14-1:0] node538;
	wire [14-1:0] node541;
	wire [14-1:0] node544;
	wire [14-1:0] node547;
	wire [14-1:0] node549;
	wire [14-1:0] node552;
	wire [14-1:0] node555;
	wire [14-1:0] node557;
	wire [14-1:0] node558;
	wire [14-1:0] node559;
	wire [14-1:0] node560;
	wire [14-1:0] node563;
	wire [14-1:0] node564;
	wire [14-1:0] node568;
	wire [14-1:0] node569;
	wire [14-1:0] node570;
	wire [14-1:0] node571;
	wire [14-1:0] node575;
	wire [14-1:0] node581;
	wire [14-1:0] node582;
	wire [14-1:0] node583;
	wire [14-1:0] node584;
	wire [14-1:0] node585;
	wire [14-1:0] node586;
	wire [14-1:0] node587;
	wire [14-1:0] node588;
	wire [14-1:0] node589;
	wire [14-1:0] node590;
	wire [14-1:0] node593;
	wire [14-1:0] node596;
	wire [14-1:0] node598;
	wire [14-1:0] node601;
	wire [14-1:0] node602;
	wire [14-1:0] node603;
	wire [14-1:0] node606;
	wire [14-1:0] node609;
	wire [14-1:0] node610;
	wire [14-1:0] node613;
	wire [14-1:0] node614;
	wire [14-1:0] node618;
	wire [14-1:0] node619;
	wire [14-1:0] node620;
	wire [14-1:0] node624;
	wire [14-1:0] node625;
	wire [14-1:0] node626;
	wire [14-1:0] node630;
	wire [14-1:0] node633;
	wire [14-1:0] node634;
	wire [14-1:0] node635;
	wire [14-1:0] node636;
	wire [14-1:0] node639;
	wire [14-1:0] node640;
	wire [14-1:0] node642;
	wire [14-1:0] node646;
	wire [14-1:0] node647;
	wire [14-1:0] node648;
	wire [14-1:0] node652;
	wire [14-1:0] node655;
	wire [14-1:0] node656;
	wire [14-1:0] node658;
	wire [14-1:0] node659;
	wire [14-1:0] node664;
	wire [14-1:0] node665;
	wire [14-1:0] node666;
	wire [14-1:0] node667;
	wire [14-1:0] node670;
	wire [14-1:0] node671;
	wire [14-1:0] node672;
	wire [14-1:0] node674;
	wire [14-1:0] node677;
	wire [14-1:0] node679;
	wire [14-1:0] node682;
	wire [14-1:0] node685;
	wire [14-1:0] node686;
	wire [14-1:0] node687;
	wire [14-1:0] node690;
	wire [14-1:0] node692;
	wire [14-1:0] node695;
	wire [14-1:0] node696;
	wire [14-1:0] node697;
	wire [14-1:0] node698;
	wire [14-1:0] node704;
	wire [14-1:0] node705;
	wire [14-1:0] node706;
	wire [14-1:0] node708;
	wire [14-1:0] node711;
	wire [14-1:0] node712;
	wire [14-1:0] node715;
	wire [14-1:0] node716;
	wire [14-1:0] node720;
	wire [14-1:0] node721;
	wire [14-1:0] node722;
	wire [14-1:0] node724;
	wire [14-1:0] node728;
	wire [14-1:0] node729;
	wire [14-1:0] node731;
	wire [14-1:0] node733;
	wire [14-1:0] node737;
	wire [14-1:0] node738;
	wire [14-1:0] node739;
	wire [14-1:0] node740;
	wire [14-1:0] node741;
	wire [14-1:0] node742;
	wire [14-1:0] node743;
	wire [14-1:0] node744;
	wire [14-1:0] node750;
	wire [14-1:0] node751;
	wire [14-1:0] node753;
	wire [14-1:0] node757;
	wire [14-1:0] node758;
	wire [14-1:0] node759;
	wire [14-1:0] node762;
	wire [14-1:0] node764;
	wire [14-1:0] node767;
	wire [14-1:0] node768;
	wire [14-1:0] node771;
	wire [14-1:0] node772;
	wire [14-1:0] node776;
	wire [14-1:0] node777;
	wire [14-1:0] node779;
	wire [14-1:0] node780;
	wire [14-1:0] node783;
	wire [14-1:0] node788;
	wire [14-1:0] node789;
	wire [14-1:0] node790;
	wire [14-1:0] node791;
	wire [14-1:0] node793;
	wire [14-1:0] node794;
	wire [14-1:0] node795;
	wire [14-1:0] node796;
	wire [14-1:0] node803;
	wire [14-1:0] node804;
	wire [14-1:0] node805;
	wire [14-1:0] node806;
	wire [14-1:0] node807;
	wire [14-1:0] node810;
	wire [14-1:0] node811;
	wire [14-1:0] node815;
	wire [14-1:0] node818;
	wire [14-1:0] node819;
	wire [14-1:0] node821;
	wire [14-1:0] node822;
	wire [14-1:0] node823;
	wire [14-1:0] node827;
	wire [14-1:0] node830;
	wire [14-1:0] node831;
	wire [14-1:0] node833;
	wire [14-1:0] node834;
	wire [14-1:0] node838;
	wire [14-1:0] node841;
	wire [14-1:0] node842;
	wire [14-1:0] node843;
	wire [14-1:0] node844;
	wire [14-1:0] node848;
	wire [14-1:0] node850;
	wire [14-1:0] node853;
	wire [14-1:0] node854;
	wire [14-1:0] node856;
	wire [14-1:0] node860;
	wire [14-1:0] node861;
	wire [14-1:0] node863;
	wire [14-1:0] node864;
	wire [14-1:0] node865;
	wire [14-1:0] node867;
	wire [14-1:0] node869;
	wire [14-1:0] node876;
	wire [14-1:0] node877;
	wire [14-1:0] node878;
	wire [14-1:0] node879;
	wire [14-1:0] node880;
	wire [14-1:0] node881;
	wire [14-1:0] node882;
	wire [14-1:0] node883;
	wire [14-1:0] node884;
	wire [14-1:0] node885;
	wire [14-1:0] node886;
	wire [14-1:0] node888;
	wire [14-1:0] node894;
	wire [14-1:0] node895;
	wire [14-1:0] node896;
	wire [14-1:0] node897;
	wire [14-1:0] node899;
	wire [14-1:0] node902;
	wire [14-1:0] node905;
	wire [14-1:0] node908;
	wire [14-1:0] node909;
	wire [14-1:0] node910;
	wire [14-1:0] node913;
	wire [14-1:0] node916;
	wire [14-1:0] node917;
	wire [14-1:0] node918;
	wire [14-1:0] node921;
	wire [14-1:0] node925;
	wire [14-1:0] node926;
	wire [14-1:0] node927;
	wire [14-1:0] node928;
	wire [14-1:0] node929;
	wire [14-1:0] node932;
	wire [14-1:0] node935;
	wire [14-1:0] node936;
	wire [14-1:0] node939;
	wire [14-1:0] node942;
	wire [14-1:0] node943;
	wire [14-1:0] node944;
	wire [14-1:0] node945;
	wire [14-1:0] node949;
	wire [14-1:0] node952;
	wire [14-1:0] node953;
	wire [14-1:0] node957;
	wire [14-1:0] node958;
	wire [14-1:0] node959;
	wire [14-1:0] node960;
	wire [14-1:0] node962;
	wire [14-1:0] node965;
	wire [14-1:0] node966;
	wire [14-1:0] node970;
	wire [14-1:0] node971;
	wire [14-1:0] node974;
	wire [14-1:0] node976;
	wire [14-1:0] node979;
	wire [14-1:0] node980;
	wire [14-1:0] node981;
	wire [14-1:0] node982;
	wire [14-1:0] node986;
	wire [14-1:0] node988;
	wire [14-1:0] node991;
	wire [14-1:0] node992;
	wire [14-1:0] node994;
	wire [14-1:0] node997;
	wire [14-1:0] node998;
	wire [14-1:0] node1001;
	wire [14-1:0] node1002;
	wire [14-1:0] node1006;
	wire [14-1:0] node1007;
	wire [14-1:0] node1008;
	wire [14-1:0] node1009;
	wire [14-1:0] node1010;
	wire [14-1:0] node1011;
	wire [14-1:0] node1013;
	wire [14-1:0] node1014;
	wire [14-1:0] node1019;
	wire [14-1:0] node1020;
	wire [14-1:0] node1024;
	wire [14-1:0] node1025;
	wire [14-1:0] node1027;
	wire [14-1:0] node1030;
	wire [14-1:0] node1031;
	wire [14-1:0] node1034;
	wire [14-1:0] node1037;
	wire [14-1:0] node1038;
	wire [14-1:0] node1039;
	wire [14-1:0] node1040;
	wire [14-1:0] node1043;
	wire [14-1:0] node1046;
	wire [14-1:0] node1047;
	wire [14-1:0] node1049;
	wire [14-1:0] node1052;
	wire [14-1:0] node1055;
	wire [14-1:0] node1056;
	wire [14-1:0] node1058;
	wire [14-1:0] node1060;
	wire [14-1:0] node1064;
	wire [14-1:0] node1065;
	wire [14-1:0] node1066;
	wire [14-1:0] node1067;
	wire [14-1:0] node1068;
	wire [14-1:0] node1070;
	wire [14-1:0] node1074;
	wire [14-1:0] node1075;
	wire [14-1:0] node1076;
	wire [14-1:0] node1080;
	wire [14-1:0] node1082;
	wire [14-1:0] node1085;
	wire [14-1:0] node1086;
	wire [14-1:0] node1087;
	wire [14-1:0] node1090;
	wire [14-1:0] node1093;
	wire [14-1:0] node1094;
	wire [14-1:0] node1097;
	wire [14-1:0] node1100;
	wire [14-1:0] node1101;
	wire [14-1:0] node1102;
	wire [14-1:0] node1103;
	wire [14-1:0] node1106;
	wire [14-1:0] node1109;
	wire [14-1:0] node1110;
	wire [14-1:0] node1111;
	wire [14-1:0] node1114;
	wire [14-1:0] node1117;
	wire [14-1:0] node1120;
	wire [14-1:0] node1121;
	wire [14-1:0] node1123;
	wire [14-1:0] node1125;
	wire [14-1:0] node1129;
	wire [14-1:0] node1130;
	wire [14-1:0] node1131;
	wire [14-1:0] node1132;
	wire [14-1:0] node1134;
	wire [14-1:0] node1135;
	wire [14-1:0] node1136;
	wire [14-1:0] node1138;
	wire [14-1:0] node1142;
	wire [14-1:0] node1143;
	wire [14-1:0] node1146;
	wire [14-1:0] node1149;
	wire [14-1:0] node1150;
	wire [14-1:0] node1151;
	wire [14-1:0] node1152;
	wire [14-1:0] node1154;
	wire [14-1:0] node1157;
	wire [14-1:0] node1158;
	wire [14-1:0] node1160;
	wire [14-1:0] node1164;
	wire [14-1:0] node1166;
	wire [14-1:0] node1169;
	wire [14-1:0] node1170;
	wire [14-1:0] node1171;
	wire [14-1:0] node1174;
	wire [14-1:0] node1176;
	wire [14-1:0] node1179;
	wire [14-1:0] node1180;
	wire [14-1:0] node1184;
	wire [14-1:0] node1185;
	wire [14-1:0] node1186;
	wire [14-1:0] node1187;
	wire [14-1:0] node1188;
	wire [14-1:0] node1189;
	wire [14-1:0] node1192;
	wire [14-1:0] node1195;
	wire [14-1:0] node1196;
	wire [14-1:0] node1200;
	wire [14-1:0] node1201;
	wire [14-1:0] node1203;
	wire [14-1:0] node1206;
	wire [14-1:0] node1209;
	wire [14-1:0] node1210;
	wire [14-1:0] node1211;
	wire [14-1:0] node1213;
	wire [14-1:0] node1216;
	wire [14-1:0] node1218;
	wire [14-1:0] node1221;
	wire [14-1:0] node1222;
	wire [14-1:0] node1223;
	wire [14-1:0] node1226;
	wire [14-1:0] node1229;
	wire [14-1:0] node1231;
	wire [14-1:0] node1234;
	wire [14-1:0] node1235;
	wire [14-1:0] node1236;
	wire [14-1:0] node1237;
	wire [14-1:0] node1240;
	wire [14-1:0] node1243;
	wire [14-1:0] node1245;
	wire [14-1:0] node1248;
	wire [14-1:0] node1249;
	wire [14-1:0] node1251;
	wire [14-1:0] node1254;
	wire [14-1:0] node1255;
	wire [14-1:0] node1258;
	wire [14-1:0] node1261;
	wire [14-1:0] node1262;
	wire [14-1:0] node1263;
	wire [14-1:0] node1264;
	wire [14-1:0] node1265;
	wire [14-1:0] node1268;
	wire [14-1:0] node1269;
	wire [14-1:0] node1273;
	wire [14-1:0] node1274;
	wire [14-1:0] node1276;
	wire [14-1:0] node1277;
	wire [14-1:0] node1281;
	wire [14-1:0] node1282;
	wire [14-1:0] node1286;
	wire [14-1:0] node1288;
	wire [14-1:0] node1289;
	wire [14-1:0] node1290;
	wire [14-1:0] node1291;
	wire [14-1:0] node1295;
	wire [14-1:0] node1297;
	wire [14-1:0] node1300;
	wire [14-1:0] node1301;
	wire [14-1:0] node1304;
	wire [14-1:0] node1306;
	wire [14-1:0] node1310;
	wire [14-1:0] node1311;
	wire [14-1:0] node1312;
	wire [14-1:0] node1313;
	wire [14-1:0] node1314;
	wire [14-1:0] node1315;
	wire [14-1:0] node1316;
	wire [14-1:0] node1318;
	wire [14-1:0] node1322;
	wire [14-1:0] node1323;
	wire [14-1:0] node1324;
	wire [14-1:0] node1327;
	wire [14-1:0] node1329;
	wire [14-1:0] node1332;
	wire [14-1:0] node1333;
	wire [14-1:0] node1336;
	wire [14-1:0] node1339;
	wire [14-1:0] node1340;
	wire [14-1:0] node1341;
	wire [14-1:0] node1344;
	wire [14-1:0] node1345;
	wire [14-1:0] node1346;
	wire [14-1:0] node1349;
	wire [14-1:0] node1352;
	wire [14-1:0] node1355;
	wire [14-1:0] node1356;
	wire [14-1:0] node1359;
	wire [14-1:0] node1360;
	wire [14-1:0] node1363;
	wire [14-1:0] node1366;
	wire [14-1:0] node1367;
	wire [14-1:0] node1368;
	wire [14-1:0] node1369;
	wire [14-1:0] node1370;
	wire [14-1:0] node1373;
	wire [14-1:0] node1376;
	wire [14-1:0] node1377;
	wire [14-1:0] node1378;
	wire [14-1:0] node1381;
	wire [14-1:0] node1384;
	wire [14-1:0] node1387;
	wire [14-1:0] node1388;
	wire [14-1:0] node1389;
	wire [14-1:0] node1393;
	wire [14-1:0] node1394;
	wire [14-1:0] node1398;
	wire [14-1:0] node1399;
	wire [14-1:0] node1400;
	wire [14-1:0] node1401;
	wire [14-1:0] node1404;
	wire [14-1:0] node1407;
	wire [14-1:0] node1408;
	wire [14-1:0] node1409;
	wire [14-1:0] node1413;
	wire [14-1:0] node1416;
	wire [14-1:0] node1417;
	wire [14-1:0] node1418;
	wire [14-1:0] node1421;
	wire [14-1:0] node1424;
	wire [14-1:0] node1425;
	wire [14-1:0] node1428;
	wire [14-1:0] node1430;
	wire [14-1:0] node1433;
	wire [14-1:0] node1434;
	wire [14-1:0] node1435;
	wire [14-1:0] node1436;
	wire [14-1:0] node1437;
	wire [14-1:0] node1438;
	wire [14-1:0] node1441;
	wire [14-1:0] node1444;
	wire [14-1:0] node1445;
	wire [14-1:0] node1446;
	wire [14-1:0] node1450;
	wire [14-1:0] node1452;
	wire [14-1:0] node1456;
	wire [14-1:0] node1457;
	wire [14-1:0] node1458;
	wire [14-1:0] node1459;
	wire [14-1:0] node1462;
	wire [14-1:0] node1465;
	wire [14-1:0] node1467;
	wire [14-1:0] node1470;
	wire [14-1:0] node1471;
	wire [14-1:0] node1473;
	wire [14-1:0] node1476;
	wire [14-1:0] node1477;
	wire [14-1:0] node1480;
	wire [14-1:0] node1483;
	wire [14-1:0] node1484;
	wire [14-1:0] node1485;
	wire [14-1:0] node1486;
	wire [14-1:0] node1488;
	wire [14-1:0] node1491;
	wire [14-1:0] node1492;
	wire [14-1:0] node1495;
	wire [14-1:0] node1497;
	wire [14-1:0] node1502;
	wire [14-1:0] node1503;
	wire [14-1:0] node1505;
	wire [14-1:0] node1506;
	wire [14-1:0] node1508;
	wire [14-1:0] node1509;
	wire [14-1:0] node1511;
	wire [14-1:0] node1514;
	wire [14-1:0] node1516;
	wire [14-1:0] node1521;
	wire [14-1:0] node1522;
	wire [14-1:0] node1523;
	wire [14-1:0] node1524;
	wire [14-1:0] node1525;
	wire [14-1:0] node1526;
	wire [14-1:0] node1527;
	wire [14-1:0] node1529;
	wire [14-1:0] node1532;
	wire [14-1:0] node1533;
	wire [14-1:0] node1534;
	wire [14-1:0] node1537;
	wire [14-1:0] node1540;
	wire [14-1:0] node1541;
	wire [14-1:0] node1544;
	wire [14-1:0] node1547;
	wire [14-1:0] node1548;
	wire [14-1:0] node1549;
	wire [14-1:0] node1550;
	wire [14-1:0] node1553;
	wire [14-1:0] node1556;
	wire [14-1:0] node1557;
	wire [14-1:0] node1561;
	wire [14-1:0] node1562;
	wire [14-1:0] node1565;
	wire [14-1:0] node1566;
	wire [14-1:0] node1569;
	wire [14-1:0] node1572;
	wire [14-1:0] node1573;
	wire [14-1:0] node1574;
	wire [14-1:0] node1575;
	wire [14-1:0] node1576;
	wire [14-1:0] node1578;
	wire [14-1:0] node1581;
	wire [14-1:0] node1584;
	wire [14-1:0] node1585;
	wire [14-1:0] node1586;
	wire [14-1:0] node1589;
	wire [14-1:0] node1593;
	wire [14-1:0] node1594;
	wire [14-1:0] node1595;
	wire [14-1:0] node1596;
	wire [14-1:0] node1599;
	wire [14-1:0] node1602;
	wire [14-1:0] node1605;
	wire [14-1:0] node1606;
	wire [14-1:0] node1609;
	wire [14-1:0] node1612;
	wire [14-1:0] node1613;
	wire [14-1:0] node1614;
	wire [14-1:0] node1615;
	wire [14-1:0] node1619;
	wire [14-1:0] node1620;
	wire [14-1:0] node1622;
	wire [14-1:0] node1625;
	wire [14-1:0] node1628;
	wire [14-1:0] node1629;
	wire [14-1:0] node1631;
	wire [14-1:0] node1633;
	wire [14-1:0] node1636;
	wire [14-1:0] node1637;
	wire [14-1:0] node1638;
	wire [14-1:0] node1642;
	wire [14-1:0] node1645;
	wire [14-1:0] node1646;
	wire [14-1:0] node1647;
	wire [14-1:0] node1648;
	wire [14-1:0] node1649;
	wire [14-1:0] node1651;
	wire [14-1:0] node1652;
	wire [14-1:0] node1655;
	wire [14-1:0] node1658;
	wire [14-1:0] node1660;
	wire [14-1:0] node1661;
	wire [14-1:0] node1664;
	wire [14-1:0] node1667;
	wire [14-1:0] node1668;
	wire [14-1:0] node1669;
	wire [14-1:0] node1670;
	wire [14-1:0] node1673;
	wire [14-1:0] node1677;
	wire [14-1:0] node1678;
	wire [14-1:0] node1679;
	wire [14-1:0] node1682;
	wire [14-1:0] node1685;
	wire [14-1:0] node1687;
	wire [14-1:0] node1690;
	wire [14-1:0] node1692;
	wire [14-1:0] node1693;
	wire [14-1:0] node1694;
	wire [14-1:0] node1697;
	wire [14-1:0] node1700;
	wire [14-1:0] node1701;
	wire [14-1:0] node1705;
	wire [14-1:0] node1706;
	wire [14-1:0] node1707;
	wire [14-1:0] node1708;
	wire [14-1:0] node1711;
	wire [14-1:0] node1712;
	wire [14-1:0] node1715;
	wire [14-1:0] node1720;
	wire [14-1:0] node1721;
	wire [14-1:0] node1722;
	wire [14-1:0] node1723;
	wire [14-1:0] node1724;
	wire [14-1:0] node1725;
	wire [14-1:0] node1731;
	wire [14-1:0] node1732;
	wire [14-1:0] node1733;
	wire [14-1:0] node1735;
	wire [14-1:0] node1736;
	wire [14-1:0] node1737;
	wire [14-1:0] node1740;
	wire [14-1:0] node1743;
	wire [14-1:0] node1746;
	wire [14-1:0] node1747;
	wire [14-1:0] node1748;
	wire [14-1:0] node1749;
	wire [14-1:0] node1753;
	wire [14-1:0] node1756;
	wire [14-1:0] node1757;
	wire [14-1:0] node1760;
	wire [14-1:0] node1763;
	wire [14-1:0] node1764;
	wire [14-1:0] node1765;
	wire [14-1:0] node1766;
	wire [14-1:0] node1770;
	wire [14-1:0] node1771;
	wire [14-1:0] node1775;
	wire [14-1:0] node1776;
	wire [14-1:0] node1781;
	wire [14-1:0] node1782;
	wire [14-1:0] node1783;
	wire [14-1:0] node1784;
	wire [14-1:0] node1785;
	wire [14-1:0] node1787;
	wire [14-1:0] node1789;
	wire [14-1:0] node1792;
	wire [14-1:0] node1793;
	wire [14-1:0] node1794;
	wire [14-1:0] node1795;
	wire [14-1:0] node1804;
	wire [14-1:0] node1805;
	wire [14-1:0] node1806;
	wire [14-1:0] node1807;
	wire [14-1:0] node1808;
	wire [14-1:0] node1809;
	wire [14-1:0] node1810;
	wire [14-1:0] node1811;
	wire [14-1:0] node1812;
	wire [14-1:0] node1815;
	wire [14-1:0] node1816;
	wire [14-1:0] node1818;
	wire [14-1:0] node1822;
	wire [14-1:0] node1823;
	wire [14-1:0] node1826;
	wire [14-1:0] node1828;
	wire [14-1:0] node1831;
	wire [14-1:0] node1832;
	wire [14-1:0] node1833;
	wire [14-1:0] node1835;
	wire [14-1:0] node1839;
	wire [14-1:0] node1841;
	wire [14-1:0] node1842;
	wire [14-1:0] node1844;
	wire [14-1:0] node1848;
	wire [14-1:0] node1849;
	wire [14-1:0] node1850;
	wire [14-1:0] node1851;
	wire [14-1:0] node1853;
	wire [14-1:0] node1856;
	wire [14-1:0] node1857;
	wire [14-1:0] node1860;
	wire [14-1:0] node1863;
	wire [14-1:0] node1864;
	wire [14-1:0] node1866;
	wire [14-1:0] node1872;
	wire [14-1:0] node1873;
	wire [14-1:0] node1874;
	wire [14-1:0] node1875;
	wire [14-1:0] node1876;
	wire [14-1:0] node1877;
	wire [14-1:0] node1879;
	wire [14-1:0] node1882;
	wire [14-1:0] node1883;
	wire [14-1:0] node1886;
	wire [14-1:0] node1889;
	wire [14-1:0] node1890;
	wire [14-1:0] node1891;
	wire [14-1:0] node1895;
	wire [14-1:0] node1896;
	wire [14-1:0] node1899;
	wire [14-1:0] node1902;
	wire [14-1:0] node1903;
	wire [14-1:0] node1904;
	wire [14-1:0] node1907;
	wire [14-1:0] node1908;
	wire [14-1:0] node1911;
	wire [14-1:0] node1914;
	wire [14-1:0] node1915;
	wire [14-1:0] node1917;
	wire [14-1:0] node1920;
	wire [14-1:0] node1921;
	wire [14-1:0] node1924;
	wire [14-1:0] node1927;
	wire [14-1:0] node1928;
	wire [14-1:0] node1929;
	wire [14-1:0] node1930;
	wire [14-1:0] node1931;
	wire [14-1:0] node1934;
	wire [14-1:0] node1937;
	wire [14-1:0] node1938;
	wire [14-1:0] node1943;
	wire [14-1:0] node1945;
	wire [14-1:0] node1946;
	wire [14-1:0] node1947;
	wire [14-1:0] node1950;
	wire [14-1:0] node1954;
	wire [14-1:0] node1955;
	wire [14-1:0] node1956;
	wire [14-1:0] node1957;
	wire [14-1:0] node1958;
	wire [14-1:0] node1960;
	wire [14-1:0] node1963;
	wire [14-1:0] node1964;
	wire [14-1:0] node1967;
	wire [14-1:0] node1970;
	wire [14-1:0] node1971;
	wire [14-1:0] node1974;
	wire [14-1:0] node1975;
	wire [14-1:0] node1979;
	wire [14-1:0] node1980;
	wire [14-1:0] node1981;
	wire [14-1:0] node1984;
	wire [14-1:0] node1985;
	wire [14-1:0] node1991;
	wire [14-1:0] node1992;
	wire [14-1:0] node1993;
	wire [14-1:0] node1994;
	wire [14-1:0] node1995;
	wire [14-1:0] node1996;
	wire [14-1:0] node1997;
	wire [14-1:0] node2000;
	wire [14-1:0] node2001;
	wire [14-1:0] node2003;
	wire [14-1:0] node2006;
	wire [14-1:0] node2008;
	wire [14-1:0] node2011;
	wire [14-1:0] node2012;
	wire [14-1:0] node2013;
	wire [14-1:0] node2015;
	wire [14-1:0] node2018;
	wire [14-1:0] node2019;
	wire [14-1:0] node2022;
	wire [14-1:0] node2026;
	wire [14-1:0] node2027;
	wire [14-1:0] node2028;
	wire [14-1:0] node2029;
	wire [14-1:0] node2031;
	wire [14-1:0] node2034;
	wire [14-1:0] node2037;
	wire [14-1:0] node2038;
	wire [14-1:0] node2042;
	wire [14-1:0] node2043;
	wire [14-1:0] node2044;
	wire [14-1:0] node2046;
	wire [14-1:0] node2051;
	wire [14-1:0] node2052;
	wire [14-1:0] node2053;
	wire [14-1:0] node2054;
	wire [14-1:0] node2056;
	wire [14-1:0] node2060;
	wire [14-1:0] node2061;
	wire [14-1:0] node2062;
	wire [14-1:0] node2065;
	wire [14-1:0] node2068;
	wire [14-1:0] node2069;
	wire [14-1:0] node2072;
	wire [14-1:0] node2075;
	wire [14-1:0] node2076;
	wire [14-1:0] node2077;
	wire [14-1:0] node2082;
	wire [14-1:0] node2084;
	wire [14-1:0] node2086;
	wire [14-1:0] node2087;
	wire [14-1:0] node2088;
	wire [14-1:0] node2089;
	wire [14-1:0] node2090;
	wire [14-1:0] node2094;
	wire [14-1:0] node2095;
	wire [14-1:0] node2098;
	wire [14-1:0] node2101;
	wire [14-1:0] node2104;
	wire [14-1:0] node2105;
	wire [14-1:0] node2106;
	wire [14-1:0] node2109;
	wire [14-1:0] node2112;
	wire [14-1:0] node2114;
	wire [14-1:0] node2118;
	wire [14-1:0] node2119;
	wire [14-1:0] node2120;
	wire [14-1:0] node2121;
	wire [14-1:0] node2122;
	wire [14-1:0] node2123;
	wire [14-1:0] node2124;
	wire [14-1:0] node2125;
	wire [14-1:0] node2127;
	wire [14-1:0] node2131;
	wire [14-1:0] node2132;
	wire [14-1:0] node2136;
	wire [14-1:0] node2138;
	wire [14-1:0] node2139;
	wire [14-1:0] node2140;
	wire [14-1:0] node2143;
	wire [14-1:0] node2146;
	wire [14-1:0] node2148;
	wire [14-1:0] node2151;
	wire [14-1:0] node2153;
	wire [14-1:0] node2154;
	wire [14-1:0] node2155;
	wire [14-1:0] node2157;
	wire [14-1:0] node2160;
	wire [14-1:0] node2161;
	wire [14-1:0] node2165;
	wire [14-1:0] node2166;
	wire [14-1:0] node2167;
	wire [14-1:0] node2172;
	wire [14-1:0] node2173;
	wire [14-1:0] node2174;
	wire [14-1:0] node2175;
	wire [14-1:0] node2176;
	wire [14-1:0] node2178;
	wire [14-1:0] node2180;
	wire [14-1:0] node2184;
	wire [14-1:0] node2185;
	wire [14-1:0] node2186;
	wire [14-1:0] node2189;
	wire [14-1:0] node2196;
	wire [14-1:0] node2197;
	wire [14-1:0] node2198;
	wire [14-1:0] node2199;
	wire [14-1:0] node2200;
	wire [14-1:0] node2201;
	wire [14-1:0] node2202;
	wire [14-1:0] node2206;
	wire [14-1:0] node2207;
	wire [14-1:0] node2209;
	wire [14-1:0] node2210;
	wire [14-1:0] node2214;
	wire [14-1:0] node2215;
	wire [14-1:0] node2220;
	wire [14-1:0] node2222;
	wire [14-1:0] node2224;
	wire [14-1:0] node2226;
	wire [14-1:0] node2228;
	wire [14-1:0] node2231;
	wire [14-1:0] node2233;
	wire [14-1:0] node2235;
	wire [14-1:0] node2237;
	wire [14-1:0] node2239;
	wire [14-1:0] node2242;
	wire [14-1:0] node2243;
	wire [14-1:0] node2245;
	wire [14-1:0] node2247;
	wire [14-1:0] node2249;
	wire [14-1:0] node2251;

	assign outp = (inp[13]) ? node876 : node1;
		assign node1 = (inp[8]) ? node3 : 14'b00000000000000;
			assign node3 = (inp[11]) ? node581 : node4;
				assign node4 = (inp[0]) ? node394 : node5;
					assign node5 = (inp[3]) ? node267 : node6;
						assign node6 = (inp[4]) ? node164 : node7;
							assign node7 = (inp[5]) ? node93 : node8;
								assign node8 = (inp[10]) ? node46 : node9;
									assign node9 = (inp[12]) ? node19 : node10;
										assign node10 = (inp[2]) ? node12 : 14'b00000000000001;
											assign node12 = (inp[9]) ? node14 : 14'b00001010110000;
												assign node14 = (inp[1]) ? node16 : 14'b00011100010000;
													assign node16 = (inp[6]) ? 14'b00001000010000 : 14'b00001000000000;
										assign node19 = (inp[1]) ? node37 : node20;
											assign node20 = (inp[6]) ? node28 : node21;
												assign node21 = (inp[7]) ? 14'b00001110110110 : node22;
													assign node22 = (inp[9]) ? node24 : 14'b00000000000001;
														assign node24 = (inp[2]) ? 14'b00001100000110 : 14'b01001100000110;
												assign node28 = (inp[9]) ? node32 : node29;
													assign node29 = (inp[7]) ? 14'b00001100110110 : 14'b00011100110110;
													assign node32 = (inp[7]) ? 14'b00001100010110 : node33;
														assign node33 = (inp[2]) ? 14'b00011100010110 : 14'b01011100010110;
											assign node37 = (inp[6]) ? node43 : node38;
												assign node38 = (inp[7]) ? node40 : 14'b01011010000110;
													assign node40 = (inp[9]) ? 14'b01001010010110 : 14'b01001010110110;
												assign node43 = (inp[2]) ? 14'b00001000110110 : 14'b01001000110110;
									assign node46 = (inp[7]) ? node70 : node47;
										assign node47 = (inp[6]) ? node53 : node48;
											assign node48 = (inp[1]) ? node50 : 14'b00000000000001;
												assign node50 = (inp[12]) ? 14'b01001000000010 : 14'b00101000000010;
											assign node53 = (inp[9]) ? node59 : node54;
												assign node54 = (inp[2]) ? node56 : 14'b01011000110010;
													assign node56 = (inp[12]) ? 14'b00011000110010 : 14'b00111000110010;
												assign node59 = (inp[2]) ? node65 : node60;
													assign node60 = (inp[12]) ? 14'b01011100010010 : node61;
														assign node61 = (inp[1]) ? 14'b01111000010010 : 14'b01111100010010;
													assign node65 = (inp[12]) ? 14'b00011000010010 : node66;
														assign node66 = (inp[1]) ? 14'b00111000010010 : 14'b00111100010010;
										assign node70 = (inp[2]) ? node82 : node71;
											assign node71 = (inp[12]) ? node77 : node72;
												assign node72 = (inp[6]) ? node74 : 14'b01101110010010;
													assign node74 = (inp[9]) ? 14'b01101100010010 : 14'b01101100110010;
												assign node77 = (inp[1]) ? 14'b01001000010010 : node78;
													assign node78 = (inp[6]) ? 14'b01001100110010 : 14'b01001110110010;
											assign node82 = (inp[6]) ? node90 : node83;
												assign node83 = (inp[9]) ? node85 : 14'b00101110110010;
													assign node85 = (inp[1]) ? node87 : 14'b00001110010010;
														assign node87 = (inp[12]) ? 14'b00001010010010 : 14'b00101010010010;
												assign node90 = (inp[1]) ? 14'b00001000110010 : 14'b00001100110010;
								assign node93 = (inp[10]) ? node137 : node94;
									assign node94 = (inp[12]) ? node110 : node95;
										assign node95 = (inp[2]) ? node103 : node96;
											assign node96 = (inp[7]) ? node100 : node97;
												assign node97 = (inp[9]) ? 14'b00100000000010 : 14'b00110010000010;
												assign node100 = (inp[9]) ? 14'b00100110010010 : 14'b00100000110010;
											assign node103 = (inp[1]) ? node107 : node104;
												assign node104 = (inp[9]) ? 14'b00000110010000 : 14'b00000110110000;
												assign node107 = (inp[6]) ? 14'b00000000110000 : 14'b00000000000000;
										assign node110 = (inp[1]) ? node122 : node111;
											assign node111 = (inp[9]) ? node115 : node112;
												assign node112 = (inp[2]) ? 14'b00010100110110 : 14'b01010100110110;
												assign node115 = (inp[6]) ? node119 : node116;
													assign node116 = (inp[2]) ? 14'b00000100000110 : 14'b01000100000110;
													assign node119 = (inp[7]) ? 14'b00000100010110 : 14'b00010100010110;
											assign node122 = (inp[7]) ? node130 : node123;
												assign node123 = (inp[6]) ? node125 : 14'b01010010000110;
													assign node125 = (inp[9]) ? 14'b01010000010110 : node126;
														assign node126 = (inp[2]) ? 14'b00010000110110 : 14'b01010000110110;
												assign node130 = (inp[2]) ? node134 : node131;
													assign node131 = (inp[9]) ? 14'b01000010010110 : 14'b01000010110110;
													assign node134 = (inp[9]) ? 14'b00000010010110 : 14'b00000010110110;
									assign node137 = (inp[12]) ? node149 : node138;
										assign node138 = (inp[2]) ? 14'b00000000000001 : node139;
											assign node139 = (inp[9]) ? node145 : node140;
												assign node140 = (inp[7]) ? node142 : 14'b01110000110010;
													assign node142 = (inp[1]) ? 14'b01100010110010 : 14'b01100110110010;
												assign node145 = (inp[1]) ? 14'b01100000000010 : 14'b01100100000010;
										assign node149 = (inp[2]) ? node151 : 14'b00000000000001;
											assign node151 = (inp[7]) ? node159 : node152;
												assign node152 = (inp[1]) ? node156 : node153;
													assign node153 = (inp[9]) ? 14'b00000100000010 : 14'b00000000000001;
													assign node156 = (inp[9]) ? 14'b00000000000010 : 14'b00010010000010;
												assign node159 = (inp[6]) ? node161 : 14'b00000010110010;
													assign node161 = (inp[1]) ? 14'b00000000010010 : 14'b00000100110010;
							assign node164 = (inp[12]) ? node242 : node165;
								assign node165 = (inp[10]) ? node203 : node166;
									assign node166 = (inp[6]) ? node182 : node167;
										assign node167 = (inp[7]) ? node173 : node168;
											assign node168 = (inp[9]) ? 14'b01101100000110 : node169;
												assign node169 = (inp[1]) ? 14'b00110010000110 : 14'b00000000000001;
											assign node173 = (inp[2]) ? node177 : node174;
												assign node174 = (inp[9]) ? 14'b01100110010110 : 14'b01100010110110;
												assign node177 = (inp[1]) ? node179 : 14'b00101110110110;
													assign node179 = (inp[5]) ? 14'b00100010110110 : 14'b00101010110110;
										assign node182 = (inp[2]) ? node192 : node183;
											assign node183 = (inp[1]) ? 14'b01111000110110 : node184;
												assign node184 = (inp[5]) ? node186 : 14'b01101100110110;
													assign node186 = (inp[7]) ? node188 : 14'b01110100110110;
														assign node188 = (inp[9]) ? 14'b01100100010110 : 14'b01100100110110;
											assign node192 = (inp[7]) ? node198 : node193;
												assign node193 = (inp[9]) ? node195 : 14'b00110100110110;
													assign node195 = (inp[1]) ? 14'b00110000010110 : 14'b00110100010110;
												assign node198 = (inp[9]) ? node200 : 14'b00100000110110;
													assign node200 = (inp[1]) ? 14'b00100000010110 : 14'b00100100010110;
									assign node203 = (inp[2]) ? node227 : node204;
										assign node204 = (inp[7]) ? node212 : node205;
											assign node205 = (inp[6]) ? 14'b01111100110000 : node206;
												assign node206 = (inp[1]) ? 14'b01110010000000 : node207;
													assign node207 = (inp[9]) ? 14'b01100100000000 : 14'b00000000000001;
											assign node212 = (inp[1]) ? node220 : node213;
												assign node213 = (inp[9]) ? node217 : node214;
													assign node214 = (inp[6]) ? 14'b01101100110000 : 14'b01101110110000;
													assign node217 = (inp[6]) ? 14'b01101100010000 : 14'b01101110010000;
												assign node220 = (inp[6]) ? node222 : 14'b01100010110000;
													assign node222 = (inp[5]) ? node224 : 14'b01101000110000;
														assign node224 = (inp[9]) ? 14'b01100000010000 : 14'b01100000110000;
										assign node227 = (inp[5]) ? node229 : 14'b00000000000001;
											assign node229 = (inp[9]) ? node231 : 14'b00000000000001;
												assign node231 = (inp[6]) ? node237 : node232;
													assign node232 = (inp[7]) ? node234 : 14'b00100100000000;
														assign node234 = (inp[1]) ? 14'b00100010010000 : 14'b00100110010000;
													assign node237 = (inp[7]) ? 14'b00100000010000 : node238;
														assign node238 = (inp[1]) ? 14'b00110000010000 : 14'b00110100010000;
								assign node242 = (inp[2]) ? 14'b00000000000001 : node243;
									assign node243 = (inp[5]) ? node259 : node244;
										assign node244 = (inp[10]) ? node246 : 14'b00000000000001;
											assign node246 = (inp[9]) ? node252 : node247;
												assign node247 = (inp[1]) ? node249 : 14'b00111100110000;
													assign node249 = (inp[7]) ? 14'b00101000110000 : 14'b00111000110000;
												assign node252 = (inp[1]) ? node256 : node253;
													assign node253 = (inp[7]) ? 14'b00101100010000 : 14'b00111100010000;
													assign node256 = (inp[6]) ? 14'b00101000010000 : 14'b00101000000000;
										assign node259 = (inp[10]) ? 14'b00000000000001 : node260;
											assign node260 = (inp[7]) ? node262 : 14'b01010100110010;
												assign node262 = (inp[6]) ? 14'b01000000010010 : 14'b01000010110010;
						assign node267 = (inp[7]) ? node361 : node268;
							assign node268 = (inp[6]) ? node334 : node269;
								assign node269 = (inp[12]) ? node311 : node270;
									assign node270 = (inp[5]) ? node288 : node271;
										assign node271 = (inp[1]) ? node279 : node272;
											assign node272 = (inp[4]) ? 14'b00000000000001 : node273;
												assign node273 = (inp[10]) ? node275 : 14'b00011110110000;
													assign node275 = (inp[9]) ? 14'b00111110010010 : 14'b00111110110010;
											assign node279 = (inp[4]) ? node281 : 14'b00000000000001;
												assign node281 = (inp[10]) ? node285 : node282;
													assign node282 = (inp[2]) ? 14'b00111010010110 : 14'b01111010110110;
													assign node285 = (inp[2]) ? 14'b00000000000001 : 14'b01111010010000;
										assign node288 = (inp[1]) ? node300 : node289;
											assign node289 = (inp[9]) ? node295 : node290;
												assign node290 = (inp[4]) ? 14'b00110110110110 : node291;
													assign node291 = (inp[10]) ? 14'b01110110110010 : 14'b00110110110010;
												assign node295 = (inp[2]) ? 14'b00110110010000 : node296;
													assign node296 = (inp[4]) ? 14'b01110110010110 : 14'b00110110010010;
											assign node300 = (inp[2]) ? node308 : node301;
												assign node301 = (inp[10]) ? node305 : node302;
													assign node302 = (inp[9]) ? 14'b01110010010110 : 14'b01110010110110;
													assign node305 = (inp[9]) ? 14'b01110010010010 : 14'b01110010110000;
												assign node308 = (inp[4]) ? 14'b00110010010000 : 14'b00010010110000;
									assign node311 = (inp[4]) ? node323 : node312;
										assign node312 = (inp[10]) ? node318 : node313;
											assign node313 = (inp[1]) ? node315 : 14'b01011110110110;
												assign node315 = (inp[5]) ? 14'b01010010010110 : 14'b01011010010110;
											assign node318 = (inp[2]) ? node320 : 14'b00000000000001;
												assign node320 = (inp[5]) ? 14'b00010010110010 : 14'b00011010110010;
										assign node323 = (inp[2]) ? 14'b00000000000001 : node324;
											assign node324 = (inp[10]) ? node328 : node325;
												assign node325 = (inp[5]) ? 14'b01010010010010 : 14'b00000000000001;
												assign node328 = (inp[5]) ? 14'b00000000000001 : node329;
													assign node329 = (inp[9]) ? 14'b00111110010000 : 14'b00111110110000;
								assign node334 = (inp[1]) ? node336 : 14'b00000000000001;
									assign node336 = (inp[9]) ? 14'b00000000000001 : node337;
										assign node337 = (inp[12]) ? node349 : node338;
											assign node338 = (inp[10]) ? node346 : node339;
												assign node339 = (inp[5]) ? node343 : node340;
													assign node340 = (inp[2]) ? 14'b00011000100000 : 14'b00000000000001;
													assign node343 = (inp[2]) ? 14'b00010000100000 : 14'b00110000100010;
												assign node346 = (inp[2]) ? 14'b00111000100010 : 14'b01111000100010;
											assign node349 = (inp[4]) ? node353 : node350;
												assign node350 = (inp[2]) ? 14'b00011000100110 : 14'b00000000000001;
												assign node353 = (inp[2]) ? 14'b00000000000001 : node354;
													assign node354 = (inp[10]) ? 14'b00111000100000 : node355;
														assign node355 = (inp[5]) ? 14'b01010000100010 : 14'b00000000000001;
							assign node361 = (inp[9]) ? 14'b00000000000001 : node362;
								assign node362 = (inp[6]) ? node364 : 14'b00000000000001;
									assign node364 = (inp[10]) ? node378 : node365;
										assign node365 = (inp[12]) ? node373 : node366;
											assign node366 = (inp[4]) ? node370 : node367;
												assign node367 = (inp[1]) ? 14'b00000000100000 : 14'b00100100100010;
												assign node370 = (inp[1]) ? 14'b01100000100110 : 14'b00101100100110;
											assign node373 = (inp[4]) ? 14'b01000100100010 : node374;
												assign node374 = (inp[5]) ? 14'b01000100100110 : 14'b01001100100110;
										assign node378 = (inp[5]) ? node388 : node379;
											assign node379 = (inp[4]) ? node385 : node380;
												assign node380 = (inp[1]) ? 14'b00001000100010 : node381;
													assign node381 = (inp[12]) ? 14'b01001100100010 : 14'b00101100100010;
												assign node385 = (inp[1]) ? 14'b00101000100000 : 14'b00000000000001;
											assign node388 = (inp[4]) ? node390 : 14'b00000000000001;
												assign node390 = (inp[1]) ? 14'b00100000100000 : 14'b00100100100000;
					assign node394 = (inp[7]) ? 14'b00000000000001 : node395;
						assign node395 = (inp[9]) ? node493 : node396;
							assign node396 = (inp[1]) ? node464 : node397;
								assign node397 = (inp[2]) ? node437 : node398;
									assign node398 = (inp[3]) ? node416 : node399;
										assign node399 = (inp[5]) ? node409 : node400;
											assign node400 = (inp[10]) ? node402 : 14'b01111110100110;
												assign node402 = (inp[6]) ? node404 : 14'b01111110100000;
													assign node404 = (inp[12]) ? 14'b00111100100000 : node405;
														assign node405 = (inp[4]) ? 14'b01111100100000 : 14'b01111100100010;
											assign node409 = (inp[12]) ? 14'b01010100100110 : node410;
												assign node410 = (inp[6]) ? node412 : 14'b01110110100010;
													assign node412 = (inp[10]) ? 14'b01110100100000 : 14'b00110100100010;
										assign node416 = (inp[12]) ? node432 : node417;
											assign node417 = (inp[6]) ? node427 : node418;
												assign node418 = (inp[5]) ? node420 : 14'b01101110100000;
													assign node420 = (inp[10]) ? node424 : node421;
														assign node421 = (inp[4]) ? 14'b01100110100110 : 14'b00100110100010;
														assign node424 = (inp[4]) ? 14'b01100110100000 : 14'b01100110100010;
												assign node427 = (inp[4]) ? 14'b01101110000110 : node428;
													assign node428 = (inp[10]) ? 14'b01100110000010 : 14'b00100110000010;
											assign node432 = (inp[5]) ? 14'b00000000000001 : node433;
												assign node433 = (inp[6]) ? 14'b01001110000010 : 14'b01001110100010;
									assign node437 = (inp[4]) ? node453 : node438;
										assign node438 = (inp[12]) ? node444 : node439;
											assign node439 = (inp[10]) ? 14'b00000000000001 : node440;
												assign node440 = (inp[3]) ? 14'b00001110100000 : 14'b00010110100000;
											assign node444 = (inp[5]) ? node448 : node445;
												assign node445 = (inp[6]) ? 14'b00011100100110 : 14'b00011110100010;
												assign node448 = (inp[10]) ? node450 : 14'b00000110100110;
													assign node450 = (inp[3]) ? 14'b00000110100010 : 14'b00010110100010;
										assign node453 = (inp[12]) ? 14'b00000000000001 : node454;
											assign node454 = (inp[10]) ? node460 : node455;
												assign node455 = (inp[3]) ? 14'b00100110000110 : node456;
													assign node456 = (inp[6]) ? 14'b00110100100110 : 14'b00111110100110;
												assign node460 = (inp[3]) ? 14'b00100110000000 : 14'b00000000000001;
								assign node464 = (inp[6]) ? 14'b00000000000001 : node465;
									assign node465 = (inp[3]) ? node483 : node466;
										assign node466 = (inp[4]) ? node480 : node467;
											assign node467 = (inp[2]) ? node477 : node468;
												assign node468 = (inp[12]) ? node472 : node469;
													assign node469 = (inp[5]) ? 14'b01110010100010 : 14'b00000000000001;
													assign node472 = (inp[10]) ? 14'b00000000000001 : node473;
														assign node473 = (inp[5]) ? 14'b01010010100110 : 14'b01011010100110;
												assign node477 = (inp[5]) ? 14'b00010010100110 : 14'b00011010100010;
											assign node480 = (inp[2]) ? 14'b00110010100110 : 14'b01110010100110;
										assign node483 = (inp[12]) ? node487 : node484;
											assign node484 = (inp[4]) ? 14'b01101010100000 : 14'b00101010100010;
											assign node487 = (inp[5]) ? node489 : 14'b00000000000001;
												assign node489 = (inp[10]) ? 14'b00000000000001 : 14'b01000010100010;
							assign node493 = (inp[3]) ? node555 : node494;
								assign node494 = (inp[1]) ? node532 : node495;
									assign node495 = (inp[5]) ? node515 : node496;
										assign node496 = (inp[6]) ? node506 : node497;
											assign node497 = (inp[10]) ? node501 : node498;
												assign node498 = (inp[12]) ? 14'b01011110000110 : 14'b00111110000110;
												assign node501 = (inp[2]) ? 14'b00111110000010 : node502;
													assign node502 = (inp[12]) ? 14'b00111110000000 : 14'b01111110000000;
											assign node506 = (inp[4]) ? 14'b00000000000001 : node507;
												assign node507 = (inp[10]) ? node511 : node508;
													assign node508 = (inp[2]) ? 14'b00011100000110 : 14'b00000000000001;
													assign node511 = (inp[2]) ? 14'b00011100000010 : 14'b01111100000010;
										assign node515 = (inp[12]) ? node527 : node516;
											assign node516 = (inp[6]) ? node520 : node517;
												assign node517 = (inp[10]) ? 14'b00000000000001 : 14'b00110110000010;
												assign node520 = (inp[10]) ? node524 : node521;
													assign node521 = (inp[2]) ? 14'b00110100000110 : 14'b01110100000110;
													assign node524 = (inp[4]) ? 14'b00110100000000 : 14'b01110100000010;
											assign node527 = (inp[4]) ? 14'b00000000000001 : node528;
												assign node528 = (inp[2]) ? 14'b00010100000010 : 14'b00000000000001;
									assign node532 = (inp[6]) ? node534 : 14'b00000000000001;
										assign node534 = (inp[12]) ? node552 : node535;
											assign node535 = (inp[10]) ? node547 : node536;
												assign node536 = (inp[4]) ? node544 : node537;
													assign node537 = (inp[2]) ? node541 : node538;
														assign node538 = (inp[5]) ? 14'b00110000000010 : 14'b00000000000001;
														assign node541 = (inp[5]) ? 14'b00010000000000 : 14'b00011000000000;
													assign node544 = (inp[5]) ? 14'b01110000000110 : 14'b00111000000110;
												assign node547 = (inp[5]) ? node549 : 14'b00000000000001;
													assign node549 = (inp[4]) ? 14'b00110000000000 : 14'b00000000000001;
											assign node552 = (inp[4]) ? 14'b00000000000001 : 14'b01011000000110;
								assign node555 = (inp[1]) ? node557 : 14'b00000000000001;
									assign node557 = (inp[6]) ? 14'b00000000000001 : node558;
										assign node558 = (inp[12]) ? node568 : node559;
											assign node559 = (inp[2]) ? node563 : node560;
												assign node560 = (inp[10]) ? 14'b01100010000000 : 14'b01100010000110;
												assign node563 = (inp[10]) ? 14'b00101010000010 : node564;
													assign node564 = (inp[5]) ? 14'b00100010000110 : 14'b00101010000110;
											assign node568 = (inp[4]) ? 14'b00000000000001 : node569;
												assign node569 = (inp[10]) ? node575 : node570;
													assign node570 = (inp[2]) ? 14'b00000010000110 : node571;
														assign node571 = (inp[5]) ? 14'b01000010000110 : 14'b01001010000110;
													assign node575 = (inp[5]) ? 14'b00000000000001 : 14'b00001010000010;
				assign node581 = (inp[10]) ? 14'b00000000000001 : node582;
					assign node582 = (inp[4]) ? node788 : node583;
						assign node583 = (inp[7]) ? node737 : node584;
							assign node584 = (inp[12]) ? node664 : node585;
								assign node585 = (inp[3]) ? node633 : node586;
									assign node586 = (inp[1]) ? node618 : node587;
										assign node587 = (inp[2]) ? node601 : node588;
											assign node588 = (inp[5]) ? node596 : node589;
												assign node589 = (inp[0]) ? node593 : node590;
													assign node590 = (inp[6]) ? 14'b01111100010100 : 14'b01101100000100;
													assign node593 = (inp[6]) ? 14'b01111100000100 : 14'b01111110000100;
												assign node596 = (inp[9]) ? node598 : 14'b01110100110100;
													assign node598 = (inp[6]) ? 14'b01110100000100 : 14'b01110110000100;
											assign node601 = (inp[6]) ? node609 : node602;
												assign node602 = (inp[0]) ? node606 : node603;
													assign node603 = (inp[5]) ? 14'b00100100000100 : 14'b00000000000001;
													assign node606 = (inp[9]) ? 14'b00110110000100 : 14'b00111110100100;
												assign node609 = (inp[9]) ? node613 : node610;
													assign node610 = (inp[0]) ? 14'b00110100100100 : 14'b00110100110100;
													assign node613 = (inp[5]) ? 14'b00110100010100 : node614;
														assign node614 = (inp[0]) ? 14'b00111100000100 : 14'b00111100010100;
										assign node618 = (inp[0]) ? node624 : node619;
											assign node619 = (inp[6]) ? 14'b01110000110100 : node620;
												assign node620 = (inp[2]) ? 14'b00101000000100 : 14'b01101000000100;
											assign node624 = (inp[6]) ? node630 : node625;
												assign node625 = (inp[5]) ? 14'b00000000000001 : node626;
													assign node626 = (inp[2]) ? 14'b00111010100100 : 14'b01111010100100;
												assign node630 = (inp[5]) ? 14'b00110000000100 : 14'b00000000000001;
									assign node633 = (inp[9]) ? node655 : node634;
										assign node634 = (inp[5]) ? node646 : node635;
											assign node635 = (inp[6]) ? node639 : node636;
												assign node636 = (inp[1]) ? 14'b01101010100100 : 14'b01111110110100;
												assign node639 = (inp[1]) ? 14'b00000000000001 : node640;
													assign node640 = (inp[0]) ? node642 : 14'b00000000000001;
														assign node642 = (inp[2]) ? 14'b00101110000100 : 14'b01101110000100;
											assign node646 = (inp[6]) ? node652 : node647;
												assign node647 = (inp[0]) ? 14'b00100010100100 : node648;
													assign node648 = (inp[2]) ? 14'b00110110110100 : 14'b01110010110100;
												assign node652 = (inp[2]) ? 14'b00110000100100 : 14'b01110000100100;
										assign node655 = (inp[6]) ? 14'b00000000000001 : node656;
											assign node656 = (inp[1]) ? node658 : 14'b00000000000001;
												assign node658 = (inp[0]) ? 14'b00101010000100 : node659;
													assign node659 = (inp[5]) ? 14'b01110010010100 : 14'b01111010010100;
								assign node664 = (inp[5]) ? node704 : node665;
									assign node665 = (inp[3]) ? node685 : node666;
										assign node666 = (inp[9]) ? node670 : node667;
											assign node667 = (inp[1]) ? 14'b01011010000100 : 14'b00000000000001;
											assign node670 = (inp[1]) ? node682 : node671;
												assign node671 = (inp[2]) ? node677 : node672;
													assign node672 = (inp[6]) ? node674 : 14'b01011110000100;
														assign node674 = (inp[0]) ? 14'b01011100000100 : 14'b01011100010100;
													assign node677 = (inp[0]) ? node679 : 14'b00001100000100;
														assign node679 = (inp[6]) ? 14'b00011100000100 : 14'b00011110000100;
												assign node682 = (inp[2]) ? 14'b00011000000100 : 14'b00000000000001;
										assign node685 = (inp[6]) ? node695 : node686;
											assign node686 = (inp[0]) ? node690 : node687;
												assign node687 = (inp[1]) ? 14'b00011010110100 : 14'b01011110110100;
												assign node690 = (inp[1]) ? node692 : 14'b00001110100100;
													assign node692 = (inp[2]) ? 14'b00001010100100 : 14'b01001010100100;
											assign node695 = (inp[9]) ? 14'b00000000000001 : node696;
												assign node696 = (inp[2]) ? 14'b00000000000001 : node697;
													assign node697 = (inp[1]) ? 14'b01011000100100 : node698;
														assign node698 = (inp[0]) ? 14'b01001110000100 : 14'b00000000000001;
									assign node704 = (inp[1]) ? node720 : node705;
										assign node705 = (inp[9]) ? node711 : node706;
											assign node706 = (inp[0]) ? node708 : 14'b00000000000001;
												assign node708 = (inp[2]) ? 14'b00000110000100 : 14'b01000110000100;
											assign node711 = (inp[0]) ? node715 : node712;
												assign node712 = (inp[2]) ? 14'b00010110010100 : 14'b01010110010100;
												assign node715 = (inp[3]) ? 14'b00000000000001 : node716;
													assign node716 = (inp[6]) ? 14'b01010100000100 : 14'b01010110000100;
										assign node720 = (inp[6]) ? node728 : node721;
											assign node721 = (inp[0]) ? 14'b00000000000001 : node722;
												assign node722 = (inp[3]) ? node724 : 14'b00010010000100;
													assign node724 = (inp[2]) ? 14'b00010010110100 : 14'b01010010010100;
											assign node728 = (inp[3]) ? 14'b00000000000001 : node729;
												assign node729 = (inp[0]) ? node731 : 14'b00010000110100;
													assign node731 = (inp[9]) ? node733 : 14'b00000000000001;
														assign node733 = (inp[2]) ? 14'b00010000000100 : 14'b01010000000100;
							assign node737 = (inp[0]) ? 14'b00000000000001 : node738;
								assign node738 = (inp[3]) ? node776 : node739;
									assign node739 = (inp[6]) ? node757 : node740;
										assign node740 = (inp[12]) ? node750 : node741;
											assign node741 = (inp[1]) ? 14'b00101010110100 : node742;
												assign node742 = (inp[5]) ? 14'b01100110010100 : node743;
													assign node743 = (inp[2]) ? 14'b00101110010100 : node744;
														assign node744 = (inp[9]) ? 14'b01101110010100 : 14'b01101110110100;
											assign node750 = (inp[5]) ? 14'b01000110110100 : node751;
												assign node751 = (inp[9]) ? node753 : 14'b01001010110100;
													assign node753 = (inp[1]) ? 14'b01001010010100 : 14'b01001110010100;
										assign node757 = (inp[9]) ? node767 : node758;
											assign node758 = (inp[12]) ? node762 : node759;
												assign node759 = (inp[2]) ? 14'b00101000110100 : 14'b01101100110100;
												assign node762 = (inp[5]) ? node764 : 14'b00001100110100;
													assign node764 = (inp[1]) ? 14'b00000000110100 : 14'b00000100110100;
											assign node767 = (inp[1]) ? node771 : node768;
												assign node768 = (inp[12]) ? 14'b00000100010100 : 14'b00100100010100;
												assign node771 = (inp[5]) ? 14'b01100000010100 : node772;
													assign node772 = (inp[2]) ? 14'b00001000010100 : 14'b01001000010100;
									assign node776 = (inp[9]) ? 14'b00000000000001 : node777;
										assign node777 = (inp[6]) ? node779 : 14'b00000000000001;
											assign node779 = (inp[1]) ? node783 : node780;
												assign node780 = (inp[2]) ? 14'b00001100100100 : 14'b01000100100100;
												assign node783 = (inp[2]) ? 14'b00000000100100 : 14'b01100000100100;
						assign node788 = (inp[2]) ? node860 : node789;
							assign node789 = (inp[12]) ? node803 : node790;
								assign node790 = (inp[9]) ? 14'b00000000000001 : node791;
									assign node791 = (inp[3]) ? node793 : 14'b00000000000001;
										assign node793 = (inp[1]) ? 14'b00000000000001 : node794;
											assign node794 = (inp[5]) ? 14'b00000000000001 : node795;
												assign node795 = (inp[0]) ? 14'b00000000000001 : node796;
													assign node796 = (inp[6]) ? 14'b10000001001000 : 14'b10000001000000;
								assign node803 = (inp[9]) ? node841 : node804;
									assign node804 = (inp[5]) ? node818 : node805;
										assign node805 = (inp[7]) ? node815 : node806;
											assign node806 = (inp[1]) ? node810 : node807;
												assign node807 = (inp[0]) ? 14'b01011110100000 : 14'b01011110110000;
												assign node810 = (inp[6]) ? 14'b01011000110000 : node811;
													assign node811 = (inp[0]) ? 14'b01011010100000 : 14'b01011010110000;
											assign node815 = (inp[1]) ? 14'b01001000100000 : 14'b01001100100000;
										assign node818 = (inp[3]) ? node830 : node819;
											assign node819 = (inp[1]) ? node821 : 14'b00000000000001;
												assign node821 = (inp[6]) ? node827 : node822;
													assign node822 = (inp[7]) ? 14'b01000010110000 : node823;
														assign node823 = (inp[0]) ? 14'b01010010100000 : 14'b01010010000000;
													assign node827 = (inp[0]) ? 14'b00000000000001 : 14'b01010000110000;
											assign node830 = (inp[7]) ? node838 : node831;
												assign node831 = (inp[0]) ? node833 : 14'b01010010110000;
													assign node833 = (inp[1]) ? 14'b01000010100000 : node834;
														assign node834 = (inp[6]) ? 14'b01000110000000 : 14'b01000110100000;
												assign node838 = (inp[6]) ? 14'b01000100100000 : 14'b00000000000001;
									assign node841 = (inp[3]) ? node853 : node842;
										assign node842 = (inp[0]) ? node848 : node843;
											assign node843 = (inp[7]) ? 14'b01000010010000 : node844;
												assign node844 = (inp[5]) ? 14'b01010000010000 : 14'b01011000010000;
											assign node848 = (inp[1]) ? node850 : 14'b00000000000001;
												assign node850 = (inp[6]) ? 14'b01010000000000 : 14'b00000000000001;
										assign node853 = (inp[6]) ? 14'b00000000000001 : node854;
											assign node854 = (inp[1]) ? node856 : 14'b00000000000001;
												assign node856 = (inp[7]) ? 14'b00000000000001 : 14'b01001010000000;
							assign node860 = (inp[5]) ? 14'b00000000000001 : node861;
								assign node861 = (inp[0]) ? node863 : 14'b00000000000001;
									assign node863 = (inp[9]) ? 14'b00000000000001 : node864;
										assign node864 = (inp[7]) ? 14'b00000000000001 : node865;
											assign node865 = (inp[1]) ? node867 : 14'b00000000000001;
												assign node867 = (inp[6]) ? node869 : 14'b00000000000001;
													assign node869 = (inp[3]) ? 14'b00000000000001 : 14'b10000000000000;
		assign node876 = (inp[5]) ? node1804 : node877;
			assign node877 = (inp[0]) ? node1521 : node878;
				assign node878 = (inp[6]) ? node1310 : node879;
					assign node879 = (inp[7]) ? node1129 : node880;
						assign node880 = (inp[1]) ? node1006 : node881;
							assign node881 = (inp[3]) ? node925 : node882;
								assign node882 = (inp[9]) ? node894 : node883;
									assign node883 = (inp[2]) ? 14'b00000000000001 : node884;
										assign node884 = (inp[12]) ? 14'b00000000000001 : node885;
											assign node885 = (inp[4]) ? 14'b00000000000001 : node886;
												assign node886 = (inp[10]) ? node888 : 14'b10000000001000;
													assign node888 = (inp[8]) ? 14'b10000000001000 : 14'b00000000000001;
									assign node894 = (inp[4]) ? node908 : node895;
										assign node895 = (inp[8]) ? node905 : node896;
											assign node896 = (inp[12]) ? node902 : node897;
												assign node897 = (inp[2]) ? node899 : 14'b00000000000001;
													assign node899 = (inp[10]) ? 14'b00000000000001 : 14'b01100100000110;
												assign node902 = (inp[10]) ? 14'b01100100000000 : 14'b01100100000100;
											assign node905 = (inp[11]) ? 14'b01100100000100 : 14'b01000100000100;
										assign node908 = (inp[2]) ? node916 : node909;
											assign node909 = (inp[8]) ? node913 : node910;
												assign node910 = (inp[10]) ? 14'b00100100000000 : 14'b00100100000100;
												assign node913 = (inp[12]) ? 14'b00000100000100 : 14'b00100100000100;
											assign node916 = (inp[8]) ? 14'b00000000000001 : node917;
												assign node917 = (inp[12]) ? node921 : node918;
													assign node918 = (inp[10]) ? 14'b00000100000010 : 14'b00000000000001;
													assign node921 = (inp[10]) ? 14'b00000100000000 : 14'b00000100000100;
								assign node925 = (inp[9]) ? node957 : node926;
									assign node926 = (inp[12]) ? node942 : node927;
										assign node927 = (inp[8]) ? node935 : node928;
											assign node928 = (inp[10]) ? node932 : node929;
												assign node929 = (inp[4]) ? 14'b00110110110110 : 14'b00000000000001;
												assign node932 = (inp[2]) ? 14'b00010110110010 : 14'b01110110110010;
											assign node935 = (inp[4]) ? node939 : node936;
												assign node936 = (inp[2]) ? 14'b01110110110100 : 14'b00000000000001;
												assign node939 = (inp[2]) ? 14'b00000000000001 : 14'b00110110110100;
										assign node942 = (inp[4]) ? node952 : node943;
											assign node943 = (inp[8]) ? node949 : node944;
												assign node944 = (inp[10]) ? 14'b01110110110000 : node945;
													assign node945 = (inp[2]) ? 14'b01110110110100 : 14'b01010010110100;
												assign node949 = (inp[2]) ? 14'b01010110110000 : 14'b01010110110100;
											assign node952 = (inp[8]) ? 14'b00010110110100 : node953;
												assign node953 = (inp[2]) ? 14'b00010110110100 : 14'b00110110110100;
									assign node957 = (inp[10]) ? node979 : node958;
										assign node958 = (inp[12]) ? node970 : node959;
											assign node959 = (inp[2]) ? node965 : node960;
												assign node960 = (inp[4]) ? node962 : 14'b00000000000001;
													assign node962 = (inp[8]) ? 14'b00110110010100 : 14'b00110110010110;
												assign node965 = (inp[4]) ? 14'b00000000000001 : node966;
													assign node966 = (inp[8]) ? 14'b01110110010100 : 14'b01110110010110;
											assign node970 = (inp[4]) ? node974 : node971;
												assign node971 = (inp[2]) ? 14'b01010110010000 : 14'b01010010010100;
												assign node974 = (inp[2]) ? node976 : 14'b00010110010100;
													assign node976 = (inp[8]) ? 14'b00000000000001 : 14'b00010110010100;
										assign node979 = (inp[2]) ? node991 : node980;
											assign node980 = (inp[8]) ? node986 : node981;
												assign node981 = (inp[12]) ? 14'b01110110010000 : node982;
													assign node982 = (inp[11]) ? 14'b01110110010010 : 14'b00110110010010;
												assign node986 = (inp[12]) ? node988 : 14'b00110110010100;
													assign node988 = (inp[4]) ? 14'b00010110010100 : 14'b01010110010100;
											assign node991 = (inp[11]) ? node997 : node992;
												assign node992 = (inp[12]) ? node994 : 14'b00010110010010;
													assign node994 = (inp[4]) ? 14'b00010110010000 : 14'b01010110010000;
												assign node997 = (inp[4]) ? node1001 : node998;
													assign node998 = (inp[8]) ? 14'b01010110010000 : 14'b00000000000001;
													assign node1001 = (inp[8]) ? 14'b00000000000001 : node1002;
														assign node1002 = (inp[12]) ? 14'b00010110010000 : 14'b00010110010010;
							assign node1006 = (inp[3]) ? node1064 : node1007;
								assign node1007 = (inp[4]) ? node1037 : node1008;
									assign node1008 = (inp[9]) ? node1024 : node1009;
										assign node1009 = (inp[12]) ? node1019 : node1010;
											assign node1010 = (inp[11]) ? 14'b01110110100110 : node1011;
												assign node1011 = (inp[10]) ? node1013 : 14'b00000000000001;
													assign node1013 = (inp[8]) ? 14'b01110110100100 : node1014;
														assign node1014 = (inp[2]) ? 14'b00000000000001 : 14'b01110110100010;
											assign node1019 = (inp[10]) ? 14'b00000000000001 : node1020;
												assign node1020 = (inp[2]) ? 14'b01110110100100 : 14'b01010110100100;
										assign node1024 = (inp[2]) ? node1030 : node1025;
											assign node1025 = (inp[12]) ? node1027 : 14'b00000000000001;
												assign node1027 = (inp[10]) ? 14'b01110110000000 : 14'b01010010000100;
											assign node1030 = (inp[12]) ? node1034 : node1031;
												assign node1031 = (inp[8]) ? 14'b01110110000100 : 14'b01110110000110;
												assign node1034 = (inp[11]) ? 14'b01010110000000 : 14'b01110110000100;
									assign node1037 = (inp[2]) ? node1055 : node1038;
										assign node1038 = (inp[9]) ? node1046 : node1039;
											assign node1039 = (inp[8]) ? node1043 : node1040;
												assign node1040 = (inp[10]) ? 14'b00110110100000 : 14'b00110110100110;
												assign node1043 = (inp[12]) ? 14'b00010110100100 : 14'b00110110100100;
											assign node1046 = (inp[8]) ? node1052 : node1047;
												assign node1047 = (inp[10]) ? node1049 : 14'b00110110000110;
													assign node1049 = (inp[11]) ? 14'b00110110000010 : 14'b00110110000000;
												assign node1052 = (inp[12]) ? 14'b00010110000100 : 14'b00110110000100;
										assign node1055 = (inp[8]) ? 14'b00000000000001 : node1056;
											assign node1056 = (inp[12]) ? node1058 : 14'b00000000000001;
												assign node1058 = (inp[10]) ? node1060 : 14'b00010110000100;
													assign node1060 = (inp[9]) ? 14'b00010110000000 : 14'b00010110100000;
								assign node1064 = (inp[4]) ? node1100 : node1065;
									assign node1065 = (inp[12]) ? node1085 : node1066;
										assign node1066 = (inp[2]) ? node1074 : node1067;
											assign node1067 = (inp[8]) ? 14'b00000000000001 : node1068;
												assign node1068 = (inp[10]) ? node1070 : 14'b00000000000001;
													assign node1070 = (inp[11]) ? 14'b01100110100010 : 14'b01100110000010;
											assign node1074 = (inp[10]) ? node1080 : node1075;
												assign node1075 = (inp[8]) ? 14'b01100110100100 : node1076;
													assign node1076 = (inp[11]) ? 14'b01100110000110 : 14'b01100110100110;
												assign node1080 = (inp[8]) ? node1082 : 14'b00000000000001;
													assign node1082 = (inp[11]) ? 14'b01100110100100 : 14'b01100110000100;
										assign node1085 = (inp[9]) ? node1093 : node1086;
											assign node1086 = (inp[10]) ? node1090 : node1087;
												assign node1087 = (inp[8]) ? 14'b01000110100000 : 14'b01000010100100;
												assign node1090 = (inp[2]) ? 14'b00000000000001 : 14'b01100110100000;
											assign node1093 = (inp[8]) ? node1097 : node1094;
												assign node1094 = (inp[10]) ? 14'b01100110000000 : 14'b01100110000100;
												assign node1097 = (inp[11]) ? 14'b01000110000000 : 14'b01000110000100;
									assign node1100 = (inp[2]) ? node1120 : node1101;
										assign node1101 = (inp[9]) ? node1109 : node1102;
											assign node1102 = (inp[12]) ? node1106 : node1103;
												assign node1103 = (inp[8]) ? 14'b00100110100100 : 14'b00100110100110;
												assign node1106 = (inp[10]) ? 14'b00100110100000 : 14'b00100110100100;
											assign node1109 = (inp[8]) ? node1117 : node1110;
												assign node1110 = (inp[10]) ? node1114 : node1111;
													assign node1111 = (inp[12]) ? 14'b00100110000100 : 14'b00100110000110;
													assign node1114 = (inp[12]) ? 14'b00100110000000 : 14'b00100110000010;
												assign node1117 = (inp[12]) ? 14'b00000110000100 : 14'b00100110000100;
										assign node1120 = (inp[8]) ? 14'b00000000000001 : node1121;
											assign node1121 = (inp[10]) ? node1123 : 14'b00000000000001;
												assign node1123 = (inp[12]) ? node1125 : 14'b00000110000010;
													assign node1125 = (inp[9]) ? 14'b00000110000000 : 14'b00000110100000;
						assign node1129 = (inp[2]) ? node1261 : node1130;
							assign node1130 = (inp[9]) ? node1184 : node1131;
								assign node1131 = (inp[3]) ? node1149 : node1132;
									assign node1132 = (inp[1]) ? node1134 : 14'b00000000000001;
										assign node1134 = (inp[8]) ? node1142 : node1135;
											assign node1135 = (inp[12]) ? 14'b00110010100100 : node1136;
												assign node1136 = (inp[10]) ? node1138 : 14'b00010010100010;
													assign node1138 = (inp[4]) ? 14'b00110010100010 : 14'b01110010100010;
											assign node1142 = (inp[12]) ? node1146 : node1143;
												assign node1143 = (inp[4]) ? 14'b00110010100100 : 14'b00010010100000;
												assign node1146 = (inp[4]) ? 14'b00010010100100 : 14'b01010010100100;
									assign node1149 = (inp[1]) ? node1169 : node1150;
										assign node1150 = (inp[8]) ? node1164 : node1151;
											assign node1151 = (inp[12]) ? node1157 : node1152;
												assign node1152 = (inp[10]) ? node1154 : 14'b00010010110010;
													assign node1154 = (inp[4]) ? 14'b00110010110010 : 14'b01110010110010;
												assign node1157 = (inp[11]) ? 14'b01110010110000 : node1158;
													assign node1158 = (inp[4]) ? node1160 : 14'b00010010110000;
														assign node1160 = (inp[10]) ? 14'b00110010110000 : 14'b00110010110100;
											assign node1164 = (inp[12]) ? node1166 : 14'b00110010110100;
												assign node1166 = (inp[4]) ? 14'b00010010110100 : 14'b01010010110100;
										assign node1169 = (inp[4]) ? node1179 : node1170;
											assign node1170 = (inp[12]) ? node1174 : node1171;
												assign node1171 = (inp[8]) ? 14'b00000010100000 : 14'b00000010100010;
												assign node1174 = (inp[11]) ? node1176 : 14'b01100010100000;
													assign node1176 = (inp[8]) ? 14'b01000010100100 : 14'b00000010100000;
											assign node1179 = (inp[11]) ? 14'b00100010100100 : node1180;
												assign node1180 = (inp[12]) ? 14'b00000010100100 : 14'b00100010100110;
								assign node1184 = (inp[8]) ? node1234 : node1185;
									assign node1185 = (inp[12]) ? node1209 : node1186;
										assign node1186 = (inp[3]) ? node1200 : node1187;
											assign node1187 = (inp[1]) ? node1195 : node1188;
												assign node1188 = (inp[4]) ? node1192 : node1189;
													assign node1189 = (inp[10]) ? 14'b01100000000010 : 14'b00000000000010;
													assign node1192 = (inp[10]) ? 14'b00100000000010 : 14'b00100000000110;
												assign node1195 = (inp[10]) ? 14'b01110010000010 : node1196;
													assign node1196 = (inp[4]) ? 14'b00110010000110 : 14'b00010010000010;
											assign node1200 = (inp[1]) ? node1206 : node1201;
												assign node1201 = (inp[10]) ? node1203 : 14'b00010010010010;
													assign node1203 = (inp[4]) ? 14'b00110010010010 : 14'b01110010010010;
												assign node1206 = (inp[10]) ? 14'b01100010000010 : 14'b00000010000010;
										assign node1209 = (inp[10]) ? node1221 : node1210;
											assign node1210 = (inp[4]) ? node1216 : node1211;
												assign node1211 = (inp[1]) ? node1213 : 14'b00000000000000;
													assign node1213 = (inp[3]) ? 14'b00000010000000 : 14'b00010010000000;
												assign node1216 = (inp[1]) ? node1218 : 14'b00100000000100;
													assign node1218 = (inp[3]) ? 14'b00100010000100 : 14'b00110010000100;
											assign node1221 = (inp[4]) ? node1229 : node1222;
												assign node1222 = (inp[1]) ? node1226 : node1223;
													assign node1223 = (inp[3]) ? 14'b01110010010000 : 14'b01100000000000;
													assign node1226 = (inp[3]) ? 14'b01100010000000 : 14'b01110010000000;
												assign node1229 = (inp[1]) ? node1231 : 14'b00100000000000;
													assign node1231 = (inp[3]) ? 14'b00100010000000 : 14'b00110010000000;
									assign node1234 = (inp[12]) ? node1248 : node1235;
										assign node1235 = (inp[4]) ? node1243 : node1236;
											assign node1236 = (inp[1]) ? node1240 : node1237;
												assign node1237 = (inp[3]) ? 14'b00010010010000 : 14'b00000000000000;
												assign node1240 = (inp[3]) ? 14'b00000010000000 : 14'b00010010000000;
											assign node1243 = (inp[3]) ? node1245 : 14'b00100000000100;
												assign node1245 = (inp[1]) ? 14'b00100010000100 : 14'b00110010010100;
										assign node1248 = (inp[4]) ? node1254 : node1249;
											assign node1249 = (inp[1]) ? node1251 : 14'b01010010010100;
												assign node1251 = (inp[3]) ? 14'b01000010000100 : 14'b01010010000100;
											assign node1254 = (inp[1]) ? node1258 : node1255;
												assign node1255 = (inp[3]) ? 14'b00010010010100 : 14'b00000000000100;
												assign node1258 = (inp[3]) ? 14'b00000010000100 : 14'b00010010000100;
							assign node1261 = (inp[4]) ? 14'b00000000000001 : node1262;
								assign node1262 = (inp[10]) ? node1286 : node1263;
									assign node1263 = (inp[1]) ? node1273 : node1264;
										assign node1264 = (inp[3]) ? node1268 : node1265;
											assign node1265 = (inp[9]) ? 14'b01000000000000 : 14'b00000000000001;
											assign node1268 = (inp[12]) ? 14'b01110010010100 : node1269;
												assign node1269 = (inp[8]) ? 14'b01110010010100 : 14'b01110010010110;
										assign node1273 = (inp[9]) ? node1281 : node1274;
											assign node1274 = (inp[3]) ? node1276 : 14'b01110010100100;
												assign node1276 = (inp[12]) ? 14'b01000010100000 : node1277;
													assign node1277 = (inp[8]) ? 14'b01100010100100 : 14'b01100010100110;
											assign node1281 = (inp[12]) ? 14'b01100010000100 : node1282;
												assign node1282 = (inp[8]) ? 14'b01110010000100 : 14'b01110010000110;
									assign node1286 = (inp[8]) ? node1288 : 14'b00000000000001;
										assign node1288 = (inp[12]) ? node1300 : node1289;
											assign node1289 = (inp[1]) ? node1295 : node1290;
												assign node1290 = (inp[3]) ? 14'b01110010110100 : node1291;
													assign node1291 = (inp[9]) ? 14'b01100000000100 : 14'b00000000000001;
												assign node1295 = (inp[3]) ? node1297 : 14'b01110010100100;
													assign node1297 = (inp[9]) ? 14'b01100010000100 : 14'b01100010100100;
											assign node1300 = (inp[1]) ? node1304 : node1301;
												assign node1301 = (inp[3]) ? 14'b01010010010000 : 14'b00000000000001;
												assign node1304 = (inp[9]) ? node1306 : 14'b01000010100000;
													assign node1306 = (inp[11]) ? 14'b01000010000000 : 14'b01010010000000;
					assign node1310 = (inp[3]) ? node1502 : node1311;
						assign node1311 = (inp[2]) ? node1433 : node1312;
							assign node1312 = (inp[4]) ? node1366 : node1313;
								assign node1313 = (inp[12]) ? node1339 : node1314;
									assign node1314 = (inp[7]) ? node1322 : node1315;
										assign node1315 = (inp[8]) ? 14'b00000000000001 : node1316;
											assign node1316 = (inp[10]) ? node1318 : 14'b00000000000001;
												assign node1318 = (inp[11]) ? 14'b01110100110010 : 14'b01110100000010;
										assign node1322 = (inp[8]) ? node1332 : node1323;
											assign node1323 = (inp[10]) ? node1327 : node1324;
												assign node1324 = (inp[9]) ? 14'b00010000010010 : 14'b00010000110010;
												assign node1327 = (inp[1]) ? node1329 : 14'b01110000110010;
													assign node1329 = (inp[9]) ? 14'b01110000000010 : 14'b01110000100010;
											assign node1332 = (inp[9]) ? node1336 : node1333;
												assign node1333 = (inp[1]) ? 14'b00010000100000 : 14'b00010000110000;
												assign node1336 = (inp[10]) ? 14'b00010000010000 : 14'b00010000000000;
									assign node1339 = (inp[9]) ? node1355 : node1340;
										assign node1340 = (inp[1]) ? node1344 : node1341;
											assign node1341 = (inp[8]) ? 14'b01010100110100 : 14'b01110100110000;
											assign node1344 = (inp[7]) ? node1352 : node1345;
												assign node1345 = (inp[10]) ? node1349 : node1346;
													assign node1346 = (inp[8]) ? 14'b01010100100100 : 14'b01010000100100;
													assign node1349 = (inp[11]) ? 14'b01110100100000 : 14'b01010100100100;
												assign node1352 = (inp[11]) ? 14'b01110000100000 : 14'b00010000100000;
										assign node1355 = (inp[1]) ? node1359 : node1356;
											assign node1356 = (inp[8]) ? 14'b01010100010100 : 14'b01010000010100;
											assign node1359 = (inp[8]) ? node1363 : node1360;
												assign node1360 = (inp[7]) ? 14'b01110000000000 : 14'b01010000000100;
												assign node1363 = (inp[7]) ? 14'b01010000000100 : 14'b01010100000100;
								assign node1366 = (inp[9]) ? node1398 : node1367;
									assign node1367 = (inp[7]) ? node1387 : node1368;
										assign node1368 = (inp[1]) ? node1376 : node1369;
											assign node1369 = (inp[8]) ? node1373 : node1370;
												assign node1370 = (inp[10]) ? 14'b00110100110010 : 14'b00110100110110;
												assign node1373 = (inp[12]) ? 14'b00010100110100 : 14'b00110100110100;
											assign node1376 = (inp[8]) ? node1384 : node1377;
												assign node1377 = (inp[12]) ? node1381 : node1378;
													assign node1378 = (inp[11]) ? 14'b00110100100110 : 14'b00110100100010;
													assign node1381 = (inp[10]) ? 14'b00110100100000 : 14'b00110100100100;
												assign node1384 = (inp[12]) ? 14'b00010100100100 : 14'b00110100100100;
										assign node1387 = (inp[8]) ? node1393 : node1388;
											assign node1388 = (inp[10]) ? 14'b00110000100010 : node1389;
												assign node1389 = (inp[1]) ? 14'b00110000100110 : 14'b00110000110110;
											assign node1393 = (inp[12]) ? 14'b00010000100100 : node1394;
												assign node1394 = (inp[1]) ? 14'b00110000100100 : 14'b00110000110100;
									assign node1398 = (inp[7]) ? node1416 : node1399;
										assign node1399 = (inp[1]) ? node1407 : node1400;
											assign node1400 = (inp[12]) ? node1404 : node1401;
												assign node1401 = (inp[8]) ? 14'b00110100010100 : 14'b00110100010010;
												assign node1404 = (inp[8]) ? 14'b00010100010100 : 14'b00110100010100;
											assign node1407 = (inp[8]) ? node1413 : node1408;
												assign node1408 = (inp[11]) ? 14'b00110100000000 : node1409;
													assign node1409 = (inp[10]) ? 14'b00110100000010 : 14'b00110100000110;
												assign node1413 = (inp[12]) ? 14'b00010100000100 : 14'b00110100000100;
										assign node1416 = (inp[1]) ? node1424 : node1417;
											assign node1417 = (inp[8]) ? node1421 : node1418;
												assign node1418 = (inp[12]) ? 14'b00110000010000 : 14'b00110000010010;
												assign node1421 = (inp[12]) ? 14'b00010000010100 : 14'b00110000010100;
											assign node1424 = (inp[11]) ? node1428 : node1425;
												assign node1425 = (inp[8]) ? 14'b00110000000100 : 14'b00110000000000;
												assign node1428 = (inp[12]) ? node1430 : 14'b00110000000100;
													assign node1430 = (inp[8]) ? 14'b00010000000100 : 14'b00110000000100;
							assign node1433 = (inp[4]) ? node1483 : node1434;
								assign node1434 = (inp[8]) ? node1456 : node1435;
									assign node1435 = (inp[10]) ? 14'b00000000000001 : node1436;
										assign node1436 = (inp[12]) ? node1444 : node1437;
											assign node1437 = (inp[1]) ? node1441 : node1438;
												assign node1438 = (inp[9]) ? 14'b01110000010110 : 14'b01110000110110;
												assign node1441 = (inp[9]) ? 14'b01110000000110 : 14'b01110000100110;
											assign node1444 = (inp[9]) ? node1450 : node1445;
												assign node1445 = (inp[1]) ? 14'b01110000100100 : node1446;
													assign node1446 = (inp[7]) ? 14'b01110000110100 : 14'b01110100110100;
												assign node1450 = (inp[7]) ? node1452 : 14'b01110100000100;
													assign node1452 = (inp[11]) ? 14'b01110000000100 : 14'b01110000010100;
									assign node1456 = (inp[12]) ? node1470 : node1457;
										assign node1457 = (inp[9]) ? node1465 : node1458;
											assign node1458 = (inp[1]) ? node1462 : node1459;
												assign node1459 = (inp[7]) ? 14'b01110000110100 : 14'b01110100110100;
												assign node1462 = (inp[7]) ? 14'b01110000100100 : 14'b01110100100100;
											assign node1465 = (inp[1]) ? node1467 : 14'b01110100010100;
												assign node1467 = (inp[7]) ? 14'b01110000000100 : 14'b01110100000100;
										assign node1470 = (inp[9]) ? node1476 : node1471;
											assign node1471 = (inp[7]) ? node1473 : 14'b01010100110000;
												assign node1473 = (inp[11]) ? 14'b01010000100000 : 14'b01010000110000;
											assign node1476 = (inp[1]) ? node1480 : node1477;
												assign node1477 = (inp[7]) ? 14'b01010000010000 : 14'b01010100010000;
												assign node1480 = (inp[7]) ? 14'b01010000000000 : 14'b01010100000000;
								assign node1483 = (inp[7]) ? 14'b00000000000001 : node1484;
									assign node1484 = (inp[8]) ? 14'b00000000000001 : node1485;
										assign node1485 = (inp[10]) ? node1491 : node1486;
											assign node1486 = (inp[12]) ? node1488 : 14'b00000000000001;
												assign node1488 = (inp[9]) ? 14'b00010100010100 : 14'b00010100100100;
											assign node1491 = (inp[12]) ? node1495 : node1492;
												assign node1492 = (inp[1]) ? 14'b00010100100010 : 14'b00010100110010;
												assign node1495 = (inp[9]) ? node1497 : 14'b00010100110000;
													assign node1497 = (inp[1]) ? 14'b00010100000000 : 14'b00010100010000;
						assign node1502 = (inp[12]) ? 14'b00000000000001 : node1503;
							assign node1503 = (inp[2]) ? node1505 : 14'b00000000000001;
								assign node1505 = (inp[9]) ? 14'b00000000000001 : node1506;
									assign node1506 = (inp[4]) ? node1508 : 14'b00000000000001;
										assign node1508 = (inp[10]) ? node1514 : node1509;
											assign node1509 = (inp[7]) ? node1511 : 14'b10000001001010;
												assign node1511 = (inp[1]) ? 14'b10000000000000 : 14'b00000000000001;
											assign node1514 = (inp[7]) ? node1516 : 14'b00000000000001;
												assign node1516 = (inp[1]) ? 14'b10000000000000 : 14'b00000000000001;
				assign node1521 = (inp[1]) ? node1781 : node1522;
					assign node1522 = (inp[3]) ? node1720 : node1523;
						assign node1523 = (inp[2]) ? node1645 : node1524;
							assign node1524 = (inp[4]) ? node1572 : node1525;
								assign node1525 = (inp[12]) ? node1547 : node1526;
									assign node1526 = (inp[7]) ? node1532 : node1527;
										assign node1527 = (inp[11]) ? node1529 : 14'b00000000000001;
											assign node1529 = (inp[8]) ? 14'b00000000000001 : 14'b01100100010010;
										assign node1532 = (inp[9]) ? node1540 : node1533;
											assign node1533 = (inp[8]) ? node1537 : node1534;
												assign node1534 = (inp[10]) ? 14'b01100000110010 : 14'b00000000110010;
												assign node1537 = (inp[10]) ? 14'b00000000110000 : 14'b00000010110000;
											assign node1540 = (inp[8]) ? node1544 : node1541;
												assign node1541 = (inp[6]) ? 14'b00000000010010 : 14'b00000010010010;
												assign node1544 = (inp[6]) ? 14'b00000000010000 : 14'b00000010010000;
									assign node1547 = (inp[9]) ? node1561 : node1548;
										assign node1548 = (inp[6]) ? node1556 : node1549;
											assign node1549 = (inp[8]) ? node1553 : node1550;
												assign node1550 = (inp[10]) ? 14'b01100010110000 : 14'b01000010110100;
												assign node1553 = (inp[7]) ? 14'b01000010110100 : 14'b01000110110100;
											assign node1556 = (inp[10]) ? 14'b01100000110000 : node1557;
												assign node1557 = (inp[8]) ? 14'b01000100110100 : 14'b01000000110100;
										assign node1561 = (inp[6]) ? node1565 : node1562;
											assign node1562 = (inp[10]) ? 14'b01100110010000 : 14'b01000110010100;
											assign node1565 = (inp[11]) ? node1569 : node1566;
												assign node1566 = (inp[10]) ? 14'b01100100010000 : 14'b01000000010100;
												assign node1569 = (inp[7]) ? 14'b01000000010100 : 14'b01000100010100;
								assign node1572 = (inp[7]) ? node1612 : node1573;
									assign node1573 = (inp[6]) ? node1593 : node1574;
										assign node1574 = (inp[9]) ? node1584 : node1575;
											assign node1575 = (inp[8]) ? node1581 : node1576;
												assign node1576 = (inp[12]) ? node1578 : 14'b00100110110110;
													assign node1578 = (inp[10]) ? 14'b00100110110000 : 14'b00100110110100;
												assign node1581 = (inp[12]) ? 14'b00000110110100 : 14'b00100110110100;
											assign node1584 = (inp[10]) ? 14'b00100110010010 : node1585;
												assign node1585 = (inp[8]) ? node1589 : node1586;
													assign node1586 = (inp[12]) ? 14'b00100110010100 : 14'b00100110010110;
													assign node1589 = (inp[12]) ? 14'b00000110010100 : 14'b00100110010100;
										assign node1593 = (inp[9]) ? node1605 : node1594;
											assign node1594 = (inp[8]) ? node1602 : node1595;
												assign node1595 = (inp[12]) ? node1599 : node1596;
													assign node1596 = (inp[10]) ? 14'b00100100110010 : 14'b00100100110110;
													assign node1599 = (inp[11]) ? 14'b00100100110100 : 14'b00100100110000;
												assign node1602 = (inp[12]) ? 14'b00000100110100 : 14'b00100100110100;
											assign node1605 = (inp[12]) ? node1609 : node1606;
												assign node1606 = (inp[8]) ? 14'b00100100010100 : 14'b00100100010110;
												assign node1609 = (inp[8]) ? 14'b00000100010100 : 14'b00100100010100;
									assign node1612 = (inp[9]) ? node1628 : node1613;
										assign node1613 = (inp[6]) ? node1619 : node1614;
											assign node1614 = (inp[8]) ? 14'b00000010110100 : node1615;
												assign node1615 = (inp[10]) ? 14'b00100010110000 : 14'b00100010110100;
											assign node1619 = (inp[8]) ? node1625 : node1620;
												assign node1620 = (inp[12]) ? node1622 : 14'b00100000110010;
													assign node1622 = (inp[10]) ? 14'b00100000110000 : 14'b00100000110100;
												assign node1625 = (inp[12]) ? 14'b00000000110100 : 14'b00100000110100;
										assign node1628 = (inp[6]) ? node1636 : node1629;
											assign node1629 = (inp[11]) ? node1631 : 14'b00000010010100;
												assign node1631 = (inp[10]) ? node1633 : 14'b00100010010100;
													assign node1633 = (inp[8]) ? 14'b00100010010100 : 14'b00100010010010;
											assign node1636 = (inp[8]) ? node1642 : node1637;
												assign node1637 = (inp[12]) ? 14'b00100000010100 : node1638;
													assign node1638 = (inp[10]) ? 14'b00100000010010 : 14'b00100000010110;
												assign node1642 = (inp[12]) ? 14'b00000000010100 : 14'b00100000010100;
							assign node1645 = (inp[4]) ? node1705 : node1646;
								assign node1646 = (inp[10]) ? node1690 : node1647;
									assign node1647 = (inp[9]) ? node1667 : node1648;
										assign node1648 = (inp[8]) ? node1658 : node1649;
											assign node1649 = (inp[12]) ? node1651 : 14'b01100010110110;
												assign node1651 = (inp[6]) ? node1655 : node1652;
													assign node1652 = (inp[7]) ? 14'b01100010110100 : 14'b01100110110100;
													assign node1655 = (inp[7]) ? 14'b01100000110100 : 14'b01100100110100;
											assign node1658 = (inp[12]) ? node1660 : 14'b01100100110100;
												assign node1660 = (inp[6]) ? node1664 : node1661;
													assign node1661 = (inp[7]) ? 14'b01000010110000 : 14'b01000110110000;
													assign node1664 = (inp[7]) ? 14'b01000000110000 : 14'b01000100110000;
										assign node1667 = (inp[6]) ? node1677 : node1668;
											assign node1668 = (inp[7]) ? 14'b01100010010100 : node1669;
												assign node1669 = (inp[12]) ? node1673 : node1670;
													assign node1670 = (inp[8]) ? 14'b01100110010100 : 14'b01100110010110;
													assign node1673 = (inp[8]) ? 14'b01000110010000 : 14'b01100110010100;
											assign node1677 = (inp[12]) ? node1685 : node1678;
												assign node1678 = (inp[7]) ? node1682 : node1679;
													assign node1679 = (inp[11]) ? 14'b01100100010110 : 14'b01100100010100;
													assign node1682 = (inp[8]) ? 14'b01100000010100 : 14'b01100000010110;
												assign node1685 = (inp[8]) ? node1687 : 14'b01100100010100;
													assign node1687 = (inp[7]) ? 14'b01000000010000 : 14'b01000100010000;
									assign node1690 = (inp[8]) ? node1692 : 14'b00000000000001;
										assign node1692 = (inp[12]) ? node1700 : node1693;
											assign node1693 = (inp[7]) ? node1697 : node1694;
												assign node1694 = (inp[6]) ? 14'b01100100110100 : 14'b01100110110100;
												assign node1697 = (inp[9]) ? 14'b01100000010100 : 14'b01100000110100;
											assign node1700 = (inp[7]) ? 14'b01000000010000 : node1701;
												assign node1701 = (inp[9]) ? 14'b01000110010000 : 14'b01000110110000;
								assign node1705 = (inp[8]) ? 14'b00000000000001 : node1706;
									assign node1706 = (inp[7]) ? 14'b00000000000001 : node1707;
										assign node1707 = (inp[12]) ? node1711 : node1708;
											assign node1708 = (inp[10]) ? 14'b00000100010010 : 14'b00000000000001;
											assign node1711 = (inp[9]) ? node1715 : node1712;
												assign node1712 = (inp[10]) ? 14'b00000110110000 : 14'b00000110110100;
												assign node1715 = (inp[6]) ? 14'b00000100010100 : 14'b00000110010100;
						assign node1720 = (inp[9]) ? 14'b00000000000001 : node1721;
							assign node1721 = (inp[6]) ? node1731 : node1722;
								assign node1722 = (inp[8]) ? 14'b00000000000001 : node1723;
									assign node1723 = (inp[4]) ? 14'b00000000000001 : node1724;
										assign node1724 = (inp[7]) ? 14'b00000000000001 : node1725;
											assign node1725 = (inp[2]) ? 14'b10000001000000 : 14'b00000000000001;
								assign node1731 = (inp[2]) ? node1763 : node1732;
									assign node1732 = (inp[4]) ? node1746 : node1733;
										assign node1733 = (inp[12]) ? node1735 : 14'b00000000000001;
											assign node1735 = (inp[8]) ? node1743 : node1736;
												assign node1736 = (inp[10]) ? node1740 : node1737;
													assign node1737 = (inp[7]) ? 14'b00000000100000 : 14'b01000000100100;
													assign node1740 = (inp[7]) ? 14'b01100000100000 : 14'b01100100100000;
												assign node1743 = (inp[7]) ? 14'b01000000100100 : 14'b01000100100100;
										assign node1746 = (inp[7]) ? node1756 : node1747;
											assign node1747 = (inp[8]) ? node1753 : node1748;
												assign node1748 = (inp[10]) ? 14'b00100100100010 : node1749;
													assign node1749 = (inp[11]) ? 14'b00100100100110 : 14'b00100100100100;
												assign node1753 = (inp[12]) ? 14'b00000100100100 : 14'b00100100100100;
											assign node1756 = (inp[12]) ? node1760 : node1757;
												assign node1757 = (inp[8]) ? 14'b00100000100100 : 14'b00100000100110;
												assign node1760 = (inp[8]) ? 14'b00000000100100 : 14'b00100000100100;
									assign node1763 = (inp[4]) ? node1775 : node1764;
										assign node1764 = (inp[8]) ? node1770 : node1765;
											assign node1765 = (inp[10]) ? 14'b00000000000001 : node1766;
												assign node1766 = (inp[12]) ? 14'b01100000100100 : 14'b01100100100110;
											assign node1770 = (inp[12]) ? 14'b01000000100000 : node1771;
												assign node1771 = (inp[7]) ? 14'b01100000100100 : 14'b01100100100100;
										assign node1775 = (inp[7]) ? 14'b00000000000001 : node1776;
											assign node1776 = (inp[8]) ? 14'b00000000000001 : 14'b00000100100010;
					assign node1781 = (inp[7]) ? 14'b00000000000001 : node1782;
						assign node1782 = (inp[12]) ? 14'b00000000000001 : node1783;
							assign node1783 = (inp[6]) ? 14'b00000000000001 : node1784;
								assign node1784 = (inp[2]) ? node1792 : node1785;
									assign node1785 = (inp[9]) ? node1787 : 14'b00000000000001;
										assign node1787 = (inp[3]) ? node1789 : 14'b00000000000001;
											assign node1789 = (inp[10]) ? 14'b00000000000001 : 14'b10000000000010;
									assign node1792 = (inp[9]) ? 14'b00000000000001 : node1793;
										assign node1793 = (inp[3]) ? 14'b00000000000001 : node1794;
											assign node1794 = (inp[4]) ? 14'b10000001000010 : node1795;
												assign node1795 = (inp[10]) ? 14'b10000000001010 : 14'b00000000000001;
			assign node1804 = (inp[12]) ? node2118 : node1805;
				assign node1805 = (inp[2]) ? node1991 : node1806;
					assign node1806 = (inp[8]) ? node1872 : node1807;
						assign node1807 = (inp[10]) ? 14'b00000000000001 : node1808;
							assign node1808 = (inp[1]) ? node1848 : node1809;
								assign node1809 = (inp[3]) ? node1831 : node1810;
									assign node1810 = (inp[9]) ? node1822 : node1811;
										assign node1811 = (inp[0]) ? node1815 : node1812;
											assign node1812 = (inp[7]) ? 14'b01010000110110 : 14'b01010100110110;
											assign node1815 = (inp[4]) ? 14'b00000100110110 : node1816;
												assign node1816 = (inp[7]) ? node1818 : 14'b01000110110110;
													assign node1818 = (inp[11]) ? 14'b01000010110110 : 14'b01000000110110;
										assign node1822 = (inp[4]) ? node1826 : node1823;
											assign node1823 = (inp[6]) ? 14'b01000100010110 : 14'b01000010010110;
											assign node1826 = (inp[6]) ? node1828 : 14'b00000110010110;
												assign node1828 = (inp[0]) ? 14'b00000000010110 : 14'b00010100010110;
									assign node1831 = (inp[0]) ? node1839 : node1832;
										assign node1832 = (inp[6]) ? 14'b00000000000001 : node1833;
											assign node1833 = (inp[4]) ? node1835 : 14'b01010110010110;
												assign node1835 = (inp[11]) ? 14'b00010010010110 : 14'b00010110010110;
										assign node1839 = (inp[6]) ? node1841 : 14'b00000000000001;
											assign node1841 = (inp[9]) ? 14'b00000000000001 : node1842;
												assign node1842 = (inp[4]) ? node1844 : 14'b01000000100110;
													assign node1844 = (inp[7]) ? 14'b00000000100110 : 14'b00000100100110;
								assign node1848 = (inp[0]) ? 14'b00000000000001 : node1849;
									assign node1849 = (inp[3]) ? node1863 : node1850;
										assign node1850 = (inp[6]) ? node1856 : node1851;
											assign node1851 = (inp[9]) ? node1853 : 14'b00010010100110;
												assign node1853 = (inp[4]) ? 14'b00010010000110 : 14'b01010010000110;
											assign node1856 = (inp[9]) ? node1860 : node1857;
												assign node1857 = (inp[7]) ? 14'b01010000100110 : 14'b00010100100110;
												assign node1860 = (inp[4]) ? 14'b00010000000110 : 14'b01010100000110;
										assign node1863 = (inp[6]) ? 14'b00000000000001 : node1864;
											assign node1864 = (inp[9]) ? node1866 : 14'b01000110100110;
												assign node1866 = (inp[4]) ? 14'b00000010000110 : 14'b01000010000110;
						assign node1872 = (inp[1]) ? node1954 : node1873;
							assign node1873 = (inp[3]) ? node1927 : node1874;
								assign node1874 = (inp[4]) ? node1902 : node1875;
									assign node1875 = (inp[9]) ? node1889 : node1876;
										assign node1876 = (inp[0]) ? node1882 : node1877;
											assign node1877 = (inp[6]) ? node1879 : 14'b00000000000001;
												assign node1879 = (inp[7]) ? 14'b01110000110000 : 14'b01110100110000;
											assign node1882 = (inp[7]) ? node1886 : node1883;
												assign node1883 = (inp[6]) ? 14'b01100100110000 : 14'b01100110110000;
												assign node1886 = (inp[6]) ? 14'b01100000110000 : 14'b01100010110000;
										assign node1889 = (inp[6]) ? node1895 : node1890;
											assign node1890 = (inp[0]) ? 14'b01100010010000 : node1891;
												assign node1891 = (inp[7]) ? 14'b01100000000000 : 14'b01100100000000;
											assign node1895 = (inp[7]) ? node1899 : node1896;
												assign node1896 = (inp[11]) ? 14'b01110100010000 : 14'b01100100010000;
												assign node1899 = (inp[0]) ? 14'b01100000010000 : 14'b01110000010000;
									assign node1902 = (inp[0]) ? node1914 : node1903;
										assign node1903 = (inp[6]) ? node1907 : node1904;
											assign node1904 = (inp[9]) ? 14'b00100000000000 : 14'b00000000000001;
											assign node1907 = (inp[9]) ? node1911 : node1908;
												assign node1908 = (inp[11]) ? 14'b00110100110000 : 14'b00110000110000;
												assign node1911 = (inp[7]) ? 14'b00110000010000 : 14'b00110100010000;
										assign node1914 = (inp[9]) ? node1920 : node1915;
											assign node1915 = (inp[7]) ? node1917 : 14'b00100110110000;
												assign node1917 = (inp[6]) ? 14'b00100000110000 : 14'b00100010110000;
											assign node1920 = (inp[7]) ? node1924 : node1921;
												assign node1921 = (inp[6]) ? 14'b00100100010000 : 14'b00100110010000;
												assign node1924 = (inp[6]) ? 14'b00100000010000 : 14'b00100010010000;
								assign node1927 = (inp[0]) ? node1943 : node1928;
									assign node1928 = (inp[6]) ? 14'b00000000000001 : node1929;
										assign node1929 = (inp[9]) ? node1937 : node1930;
											assign node1930 = (inp[7]) ? node1934 : node1931;
												assign node1931 = (inp[4]) ? 14'b00110110110000 : 14'b01110110110000;
												assign node1934 = (inp[4]) ? 14'b00110010110000 : 14'b01110010110000;
											assign node1937 = (inp[4]) ? 14'b00110010010000 : node1938;
												assign node1938 = (inp[7]) ? 14'b01110010010000 : 14'b01110110010000;
									assign node1943 = (inp[6]) ? node1945 : 14'b00000000000001;
										assign node1945 = (inp[9]) ? 14'b00000000000001 : node1946;
											assign node1946 = (inp[7]) ? node1950 : node1947;
												assign node1947 = (inp[4]) ? 14'b00100100100000 : 14'b01100100100000;
												assign node1950 = (inp[4]) ? 14'b00100000100000 : 14'b01100000100000;
							assign node1954 = (inp[0]) ? 14'b00000000000001 : node1955;
								assign node1955 = (inp[3]) ? node1979 : node1956;
									assign node1956 = (inp[6]) ? node1970 : node1957;
										assign node1957 = (inp[7]) ? node1963 : node1958;
											assign node1958 = (inp[4]) ? node1960 : 14'b01110110000000;
												assign node1960 = (inp[9]) ? 14'b00110110000000 : 14'b00110110100000;
											assign node1963 = (inp[11]) ? node1967 : node1964;
												assign node1964 = (inp[9]) ? 14'b01110010000000 : 14'b01110010100000;
												assign node1967 = (inp[9]) ? 14'b00110010000000 : 14'b00110010100000;
										assign node1970 = (inp[7]) ? node1974 : node1971;
											assign node1971 = (inp[9]) ? 14'b00110100000000 : 14'b01110100100000;
											assign node1974 = (inp[4]) ? 14'b00110000100000 : node1975;
												assign node1975 = (inp[9]) ? 14'b01110000000000 : 14'b01110000100000;
									assign node1979 = (inp[6]) ? 14'b00000000000001 : node1980;
										assign node1980 = (inp[4]) ? node1984 : node1981;
											assign node1981 = (inp[9]) ? 14'b01100010000000 : 14'b01100010100000;
											assign node1984 = (inp[7]) ? 14'b00100010000000 : node1985;
												assign node1985 = (inp[9]) ? 14'b00100110000000 : 14'b00100110100000;
					assign node1991 = (inp[7]) ? 14'b00000000000001 : node1992;
						assign node1992 = (inp[10]) ? node2082 : node1993;
							assign node1993 = (inp[8]) ? node2051 : node1994;
								assign node1994 = (inp[3]) ? node2026 : node1995;
									assign node1995 = (inp[1]) ? node2011 : node1996;
										assign node1996 = (inp[6]) ? node2000 : node1997;
											assign node1997 = (inp[0]) ? 14'b01000010110010 : 14'b00000000000001;
											assign node2000 = (inp[9]) ? node2006 : node2001;
												assign node2001 = (inp[4]) ? node2003 : 14'b01000100110010;
													assign node2003 = (inp[0]) ? 14'b01000000110010 : 14'b01010000110010;
												assign node2006 = (inp[0]) ? node2008 : 14'b01010100010010;
													assign node2008 = (inp[4]) ? 14'b01000000010010 : 14'b01000100010010;
										assign node2011 = (inp[0]) ? 14'b00000000000001 : node2012;
											assign node2012 = (inp[9]) ? node2018 : node2013;
												assign node2013 = (inp[6]) ? node2015 : 14'b01010010100010;
													assign node2015 = (inp[4]) ? 14'b01010000100010 : 14'b01010100100010;
												assign node2018 = (inp[4]) ? node2022 : node2019;
													assign node2019 = (inp[11]) ? 14'b01010100000010 : 14'b01010110000010;
													assign node2022 = (inp[6]) ? 14'b01010000000010 : 14'b01010010000010;
									assign node2026 = (inp[9]) ? node2042 : node2027;
										assign node2027 = (inp[4]) ? node2037 : node2028;
											assign node2028 = (inp[1]) ? node2034 : node2029;
												assign node2029 = (inp[6]) ? node2031 : 14'b00000000000001;
													assign node2031 = (inp[0]) ? 14'b01000100100010 : 14'b00000000000001;
												assign node2034 = (inp[6]) ? 14'b00000000000001 : 14'b01000110100010;
											assign node2037 = (inp[1]) ? 14'b00000000000001 : node2038;
												assign node2038 = (inp[6]) ? 14'b01000000100010 : 14'b01010010110010;
										assign node2042 = (inp[0]) ? 14'b00000000000001 : node2043;
											assign node2043 = (inp[6]) ? 14'b00000000000001 : node2044;
												assign node2044 = (inp[1]) ? node2046 : 14'b01010110010010;
													assign node2046 = (inp[11]) ? 14'b01000010000010 : 14'b01000110000010;
								assign node2051 = (inp[1]) ? node2075 : node2052;
									assign node2052 = (inp[4]) ? node2060 : node2053;
										assign node2053 = (inp[9]) ? 14'b00000000000001 : node2054;
											assign node2054 = (inp[6]) ? node2056 : 14'b00000000000001;
												assign node2056 = (inp[3]) ? 14'b10000001001000 : 14'b00000000000001;
										assign node2060 = (inp[3]) ? node2068 : node2061;
											assign node2061 = (inp[9]) ? node2065 : node2062;
												assign node2062 = (inp[6]) ? 14'b00000100110000 : 14'b00000110110000;
												assign node2065 = (inp[0]) ? 14'b00000100010000 : 14'b00010100010000;
											assign node2068 = (inp[6]) ? node2072 : node2069;
												assign node2069 = (inp[9]) ? 14'b00010110010000 : 14'b00000000000001;
												assign node2072 = (inp[0]) ? 14'b00000100100000 : 14'b00000000000001;
									assign node2075 = (inp[0]) ? 14'b00000000000001 : node2076;
										assign node2076 = (inp[6]) ? 14'b00000000000001 : node2077;
											assign node2077 = (inp[4]) ? 14'b00000110100000 : 14'b00000000000001;
							assign node2082 = (inp[8]) ? node2084 : 14'b00000000000001;
								assign node2084 = (inp[4]) ? node2086 : 14'b00000000000001;
									assign node2086 = (inp[6]) ? node2104 : node2087;
										assign node2087 = (inp[0]) ? node2101 : node2088;
											assign node2088 = (inp[3]) ? node2094 : node2089;
												assign node2089 = (inp[1]) ? 14'b00010110100000 : node2090;
													assign node2090 = (inp[9]) ? 14'b00000100000000 : 14'b00000000000001;
												assign node2094 = (inp[1]) ? node2098 : node2095;
													assign node2095 = (inp[9]) ? 14'b00010110010000 : 14'b00010110110000;
													assign node2098 = (inp[9]) ? 14'b00000110000000 : 14'b00000110100000;
											assign node2101 = (inp[1]) ? 14'b00000000000001 : 14'b00000110010000;
										assign node2104 = (inp[3]) ? node2112 : node2105;
											assign node2105 = (inp[1]) ? node2109 : node2106;
												assign node2106 = (inp[9]) ? 14'b00000100010000 : 14'b00000100110000;
												assign node2109 = (inp[0]) ? 14'b00000000000001 : 14'b00010100000000;
											assign node2112 = (inp[0]) ? node2114 : 14'b00000000000001;
												assign node2114 = (inp[1]) ? 14'b00000000000001 : 14'b00000100100000;
				assign node2118 = (inp[8]) ? node2196 : node2119;
					assign node2119 = (inp[10]) ? 14'b00000000000001 : node2120;
						assign node2120 = (inp[3]) ? node2172 : node2121;
							assign node2121 = (inp[4]) ? node2151 : node2122;
								assign node2122 = (inp[7]) ? node2136 : node2123;
									assign node2123 = (inp[2]) ? node2131 : node2124;
										assign node2124 = (inp[0]) ? 14'b01000110110100 : node2125;
											assign node2125 = (inp[6]) ? node2127 : 14'b01010110000100;
												assign node2127 = (inp[9]) ? 14'b01010100000100 : 14'b01010100100100;
										assign node2131 = (inp[1]) ? 14'b00000000000001 : node2132;
											assign node2132 = (inp[6]) ? 14'b01010100110000 : 14'b01000110110000;
									assign node2136 = (inp[2]) ? node2138 : 14'b00000000000001;
										assign node2138 = (inp[9]) ? node2146 : node2139;
											assign node2139 = (inp[0]) ? node2143 : node2140;
												assign node2140 = (inp[1]) ? 14'b01010010100000 : 14'b00000000000001;
												assign node2143 = (inp[1]) ? 14'b00000000000001 : 14'b01000000110000;
											assign node2146 = (inp[0]) ? node2148 : 14'b01010000010000;
												assign node2148 = (inp[11]) ? 14'b01000010010000 : 14'b01000000010000;
								assign node2151 = (inp[7]) ? node2153 : 14'b00000000000001;
									assign node2153 = (inp[0]) ? node2165 : node2154;
										assign node2154 = (inp[1]) ? node2160 : node2155;
											assign node2155 = (inp[9]) ? node2157 : 14'b00000000000001;
												assign node2157 = (inp[6]) ? 14'b00010000010100 : 14'b00000000000100;
											assign node2160 = (inp[9]) ? 14'b00010010000100 : node2161;
												assign node2161 = (inp[6]) ? 14'b00010000100100 : 14'b00010010100100;
										assign node2165 = (inp[1]) ? 14'b00000000000001 : node2166;
											assign node2166 = (inp[2]) ? 14'b00000000000001 : node2167;
												assign node2167 = (inp[11]) ? 14'b00000000110100 : 14'b00000010010100;
							assign node2172 = (inp[0]) ? 14'b00000000000001 : node2173;
								assign node2173 = (inp[6]) ? 14'b00000000000001 : node2174;
									assign node2174 = (inp[11]) ? node2184 : node2175;
										assign node2175 = (inp[2]) ? 14'b00000000000001 : node2176;
											assign node2176 = (inp[7]) ? node2178 : 14'b00000000000001;
												assign node2178 = (inp[4]) ? node2180 : 14'b00000000000001;
													assign node2180 = (inp[9]) ? 14'b00000010000100 : 14'b00000010100100;
										assign node2184 = (inp[1]) ? 14'b00000000000001 : node2185;
											assign node2185 = (inp[4]) ? node2189 : node2186;
												assign node2186 = (inp[9]) ? 14'b01010010010000 : 14'b01010110110000;
												assign node2189 = (inp[9]) ? 14'b00010010010100 : 14'b00010010110100;
					assign node2196 = (inp[4]) ? node2242 : node2197;
						assign node2197 = (inp[6]) ? node2231 : node2198;
							assign node2198 = (inp[9]) ? node2220 : node2199;
								assign node2199 = (inp[3]) ? 14'b00000000000001 : node2200;
									assign node2200 = (inp[11]) ? node2206 : node2201;
										assign node2201 = (inp[0]) ? 14'b00000000000001 : node2202;
											assign node2202 = (inp[7]) ? 14'b10001000001000 : 14'b00000000000001;
										assign node2206 = (inp[0]) ? node2214 : node2207;
											assign node2207 = (inp[2]) ? node2209 : 14'b00000000000001;
												assign node2209 = (inp[1]) ? 14'b00000000000001 : node2210;
													assign node2210 = (inp[7]) ? 14'b10001000001000 : 14'b00000000000001;
											assign node2214 = (inp[2]) ? 14'b00000000000001 : node2215;
												assign node2215 = (inp[7]) ? 14'b00000000000001 : 14'b10001001001000;
								assign node2220 = (inp[0]) ? node2222 : 14'b00000000000001;
									assign node2222 = (inp[2]) ? node2224 : 14'b00000000000001;
										assign node2224 = (inp[11]) ? node2226 : 14'b00000000000001;
											assign node2226 = (inp[10]) ? node2228 : 14'b00000000000001;
												assign node2228 = (inp[3]) ? 14'b10001000000000 : 14'b00000000000001;
							assign node2231 = (inp[3]) ? node2233 : 14'b00000000000001;
								assign node2233 = (inp[0]) ? node2235 : 14'b00000000000001;
									assign node2235 = (inp[1]) ? node2237 : 14'b00000000000001;
										assign node2237 = (inp[7]) ? node2239 : 14'b00000000000001;
											assign node2239 = (inp[9]) ? 14'b10001001000000 : 14'b00000000000001;
						assign node2242 = (inp[11]) ? 14'b00000000000001 : node2243;
							assign node2243 = (inp[0]) ? node2245 : 14'b00000000000001;
								assign node2245 = (inp[10]) ? node2247 : 14'b00000000000001;
									assign node2247 = (inp[7]) ? node2249 : 14'b00000000000001;
										assign node2249 = (inp[6]) ? node2251 : 14'b00000000000001;
											assign node2251 = (inp[2]) ? 14'b10001001001010 : 14'b00000000000001;

endmodule