module dtc_split5_bm86 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node15;
	wire [3-1:0] node16;
	wire [3-1:0] node19;
	wire [3-1:0] node20;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node30;
	wire [3-1:0] node32;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node39;
	wire [3-1:0] node43;
	wire [3-1:0] node44;
	wire [3-1:0] node46;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node59;
	wire [3-1:0] node62;
	wire [3-1:0] node63;
	wire [3-1:0] node67;
	wire [3-1:0] node68;
	wire [3-1:0] node70;
	wire [3-1:0] node72;
	wire [3-1:0] node75;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node81;
	wire [3-1:0] node84;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node95;
	wire [3-1:0] node96;
	wire [3-1:0] node100;
	wire [3-1:0] node101;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node108;
	wire [3-1:0] node110;
	wire [3-1:0] node112;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node120;
	wire [3-1:0] node121;
	wire [3-1:0] node122;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node128;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node134;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node145;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node160;
	wire [3-1:0] node161;
	wire [3-1:0] node163;
	wire [3-1:0] node168;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node173;
	wire [3-1:0] node174;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node188;
	wire [3-1:0] node190;
	wire [3-1:0] node193;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node200;
	wire [3-1:0] node203;
	wire [3-1:0] node207;
	wire [3-1:0] node208;
	wire [3-1:0] node209;
	wire [3-1:0] node210;
	wire [3-1:0] node214;
	wire [3-1:0] node216;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node225;
	wire [3-1:0] node228;
	wire [3-1:0] node229;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node236;
	wire [3-1:0] node237;
	wire [3-1:0] node238;
	wire [3-1:0] node241;
	wire [3-1:0] node244;
	wire [3-1:0] node246;
	wire [3-1:0] node249;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node254;
	wire [3-1:0] node255;
	wire [3-1:0] node258;
	wire [3-1:0] node261;
	wire [3-1:0] node262;
	wire [3-1:0] node263;
	wire [3-1:0] node267;
	wire [3-1:0] node269;
	wire [3-1:0] node272;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node286;
	wire [3-1:0] node288;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node292;
	wire [3-1:0] node294;
	wire [3-1:0] node295;
	wire [3-1:0] node299;
	wire [3-1:0] node300;
	wire [3-1:0] node301;
	wire [3-1:0] node304;
	wire [3-1:0] node306;
	wire [3-1:0] node309;
	wire [3-1:0] node310;
	wire [3-1:0] node311;
	wire [3-1:0] node316;
	wire [3-1:0] node317;
	wire [3-1:0] node319;
	wire [3-1:0] node322;
	wire [3-1:0] node323;
	wire [3-1:0] node326;
	wire [3-1:0] node329;
	wire [3-1:0] node331;
	wire [3-1:0] node333;
	wire [3-1:0] node334;
	wire [3-1:0] node336;
	wire [3-1:0] node337;
	wire [3-1:0] node342;
	wire [3-1:0] node344;
	wire [3-1:0] node345;
	wire [3-1:0] node347;
	wire [3-1:0] node348;
	wire [3-1:0] node350;
	wire [3-1:0] node352;
	wire [3-1:0] node355;
	wire [3-1:0] node357;
	wire [3-1:0] node359;
	wire [3-1:0] node362;
	wire [3-1:0] node363;
	wire [3-1:0] node365;
	wire [3-1:0] node367;
	wire [3-1:0] node370;
	wire [3-1:0] node371;
	wire [3-1:0] node372;
	wire [3-1:0] node374;
	wire [3-1:0] node377;
	wire [3-1:0] node380;
	wire [3-1:0] node381;
	wire [3-1:0] node384;

	assign outp = (inp[3]) ? node284 : node1;
		assign node1 = (inp[0]) ? node117 : node2;
			assign node2 = (inp[6]) ? 3'b000 : node3;
				assign node3 = (inp[4]) ? node89 : node4;
					assign node4 = (inp[9]) ? node54 : node5;
						assign node5 = (inp[7]) ? node35 : node6;
							assign node6 = (inp[1]) ? node14 : node7;
								assign node7 = (inp[2]) ? node9 : 3'b000;
									assign node9 = (inp[10]) ? node11 : 3'b000;
										assign node11 = (inp[8]) ? 3'b000 : 3'b100;
								assign node14 = (inp[5]) ? node26 : node15;
									assign node15 = (inp[2]) ? node19 : node16;
										assign node16 = (inp[10]) ? 3'b110 : 3'b100;
										assign node19 = (inp[8]) ? node23 : node20;
											assign node20 = (inp[10]) ? 3'b110 : 3'b010;
											assign node23 = (inp[11]) ? 3'b000 : 3'b010;
									assign node26 = (inp[8]) ? node30 : node27;
										assign node27 = (inp[2]) ? 3'b100 : 3'b000;
										assign node30 = (inp[11]) ? node32 : 3'b000;
											assign node32 = (inp[2]) ? 3'b010 : 3'b100;
							assign node35 = (inp[1]) ? node43 : node36;
								assign node36 = (inp[5]) ? 3'b010 : node37;
									assign node37 = (inp[2]) ? node39 : 3'b010;
										assign node39 = (inp[11]) ? 3'b000 : 3'b010;
								assign node43 = (inp[5]) ? node49 : node44;
									assign node44 = (inp[11]) ? node46 : 3'b110;
										assign node46 = (inp[2]) ? 3'b100 : 3'b110;
									assign node49 = (inp[11]) ? node51 : 3'b010;
										assign node51 = (inp[2]) ? 3'b110 : 3'b010;
						assign node54 = (inp[7]) ? node84 : node55;
							assign node55 = (inp[11]) ? node67 : node56;
								assign node56 = (inp[1]) ? node58 : 3'b110;
									assign node58 = (inp[8]) ? node62 : node59;
										assign node59 = (inp[10]) ? 3'b001 : 3'b010;
										assign node62 = (inp[2]) ? 3'b110 : node63;
											assign node63 = (inp[10]) ? 3'b000 : 3'b100;
								assign node67 = (inp[8]) ? node75 : node68;
									assign node68 = (inp[1]) ? node70 : 3'b110;
										assign node70 = (inp[2]) ? node72 : 3'b110;
											assign node72 = (inp[10]) ? 3'b001 : 3'b100;
									assign node75 = (inp[1]) ? node77 : 3'b001;
										assign node77 = (inp[2]) ? node81 : node78;
											assign node78 = (inp[10]) ? 3'b110 : 3'b010;
											assign node81 = (inp[5]) ? 3'b100 : 3'b101;
							assign node84 = (inp[11]) ? node86 : 3'b011;
								assign node86 = (inp[2]) ? 3'b111 : 3'b011;
					assign node89 = (inp[7]) ? 3'b000 : node90;
						assign node90 = (inp[9]) ? node92 : 3'b000;
							assign node92 = (inp[1]) ? node100 : node93;
								assign node93 = (inp[10]) ? node95 : 3'b000;
									assign node95 = (inp[5]) ? 3'b000 : node96;
										assign node96 = (inp[2]) ? 3'b010 : 3'b000;
								assign node100 = (inp[2]) ? node108 : node101;
									assign node101 = (inp[10]) ? node103 : 3'b000;
										assign node103 = (inp[5]) ? 3'b000 : node104;
											assign node104 = (inp[8]) ? 3'b100 : 3'b000;
									assign node108 = (inp[8]) ? node110 : 3'b100;
										assign node110 = (inp[10]) ? node112 : 3'b000;
											assign node112 = (inp[5]) ? 3'b100 : 3'b010;
			assign node117 = (inp[6]) ? node279 : node118;
				assign node118 = (inp[4]) ? node168 : node119;
					assign node119 = (inp[7]) ? 3'b111 : node120;
						assign node120 = (inp[1]) ? node152 : node121;
							assign node121 = (inp[5]) ? node139 : node122;
								assign node122 = (inp[9]) ? node132 : node123;
									assign node123 = (inp[8]) ? 3'b001 : node124;
										assign node124 = (inp[2]) ? node128 : node125;
											assign node125 = (inp[10]) ? 3'b101 : 3'b001;
											assign node128 = (inp[11]) ? 3'b011 : 3'b101;
									assign node132 = (inp[10]) ? 3'b111 : node133;
										assign node133 = (inp[8]) ? 3'b111 : node134;
											assign node134 = (inp[2]) ? 3'b011 : 3'b001;
								assign node139 = (inp[9]) ? node145 : node140;
									assign node140 = (inp[8]) ? 3'b010 : node141;
										assign node141 = (inp[10]) ? 3'b110 : 3'b010;
									assign node145 = (inp[10]) ? 3'b011 : node146;
										assign node146 = (inp[2]) ? 3'b101 : node147;
											assign node147 = (inp[8]) ? 3'b011 : 3'b001;
							assign node152 = (inp[9]) ? node160 : node153;
								assign node153 = (inp[5]) ? node155 : 3'b111;
									assign node155 = (inp[2]) ? node157 : 3'b101;
										assign node157 = (inp[11]) ? 3'b111 : 3'b101;
								assign node160 = (inp[10]) ? 3'b111 : node161;
									assign node161 = (inp[5]) ? node163 : 3'b111;
										assign node163 = (inp[2]) ? 3'b111 : 3'b011;
					assign node168 = (inp[9]) ? node228 : node169;
						assign node169 = (inp[1]) ? node193 : node170;
							assign node170 = (inp[5]) ? node178 : node171;
								assign node171 = (inp[10]) ? node173 : 3'b100;
									assign node173 = (inp[7]) ? 3'b100 : node174;
										assign node174 = (inp[2]) ? 3'b110 : 3'b100;
								assign node178 = (inp[7]) ? node188 : node179;
									assign node179 = (inp[10]) ? node183 : node180;
										assign node180 = (inp[11]) ? 3'b000 : 3'b100;
										assign node183 = (inp[2]) ? node185 : 3'b000;
											assign node185 = (inp[8]) ? 3'b100 : 3'b000;
									assign node188 = (inp[11]) ? node190 : 3'b100;
										assign node190 = (inp[2]) ? 3'b000 : 3'b100;
							assign node193 = (inp[5]) ? node207 : node194;
								assign node194 = (inp[7]) ? 3'b110 : node195;
									assign node195 = (inp[8]) ? node203 : node196;
										assign node196 = (inp[2]) ? node200 : node197;
											assign node197 = (inp[10]) ? 3'b100 : 3'b110;
											assign node200 = (inp[11]) ? 3'b110 : 3'b010;
										assign node203 = (inp[2]) ? 3'b100 : 3'b110;
								assign node207 = (inp[2]) ? node219 : node208;
									assign node208 = (inp[11]) ? node214 : node209;
										assign node209 = (inp[7]) ? 3'b100 : node210;
											assign node210 = (inp[8]) ? 3'b100 : 3'b000;
										assign node214 = (inp[8]) ? node216 : 3'b100;
											assign node216 = (inp[7]) ? 3'b100 : 3'b110;
									assign node219 = (inp[10]) ? node221 : 3'b010;
										assign node221 = (inp[11]) ? node225 : node222;
											assign node222 = (inp[7]) ? 3'b100 : 3'b110;
											assign node225 = (inp[7]) ? 3'b010 : 3'b000;
						assign node228 = (inp[7]) ? node272 : node229;
							assign node229 = (inp[1]) ? node249 : node230;
								assign node230 = (inp[5]) ? node236 : node231;
									assign node231 = (inp[10]) ? 3'b110 : node232;
										assign node232 = (inp[11]) ? 3'b101 : 3'b110;
									assign node236 = (inp[2]) ? node244 : node237;
										assign node237 = (inp[10]) ? node241 : node238;
											assign node238 = (inp[8]) ? 3'b100 : 3'b110;
											assign node241 = (inp[11]) ? 3'b010 : 3'b000;
										assign node244 = (inp[10]) ? node246 : 3'b010;
											assign node246 = (inp[11]) ? 3'b110 : 3'b010;
								assign node249 = (inp[2]) ? node261 : node250;
									assign node250 = (inp[11]) ? node254 : node251;
										assign node251 = (inp[10]) ? 3'b110 : 3'b010;
										assign node254 = (inp[10]) ? node258 : node255;
											assign node255 = (inp[5]) ? 3'b110 : 3'b101;
											assign node258 = (inp[8]) ? 3'b011 : 3'b001;
									assign node261 = (inp[8]) ? node267 : node262;
										assign node262 = (inp[11]) ? 3'b101 : node263;
											assign node263 = (inp[10]) ? 3'b011 : 3'b001;
										assign node267 = (inp[5]) ? node269 : 3'b111;
											assign node269 = (inp[11]) ? 3'b011 : 3'b001;
							assign node272 = (inp[5]) ? node274 : 3'b111;
								assign node274 = (inp[11]) ? node276 : 3'b101;
									assign node276 = (inp[2]) ? 3'b011 : 3'b101;
				assign node279 = (inp[4]) ? 3'b000 : node280;
					assign node280 = (inp[9]) ? 3'b111 : 3'b000;
		assign node284 = (inp[9]) ? node286 : 3'b000;
			assign node286 = (inp[0]) ? node288 : 3'b000;
				assign node288 = (inp[4]) ? node342 : node289;
					assign node289 = (inp[6]) ? node329 : node290;
						assign node290 = (inp[7]) ? node316 : node291;
							assign node291 = (inp[1]) ? node299 : node292;
								assign node292 = (inp[2]) ? node294 : 3'b000;
									assign node294 = (inp[5]) ? 3'b000 : node295;
										assign node295 = (inp[10]) ? 3'b100 : 3'b000;
								assign node299 = (inp[10]) ? node309 : node300;
									assign node300 = (inp[5]) ? node304 : node301;
										assign node301 = (inp[2]) ? 3'b001 : 3'b100;
										assign node304 = (inp[2]) ? node306 : 3'b000;
											assign node306 = (inp[8]) ? 3'b000 : 3'b100;
									assign node309 = (inp[5]) ? 3'b100 : node310;
										assign node310 = (inp[8]) ? 3'b110 : node311;
											assign node311 = (inp[11]) ? 3'b110 : 3'b010;
							assign node316 = (inp[2]) ? node322 : node317;
								assign node317 = (inp[1]) ? node319 : 3'b010;
									assign node319 = (inp[5]) ? 3'b010 : 3'b110;
								assign node322 = (inp[5]) ? node326 : node323;
									assign node323 = (inp[11]) ? 3'b101 : 3'b110;
									assign node326 = (inp[11]) ? 3'b110 : 3'b010;
						assign node329 = (inp[1]) ? node331 : 3'b000;
							assign node331 = (inp[5]) ? node333 : 3'b000;
								assign node333 = (inp[8]) ? 3'b000 : node334;
									assign node334 = (inp[2]) ? node336 : 3'b000;
										assign node336 = (inp[7]) ? 3'b001 : node337;
											assign node337 = (inp[11]) ? 3'b001 : 3'b000;
					assign node342 = (inp[1]) ? node344 : 3'b000;
						assign node344 = (inp[11]) ? node362 : node345;
							assign node345 = (inp[6]) ? node347 : 3'b000;
								assign node347 = (inp[8]) ? node355 : node348;
									assign node348 = (inp[5]) ? node350 : 3'b000;
										assign node350 = (inp[2]) ? node352 : 3'b000;
											assign node352 = (inp[7]) ? 3'b100 : 3'b000;
									assign node355 = (inp[7]) ? node357 : 3'b000;
										assign node357 = (inp[2]) ? node359 : 3'b000;
											assign node359 = (inp[5]) ? 3'b010 : 3'b000;
							assign node362 = (inp[2]) ? node370 : node363;
								assign node363 = (inp[8]) ? node365 : 3'b000;
									assign node365 = (inp[6]) ? node367 : 3'b000;
										assign node367 = (inp[7]) ? 3'b100 : 3'b000;
								assign node370 = (inp[7]) ? node380 : node371;
									assign node371 = (inp[5]) ? node377 : node372;
										assign node372 = (inp[8]) ? node374 : 3'b000;
											assign node374 = (inp[6]) ? 3'b000 : 3'b100;
										assign node377 = (inp[6]) ? 3'b100 : 3'b000;
									assign node380 = (inp[6]) ? node384 : node381;
										assign node381 = (inp[5]) ? 3'b000 : 3'b100;
										assign node384 = (inp[5]) ? 3'b010 : 3'b000;

endmodule