module dtc_split125_bm98 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node11;
	wire [3-1:0] node14;
	wire [3-1:0] node16;
	wire [3-1:0] node18;
	wire [3-1:0] node20;
	wire [3-1:0] node22;
	wire [3-1:0] node24;
	wire [3-1:0] node27;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node30;
	wire [3-1:0] node31;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node41;
	wire [3-1:0] node42;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node52;
	wire [3-1:0] node55;
	wire [3-1:0] node56;
	wire [3-1:0] node58;
	wire [3-1:0] node61;
	wire [3-1:0] node62;
	wire [3-1:0] node65;
	wire [3-1:0] node68;
	wire [3-1:0] node69;
	wire [3-1:0] node70;
	wire [3-1:0] node71;
	wire [3-1:0] node73;
	wire [3-1:0] node74;
	wire [3-1:0] node76;
	wire [3-1:0] node77;
	wire [3-1:0] node78;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node90;
	wire [3-1:0] node91;
	wire [3-1:0] node92;
	wire [3-1:0] node93;
	wire [3-1:0] node97;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node108;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node113;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node129;
	wire [3-1:0] node131;
	wire [3-1:0] node132;
	wire [3-1:0] node133;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node142;
	wire [3-1:0] node144;
	wire [3-1:0] node148;
	wire [3-1:0] node149;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node159;
	wire [3-1:0] node161;
	wire [3-1:0] node162;
	wire [3-1:0] node163;
	wire [3-1:0] node164;
	wire [3-1:0] node165;
	wire [3-1:0] node171;
	wire [3-1:0] node172;
	wire [3-1:0] node173;
	wire [3-1:0] node175;
	wire [3-1:0] node180;
	wire [3-1:0] node181;
	wire [3-1:0] node183;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node188;
	wire [3-1:0] node191;
	wire [3-1:0] node193;
	wire [3-1:0] node196;
	wire [3-1:0] node197;
	wire [3-1:0] node198;
	wire [3-1:0] node199;
	wire [3-1:0] node201;
	wire [3-1:0] node205;
	wire [3-1:0] node206;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node214;
	wire [3-1:0] node215;
	wire [3-1:0] node216;
	wire [3-1:0] node217;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node226;

	assign outp = (inp[0]) ? node68 : node1;
		assign node1 = (inp[6]) ? node3 : 3'b111;
			assign node3 = (inp[9]) ? node27 : node4;
				assign node4 = (inp[3]) ? node14 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b100;
						assign node7 = (inp[5]) ? node11 : node8;
							assign node8 = (inp[1]) ? 3'b101 : 3'b100;
							assign node11 = (inp[8]) ? 3'b100 : 3'b000;
					assign node14 = (inp[7]) ? node16 : 3'b010;
						assign node16 = (inp[1]) ? node18 : 3'b010;
							assign node18 = (inp[11]) ? node20 : 3'b110;
								assign node20 = (inp[2]) ? node22 : 3'b010;
									assign node22 = (inp[4]) ? node24 : 3'b010;
										assign node24 = (inp[10]) ? 3'b110 : 3'b010;
				assign node27 = (inp[1]) ? node41 : node28;
					assign node28 = (inp[3]) ? 3'b111 : node29;
						assign node29 = (inp[5]) ? node35 : node30;
							assign node30 = (inp[8]) ? 3'b101 : node31;
								assign node31 = (inp[4]) ? 3'b111 : 3'b101;
							assign node35 = (inp[4]) ? 3'b101 : node36;
								assign node36 = (inp[8]) ? 3'b001 : 3'b101;
					assign node41 = (inp[3]) ? node55 : node42;
						assign node42 = (inp[2]) ? node52 : node43;
							assign node43 = (inp[4]) ? node45 : 3'b001;
								assign node45 = (inp[7]) ? node47 : 3'b100;
									assign node47 = (inp[5]) ? 3'b001 : node48;
										assign node48 = (inp[11]) ? 3'b110 : 3'b001;
							assign node52 = (inp[8]) ? 3'b100 : 3'b110;
						assign node55 = (inp[7]) ? node61 : node56;
							assign node56 = (inp[4]) ? node58 : 3'b011;
								assign node58 = (inp[2]) ? 3'b111 : 3'b001;
							assign node61 = (inp[4]) ? node65 : node62;
								assign node62 = (inp[2]) ? 3'b001 : 3'b101;
								assign node65 = (inp[8]) ? 3'b111 : 3'b011;
		assign node68 = (inp[3]) ? node138 : node69;
			assign node69 = (inp[6]) ? node125 : node70;
				assign node70 = (inp[9]) ? node90 : node71;
					assign node71 = (inp[4]) ? node73 : 3'b010;
						assign node73 = (inp[1]) ? node87 : node74;
							assign node74 = (inp[7]) ? node76 : 3'b010;
								assign node76 = (inp[11]) ? node82 : node77;
									assign node77 = (inp[10]) ? 3'b010 : node78;
										assign node78 = (inp[8]) ? 3'b000 : 3'b010;
									assign node82 = (inp[8]) ? node84 : 3'b000;
										assign node84 = (inp[5]) ? 3'b000 : 3'b010;
							assign node87 = (inp[7]) ? 3'b010 : 3'b000;
					assign node90 = (inp[2]) ? node104 : node91;
						assign node91 = (inp[7]) ? node97 : node92;
							assign node92 = (inp[4]) ? 3'b010 : node93;
								assign node93 = (inp[10]) ? 3'b000 : 3'b010;
							assign node97 = (inp[5]) ? 3'b000 : node98;
								assign node98 = (inp[10]) ? 3'b000 : node99;
									assign node99 = (inp[4]) ? 3'b010 : 3'b000;
						assign node104 = (inp[7]) ? node118 : node105;
							assign node105 = (inp[10]) ? node111 : node106;
								assign node106 = (inp[11]) ? node108 : 3'b010;
									assign node108 = (inp[8]) ? 3'b010 : 3'b000;
								assign node111 = (inp[8]) ? 3'b000 : node112;
									assign node112 = (inp[5]) ? 3'b000 : node113;
										assign node113 = (inp[1]) ? 3'b010 : 3'b000;
							assign node118 = (inp[4]) ? node120 : 3'b010;
								assign node120 = (inp[5]) ? node122 : 3'b010;
									assign node122 = (inp[8]) ? 3'b000 : 3'b010;
				assign node125 = (inp[9]) ? node127 : 3'b000;
					assign node127 = (inp[4]) ? node129 : 3'b000;
						assign node129 = (inp[7]) ? node131 : 3'b100;
							assign node131 = (inp[1]) ? 3'b000 : node132;
								assign node132 = (inp[10]) ? 3'b010 : node133;
									assign node133 = (inp[2]) ? 3'b100 : 3'b110;
			assign node138 = (inp[9]) ? node180 : node139;
				assign node139 = (inp[1]) ? node159 : node140;
					assign node140 = (inp[6]) ? node148 : node141;
						assign node141 = (inp[2]) ? 3'b001 : node142;
							assign node142 = (inp[8]) ? node144 : 3'b111;
								assign node144 = (inp[11]) ? 3'b001 : 3'b101;
						assign node148 = (inp[7]) ? node152 : node149;
							assign node149 = (inp[4]) ? 3'b001 : 3'b000;
							assign node152 = (inp[4]) ? node154 : 3'b000;
								assign node154 = (inp[5]) ? 3'b010 : node155;
									assign node155 = (inp[2]) ? 3'b000 : 3'b100;
					assign node159 = (inp[4]) ? node161 : 3'b000;
						assign node161 = (inp[7]) ? node171 : node162;
							assign node162 = (inp[6]) ? 3'b100 : node163;
								assign node163 = (inp[8]) ? 3'b001 : node164;
									assign node164 = (inp[11]) ? 3'b110 : node165;
										assign node165 = (inp[10]) ? 3'b101 : 3'b001;
							assign node171 = (inp[6]) ? 3'b000 : node172;
								assign node172 = (inp[10]) ? 3'b010 : node173;
									assign node173 = (inp[8]) ? node175 : 3'b010;
										assign node175 = (inp[5]) ? 3'b010 : 3'b100;
				assign node180 = (inp[6]) ? node196 : node181;
					assign node181 = (inp[1]) ? node183 : 3'b111;
						assign node183 = (inp[2]) ? node185 : 3'b001;
							assign node185 = (inp[11]) ? node187 : 3'b011;
								assign node187 = (inp[8]) ? node191 : node188;
									assign node188 = (inp[5]) ? 3'b001 : 3'b101;
									assign node191 = (inp[5]) ? node193 : 3'b110;
										assign node193 = (inp[7]) ? 3'b101 : 3'b111;
					assign node196 = (inp[1]) ? node214 : node197;
						assign node197 = (inp[7]) ? node205 : node198;
							assign node198 = (inp[2]) ? 3'b101 : node199;
								assign node199 = (inp[8]) ? node201 : 3'b010;
									assign node201 = (inp[11]) ? 3'b001 : 3'b101;
							assign node205 = (inp[4]) ? node209 : node206;
								assign node206 = (inp[11]) ? 3'b110 : 3'b010;
								assign node209 = (inp[5]) ? node211 : 3'b001;
									assign node211 = (inp[2]) ? 3'b010 : 3'b001;
						assign node214 = (inp[7]) ? node222 : node215;
							assign node215 = (inp[4]) ? 3'b000 : node216;
								assign node216 = (inp[8]) ? 3'b110 : node217;
									assign node217 = (inp[5]) ? 3'b110 : 3'b010;
							assign node222 = (inp[2]) ? 3'b100 : node223;
								assign node223 = (inp[4]) ? node225 : 3'b100;
									assign node225 = (inp[8]) ? 3'b110 : node226;
										assign node226 = (inp[5]) ? 3'b010 : 3'b110;

endmodule