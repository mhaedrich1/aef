module dtc_split5_bm62 (
	input  wire [16-1:0] inp,
	output wire [4-1:0] outp
);

	wire [4-1:0] node1;
	wire [4-1:0] node2;
	wire [4-1:0] node3;
	wire [4-1:0] node4;
	wire [4-1:0] node5;
	wire [4-1:0] node6;
	wire [4-1:0] node7;
	wire [4-1:0] node8;
	wire [4-1:0] node9;
	wire [4-1:0] node10;
	wire [4-1:0] node11;
	wire [4-1:0] node12;
	wire [4-1:0] node14;
	wire [4-1:0] node15;
	wire [4-1:0] node18;
	wire [4-1:0] node21;
	wire [4-1:0] node22;
	wire [4-1:0] node25;
	wire [4-1:0] node28;
	wire [4-1:0] node29;
	wire [4-1:0] node30;
	wire [4-1:0] node32;
	wire [4-1:0] node35;
	wire [4-1:0] node37;
	wire [4-1:0] node40;
	wire [4-1:0] node41;
	wire [4-1:0] node44;
	wire [4-1:0] node47;
	wire [4-1:0] node48;
	wire [4-1:0] node49;
	wire [4-1:0] node50;
	wire [4-1:0] node51;
	wire [4-1:0] node55;
	wire [4-1:0] node57;
	wire [4-1:0] node60;
	wire [4-1:0] node61;
	wire [4-1:0] node62;
	wire [4-1:0] node64;
	wire [4-1:0] node67;
	wire [4-1:0] node69;
	wire [4-1:0] node73;
	wire [4-1:0] node74;
	wire [4-1:0] node75;
	wire [4-1:0] node78;
	wire [4-1:0] node79;
	wire [4-1:0] node82;
	wire [4-1:0] node85;
	wire [4-1:0] node86;
	wire [4-1:0] node89;
	wire [4-1:0] node92;
	wire [4-1:0] node93;
	wire [4-1:0] node94;
	wire [4-1:0] node95;
	wire [4-1:0] node96;
	wire [4-1:0] node99;
	wire [4-1:0] node102;
	wire [4-1:0] node103;
	wire [4-1:0] node106;
	wire [4-1:0] node109;
	wire [4-1:0] node110;
	wire [4-1:0] node111;
	wire [4-1:0] node114;
	wire [4-1:0] node115;
	wire [4-1:0] node119;
	wire [4-1:0] node121;
	wire [4-1:0] node124;
	wire [4-1:0] node125;
	wire [4-1:0] node126;
	wire [4-1:0] node127;
	wire [4-1:0] node128;
	wire [4-1:0] node131;
	wire [4-1:0] node134;
	wire [4-1:0] node136;
	wire [4-1:0] node139;
	wire [4-1:0] node141;
	wire [4-1:0] node144;
	wire [4-1:0] node145;
	wire [4-1:0] node148;
	wire [4-1:0] node150;
	wire [4-1:0] node151;
	wire [4-1:0] node155;
	wire [4-1:0] node156;
	wire [4-1:0] node157;
	wire [4-1:0] node158;
	wire [4-1:0] node159;
	wire [4-1:0] node160;
	wire [4-1:0] node161;
	wire [4-1:0] node164;
	wire [4-1:0] node168;
	wire [4-1:0] node169;
	wire [4-1:0] node172;
	wire [4-1:0] node174;
	wire [4-1:0] node175;
	wire [4-1:0] node178;
	wire [4-1:0] node181;
	wire [4-1:0] node182;
	wire [4-1:0] node183;
	wire [4-1:0] node184;
	wire [4-1:0] node187;
	wire [4-1:0] node190;
	wire [4-1:0] node191;
	wire [4-1:0] node194;
	wire [4-1:0] node197;
	wire [4-1:0] node198;
	wire [4-1:0] node199;
	wire [4-1:0] node201;
	wire [4-1:0] node205;
	wire [4-1:0] node206;
	wire [4-1:0] node207;
	wire [4-1:0] node210;
	wire [4-1:0] node214;
	wire [4-1:0] node215;
	wire [4-1:0] node216;
	wire [4-1:0] node217;
	wire [4-1:0] node218;
	wire [4-1:0] node222;
	wire [4-1:0] node224;
	wire [4-1:0] node227;
	wire [4-1:0] node228;
	wire [4-1:0] node230;
	wire [4-1:0] node231;
	wire [4-1:0] node235;
	wire [4-1:0] node236;
	wire [4-1:0] node240;
	wire [4-1:0] node241;
	wire [4-1:0] node242;
	wire [4-1:0] node243;
	wire [4-1:0] node245;
	wire [4-1:0] node249;
	wire [4-1:0] node251;
	wire [4-1:0] node252;
	wire [4-1:0] node256;
	wire [4-1:0] node257;
	wire [4-1:0] node258;
	wire [4-1:0] node261;
	wire [4-1:0] node264;
	wire [4-1:0] node265;
	wire [4-1:0] node266;
	wire [4-1:0] node270;
	wire [4-1:0] node272;
	wire [4-1:0] node275;
	wire [4-1:0] node276;
	wire [4-1:0] node277;
	wire [4-1:0] node278;
	wire [4-1:0] node279;
	wire [4-1:0] node280;
	wire [4-1:0] node283;
	wire [4-1:0] node287;
	wire [4-1:0] node288;
	wire [4-1:0] node289;
	wire [4-1:0] node290;
	wire [4-1:0] node293;
	wire [4-1:0] node296;
	wire [4-1:0] node298;
	wire [4-1:0] node301;
	wire [4-1:0] node303;
	wire [4-1:0] node306;
	wire [4-1:0] node307;
	wire [4-1:0] node308;
	wire [4-1:0] node309;
	wire [4-1:0] node311;
	wire [4-1:0] node314;
	wire [4-1:0] node315;
	wire [4-1:0] node319;
	wire [4-1:0] node320;
	wire [4-1:0] node323;
	wire [4-1:0] node326;
	wire [4-1:0] node329;
	wire [4-1:0] node330;
	wire [4-1:0] node331;
	wire [4-1:0] node332;
	wire [4-1:0] node333;
	wire [4-1:0] node334;
	wire [4-1:0] node337;
	wire [4-1:0] node340;
	wire [4-1:0] node343;
	wire [4-1:0] node345;
	wire [4-1:0] node347;
	wire [4-1:0] node350;
	wire [4-1:0] node351;
	wire [4-1:0] node354;
	wire [4-1:0] node357;
	wire [4-1:0] node358;
	wire [4-1:0] node359;
	wire [4-1:0] node360;
	wire [4-1:0] node363;
	wire [4-1:0] node367;
	wire [4-1:0] node368;
	wire [4-1:0] node369;
	wire [4-1:0] node370;
	wire [4-1:0] node374;
	wire [4-1:0] node376;
	wire [4-1:0] node379;
	wire [4-1:0] node381;
	wire [4-1:0] node383;
	wire [4-1:0] node386;
	wire [4-1:0] node387;
	wire [4-1:0] node388;
	wire [4-1:0] node389;
	wire [4-1:0] node390;
	wire [4-1:0] node391;
	wire [4-1:0] node392;
	wire [4-1:0] node395;
	wire [4-1:0] node396;
	wire [4-1:0] node400;
	wire [4-1:0] node401;
	wire [4-1:0] node402;
	wire [4-1:0] node403;
	wire [4-1:0] node406;
	wire [4-1:0] node409;
	wire [4-1:0] node412;
	wire [4-1:0] node413;
	wire [4-1:0] node414;
	wire [4-1:0] node418;
	wire [4-1:0] node419;
	wire [4-1:0] node423;
	wire [4-1:0] node424;
	wire [4-1:0] node425;
	wire [4-1:0] node428;
	wire [4-1:0] node430;
	wire [4-1:0] node433;
	wire [4-1:0] node434;
	wire [4-1:0] node435;
	wire [4-1:0] node436;
	wire [4-1:0] node440;
	wire [4-1:0] node441;
	wire [4-1:0] node444;
	wire [4-1:0] node447;
	wire [4-1:0] node448;
	wire [4-1:0] node452;
	wire [4-1:0] node453;
	wire [4-1:0] node454;
	wire [4-1:0] node455;
	wire [4-1:0] node457;
	wire [4-1:0] node460;
	wire [4-1:0] node461;
	wire [4-1:0] node464;
	wire [4-1:0] node466;
	wire [4-1:0] node469;
	wire [4-1:0] node470;
	wire [4-1:0] node472;
	wire [4-1:0] node473;
	wire [4-1:0] node478;
	wire [4-1:0] node479;
	wire [4-1:0] node480;
	wire [4-1:0] node481;
	wire [4-1:0] node482;
	wire [4-1:0] node485;
	wire [4-1:0] node489;
	wire [4-1:0] node491;
	wire [4-1:0] node494;
	wire [4-1:0] node495;
	wire [4-1:0] node498;
	wire [4-1:0] node500;
	wire [4-1:0] node501;
	wire [4-1:0] node504;
	wire [4-1:0] node507;
	wire [4-1:0] node508;
	wire [4-1:0] node509;
	wire [4-1:0] node510;
	wire [4-1:0] node513;
	wire [4-1:0] node514;
	wire [4-1:0] node515;
	wire [4-1:0] node518;
	wire [4-1:0] node521;
	wire [4-1:0] node522;
	wire [4-1:0] node523;
	wire [4-1:0] node528;
	wire [4-1:0] node529;
	wire [4-1:0] node530;
	wire [4-1:0] node531;
	wire [4-1:0] node534;
	wire [4-1:0] node537;
	wire [4-1:0] node539;
	wire [4-1:0] node542;
	wire [4-1:0] node543;
	wire [4-1:0] node546;
	wire [4-1:0] node547;
	wire [4-1:0] node551;
	wire [4-1:0] node552;
	wire [4-1:0] node553;
	wire [4-1:0] node554;
	wire [4-1:0] node555;
	wire [4-1:0] node558;
	wire [4-1:0] node561;
	wire [4-1:0] node564;
	wire [4-1:0] node565;
	wire [4-1:0] node568;
	wire [4-1:0] node569;
	wire [4-1:0] node572;
	wire [4-1:0] node573;
	wire [4-1:0] node576;
	wire [4-1:0] node579;
	wire [4-1:0] node580;
	wire [4-1:0] node581;
	wire [4-1:0] node582;
	wire [4-1:0] node583;
	wire [4-1:0] node586;
	wire [4-1:0] node590;
	wire [4-1:0] node592;
	wire [4-1:0] node593;
	wire [4-1:0] node596;
	wire [4-1:0] node599;
	wire [4-1:0] node600;
	wire [4-1:0] node603;
	wire [4-1:0] node605;
	wire [4-1:0] node607;
	wire [4-1:0] node610;
	wire [4-1:0] node611;
	wire [4-1:0] node612;
	wire [4-1:0] node613;
	wire [4-1:0] node614;
	wire [4-1:0] node615;
	wire [4-1:0] node617;
	wire [4-1:0] node620;
	wire [4-1:0] node621;
	wire [4-1:0] node625;
	wire [4-1:0] node626;
	wire [4-1:0] node628;
	wire [4-1:0] node631;
	wire [4-1:0] node632;
	wire [4-1:0] node636;
	wire [4-1:0] node637;
	wire [4-1:0] node638;
	wire [4-1:0] node639;
	wire [4-1:0] node644;
	wire [4-1:0] node646;
	wire [4-1:0] node648;
	wire [4-1:0] node649;
	wire [4-1:0] node653;
	wire [4-1:0] node654;
	wire [4-1:0] node655;
	wire [4-1:0] node656;
	wire [4-1:0] node659;
	wire [4-1:0] node660;
	wire [4-1:0] node663;
	wire [4-1:0] node666;
	wire [4-1:0] node667;
	wire [4-1:0] node669;
	wire [4-1:0] node672;
	wire [4-1:0] node675;
	wire [4-1:0] node676;
	wire [4-1:0] node678;
	wire [4-1:0] node679;
	wire [4-1:0] node680;
	wire [4-1:0] node683;
	wire [4-1:0] node687;
	wire [4-1:0] node688;
	wire [4-1:0] node691;
	wire [4-1:0] node693;
	wire [4-1:0] node696;
	wire [4-1:0] node697;
	wire [4-1:0] node698;
	wire [4-1:0] node699;
	wire [4-1:0] node700;
	wire [4-1:0] node701;
	wire [4-1:0] node704;
	wire [4-1:0] node707;
	wire [4-1:0] node708;
	wire [4-1:0] node712;
	wire [4-1:0] node714;
	wire [4-1:0] node715;
	wire [4-1:0] node718;
	wire [4-1:0] node721;
	wire [4-1:0] node722;
	wire [4-1:0] node723;
	wire [4-1:0] node724;
	wire [4-1:0] node727;
	wire [4-1:0] node730;
	wire [4-1:0] node732;
	wire [4-1:0] node735;
	wire [4-1:0] node736;
	wire [4-1:0] node737;
	wire [4-1:0] node740;
	wire [4-1:0] node743;
	wire [4-1:0] node746;
	wire [4-1:0] node747;
	wire [4-1:0] node748;
	wire [4-1:0] node749;
	wire [4-1:0] node753;
	wire [4-1:0] node755;
	wire [4-1:0] node757;
	wire [4-1:0] node760;
	wire [4-1:0] node761;
	wire [4-1:0] node762;
	wire [4-1:0] node765;
	wire [4-1:0] node767;
	wire [4-1:0] node770;
	wire [4-1:0] node771;
	wire [4-1:0] node773;
	wire [4-1:0] node776;
	wire [4-1:0] node779;
	wire [4-1:0] node780;
	wire [4-1:0] node781;
	wire [4-1:0] node782;
	wire [4-1:0] node783;
	wire [4-1:0] node784;
	wire [4-1:0] node785;
	wire [4-1:0] node786;
	wire [4-1:0] node791;
	wire [4-1:0] node792;
	wire [4-1:0] node793;
	wire [4-1:0] node796;
	wire [4-1:0] node799;
	wire [4-1:0] node800;
	wire [4-1:0] node801;
	wire [4-1:0] node802;
	wire [4-1:0] node805;
	wire [4-1:0] node808;
	wire [4-1:0] node811;
	wire [4-1:0] node812;
	wire [4-1:0] node816;
	wire [4-1:0] node817;
	wire [4-1:0] node818;
	wire [4-1:0] node819;
	wire [4-1:0] node820;
	wire [4-1:0] node823;
	wire [4-1:0] node827;
	wire [4-1:0] node828;
	wire [4-1:0] node830;
	wire [4-1:0] node831;
	wire [4-1:0] node834;
	wire [4-1:0] node837;
	wire [4-1:0] node840;
	wire [4-1:0] node841;
	wire [4-1:0] node842;
	wire [4-1:0] node844;
	wire [4-1:0] node845;
	wire [4-1:0] node848;
	wire [4-1:0] node851;
	wire [4-1:0] node852;
	wire [4-1:0] node853;
	wire [4-1:0] node856;
	wire [4-1:0] node860;
	wire [4-1:0] node861;
	wire [4-1:0] node862;
	wire [4-1:0] node866;
	wire [4-1:0] node867;
	wire [4-1:0] node869;
	wire [4-1:0] node872;
	wire [4-1:0] node873;
	wire [4-1:0] node877;
	wire [4-1:0] node878;
	wire [4-1:0] node879;
	wire [4-1:0] node880;
	wire [4-1:0] node881;
	wire [4-1:0] node882;
	wire [4-1:0] node883;
	wire [4-1:0] node887;
	wire [4-1:0] node890;
	wire [4-1:0] node891;
	wire [4-1:0] node895;
	wire [4-1:0] node896;
	wire [4-1:0] node898;
	wire [4-1:0] node899;
	wire [4-1:0] node902;
	wire [4-1:0] node905;
	wire [4-1:0] node908;
	wire [4-1:0] node909;
	wire [4-1:0] node910;
	wire [4-1:0] node911;
	wire [4-1:0] node914;
	wire [4-1:0] node918;
	wire [4-1:0] node919;
	wire [4-1:0] node920;
	wire [4-1:0] node924;
	wire [4-1:0] node927;
	wire [4-1:0] node928;
	wire [4-1:0] node929;
	wire [4-1:0] node930;
	wire [4-1:0] node931;
	wire [4-1:0] node932;
	wire [4-1:0] node938;
	wire [4-1:0] node939;
	wire [4-1:0] node940;
	wire [4-1:0] node942;
	wire [4-1:0] node946;
	wire [4-1:0] node947;
	wire [4-1:0] node948;
	wire [4-1:0] node953;
	wire [4-1:0] node954;
	wire [4-1:0] node955;
	wire [4-1:0] node956;
	wire [4-1:0] node959;
	wire [4-1:0] node963;
	wire [4-1:0] node965;
	wire [4-1:0] node966;
	wire [4-1:0] node969;
	wire [4-1:0] node971;
	wire [4-1:0] node974;
	wire [4-1:0] node975;
	wire [4-1:0] node976;
	wire [4-1:0] node977;
	wire [4-1:0] node978;
	wire [4-1:0] node979;
	wire [4-1:0] node983;
	wire [4-1:0] node985;
	wire [4-1:0] node986;
	wire [4-1:0] node990;
	wire [4-1:0] node991;
	wire [4-1:0] node992;
	wire [4-1:0] node993;
	wire [4-1:0] node997;
	wire [4-1:0] node998;
	wire [4-1:0] node1001;
	wire [4-1:0] node1004;
	wire [4-1:0] node1005;
	wire [4-1:0] node1006;
	wire [4-1:0] node1007;
	wire [4-1:0] node1010;
	wire [4-1:0] node1014;
	wire [4-1:0] node1015;
	wire [4-1:0] node1016;
	wire [4-1:0] node1021;
	wire [4-1:0] node1022;
	wire [4-1:0] node1023;
	wire [4-1:0] node1024;
	wire [4-1:0] node1026;
	wire [4-1:0] node1027;
	wire [4-1:0] node1031;
	wire [4-1:0] node1034;
	wire [4-1:0] node1035;
	wire [4-1:0] node1036;
	wire [4-1:0] node1040;
	wire [4-1:0] node1042;
	wire [4-1:0] node1045;
	wire [4-1:0] node1046;
	wire [4-1:0] node1047;
	wire [4-1:0] node1049;
	wire [4-1:0] node1052;
	wire [4-1:0] node1053;
	wire [4-1:0] node1056;
	wire [4-1:0] node1059;
	wire [4-1:0] node1060;
	wire [4-1:0] node1061;
	wire [4-1:0] node1062;
	wire [4-1:0] node1067;
	wire [4-1:0] node1070;
	wire [4-1:0] node1071;
	wire [4-1:0] node1072;
	wire [4-1:0] node1073;
	wire [4-1:0] node1076;
	wire [4-1:0] node1077;
	wire [4-1:0] node1079;
	wire [4-1:0] node1082;
	wire [4-1:0] node1083;
	wire [4-1:0] node1084;
	wire [4-1:0] node1087;
	wire [4-1:0] node1091;
	wire [4-1:0] node1092;
	wire [4-1:0] node1093;
	wire [4-1:0] node1094;
	wire [4-1:0] node1099;
	wire [4-1:0] node1101;
	wire [4-1:0] node1102;
	wire [4-1:0] node1105;
	wire [4-1:0] node1107;
	wire [4-1:0] node1110;
	wire [4-1:0] node1111;
	wire [4-1:0] node1112;
	wire [4-1:0] node1113;
	wire [4-1:0] node1117;
	wire [4-1:0] node1119;
	wire [4-1:0] node1121;
	wire [4-1:0] node1123;
	wire [4-1:0] node1126;
	wire [4-1:0] node1127;
	wire [4-1:0] node1128;
	wire [4-1:0] node1130;
	wire [4-1:0] node1133;
	wire [4-1:0] node1134;
	wire [4-1:0] node1138;
	wire [4-1:0] node1139;
	wire [4-1:0] node1140;
	wire [4-1:0] node1142;
	wire [4-1:0] node1145;
	wire [4-1:0] node1146;
	wire [4-1:0] node1149;
	wire [4-1:0] node1152;
	wire [4-1:0] node1154;
	wire [4-1:0] node1157;
	wire [4-1:0] node1158;
	wire [4-1:0] node1159;
	wire [4-1:0] node1160;
	wire [4-1:0] node1161;
	wire [4-1:0] node1162;
	wire [4-1:0] node1163;
	wire [4-1:0] node1165;
	wire [4-1:0] node1167;
	wire [4-1:0] node1171;
	wire [4-1:0] node1172;
	wire [4-1:0] node1173;
	wire [4-1:0] node1175;
	wire [4-1:0] node1178;
	wire [4-1:0] node1179;
	wire [4-1:0] node1183;
	wire [4-1:0] node1185;
	wire [4-1:0] node1188;
	wire [4-1:0] node1189;
	wire [4-1:0] node1190;
	wire [4-1:0] node1191;
	wire [4-1:0] node1195;
	wire [4-1:0] node1196;
	wire [4-1:0] node1200;
	wire [4-1:0] node1201;
	wire [4-1:0] node1204;
	wire [4-1:0] node1207;
	wire [4-1:0] node1208;
	wire [4-1:0] node1209;
	wire [4-1:0] node1210;
	wire [4-1:0] node1213;
	wire [4-1:0] node1216;
	wire [4-1:0] node1218;
	wire [4-1:0] node1221;
	wire [4-1:0] node1222;
	wire [4-1:0] node1223;
	wire [4-1:0] node1226;
	wire [4-1:0] node1229;
	wire [4-1:0] node1230;
	wire [4-1:0] node1233;
	wire [4-1:0] node1236;
	wire [4-1:0] node1237;
	wire [4-1:0] node1238;
	wire [4-1:0] node1239;
	wire [4-1:0] node1241;
	wire [4-1:0] node1243;
	wire [4-1:0] node1246;
	wire [4-1:0] node1247;
	wire [4-1:0] node1250;
	wire [4-1:0] node1253;
	wire [4-1:0] node1254;
	wire [4-1:0] node1255;
	wire [4-1:0] node1257;
	wire [4-1:0] node1259;
	wire [4-1:0] node1264;
	wire [4-1:0] node1265;
	wire [4-1:0] node1266;
	wire [4-1:0] node1267;
	wire [4-1:0] node1268;
	wire [4-1:0] node1271;
	wire [4-1:0] node1275;
	wire [4-1:0] node1276;
	wire [4-1:0] node1278;
	wire [4-1:0] node1279;
	wire [4-1:0] node1282;
	wire [4-1:0] node1285;
	wire [4-1:0] node1286;
	wire [4-1:0] node1289;
	wire [4-1:0] node1292;
	wire [4-1:0] node1293;
	wire [4-1:0] node1294;
	wire [4-1:0] node1295;
	wire [4-1:0] node1296;
	wire [4-1:0] node1300;
	wire [4-1:0] node1302;
	wire [4-1:0] node1305;
	wire [4-1:0] node1306;
	wire [4-1:0] node1309;
	wire [4-1:0] node1312;
	wire [4-1:0] node1313;
	wire [4-1:0] node1314;
	wire [4-1:0] node1318;
	wire [4-1:0] node1319;
	wire [4-1:0] node1322;
	wire [4-1:0] node1325;
	wire [4-1:0] node1326;
	wire [4-1:0] node1327;
	wire [4-1:0] node1328;
	wire [4-1:0] node1329;
	wire [4-1:0] node1330;
	wire [4-1:0] node1331;
	wire [4-1:0] node1332;
	wire [4-1:0] node1337;
	wire [4-1:0] node1338;
	wire [4-1:0] node1339;
	wire [4-1:0] node1342;
	wire [4-1:0] node1346;
	wire [4-1:0] node1347;
	wire [4-1:0] node1348;
	wire [4-1:0] node1349;
	wire [4-1:0] node1353;
	wire [4-1:0] node1356;
	wire [4-1:0] node1359;
	wire [4-1:0] node1360;
	wire [4-1:0] node1361;
	wire [4-1:0] node1362;
	wire [4-1:0] node1364;
	wire [4-1:0] node1367;
	wire [4-1:0] node1368;
	wire [4-1:0] node1372;
	wire [4-1:0] node1374;
	wire [4-1:0] node1375;
	wire [4-1:0] node1378;
	wire [4-1:0] node1381;
	wire [4-1:0] node1382;
	wire [4-1:0] node1385;
	wire [4-1:0] node1387;
	wire [4-1:0] node1389;
	wire [4-1:0] node1392;
	wire [4-1:0] node1393;
	wire [4-1:0] node1394;
	wire [4-1:0] node1397;
	wire [4-1:0] node1398;
	wire [4-1:0] node1401;
	wire [4-1:0] node1402;
	wire [4-1:0] node1403;
	wire [4-1:0] node1407;
	wire [4-1:0] node1409;
	wire [4-1:0] node1412;
	wire [4-1:0] node1413;
	wire [4-1:0] node1414;
	wire [4-1:0] node1417;
	wire [4-1:0] node1418;
	wire [4-1:0] node1420;
	wire [4-1:0] node1424;
	wire [4-1:0] node1425;
	wire [4-1:0] node1427;
	wire [4-1:0] node1428;
	wire [4-1:0] node1432;
	wire [4-1:0] node1433;
	wire [4-1:0] node1435;
	wire [4-1:0] node1438;
	wire [4-1:0] node1440;
	wire [4-1:0] node1443;
	wire [4-1:0] node1444;
	wire [4-1:0] node1445;
	wire [4-1:0] node1446;
	wire [4-1:0] node1447;
	wire [4-1:0] node1451;
	wire [4-1:0] node1452;
	wire [4-1:0] node1454;
	wire [4-1:0] node1455;
	wire [4-1:0] node1458;
	wire [4-1:0] node1461;
	wire [4-1:0] node1464;
	wire [4-1:0] node1465;
	wire [4-1:0] node1466;
	wire [4-1:0] node1467;
	wire [4-1:0] node1468;
	wire [4-1:0] node1472;
	wire [4-1:0] node1475;
	wire [4-1:0] node1478;
	wire [4-1:0] node1479;
	wire [4-1:0] node1482;
	wire [4-1:0] node1483;
	wire [4-1:0] node1487;
	wire [4-1:0] node1488;
	wire [4-1:0] node1489;
	wire [4-1:0] node1490;
	wire [4-1:0] node1491;
	wire [4-1:0] node1495;
	wire [4-1:0] node1496;
	wire [4-1:0] node1497;
	wire [4-1:0] node1500;
	wire [4-1:0] node1504;
	wire [4-1:0] node1505;
	wire [4-1:0] node1506;
	wire [4-1:0] node1510;
	wire [4-1:0] node1513;
	wire [4-1:0] node1514;
	wire [4-1:0] node1515;
	wire [4-1:0] node1516;
	wire [4-1:0] node1517;
	wire [4-1:0] node1521;
	wire [4-1:0] node1523;
	wire [4-1:0] node1526;
	wire [4-1:0] node1527;
	wire [4-1:0] node1528;
	wire [4-1:0] node1533;
	wire [4-1:0] node1535;
	wire [4-1:0] node1536;
	wire [4-1:0] node1539;
	wire [4-1:0] node1542;
	wire [4-1:0] node1543;
	wire [4-1:0] node1544;
	wire [4-1:0] node1545;
	wire [4-1:0] node1546;
	wire [4-1:0] node1547;
	wire [4-1:0] node1548;
	wire [4-1:0] node1549;
	wire [4-1:0] node1551;
	wire [4-1:0] node1554;
	wire [4-1:0] node1556;
	wire [4-1:0] node1559;
	wire [4-1:0] node1560;
	wire [4-1:0] node1562;
	wire [4-1:0] node1565;
	wire [4-1:0] node1566;
	wire [4-1:0] node1568;
	wire [4-1:0] node1571;
	wire [4-1:0] node1574;
	wire [4-1:0] node1575;
	wire [4-1:0] node1576;
	wire [4-1:0] node1577;
	wire [4-1:0] node1578;
	wire [4-1:0] node1579;
	wire [4-1:0] node1582;
	wire [4-1:0] node1585;
	wire [4-1:0] node1586;
	wire [4-1:0] node1589;
	wire [4-1:0] node1592;
	wire [4-1:0] node1593;
	wire [4-1:0] node1595;
	wire [4-1:0] node1598;
	wire [4-1:0] node1601;
	wire [4-1:0] node1603;
	wire [4-1:0] node1605;
	wire [4-1:0] node1608;
	wire [4-1:0] node1609;
	wire [4-1:0] node1612;
	wire [4-1:0] node1614;
	wire [4-1:0] node1616;
	wire [4-1:0] node1619;
	wire [4-1:0] node1620;
	wire [4-1:0] node1621;
	wire [4-1:0] node1622;
	wire [4-1:0] node1623;
	wire [4-1:0] node1626;
	wire [4-1:0] node1628;
	wire [4-1:0] node1631;
	wire [4-1:0] node1633;
	wire [4-1:0] node1635;
	wire [4-1:0] node1638;
	wire [4-1:0] node1639;
	wire [4-1:0] node1640;
	wire [4-1:0] node1644;
	wire [4-1:0] node1645;
	wire [4-1:0] node1646;
	wire [4-1:0] node1647;
	wire [4-1:0] node1652;
	wire [4-1:0] node1653;
	wire [4-1:0] node1656;
	wire [4-1:0] node1659;
	wire [4-1:0] node1660;
	wire [4-1:0] node1661;
	wire [4-1:0] node1662;
	wire [4-1:0] node1666;
	wire [4-1:0] node1667;
	wire [4-1:0] node1669;
	wire [4-1:0] node1670;
	wire [4-1:0] node1674;
	wire [4-1:0] node1675;
	wire [4-1:0] node1679;
	wire [4-1:0] node1680;
	wire [4-1:0] node1682;
	wire [4-1:0] node1683;
	wire [4-1:0] node1686;
	wire [4-1:0] node1689;
	wire [4-1:0] node1690;
	wire [4-1:0] node1692;
	wire [4-1:0] node1696;
	wire [4-1:0] node1697;
	wire [4-1:0] node1698;
	wire [4-1:0] node1699;
	wire [4-1:0] node1700;
	wire [4-1:0] node1702;
	wire [4-1:0] node1704;
	wire [4-1:0] node1705;
	wire [4-1:0] node1708;
	wire [4-1:0] node1711;
	wire [4-1:0] node1712;
	wire [4-1:0] node1713;
	wire [4-1:0] node1716;
	wire [4-1:0] node1719;
	wire [4-1:0] node1721;
	wire [4-1:0] node1724;
	wire [4-1:0] node1725;
	wire [4-1:0] node1726;
	wire [4-1:0] node1729;
	wire [4-1:0] node1731;
	wire [4-1:0] node1733;
	wire [4-1:0] node1736;
	wire [4-1:0] node1737;
	wire [4-1:0] node1738;
	wire [4-1:0] node1741;
	wire [4-1:0] node1744;
	wire [4-1:0] node1746;
	wire [4-1:0] node1749;
	wire [4-1:0] node1750;
	wire [4-1:0] node1751;
	wire [4-1:0] node1752;
	wire [4-1:0] node1754;
	wire [4-1:0] node1756;
	wire [4-1:0] node1759;
	wire [4-1:0] node1760;
	wire [4-1:0] node1763;
	wire [4-1:0] node1766;
	wire [4-1:0] node1768;
	wire [4-1:0] node1771;
	wire [4-1:0] node1772;
	wire [4-1:0] node1773;
	wire [4-1:0] node1774;
	wire [4-1:0] node1777;
	wire [4-1:0] node1781;
	wire [4-1:0] node1782;
	wire [4-1:0] node1783;
	wire [4-1:0] node1784;
	wire [4-1:0] node1790;
	wire [4-1:0] node1791;
	wire [4-1:0] node1792;
	wire [4-1:0] node1793;
	wire [4-1:0] node1796;
	wire [4-1:0] node1799;
	wire [4-1:0] node1800;
	wire [4-1:0] node1802;
	wire [4-1:0] node1803;
	wire [4-1:0] node1806;
	wire [4-1:0] node1808;
	wire [4-1:0] node1811;
	wire [4-1:0] node1812;
	wire [4-1:0] node1813;
	wire [4-1:0] node1815;
	wire [4-1:0] node1818;
	wire [4-1:0] node1820;
	wire [4-1:0] node1823;
	wire [4-1:0] node1825;
	wire [4-1:0] node1826;
	wire [4-1:0] node1830;
	wire [4-1:0] node1831;
	wire [4-1:0] node1832;
	wire [4-1:0] node1833;
	wire [4-1:0] node1834;
	wire [4-1:0] node1837;
	wire [4-1:0] node1840;
	wire [4-1:0] node1841;
	wire [4-1:0] node1845;
	wire [4-1:0] node1846;
	wire [4-1:0] node1849;
	wire [4-1:0] node1852;
	wire [4-1:0] node1853;
	wire [4-1:0] node1855;
	wire [4-1:0] node1857;
	wire [4-1:0] node1859;
	wire [4-1:0] node1862;
	wire [4-1:0] node1863;
	wire [4-1:0] node1864;
	wire [4-1:0] node1868;
	wire [4-1:0] node1870;
	wire [4-1:0] node1871;
	wire [4-1:0] node1875;
	wire [4-1:0] node1876;
	wire [4-1:0] node1877;
	wire [4-1:0] node1878;
	wire [4-1:0] node1879;
	wire [4-1:0] node1880;
	wire [4-1:0] node1881;
	wire [4-1:0] node1883;
	wire [4-1:0] node1886;
	wire [4-1:0] node1888;
	wire [4-1:0] node1891;
	wire [4-1:0] node1892;
	wire [4-1:0] node1893;
	wire [4-1:0] node1898;
	wire [4-1:0] node1899;
	wire [4-1:0] node1900;
	wire [4-1:0] node1902;
	wire [4-1:0] node1906;
	wire [4-1:0] node1907;
	wire [4-1:0] node1908;
	wire [4-1:0] node1912;
	wire [4-1:0] node1914;
	wire [4-1:0] node1917;
	wire [4-1:0] node1918;
	wire [4-1:0] node1919;
	wire [4-1:0] node1921;
	wire [4-1:0] node1924;
	wire [4-1:0] node1926;
	wire [4-1:0] node1927;
	wire [4-1:0] node1930;
	wire [4-1:0] node1933;
	wire [4-1:0] node1934;
	wire [4-1:0] node1935;
	wire [4-1:0] node1938;
	wire [4-1:0] node1941;
	wire [4-1:0] node1942;
	wire [4-1:0] node1944;
	wire [4-1:0] node1947;
	wire [4-1:0] node1950;
	wire [4-1:0] node1951;
	wire [4-1:0] node1952;
	wire [4-1:0] node1953;
	wire [4-1:0] node1954;
	wire [4-1:0] node1957;
	wire [4-1:0] node1958;
	wire [4-1:0] node1961;
	wire [4-1:0] node1964;
	wire [4-1:0] node1965;
	wire [4-1:0] node1968;
	wire [4-1:0] node1970;
	wire [4-1:0] node1973;
	wire [4-1:0] node1974;
	wire [4-1:0] node1975;
	wire [4-1:0] node1977;
	wire [4-1:0] node1979;
	wire [4-1:0] node1982;
	wire [4-1:0] node1984;
	wire [4-1:0] node1987;
	wire [4-1:0] node1989;
	wire [4-1:0] node1992;
	wire [4-1:0] node1993;
	wire [4-1:0] node1994;
	wire [4-1:0] node1995;
	wire [4-1:0] node1998;
	wire [4-1:0] node2001;
	wire [4-1:0] node2002;
	wire [4-1:0] node2004;
	wire [4-1:0] node2008;
	wire [4-1:0] node2009;
	wire [4-1:0] node2010;
	wire [4-1:0] node2011;
	wire [4-1:0] node2016;
	wire [4-1:0] node2018;
	wire [4-1:0] node2020;
	wire [4-1:0] node2023;
	wire [4-1:0] node2024;
	wire [4-1:0] node2025;
	wire [4-1:0] node2026;
	wire [4-1:0] node2027;
	wire [4-1:0] node2028;
	wire [4-1:0] node2029;
	wire [4-1:0] node2033;
	wire [4-1:0] node2036;
	wire [4-1:0] node2038;
	wire [4-1:0] node2040;
	wire [4-1:0] node2043;
	wire [4-1:0] node2044;
	wire [4-1:0] node2045;
	wire [4-1:0] node2046;
	wire [4-1:0] node2049;
	wire [4-1:0] node2050;
	wire [4-1:0] node2054;
	wire [4-1:0] node2055;
	wire [4-1:0] node2057;
	wire [4-1:0] node2060;
	wire [4-1:0] node2061;
	wire [4-1:0] node2065;
	wire [4-1:0] node2066;
	wire [4-1:0] node2067;
	wire [4-1:0] node2068;
	wire [4-1:0] node2073;
	wire [4-1:0] node2076;
	wire [4-1:0] node2077;
	wire [4-1:0] node2078;
	wire [4-1:0] node2079;
	wire [4-1:0] node2082;
	wire [4-1:0] node2085;
	wire [4-1:0] node2086;
	wire [4-1:0] node2087;
	wire [4-1:0] node2088;
	wire [4-1:0] node2093;
	wire [4-1:0] node2094;
	wire [4-1:0] node2095;
	wire [4-1:0] node2100;
	wire [4-1:0] node2101;
	wire [4-1:0] node2102;
	wire [4-1:0] node2105;
	wire [4-1:0] node2106;
	wire [4-1:0] node2109;
	wire [4-1:0] node2112;
	wire [4-1:0] node2113;
	wire [4-1:0] node2115;
	wire [4-1:0] node2116;
	wire [4-1:0] node2120;
	wire [4-1:0] node2121;
	wire [4-1:0] node2124;
	wire [4-1:0] node2127;
	wire [4-1:0] node2128;
	wire [4-1:0] node2129;
	wire [4-1:0] node2130;
	wire [4-1:0] node2131;
	wire [4-1:0] node2134;
	wire [4-1:0] node2135;
	wire [4-1:0] node2138;
	wire [4-1:0] node2141;
	wire [4-1:0] node2142;
	wire [4-1:0] node2143;
	wire [4-1:0] node2146;
	wire [4-1:0] node2149;
	wire [4-1:0] node2150;
	wire [4-1:0] node2152;
	wire [4-1:0] node2155;
	wire [4-1:0] node2156;
	wire [4-1:0] node2160;
	wire [4-1:0] node2161;
	wire [4-1:0] node2162;
	wire [4-1:0] node2165;
	wire [4-1:0] node2166;
	wire [4-1:0] node2168;
	wire [4-1:0] node2171;
	wire [4-1:0] node2174;
	wire [4-1:0] node2175;
	wire [4-1:0] node2178;
	wire [4-1:0] node2181;
	wire [4-1:0] node2182;
	wire [4-1:0] node2183;
	wire [4-1:0] node2184;
	wire [4-1:0] node2185;
	wire [4-1:0] node2188;
	wire [4-1:0] node2191;
	wire [4-1:0] node2193;
	wire [4-1:0] node2194;
	wire [4-1:0] node2197;
	wire [4-1:0] node2200;
	wire [4-1:0] node2201;
	wire [4-1:0] node2202;
	wire [4-1:0] node2205;
	wire [4-1:0] node2209;
	wire [4-1:0] node2210;
	wire [4-1:0] node2211;
	wire [4-1:0] node2214;
	wire [4-1:0] node2216;
	wire [4-1:0] node2219;
	wire [4-1:0] node2220;
	wire [4-1:0] node2221;
	wire [4-1:0] node2226;
	wire [4-1:0] node2227;
	wire [4-1:0] node2228;
	wire [4-1:0] node2229;
	wire [4-1:0] node2230;
	wire [4-1:0] node2231;
	wire [4-1:0] node2232;
	wire [4-1:0] node2234;
	wire [4-1:0] node2235;
	wire [4-1:0] node2238;
	wire [4-1:0] node2241;
	wire [4-1:0] node2243;
	wire [4-1:0] node2246;
	wire [4-1:0] node2247;
	wire [4-1:0] node2248;
	wire [4-1:0] node2250;
	wire [4-1:0] node2253;
	wire [4-1:0] node2255;
	wire [4-1:0] node2258;
	wire [4-1:0] node2260;
	wire [4-1:0] node2263;
	wire [4-1:0] node2264;
	wire [4-1:0] node2265;
	wire [4-1:0] node2266;
	wire [4-1:0] node2270;
	wire [4-1:0] node2271;
	wire [4-1:0] node2272;
	wire [4-1:0] node2276;
	wire [4-1:0] node2278;
	wire [4-1:0] node2280;
	wire [4-1:0] node2283;
	wire [4-1:0] node2284;
	wire [4-1:0] node2285;
	wire [4-1:0] node2287;
	wire [4-1:0] node2290;
	wire [4-1:0] node2292;
	wire [4-1:0] node2294;
	wire [4-1:0] node2297;
	wire [4-1:0] node2299;
	wire [4-1:0] node2301;
	wire [4-1:0] node2304;
	wire [4-1:0] node2305;
	wire [4-1:0] node2306;
	wire [4-1:0] node2307;
	wire [4-1:0] node2308;
	wire [4-1:0] node2311;
	wire [4-1:0] node2313;
	wire [4-1:0] node2316;
	wire [4-1:0] node2317;
	wire [4-1:0] node2318;
	wire [4-1:0] node2321;
	wire [4-1:0] node2325;
	wire [4-1:0] node2326;
	wire [4-1:0] node2327;
	wire [4-1:0] node2328;
	wire [4-1:0] node2332;
	wire [4-1:0] node2333;
	wire [4-1:0] node2335;
	wire [4-1:0] node2339;
	wire [4-1:0] node2340;
	wire [4-1:0] node2341;
	wire [4-1:0] node2343;
	wire [4-1:0] node2346;
	wire [4-1:0] node2348;
	wire [4-1:0] node2351;
	wire [4-1:0] node2354;
	wire [4-1:0] node2355;
	wire [4-1:0] node2356;
	wire [4-1:0] node2358;
	wire [4-1:0] node2359;
	wire [4-1:0] node2361;
	wire [4-1:0] node2365;
	wire [4-1:0] node2366;
	wire [4-1:0] node2367;
	wire [4-1:0] node2370;
	wire [4-1:0] node2373;
	wire [4-1:0] node2374;
	wire [4-1:0] node2377;
	wire [4-1:0] node2380;
	wire [4-1:0] node2381;
	wire [4-1:0] node2382;
	wire [4-1:0] node2383;
	wire [4-1:0] node2385;
	wire [4-1:0] node2388;
	wire [4-1:0] node2390;
	wire [4-1:0] node2393;
	wire [4-1:0] node2395;
	wire [4-1:0] node2396;
	wire [4-1:0] node2400;
	wire [4-1:0] node2401;
	wire [4-1:0] node2402;
	wire [4-1:0] node2405;
	wire [4-1:0] node2407;
	wire [4-1:0] node2410;
	wire [4-1:0] node2412;
	wire [4-1:0] node2414;
	wire [4-1:0] node2417;
	wire [4-1:0] node2418;
	wire [4-1:0] node2419;
	wire [4-1:0] node2420;
	wire [4-1:0] node2421;
	wire [4-1:0] node2423;
	wire [4-1:0] node2424;
	wire [4-1:0] node2426;
	wire [4-1:0] node2429;
	wire [4-1:0] node2432;
	wire [4-1:0] node2434;
	wire [4-1:0] node2436;
	wire [4-1:0] node2439;
	wire [4-1:0] node2440;
	wire [4-1:0] node2442;
	wire [4-1:0] node2444;
	wire [4-1:0] node2447;
	wire [4-1:0] node2448;
	wire [4-1:0] node2450;
	wire [4-1:0] node2453;
	wire [4-1:0] node2456;
	wire [4-1:0] node2457;
	wire [4-1:0] node2458;
	wire [4-1:0] node2459;
	wire [4-1:0] node2461;
	wire [4-1:0] node2462;
	wire [4-1:0] node2466;
	wire [4-1:0] node2468;
	wire [4-1:0] node2471;
	wire [4-1:0] node2472;
	wire [4-1:0] node2475;
	wire [4-1:0] node2476;
	wire [4-1:0] node2477;
	wire [4-1:0] node2482;
	wire [4-1:0] node2483;
	wire [4-1:0] node2485;
	wire [4-1:0] node2486;
	wire [4-1:0] node2489;
	wire [4-1:0] node2492;
	wire [4-1:0] node2493;
	wire [4-1:0] node2496;
	wire [4-1:0] node2498;
	wire [4-1:0] node2500;
	wire [4-1:0] node2503;
	wire [4-1:0] node2504;
	wire [4-1:0] node2505;
	wire [4-1:0] node2506;
	wire [4-1:0] node2507;
	wire [4-1:0] node2510;
	wire [4-1:0] node2511;
	wire [4-1:0] node2515;
	wire [4-1:0] node2517;
	wire [4-1:0] node2518;
	wire [4-1:0] node2521;
	wire [4-1:0] node2524;
	wire [4-1:0] node2525;
	wire [4-1:0] node2526;
	wire [4-1:0] node2527;
	wire [4-1:0] node2528;
	wire [4-1:0] node2532;
	wire [4-1:0] node2533;
	wire [4-1:0] node2537;
	wire [4-1:0] node2538;
	wire [4-1:0] node2539;
	wire [4-1:0] node2542;
	wire [4-1:0] node2545;
	wire [4-1:0] node2547;
	wire [4-1:0] node2550;
	wire [4-1:0] node2551;
	wire [4-1:0] node2552;
	wire [4-1:0] node2557;
	wire [4-1:0] node2558;
	wire [4-1:0] node2559;
	wire [4-1:0] node2561;
	wire [4-1:0] node2562;
	wire [4-1:0] node2564;
	wire [4-1:0] node2568;
	wire [4-1:0] node2569;
	wire [4-1:0] node2571;
	wire [4-1:0] node2573;
	wire [4-1:0] node2576;
	wire [4-1:0] node2578;
	wire [4-1:0] node2581;
	wire [4-1:0] node2582;
	wire [4-1:0] node2583;
	wire [4-1:0] node2584;
	wire [4-1:0] node2586;
	wire [4-1:0] node2590;
	wire [4-1:0] node2592;
	wire [4-1:0] node2595;
	wire [4-1:0] node2596;
	wire [4-1:0] node2600;
	wire [4-1:0] node2601;
	wire [4-1:0] node2602;
	wire [4-1:0] node2603;
	wire [4-1:0] node2604;
	wire [4-1:0] node2605;
	wire [4-1:0] node2607;
	wire [4-1:0] node2608;
	wire [4-1:0] node2612;
	wire [4-1:0] node2613;
	wire [4-1:0] node2614;
	wire [4-1:0] node2617;
	wire [4-1:0] node2620;
	wire [4-1:0] node2621;
	wire [4-1:0] node2622;
	wire [4-1:0] node2625;
	wire [4-1:0] node2629;
	wire [4-1:0] node2630;
	wire [4-1:0] node2631;
	wire [4-1:0] node2632;
	wire [4-1:0] node2635;
	wire [4-1:0] node2638;
	wire [4-1:0] node2640;
	wire [4-1:0] node2641;
	wire [4-1:0] node2645;
	wire [4-1:0] node2646;
	wire [4-1:0] node2647;
	wire [4-1:0] node2648;
	wire [4-1:0] node2651;
	wire [4-1:0] node2654;
	wire [4-1:0] node2655;
	wire [4-1:0] node2658;
	wire [4-1:0] node2661;
	wire [4-1:0] node2662;
	wire [4-1:0] node2663;
	wire [4-1:0] node2667;
	wire [4-1:0] node2670;
	wire [4-1:0] node2671;
	wire [4-1:0] node2672;
	wire [4-1:0] node2673;
	wire [4-1:0] node2675;
	wire [4-1:0] node2676;
	wire [4-1:0] node2680;
	wire [4-1:0] node2681;
	wire [4-1:0] node2684;
	wire [4-1:0] node2687;
	wire [4-1:0] node2688;
	wire [4-1:0] node2689;
	wire [4-1:0] node2690;
	wire [4-1:0] node2693;
	wire [4-1:0] node2696;
	wire [4-1:0] node2698;
	wire [4-1:0] node2701;
	wire [4-1:0] node2702;
	wire [4-1:0] node2703;
	wire [4-1:0] node2706;
	wire [4-1:0] node2709;
	wire [4-1:0] node2712;
	wire [4-1:0] node2713;
	wire [4-1:0] node2714;
	wire [4-1:0] node2717;
	wire [4-1:0] node2718;
	wire [4-1:0] node2719;
	wire [4-1:0] node2722;
	wire [4-1:0] node2726;
	wire [4-1:0] node2727;
	wire [4-1:0] node2730;
	wire [4-1:0] node2731;
	wire [4-1:0] node2732;
	wire [4-1:0] node2737;
	wire [4-1:0] node2738;
	wire [4-1:0] node2739;
	wire [4-1:0] node2740;
	wire [4-1:0] node2741;
	wire [4-1:0] node2742;
	wire [4-1:0] node2745;
	wire [4-1:0] node2747;
	wire [4-1:0] node2750;
	wire [4-1:0] node2753;
	wire [4-1:0] node2755;
	wire [4-1:0] node2756;
	wire [4-1:0] node2760;
	wire [4-1:0] node2761;
	wire [4-1:0] node2762;
	wire [4-1:0] node2765;
	wire [4-1:0] node2766;
	wire [4-1:0] node2771;
	wire [4-1:0] node2772;
	wire [4-1:0] node2773;
	wire [4-1:0] node2775;
	wire [4-1:0] node2776;
	wire [4-1:0] node2780;
	wire [4-1:0] node2781;
	wire [4-1:0] node2783;
	wire [4-1:0] node2786;
	wire [4-1:0] node2787;
	wire [4-1:0] node2790;
	wire [4-1:0] node2793;
	wire [4-1:0] node2794;
	wire [4-1:0] node2795;
	wire [4-1:0] node2796;
	wire [4-1:0] node2799;
	wire [4-1:0] node2800;
	wire [4-1:0] node2803;
	wire [4-1:0] node2806;
	wire [4-1:0] node2809;
	wire [4-1:0] node2810;
	wire [4-1:0] node2813;
	wire [4-1:0] node2816;
	wire [4-1:0] node2817;
	wire [4-1:0] node2818;
	wire [4-1:0] node2819;
	wire [4-1:0] node2820;
	wire [4-1:0] node2821;
	wire [4-1:0] node2822;
	wire [4-1:0] node2823;
	wire [4-1:0] node2828;
	wire [4-1:0] node2829;
	wire [4-1:0] node2830;
	wire [4-1:0] node2835;
	wire [4-1:0] node2836;
	wire [4-1:0] node2837;
	wire [4-1:0] node2841;
	wire [4-1:0] node2844;
	wire [4-1:0] node2845;
	wire [4-1:0] node2847;
	wire [4-1:0] node2848;
	wire [4-1:0] node2849;
	wire [4-1:0] node2852;
	wire [4-1:0] node2856;
	wire [4-1:0] node2857;
	wire [4-1:0] node2858;
	wire [4-1:0] node2859;
	wire [4-1:0] node2863;
	wire [4-1:0] node2866;
	wire [4-1:0] node2867;
	wire [4-1:0] node2868;
	wire [4-1:0] node2872;
	wire [4-1:0] node2873;
	wire [4-1:0] node2877;
	wire [4-1:0] node2878;
	wire [4-1:0] node2879;
	wire [4-1:0] node2881;
	wire [4-1:0] node2882;
	wire [4-1:0] node2884;
	wire [4-1:0] node2888;
	wire [4-1:0] node2889;
	wire [4-1:0] node2890;
	wire [4-1:0] node2895;
	wire [4-1:0] node2896;
	wire [4-1:0] node2898;
	wire [4-1:0] node2899;
	wire [4-1:0] node2903;
	wire [4-1:0] node2904;
	wire [4-1:0] node2907;
	wire [4-1:0] node2910;
	wire [4-1:0] node2911;
	wire [4-1:0] node2912;
	wire [4-1:0] node2913;
	wire [4-1:0] node2914;
	wire [4-1:0] node2915;
	wire [4-1:0] node2919;
	wire [4-1:0] node2922;
	wire [4-1:0] node2923;
	wire [4-1:0] node2925;
	wire [4-1:0] node2928;
	wire [4-1:0] node2929;
	wire [4-1:0] node2933;
	wire [4-1:0] node2934;
	wire [4-1:0] node2935;
	wire [4-1:0] node2936;
	wire [4-1:0] node2939;
	wire [4-1:0] node2942;
	wire [4-1:0] node2945;
	wire [4-1:0] node2946;
	wire [4-1:0] node2948;
	wire [4-1:0] node2951;
	wire [4-1:0] node2953;
	wire [4-1:0] node2956;
	wire [4-1:0] node2957;
	wire [4-1:0] node2958;
	wire [4-1:0] node2960;
	wire [4-1:0] node2962;
	wire [4-1:0] node2965;
	wire [4-1:0] node2966;
	wire [4-1:0] node2967;
	wire [4-1:0] node2970;
	wire [4-1:0] node2973;
	wire [4-1:0] node2974;
	wire [4-1:0] node2978;
	wire [4-1:0] node2979;
	wire [4-1:0] node2980;
	wire [4-1:0] node2982;
	wire [4-1:0] node2984;
	wire [4-1:0] node2987;
	wire [4-1:0] node2988;
	wire [4-1:0] node2991;
	wire [4-1:0] node2994;
	wire [4-1:0] node2996;
	wire [4-1:0] node2999;
	wire [4-1:0] node3000;
	wire [4-1:0] node3001;
	wire [4-1:0] node3002;
	wire [4-1:0] node3003;
	wire [4-1:0] node3004;
	wire [4-1:0] node3005;
	wire [4-1:0] node3006;
	wire [4-1:0] node3007;
	wire [4-1:0] node3008;
	wire [4-1:0] node3009;
	wire [4-1:0] node3010;
	wire [4-1:0] node3015;
	wire [4-1:0] node3016;
	wire [4-1:0] node3020;
	wire [4-1:0] node3021;
	wire [4-1:0] node3024;
	wire [4-1:0] node3026;
	wire [4-1:0] node3029;
	wire [4-1:0] node3030;
	wire [4-1:0] node3032;
	wire [4-1:0] node3033;
	wire [4-1:0] node3034;
	wire [4-1:0] node3037;
	wire [4-1:0] node3040;
	wire [4-1:0] node3041;
	wire [4-1:0] node3044;
	wire [4-1:0] node3047;
	wire [4-1:0] node3048;
	wire [4-1:0] node3050;
	wire [4-1:0] node3053;
	wire [4-1:0] node3055;
	wire [4-1:0] node3058;
	wire [4-1:0] node3059;
	wire [4-1:0] node3060;
	wire [4-1:0] node3061;
	wire [4-1:0] node3062;
	wire [4-1:0] node3066;
	wire [4-1:0] node3068;
	wire [4-1:0] node3069;
	wire [4-1:0] node3073;
	wire [4-1:0] node3074;
	wire [4-1:0] node3075;
	wire [4-1:0] node3078;
	wire [4-1:0] node3079;
	wire [4-1:0] node3083;
	wire [4-1:0] node3084;
	wire [4-1:0] node3087;
	wire [4-1:0] node3090;
	wire [4-1:0] node3091;
	wire [4-1:0] node3092;
	wire [4-1:0] node3093;
	wire [4-1:0] node3097;
	wire [4-1:0] node3100;
	wire [4-1:0] node3101;
	wire [4-1:0] node3102;
	wire [4-1:0] node3104;
	wire [4-1:0] node3107;
	wire [4-1:0] node3110;
	wire [4-1:0] node3113;
	wire [4-1:0] node3114;
	wire [4-1:0] node3115;
	wire [4-1:0] node3116;
	wire [4-1:0] node3117;
	wire [4-1:0] node3119;
	wire [4-1:0] node3121;
	wire [4-1:0] node3124;
	wire [4-1:0] node3127;
	wire [4-1:0] node3128;
	wire [4-1:0] node3130;
	wire [4-1:0] node3131;
	wire [4-1:0] node3134;
	wire [4-1:0] node3137;
	wire [4-1:0] node3138;
	wire [4-1:0] node3140;
	wire [4-1:0] node3143;
	wire [4-1:0] node3145;
	wire [4-1:0] node3148;
	wire [4-1:0] node3149;
	wire [4-1:0] node3150;
	wire [4-1:0] node3152;
	wire [4-1:0] node3155;
	wire [4-1:0] node3157;
	wire [4-1:0] node3160;
	wire [4-1:0] node3161;
	wire [4-1:0] node3162;
	wire [4-1:0] node3165;
	wire [4-1:0] node3168;
	wire [4-1:0] node3170;
	wire [4-1:0] node3171;
	wire [4-1:0] node3174;
	wire [4-1:0] node3177;
	wire [4-1:0] node3178;
	wire [4-1:0] node3179;
	wire [4-1:0] node3180;
	wire [4-1:0] node3184;
	wire [4-1:0] node3185;
	wire [4-1:0] node3188;
	wire [4-1:0] node3191;
	wire [4-1:0] node3192;
	wire [4-1:0] node3193;
	wire [4-1:0] node3196;
	wire [4-1:0] node3197;
	wire [4-1:0] node3199;
	wire [4-1:0] node3203;
	wire [4-1:0] node3204;
	wire [4-1:0] node3205;
	wire [4-1:0] node3209;
	wire [4-1:0] node3211;
	wire [4-1:0] node3213;
	wire [4-1:0] node3216;
	wire [4-1:0] node3217;
	wire [4-1:0] node3218;
	wire [4-1:0] node3219;
	wire [4-1:0] node3220;
	wire [4-1:0] node3221;
	wire [4-1:0] node3223;
	wire [4-1:0] node3227;
	wire [4-1:0] node3229;
	wire [4-1:0] node3230;
	wire [4-1:0] node3233;
	wire [4-1:0] node3236;
	wire [4-1:0] node3237;
	wire [4-1:0] node3238;
	wire [4-1:0] node3239;
	wire [4-1:0] node3243;
	wire [4-1:0] node3244;
	wire [4-1:0] node3248;
	wire [4-1:0] node3249;
	wire [4-1:0] node3252;
	wire [4-1:0] node3253;
	wire [4-1:0] node3256;
	wire [4-1:0] node3259;
	wire [4-1:0] node3260;
	wire [4-1:0] node3261;
	wire [4-1:0] node3262;
	wire [4-1:0] node3264;
	wire [4-1:0] node3267;
	wire [4-1:0] node3268;
	wire [4-1:0] node3272;
	wire [4-1:0] node3273;
	wire [4-1:0] node3274;
	wire [4-1:0] node3277;
	wire [4-1:0] node3280;
	wire [4-1:0] node3281;
	wire [4-1:0] node3285;
	wire [4-1:0] node3286;
	wire [4-1:0] node3287;
	wire [4-1:0] node3288;
	wire [4-1:0] node3291;
	wire [4-1:0] node3294;
	wire [4-1:0] node3296;
	wire [4-1:0] node3297;
	wire [4-1:0] node3301;
	wire [4-1:0] node3302;
	wire [4-1:0] node3303;
	wire [4-1:0] node3306;
	wire [4-1:0] node3309;
	wire [4-1:0] node3311;
	wire [4-1:0] node3312;
	wire [4-1:0] node3316;
	wire [4-1:0] node3317;
	wire [4-1:0] node3318;
	wire [4-1:0] node3319;
	wire [4-1:0] node3320;
	wire [4-1:0] node3321;
	wire [4-1:0] node3322;
	wire [4-1:0] node3325;
	wire [4-1:0] node3328;
	wire [4-1:0] node3329;
	wire [4-1:0] node3333;
	wire [4-1:0] node3335;
	wire [4-1:0] node3337;
	wire [4-1:0] node3340;
	wire [4-1:0] node3341;
	wire [4-1:0] node3342;
	wire [4-1:0] node3346;
	wire [4-1:0] node3348;
	wire [4-1:0] node3349;
	wire [4-1:0] node3353;
	wire [4-1:0] node3354;
	wire [4-1:0] node3355;
	wire [4-1:0] node3356;
	wire [4-1:0] node3359;
	wire [4-1:0] node3362;
	wire [4-1:0] node3363;
	wire [4-1:0] node3365;
	wire [4-1:0] node3369;
	wire [4-1:0] node3370;
	wire [4-1:0] node3371;
	wire [4-1:0] node3374;
	wire [4-1:0] node3378;
	wire [4-1:0] node3379;
	wire [4-1:0] node3380;
	wire [4-1:0] node3381;
	wire [4-1:0] node3383;
	wire [4-1:0] node3384;
	wire [4-1:0] node3387;
	wire [4-1:0] node3390;
	wire [4-1:0] node3391;
	wire [4-1:0] node3392;
	wire [4-1:0] node3395;
	wire [4-1:0] node3398;
	wire [4-1:0] node3399;
	wire [4-1:0] node3402;
	wire [4-1:0] node3405;
	wire [4-1:0] node3406;
	wire [4-1:0] node3407;
	wire [4-1:0] node3411;
	wire [4-1:0] node3413;
	wire [4-1:0] node3416;
	wire [4-1:0] node3417;
	wire [4-1:0] node3418;
	wire [4-1:0] node3420;
	wire [4-1:0] node3423;
	wire [4-1:0] node3425;
	wire [4-1:0] node3427;
	wire [4-1:0] node3430;
	wire [4-1:0] node3431;
	wire [4-1:0] node3432;
	wire [4-1:0] node3433;
	wire [4-1:0] node3436;
	wire [4-1:0] node3440;
	wire [4-1:0] node3443;
	wire [4-1:0] node3444;
	wire [4-1:0] node3445;
	wire [4-1:0] node3446;
	wire [4-1:0] node3447;
	wire [4-1:0] node3448;
	wire [4-1:0] node3449;
	wire [4-1:0] node3452;
	wire [4-1:0] node3455;
	wire [4-1:0] node3456;
	wire [4-1:0] node3457;
	wire [4-1:0] node3460;
	wire [4-1:0] node3464;
	wire [4-1:0] node3465;
	wire [4-1:0] node3467;
	wire [4-1:0] node3470;
	wire [4-1:0] node3471;
	wire [4-1:0] node3472;
	wire [4-1:0] node3475;
	wire [4-1:0] node3478;
	wire [4-1:0] node3481;
	wire [4-1:0] node3482;
	wire [4-1:0] node3483;
	wire [4-1:0] node3484;
	wire [4-1:0] node3485;
	wire [4-1:0] node3487;
	wire [4-1:0] node3490;
	wire [4-1:0] node3492;
	wire [4-1:0] node3495;
	wire [4-1:0] node3496;
	wire [4-1:0] node3497;
	wire [4-1:0] node3500;
	wire [4-1:0] node3504;
	wire [4-1:0] node3505;
	wire [4-1:0] node3508;
	wire [4-1:0] node3511;
	wire [4-1:0] node3512;
	wire [4-1:0] node3514;
	wire [4-1:0] node3515;
	wire [4-1:0] node3518;
	wire [4-1:0] node3520;
	wire [4-1:0] node3523;
	wire [4-1:0] node3524;
	wire [4-1:0] node3525;
	wire [4-1:0] node3526;
	wire [4-1:0] node3529;
	wire [4-1:0] node3532;
	wire [4-1:0] node3533;
	wire [4-1:0] node3536;
	wire [4-1:0] node3539;
	wire [4-1:0] node3540;
	wire [4-1:0] node3541;
	wire [4-1:0] node3545;
	wire [4-1:0] node3548;
	wire [4-1:0] node3549;
	wire [4-1:0] node3550;
	wire [4-1:0] node3551;
	wire [4-1:0] node3552;
	wire [4-1:0] node3555;
	wire [4-1:0] node3558;
	wire [4-1:0] node3559;
	wire [4-1:0] node3561;
	wire [4-1:0] node3564;
	wire [4-1:0] node3567;
	wire [4-1:0] node3568;
	wire [4-1:0] node3569;
	wire [4-1:0] node3570;
	wire [4-1:0] node3571;
	wire [4-1:0] node3575;
	wire [4-1:0] node3577;
	wire [4-1:0] node3580;
	wire [4-1:0] node3582;
	wire [4-1:0] node3585;
	wire [4-1:0] node3586;
	wire [4-1:0] node3590;
	wire [4-1:0] node3591;
	wire [4-1:0] node3592;
	wire [4-1:0] node3593;
	wire [4-1:0] node3595;
	wire [4-1:0] node3598;
	wire [4-1:0] node3599;
	wire [4-1:0] node3603;
	wire [4-1:0] node3604;
	wire [4-1:0] node3606;
	wire [4-1:0] node3608;
	wire [4-1:0] node3611;
	wire [4-1:0] node3612;
	wire [4-1:0] node3613;
	wire [4-1:0] node3618;
	wire [4-1:0] node3619;
	wire [4-1:0] node3620;
	wire [4-1:0] node3621;
	wire [4-1:0] node3624;
	wire [4-1:0] node3627;
	wire [4-1:0] node3629;
	wire [4-1:0] node3632;
	wire [4-1:0] node3633;
	wire [4-1:0] node3634;
	wire [4-1:0] node3637;
	wire [4-1:0] node3641;
	wire [4-1:0] node3642;
	wire [4-1:0] node3643;
	wire [4-1:0] node3644;
	wire [4-1:0] node3645;
	wire [4-1:0] node3647;
	wire [4-1:0] node3648;
	wire [4-1:0] node3652;
	wire [4-1:0] node3653;
	wire [4-1:0] node3654;
	wire [4-1:0] node3657;
	wire [4-1:0] node3661;
	wire [4-1:0] node3662;
	wire [4-1:0] node3663;
	wire [4-1:0] node3666;
	wire [4-1:0] node3668;
	wire [4-1:0] node3671;
	wire [4-1:0] node3672;
	wire [4-1:0] node3675;
	wire [4-1:0] node3677;
	wire [4-1:0] node3680;
	wire [4-1:0] node3681;
	wire [4-1:0] node3682;
	wire [4-1:0] node3683;
	wire [4-1:0] node3684;
	wire [4-1:0] node3688;
	wire [4-1:0] node3689;
	wire [4-1:0] node3690;
	wire [4-1:0] node3695;
	wire [4-1:0] node3696;
	wire [4-1:0] node3698;
	wire [4-1:0] node3701;
	wire [4-1:0] node3704;
	wire [4-1:0] node3705;
	wire [4-1:0] node3706;
	wire [4-1:0] node3707;
	wire [4-1:0] node3708;
	wire [4-1:0] node3711;
	wire [4-1:0] node3715;
	wire [4-1:0] node3718;
	wire [4-1:0] node3719;
	wire [4-1:0] node3720;
	wire [4-1:0] node3722;
	wire [4-1:0] node3725;
	wire [4-1:0] node3727;
	wire [4-1:0] node3730;
	wire [4-1:0] node3731;
	wire [4-1:0] node3732;
	wire [4-1:0] node3735;
	wire [4-1:0] node3739;
	wire [4-1:0] node3740;
	wire [4-1:0] node3741;
	wire [4-1:0] node3742;
	wire [4-1:0] node3743;
	wire [4-1:0] node3745;
	wire [4-1:0] node3748;
	wire [4-1:0] node3749;
	wire [4-1:0] node3753;
	wire [4-1:0] node3754;
	wire [4-1:0] node3756;
	wire [4-1:0] node3759;
	wire [4-1:0] node3760;
	wire [4-1:0] node3762;
	wire [4-1:0] node3766;
	wire [4-1:0] node3767;
	wire [4-1:0] node3768;
	wire [4-1:0] node3770;
	wire [4-1:0] node3773;
	wire [4-1:0] node3775;
	wire [4-1:0] node3776;
	wire [4-1:0] node3779;
	wire [4-1:0] node3782;
	wire [4-1:0] node3783;
	wire [4-1:0] node3784;
	wire [4-1:0] node3789;
	wire [4-1:0] node3790;
	wire [4-1:0] node3791;
	wire [4-1:0] node3792;
	wire [4-1:0] node3795;
	wire [4-1:0] node3797;
	wire [4-1:0] node3800;
	wire [4-1:0] node3801;
	wire [4-1:0] node3803;
	wire [4-1:0] node3807;
	wire [4-1:0] node3809;
	wire [4-1:0] node3810;
	wire [4-1:0] node3812;
	wire [4-1:0] node3814;
	wire [4-1:0] node3818;
	wire [4-1:0] node3819;
	wire [4-1:0] node3820;
	wire [4-1:0] node3821;
	wire [4-1:0] node3822;
	wire [4-1:0] node3823;
	wire [4-1:0] node3824;
	wire [4-1:0] node3825;
	wire [4-1:0] node3828;
	wire [4-1:0] node3831;
	wire [4-1:0] node3832;
	wire [4-1:0] node3836;
	wire [4-1:0] node3837;
	wire [4-1:0] node3838;
	wire [4-1:0] node3842;
	wire [4-1:0] node3843;
	wire [4-1:0] node3845;
	wire [4-1:0] node3848;
	wire [4-1:0] node3849;
	wire [4-1:0] node3850;
	wire [4-1:0] node3855;
	wire [4-1:0] node3856;
	wire [4-1:0] node3857;
	wire [4-1:0] node3859;
	wire [4-1:0] node3860;
	wire [4-1:0] node3863;
	wire [4-1:0] node3864;
	wire [4-1:0] node3868;
	wire [4-1:0] node3869;
	wire [4-1:0] node3870;
	wire [4-1:0] node3874;
	wire [4-1:0] node3877;
	wire [4-1:0] node3878;
	wire [4-1:0] node3879;
	wire [4-1:0] node3881;
	wire [4-1:0] node3884;
	wire [4-1:0] node3885;
	wire [4-1:0] node3889;
	wire [4-1:0] node3890;
	wire [4-1:0] node3892;
	wire [4-1:0] node3893;
	wire [4-1:0] node3897;
	wire [4-1:0] node3898;
	wire [4-1:0] node3902;
	wire [4-1:0] node3903;
	wire [4-1:0] node3904;
	wire [4-1:0] node3905;
	wire [4-1:0] node3906;
	wire [4-1:0] node3908;
	wire [4-1:0] node3909;
	wire [4-1:0] node3914;
	wire [4-1:0] node3915;
	wire [4-1:0] node3916;
	wire [4-1:0] node3919;
	wire [4-1:0] node3922;
	wire [4-1:0] node3924;
	wire [4-1:0] node3927;
	wire [4-1:0] node3928;
	wire [4-1:0] node3929;
	wire [4-1:0] node3932;
	wire [4-1:0] node3935;
	wire [4-1:0] node3936;
	wire [4-1:0] node3937;
	wire [4-1:0] node3939;
	wire [4-1:0] node3944;
	wire [4-1:0] node3945;
	wire [4-1:0] node3946;
	wire [4-1:0] node3947;
	wire [4-1:0] node3949;
	wire [4-1:0] node3950;
	wire [4-1:0] node3953;
	wire [4-1:0] node3956;
	wire [4-1:0] node3957;
	wire [4-1:0] node3958;
	wire [4-1:0] node3961;
	wire [4-1:0] node3964;
	wire [4-1:0] node3966;
	wire [4-1:0] node3969;
	wire [4-1:0] node3970;
	wire [4-1:0] node3971;
	wire [4-1:0] node3972;
	wire [4-1:0] node3976;
	wire [4-1:0] node3979;
	wire [4-1:0] node3981;
	wire [4-1:0] node3984;
	wire [4-1:0] node3985;
	wire [4-1:0] node3987;
	wire [4-1:0] node3989;
	wire [4-1:0] node3992;
	wire [4-1:0] node3993;
	wire [4-1:0] node3994;
	wire [4-1:0] node3995;
	wire [4-1:0] node3999;
	wire [4-1:0] node4002;
	wire [4-1:0] node4005;
	wire [4-1:0] node4006;
	wire [4-1:0] node4007;
	wire [4-1:0] node4008;
	wire [4-1:0] node4009;
	wire [4-1:0] node4010;
	wire [4-1:0] node4014;
	wire [4-1:0] node4016;
	wire [4-1:0] node4017;
	wire [4-1:0] node4019;
	wire [4-1:0] node4022;
	wire [4-1:0] node4025;
	wire [4-1:0] node4026;
	wire [4-1:0] node4027;
	wire [4-1:0] node4031;
	wire [4-1:0] node4032;
	wire [4-1:0] node4033;
	wire [4-1:0] node4037;
	wire [4-1:0] node4039;
	wire [4-1:0] node4042;
	wire [4-1:0] node4043;
	wire [4-1:0] node4044;
	wire [4-1:0] node4045;
	wire [4-1:0] node4046;
	wire [4-1:0] node4047;
	wire [4-1:0] node4051;
	wire [4-1:0] node4052;
	wire [4-1:0] node4057;
	wire [4-1:0] node4058;
	wire [4-1:0] node4059;
	wire [4-1:0] node4061;
	wire [4-1:0] node4064;
	wire [4-1:0] node4067;
	wire [4-1:0] node4068;
	wire [4-1:0] node4072;
	wire [4-1:0] node4073;
	wire [4-1:0] node4074;
	wire [4-1:0] node4076;
	wire [4-1:0] node4078;
	wire [4-1:0] node4081;
	wire [4-1:0] node4083;
	wire [4-1:0] node4086;
	wire [4-1:0] node4087;
	wire [4-1:0] node4090;
	wire [4-1:0] node4092;
	wire [4-1:0] node4093;
	wire [4-1:0] node4096;
	wire [4-1:0] node4099;
	wire [4-1:0] node4100;
	wire [4-1:0] node4101;
	wire [4-1:0] node4102;
	wire [4-1:0] node4104;
	wire [4-1:0] node4105;
	wire [4-1:0] node4109;
	wire [4-1:0] node4110;
	wire [4-1:0] node4112;
	wire [4-1:0] node4113;
	wire [4-1:0] node4116;
	wire [4-1:0] node4119;
	wire [4-1:0] node4120;
	wire [4-1:0] node4124;
	wire [4-1:0] node4125;
	wire [4-1:0] node4126;
	wire [4-1:0] node4129;
	wire [4-1:0] node4132;
	wire [4-1:0] node4133;
	wire [4-1:0] node4136;
	wire [4-1:0] node4139;
	wire [4-1:0] node4140;
	wire [4-1:0] node4141;
	wire [4-1:0] node4142;
	wire [4-1:0] node4144;
	wire [4-1:0] node4148;
	wire [4-1:0] node4149;
	wire [4-1:0] node4152;
	wire [4-1:0] node4153;
	wire [4-1:0] node4155;
	wire [4-1:0] node4158;
	wire [4-1:0] node4161;
	wire [4-1:0] node4162;
	wire [4-1:0] node4164;
	wire [4-1:0] node4166;
	wire [4-1:0] node4167;
	wire [4-1:0] node4170;
	wire [4-1:0] node4173;
	wire [4-1:0] node4175;
	wire [4-1:0] node4178;
	wire [4-1:0] node4179;
	wire [4-1:0] node4180;
	wire [4-1:0] node4181;
	wire [4-1:0] node4182;
	wire [4-1:0] node4183;
	wire [4-1:0] node4184;
	wire [4-1:0] node4185;
	wire [4-1:0] node4188;
	wire [4-1:0] node4191;
	wire [4-1:0] node4193;
	wire [4-1:0] node4196;
	wire [4-1:0] node4198;
	wire [4-1:0] node4199;
	wire [4-1:0] node4203;
	wire [4-1:0] node4204;
	wire [4-1:0] node4205;
	wire [4-1:0] node4206;
	wire [4-1:0] node4209;
	wire [4-1:0] node4212;
	wire [4-1:0] node4213;
	wire [4-1:0] node4216;
	wire [4-1:0] node4219;
	wire [4-1:0] node4222;
	wire [4-1:0] node4223;
	wire [4-1:0] node4224;
	wire [4-1:0] node4225;
	wire [4-1:0] node4228;
	wire [4-1:0] node4230;
	wire [4-1:0] node4233;
	wire [4-1:0] node4234;
	wire [4-1:0] node4235;
	wire [4-1:0] node4237;
	wire [4-1:0] node4241;
	wire [4-1:0] node4244;
	wire [4-1:0] node4245;
	wire [4-1:0] node4246;
	wire [4-1:0] node4247;
	wire [4-1:0] node4249;
	wire [4-1:0] node4253;
	wire [4-1:0] node4254;
	wire [4-1:0] node4256;
	wire [4-1:0] node4259;
	wire [4-1:0] node4262;
	wire [4-1:0] node4263;
	wire [4-1:0] node4264;
	wire [4-1:0] node4266;
	wire [4-1:0] node4269;
	wire [4-1:0] node4271;
	wire [4-1:0] node4274;
	wire [4-1:0] node4277;
	wire [4-1:0] node4278;
	wire [4-1:0] node4279;
	wire [4-1:0] node4280;
	wire [4-1:0] node4281;
	wire [4-1:0] node4283;
	wire [4-1:0] node4287;
	wire [4-1:0] node4288;
	wire [4-1:0] node4290;
	wire [4-1:0] node4293;
	wire [4-1:0] node4294;
	wire [4-1:0] node4298;
	wire [4-1:0] node4299;
	wire [4-1:0] node4300;
	wire [4-1:0] node4302;
	wire [4-1:0] node4306;
	wire [4-1:0] node4307;
	wire [4-1:0] node4308;
	wire [4-1:0] node4312;
	wire [4-1:0] node4314;
	wire [4-1:0] node4315;
	wire [4-1:0] node4318;
	wire [4-1:0] node4321;
	wire [4-1:0] node4322;
	wire [4-1:0] node4323;
	wire [4-1:0] node4324;
	wire [4-1:0] node4325;
	wire [4-1:0] node4328;
	wire [4-1:0] node4331;
	wire [4-1:0] node4332;
	wire [4-1:0] node4336;
	wire [4-1:0] node4337;
	wire [4-1:0] node4340;
	wire [4-1:0] node4343;
	wire [4-1:0] node4344;
	wire [4-1:0] node4345;
	wire [4-1:0] node4346;
	wire [4-1:0] node4350;
	wire [4-1:0] node4353;
	wire [4-1:0] node4354;
	wire [4-1:0] node4357;
	wire [4-1:0] node4358;
	wire [4-1:0] node4361;
	wire [4-1:0] node4363;
	wire [4-1:0] node4366;
	wire [4-1:0] node4367;
	wire [4-1:0] node4368;
	wire [4-1:0] node4369;
	wire [4-1:0] node4370;
	wire [4-1:0] node4372;
	wire [4-1:0] node4375;
	wire [4-1:0] node4376;
	wire [4-1:0] node4377;
	wire [4-1:0] node4381;
	wire [4-1:0] node4382;
	wire [4-1:0] node4386;
	wire [4-1:0] node4387;
	wire [4-1:0] node4388;
	wire [4-1:0] node4390;
	wire [4-1:0] node4394;
	wire [4-1:0] node4395;
	wire [4-1:0] node4396;
	wire [4-1:0] node4398;
	wire [4-1:0] node4401;
	wire [4-1:0] node4404;
	wire [4-1:0] node4406;
	wire [4-1:0] node4409;
	wire [4-1:0] node4410;
	wire [4-1:0] node4411;
	wire [4-1:0] node4412;
	wire [4-1:0] node4413;
	wire [4-1:0] node4418;
	wire [4-1:0] node4420;
	wire [4-1:0] node4421;
	wire [4-1:0] node4425;
	wire [4-1:0] node4426;
	wire [4-1:0] node4427;
	wire [4-1:0] node4429;
	wire [4-1:0] node4433;
	wire [4-1:0] node4434;
	wire [4-1:0] node4436;
	wire [4-1:0] node4439;
	wire [4-1:0] node4442;
	wire [4-1:0] node4443;
	wire [4-1:0] node4444;
	wire [4-1:0] node4445;
	wire [4-1:0] node4446;
	wire [4-1:0] node4449;
	wire [4-1:0] node4452;
	wire [4-1:0] node4453;
	wire [4-1:0] node4454;
	wire [4-1:0] node4458;
	wire [4-1:0] node4459;
	wire [4-1:0] node4460;
	wire [4-1:0] node4464;
	wire [4-1:0] node4467;
	wire [4-1:0] node4468;
	wire [4-1:0] node4470;
	wire [4-1:0] node4472;
	wire [4-1:0] node4475;
	wire [4-1:0] node4477;
	wire [4-1:0] node4479;
	wire [4-1:0] node4482;
	wire [4-1:0] node4483;
	wire [4-1:0] node4484;
	wire [4-1:0] node4485;
	wire [4-1:0] node4486;
	wire [4-1:0] node4490;
	wire [4-1:0] node4492;
	wire [4-1:0] node4495;
	wire [4-1:0] node4496;
	wire [4-1:0] node4498;
	wire [4-1:0] node4501;
	wire [4-1:0] node4503;
	wire [4-1:0] node4506;
	wire [4-1:0] node4507;
	wire [4-1:0] node4508;
	wire [4-1:0] node4510;
	wire [4-1:0] node4513;
	wire [4-1:0] node4515;
	wire [4-1:0] node4516;
	wire [4-1:0] node4520;
	wire [4-1:0] node4523;
	wire [4-1:0] node4524;
	wire [4-1:0] node4525;
	wire [4-1:0] node4526;
	wire [4-1:0] node4527;
	wire [4-1:0] node4528;
	wire [4-1:0] node4529;
	wire [4-1:0] node4530;
	wire [4-1:0] node4531;
	wire [4-1:0] node4534;
	wire [4-1:0] node4537;
	wire [4-1:0] node4539;
	wire [4-1:0] node4540;
	wire [4-1:0] node4544;
	wire [4-1:0] node4545;
	wire [4-1:0] node4546;
	wire [4-1:0] node4547;
	wire [4-1:0] node4551;
	wire [4-1:0] node4553;
	wire [4-1:0] node4554;
	wire [4-1:0] node4557;
	wire [4-1:0] node4560;
	wire [4-1:0] node4561;
	wire [4-1:0] node4564;
	wire [4-1:0] node4567;
	wire [4-1:0] node4568;
	wire [4-1:0] node4569;
	wire [4-1:0] node4570;
	wire [4-1:0] node4571;
	wire [4-1:0] node4574;
	wire [4-1:0] node4577;
	wire [4-1:0] node4578;
	wire [4-1:0] node4582;
	wire [4-1:0] node4583;
	wire [4-1:0] node4584;
	wire [4-1:0] node4587;
	wire [4-1:0] node4590;
	wire [4-1:0] node4593;
	wire [4-1:0] node4594;
	wire [4-1:0] node4595;
	wire [4-1:0] node4596;
	wire [4-1:0] node4599;
	wire [4-1:0] node4603;
	wire [4-1:0] node4604;
	wire [4-1:0] node4605;
	wire [4-1:0] node4606;
	wire [4-1:0] node4609;
	wire [4-1:0] node4613;
	wire [4-1:0] node4615;
	wire [4-1:0] node4618;
	wire [4-1:0] node4619;
	wire [4-1:0] node4620;
	wire [4-1:0] node4621;
	wire [4-1:0] node4622;
	wire [4-1:0] node4625;
	wire [4-1:0] node4626;
	wire [4-1:0] node4629;
	wire [4-1:0] node4632;
	wire [4-1:0] node4634;
	wire [4-1:0] node4635;
	wire [4-1:0] node4639;
	wire [4-1:0] node4640;
	wire [4-1:0] node4641;
	wire [4-1:0] node4644;
	wire [4-1:0] node4645;
	wire [4-1:0] node4648;
	wire [4-1:0] node4651;
	wire [4-1:0] node4652;
	wire [4-1:0] node4653;
	wire [4-1:0] node4654;
	wire [4-1:0] node4658;
	wire [4-1:0] node4660;
	wire [4-1:0] node4664;
	wire [4-1:0] node4665;
	wire [4-1:0] node4666;
	wire [4-1:0] node4667;
	wire [4-1:0] node4670;
	wire [4-1:0] node4673;
	wire [4-1:0] node4674;
	wire [4-1:0] node4677;
	wire [4-1:0] node4680;
	wire [4-1:0] node4681;
	wire [4-1:0] node4683;
	wire [4-1:0] node4686;
	wire [4-1:0] node4687;
	wire [4-1:0] node4689;
	wire [4-1:0] node4692;
	wire [4-1:0] node4693;
	wire [4-1:0] node4696;
	wire [4-1:0] node4699;
	wire [4-1:0] node4700;
	wire [4-1:0] node4701;
	wire [4-1:0] node4702;
	wire [4-1:0] node4703;
	wire [4-1:0] node4704;
	wire [4-1:0] node4706;
	wire [4-1:0] node4707;
	wire [4-1:0] node4710;
	wire [4-1:0] node4713;
	wire [4-1:0] node4715;
	wire [4-1:0] node4718;
	wire [4-1:0] node4719;
	wire [4-1:0] node4720;
	wire [4-1:0] node4721;
	wire [4-1:0] node4724;
	wire [4-1:0] node4727;
	wire [4-1:0] node4730;
	wire [4-1:0] node4731;
	wire [4-1:0] node4735;
	wire [4-1:0] node4736;
	wire [4-1:0] node4737;
	wire [4-1:0] node4738;
	wire [4-1:0] node4739;
	wire [4-1:0] node4744;
	wire [4-1:0] node4745;
	wire [4-1:0] node4746;
	wire [4-1:0] node4749;
	wire [4-1:0] node4753;
	wire [4-1:0] node4754;
	wire [4-1:0] node4756;
	wire [4-1:0] node4759;
	wire [4-1:0] node4760;
	wire [4-1:0] node4761;
	wire [4-1:0] node4766;
	wire [4-1:0] node4767;
	wire [4-1:0] node4768;
	wire [4-1:0] node4769;
	wire [4-1:0] node4770;
	wire [4-1:0] node4771;
	wire [4-1:0] node4774;
	wire [4-1:0] node4777;
	wire [4-1:0] node4778;
	wire [4-1:0] node4781;
	wire [4-1:0] node4785;
	wire [4-1:0] node4786;
	wire [4-1:0] node4787;
	wire [4-1:0] node4788;
	wire [4-1:0] node4791;
	wire [4-1:0] node4794;
	wire [4-1:0] node4795;
	wire [4-1:0] node4799;
	wire [4-1:0] node4800;
	wire [4-1:0] node4801;
	wire [4-1:0] node4806;
	wire [4-1:0] node4807;
	wire [4-1:0] node4808;
	wire [4-1:0] node4809;
	wire [4-1:0] node4810;
	wire [4-1:0] node4813;
	wire [4-1:0] node4816;
	wire [4-1:0] node4819;
	wire [4-1:0] node4822;
	wire [4-1:0] node4823;
	wire [4-1:0] node4824;
	wire [4-1:0] node4825;
	wire [4-1:0] node4829;
	wire [4-1:0] node4833;
	wire [4-1:0] node4834;
	wire [4-1:0] node4835;
	wire [4-1:0] node4836;
	wire [4-1:0] node4837;
	wire [4-1:0] node4838;
	wire [4-1:0] node4840;
	wire [4-1:0] node4843;
	wire [4-1:0] node4845;
	wire [4-1:0] node4848;
	wire [4-1:0] node4851;
	wire [4-1:0] node4852;
	wire [4-1:0] node4854;
	wire [4-1:0] node4856;
	wire [4-1:0] node4859;
	wire [4-1:0] node4860;
	wire [4-1:0] node4864;
	wire [4-1:0] node4865;
	wire [4-1:0] node4867;
	wire [4-1:0] node4868;
	wire [4-1:0] node4870;
	wire [4-1:0] node4873;
	wire [4-1:0] node4876;
	wire [4-1:0] node4877;
	wire [4-1:0] node4878;
	wire [4-1:0] node4883;
	wire [4-1:0] node4884;
	wire [4-1:0] node4885;
	wire [4-1:0] node4886;
	wire [4-1:0] node4889;
	wire [4-1:0] node4890;
	wire [4-1:0] node4893;
	wire [4-1:0] node4896;
	wire [4-1:0] node4897;
	wire [4-1:0] node4898;
	wire [4-1:0] node4902;
	wire [4-1:0] node4903;
	wire [4-1:0] node4906;
	wire [4-1:0] node4907;
	wire [4-1:0] node4911;
	wire [4-1:0] node4912;
	wire [4-1:0] node4914;
	wire [4-1:0] node4915;
	wire [4-1:0] node4916;
	wire [4-1:0] node4919;
	wire [4-1:0] node4923;
	wire [4-1:0] node4924;
	wire [4-1:0] node4926;
	wire [4-1:0] node4929;
	wire [4-1:0] node4932;
	wire [4-1:0] node4933;
	wire [4-1:0] node4934;
	wire [4-1:0] node4935;
	wire [4-1:0] node4936;
	wire [4-1:0] node4937;
	wire [4-1:0] node4938;
	wire [4-1:0] node4940;
	wire [4-1:0] node4941;
	wire [4-1:0] node4944;
	wire [4-1:0] node4947;
	wire [4-1:0] node4950;
	wire [4-1:0] node4952;
	wire [4-1:0] node4953;
	wire [4-1:0] node4955;
	wire [4-1:0] node4959;
	wire [4-1:0] node4960;
	wire [4-1:0] node4961;
	wire [4-1:0] node4965;
	wire [4-1:0] node4966;
	wire [4-1:0] node4969;
	wire [4-1:0] node4972;
	wire [4-1:0] node4973;
	wire [4-1:0] node4974;
	wire [4-1:0] node4975;
	wire [4-1:0] node4976;
	wire [4-1:0] node4978;
	wire [4-1:0] node4982;
	wire [4-1:0] node4983;
	wire [4-1:0] node4985;
	wire [4-1:0] node4990;
	wire [4-1:0] node4991;
	wire [4-1:0] node4993;
	wire [4-1:0] node4994;
	wire [4-1:0] node4995;
	wire [4-1:0] node4999;
	wire [4-1:0] node5000;
	wire [4-1:0] node5004;
	wire [4-1:0] node5005;
	wire [4-1:0] node5006;
	wire [4-1:0] node5010;
	wire [4-1:0] node5011;
	wire [4-1:0] node5012;
	wire [4-1:0] node5016;
	wire [4-1:0] node5018;
	wire [4-1:0] node5021;
	wire [4-1:0] node5022;
	wire [4-1:0] node5023;
	wire [4-1:0] node5024;
	wire [4-1:0] node5025;
	wire [4-1:0] node5027;
	wire [4-1:0] node5028;
	wire [4-1:0] node5032;
	wire [4-1:0] node5035;
	wire [4-1:0] node5036;
	wire [4-1:0] node5039;
	wire [4-1:0] node5041;
	wire [4-1:0] node5044;
	wire [4-1:0] node5045;
	wire [4-1:0] node5047;
	wire [4-1:0] node5048;
	wire [4-1:0] node5051;
	wire [4-1:0] node5052;
	wire [4-1:0] node5056;
	wire [4-1:0] node5057;
	wire [4-1:0] node5058;
	wire [4-1:0] node5059;
	wire [4-1:0] node5062;
	wire [4-1:0] node5065;
	wire [4-1:0] node5066;
	wire [4-1:0] node5070;
	wire [4-1:0] node5073;
	wire [4-1:0] node5074;
	wire [4-1:0] node5076;
	wire [4-1:0] node5077;
	wire [4-1:0] node5079;
	wire [4-1:0] node5080;
	wire [4-1:0] node5084;
	wire [4-1:0] node5086;
	wire [4-1:0] node5087;
	wire [4-1:0] node5090;
	wire [4-1:0] node5093;
	wire [4-1:0] node5094;
	wire [4-1:0] node5095;
	wire [4-1:0] node5097;
	wire [4-1:0] node5100;
	wire [4-1:0] node5102;
	wire [4-1:0] node5105;
	wire [4-1:0] node5108;
	wire [4-1:0] node5109;
	wire [4-1:0] node5110;
	wire [4-1:0] node5111;
	wire [4-1:0] node5112;
	wire [4-1:0] node5113;
	wire [4-1:0] node5115;
	wire [4-1:0] node5116;
	wire [4-1:0] node5119;
	wire [4-1:0] node5122;
	wire [4-1:0] node5123;
	wire [4-1:0] node5127;
	wire [4-1:0] node5128;
	wire [4-1:0] node5129;
	wire [4-1:0] node5130;
	wire [4-1:0] node5135;
	wire [4-1:0] node5136;
	wire [4-1:0] node5139;
	wire [4-1:0] node5142;
	wire [4-1:0] node5144;
	wire [4-1:0] node5145;
	wire [4-1:0] node5146;
	wire [4-1:0] node5148;
	wire [4-1:0] node5152;
	wire [4-1:0] node5154;
	wire [4-1:0] node5155;
	wire [4-1:0] node5159;
	wire [4-1:0] node5160;
	wire [4-1:0] node5161;
	wire [4-1:0] node5162;
	wire [4-1:0] node5164;
	wire [4-1:0] node5165;
	wire [4-1:0] node5169;
	wire [4-1:0] node5172;
	wire [4-1:0] node5173;
	wire [4-1:0] node5174;
	wire [4-1:0] node5178;
	wire [4-1:0] node5181;
	wire [4-1:0] node5182;
	wire [4-1:0] node5183;
	wire [4-1:0] node5185;
	wire [4-1:0] node5186;
	wire [4-1:0] node5189;
	wire [4-1:0] node5192;
	wire [4-1:0] node5193;
	wire [4-1:0] node5196;
	wire [4-1:0] node5199;
	wire [4-1:0] node5200;
	wire [4-1:0] node5201;
	wire [4-1:0] node5202;
	wire [4-1:0] node5205;
	wire [4-1:0] node5209;
	wire [4-1:0] node5210;
	wire [4-1:0] node5213;
	wire [4-1:0] node5214;
	wire [4-1:0] node5218;
	wire [4-1:0] node5219;
	wire [4-1:0] node5220;
	wire [4-1:0] node5221;
	wire [4-1:0] node5223;
	wire [4-1:0] node5226;
	wire [4-1:0] node5227;
	wire [4-1:0] node5228;
	wire [4-1:0] node5232;
	wire [4-1:0] node5234;
	wire [4-1:0] node5237;
	wire [4-1:0] node5238;
	wire [4-1:0] node5239;
	wire [4-1:0] node5241;
	wire [4-1:0] node5245;
	wire [4-1:0] node5248;
	wire [4-1:0] node5249;
	wire [4-1:0] node5250;
	wire [4-1:0] node5251;
	wire [4-1:0] node5252;
	wire [4-1:0] node5254;
	wire [4-1:0] node5257;
	wire [4-1:0] node5259;
	wire [4-1:0] node5262;
	wire [4-1:0] node5263;
	wire [4-1:0] node5265;
	wire [4-1:0] node5269;
	wire [4-1:0] node5270;
	wire [4-1:0] node5272;
	wire [4-1:0] node5275;
	wire [4-1:0] node5277;
	wire [4-1:0] node5280;
	wire [4-1:0] node5281;
	wire [4-1:0] node5282;
	wire [4-1:0] node5283;
	wire [4-1:0] node5284;
	wire [4-1:0] node5288;
	wire [4-1:0] node5291;
	wire [4-1:0] node5294;
	wire [4-1:0] node5295;
	wire [4-1:0] node5298;
	wire [4-1:0] node5301;
	wire [4-1:0] node5302;
	wire [4-1:0] node5303;
	wire [4-1:0] node5304;
	wire [4-1:0] node5305;
	wire [4-1:0] node5306;
	wire [4-1:0] node5307;
	wire [4-1:0] node5308;
	wire [4-1:0] node5311;
	wire [4-1:0] node5314;
	wire [4-1:0] node5315;
	wire [4-1:0] node5316;
	wire [4-1:0] node5319;
	wire [4-1:0] node5322;
	wire [4-1:0] node5323;
	wire [4-1:0] node5326;
	wire [4-1:0] node5327;
	wire [4-1:0] node5331;
	wire [4-1:0] node5332;
	wire [4-1:0] node5334;
	wire [4-1:0] node5335;
	wire [4-1:0] node5338;
	wire [4-1:0] node5341;
	wire [4-1:0] node5342;
	wire [4-1:0] node5343;
	wire [4-1:0] node5347;
	wire [4-1:0] node5349;
	wire [4-1:0] node5352;
	wire [4-1:0] node5353;
	wire [4-1:0] node5355;
	wire [4-1:0] node5356;
	wire [4-1:0] node5357;
	wire [4-1:0] node5361;
	wire [4-1:0] node5362;
	wire [4-1:0] node5366;
	wire [4-1:0] node5367;
	wire [4-1:0] node5369;
	wire [4-1:0] node5372;
	wire [4-1:0] node5373;
	wire [4-1:0] node5375;
	wire [4-1:0] node5378;
	wire [4-1:0] node5381;
	wire [4-1:0] node5382;
	wire [4-1:0] node5383;
	wire [4-1:0] node5384;
	wire [4-1:0] node5387;
	wire [4-1:0] node5388;
	wire [4-1:0] node5389;
	wire [4-1:0] node5393;
	wire [4-1:0] node5395;
	wire [4-1:0] node5396;
	wire [4-1:0] node5400;
	wire [4-1:0] node5401;
	wire [4-1:0] node5403;
	wire [4-1:0] node5405;
	wire [4-1:0] node5408;
	wire [4-1:0] node5410;
	wire [4-1:0] node5412;
	wire [4-1:0] node5415;
	wire [4-1:0] node5416;
	wire [4-1:0] node5417;
	wire [4-1:0] node5418;
	wire [4-1:0] node5419;
	wire [4-1:0] node5423;
	wire [4-1:0] node5425;
	wire [4-1:0] node5427;
	wire [4-1:0] node5430;
	wire [4-1:0] node5431;
	wire [4-1:0] node5432;
	wire [4-1:0] node5434;
	wire [4-1:0] node5437;
	wire [4-1:0] node5439;
	wire [4-1:0] node5442;
	wire [4-1:0] node5445;
	wire [4-1:0] node5446;
	wire [4-1:0] node5447;
	wire [4-1:0] node5448;
	wire [4-1:0] node5453;
	wire [4-1:0] node5454;
	wire [4-1:0] node5456;
	wire [4-1:0] node5459;
	wire [4-1:0] node5461;
	wire [4-1:0] node5464;
	wire [4-1:0] node5465;
	wire [4-1:0] node5466;
	wire [4-1:0] node5467;
	wire [4-1:0] node5468;
	wire [4-1:0] node5469;
	wire [4-1:0] node5470;
	wire [4-1:0] node5474;
	wire [4-1:0] node5476;
	wire [4-1:0] node5479;
	wire [4-1:0] node5480;
	wire [4-1:0] node5481;
	wire [4-1:0] node5485;
	wire [4-1:0] node5486;
	wire [4-1:0] node5487;
	wire [4-1:0] node5490;
	wire [4-1:0] node5494;
	wire [4-1:0] node5495;
	wire [4-1:0] node5496;
	wire [4-1:0] node5500;
	wire [4-1:0] node5501;
	wire [4-1:0] node5502;
	wire [4-1:0] node5503;
	wire [4-1:0] node5506;
	wire [4-1:0] node5510;
	wire [4-1:0] node5512;
	wire [4-1:0] node5515;
	wire [4-1:0] node5516;
	wire [4-1:0] node5517;
	wire [4-1:0] node5518;
	wire [4-1:0] node5519;
	wire [4-1:0] node5524;
	wire [4-1:0] node5525;
	wire [4-1:0] node5526;
	wire [4-1:0] node5530;
	wire [4-1:0] node5533;
	wire [4-1:0] node5534;
	wire [4-1:0] node5535;
	wire [4-1:0] node5539;
	wire [4-1:0] node5540;
	wire [4-1:0] node5541;
	wire [4-1:0] node5545;
	wire [4-1:0] node5548;
	wire [4-1:0] node5549;
	wire [4-1:0] node5550;
	wire [4-1:0] node5551;
	wire [4-1:0] node5552;
	wire [4-1:0] node5555;
	wire [4-1:0] node5558;
	wire [4-1:0] node5559;
	wire [4-1:0] node5560;
	wire [4-1:0] node5563;
	wire [4-1:0] node5566;
	wire [4-1:0] node5568;
	wire [4-1:0] node5571;
	wire [4-1:0] node5572;
	wire [4-1:0] node5573;
	wire [4-1:0] node5574;
	wire [4-1:0] node5577;
	wire [4-1:0] node5581;
	wire [4-1:0] node5583;
	wire [4-1:0] node5584;
	wire [4-1:0] node5587;
	wire [4-1:0] node5590;
	wire [4-1:0] node5591;
	wire [4-1:0] node5592;
	wire [4-1:0] node5593;
	wire [4-1:0] node5595;
	wire [4-1:0] node5598;
	wire [4-1:0] node5600;
	wire [4-1:0] node5601;
	wire [4-1:0] node5604;
	wire [4-1:0] node5607;
	wire [4-1:0] node5608;
	wire [4-1:0] node5610;
	wire [4-1:0] node5613;
	wire [4-1:0] node5614;
	wire [4-1:0] node5617;
	wire [4-1:0] node5620;
	wire [4-1:0] node5621;
	wire [4-1:0] node5622;
	wire [4-1:0] node5623;
	wire [4-1:0] node5624;
	wire [4-1:0] node5628;
	wire [4-1:0] node5629;
	wire [4-1:0] node5633;
	wire [4-1:0] node5636;
	wire [4-1:0] node5637;
	wire [4-1:0] node5639;
	wire [4-1:0] node5642;
	wire [4-1:0] node5643;
	wire [4-1:0] node5646;
	wire [4-1:0] node5649;
	wire [4-1:0] node5650;
	wire [4-1:0] node5651;
	wire [4-1:0] node5652;
	wire [4-1:0] node5653;
	wire [4-1:0] node5654;
	wire [4-1:0] node5655;
	wire [4-1:0] node5656;
	wire [4-1:0] node5657;
	wire [4-1:0] node5660;
	wire [4-1:0] node5664;
	wire [4-1:0] node5665;
	wire [4-1:0] node5666;
	wire [4-1:0] node5669;
	wire [4-1:0] node5672;
	wire [4-1:0] node5673;
	wire [4-1:0] node5677;
	wire [4-1:0] node5678;
	wire [4-1:0] node5680;
	wire [4-1:0] node5681;
	wire [4-1:0] node5684;
	wire [4-1:0] node5687;
	wire [4-1:0] node5690;
	wire [4-1:0] node5691;
	wire [4-1:0] node5692;
	wire [4-1:0] node5694;
	wire [4-1:0] node5695;
	wire [4-1:0] node5698;
	wire [4-1:0] node5701;
	wire [4-1:0] node5703;
	wire [4-1:0] node5706;
	wire [4-1:0] node5707;
	wire [4-1:0] node5708;
	wire [4-1:0] node5711;
	wire [4-1:0] node5714;
	wire [4-1:0] node5715;
	wire [4-1:0] node5719;
	wire [4-1:0] node5720;
	wire [4-1:0] node5721;
	wire [4-1:0] node5723;
	wire [4-1:0] node5724;
	wire [4-1:0] node5725;
	wire [4-1:0] node5730;
	wire [4-1:0] node5731;
	wire [4-1:0] node5735;
	wire [4-1:0] node5736;
	wire [4-1:0] node5737;
	wire [4-1:0] node5738;
	wire [4-1:0] node5741;
	wire [4-1:0] node5744;
	wire [4-1:0] node5747;
	wire [4-1:0] node5748;
	wire [4-1:0] node5751;
	wire [4-1:0] node5752;
	wire [4-1:0] node5755;
	wire [4-1:0] node5756;
	wire [4-1:0] node5760;
	wire [4-1:0] node5761;
	wire [4-1:0] node5762;
	wire [4-1:0] node5763;
	wire [4-1:0] node5764;
	wire [4-1:0] node5766;
	wire [4-1:0] node5767;
	wire [4-1:0] node5770;
	wire [4-1:0] node5774;
	wire [4-1:0] node5775;
	wire [4-1:0] node5777;
	wire [4-1:0] node5779;
	wire [4-1:0] node5782;
	wire [4-1:0] node5784;
	wire [4-1:0] node5787;
	wire [4-1:0] node5788;
	wire [4-1:0] node5789;
	wire [4-1:0] node5790;
	wire [4-1:0] node5793;
	wire [4-1:0] node5795;
	wire [4-1:0] node5798;
	wire [4-1:0] node5799;
	wire [4-1:0] node5803;
	wire [4-1:0] node5804;
	wire [4-1:0] node5805;
	wire [4-1:0] node5808;
	wire [4-1:0] node5810;
	wire [4-1:0] node5813;
	wire [4-1:0] node5814;
	wire [4-1:0] node5815;
	wire [4-1:0] node5818;
	wire [4-1:0] node5821;
	wire [4-1:0] node5824;
	wire [4-1:0] node5825;
	wire [4-1:0] node5826;
	wire [4-1:0] node5827;
	wire [4-1:0] node5830;
	wire [4-1:0] node5832;
	wire [4-1:0] node5835;
	wire [4-1:0] node5836;
	wire [4-1:0] node5838;
	wire [4-1:0] node5840;
	wire [4-1:0] node5844;
	wire [4-1:0] node5845;
	wire [4-1:0] node5846;
	wire [4-1:0] node5847;
	wire [4-1:0] node5848;
	wire [4-1:0] node5851;
	wire [4-1:0] node5854;
	wire [4-1:0] node5855;
	wire [4-1:0] node5859;
	wire [4-1:0] node5862;
	wire [4-1:0] node5863;
	wire [4-1:0] node5864;
	wire [4-1:0] node5868;
	wire [4-1:0] node5869;
	wire [4-1:0] node5870;
	wire [4-1:0] node5873;
	wire [4-1:0] node5876;
	wire [4-1:0] node5879;
	wire [4-1:0] node5880;
	wire [4-1:0] node5881;
	wire [4-1:0] node5882;
	wire [4-1:0] node5883;
	wire [4-1:0] node5884;
	wire [4-1:0] node5888;
	wire [4-1:0] node5889;
	wire [4-1:0] node5891;
	wire [4-1:0] node5892;
	wire [4-1:0] node5895;
	wire [4-1:0] node5898;
	wire [4-1:0] node5899;
	wire [4-1:0] node5902;
	wire [4-1:0] node5905;
	wire [4-1:0] node5906;
	wire [4-1:0] node5907;
	wire [4-1:0] node5908;
	wire [4-1:0] node5911;
	wire [4-1:0] node5914;
	wire [4-1:0] node5915;
	wire [4-1:0] node5918;
	wire [4-1:0] node5921;
	wire [4-1:0] node5922;
	wire [4-1:0] node5924;
	wire [4-1:0] node5925;
	wire [4-1:0] node5928;
	wire [4-1:0] node5932;
	wire [4-1:0] node5933;
	wire [4-1:0] node5934;
	wire [4-1:0] node5935;
	wire [4-1:0] node5937;
	wire [4-1:0] node5938;
	wire [4-1:0] node5942;
	wire [4-1:0] node5943;
	wire [4-1:0] node5946;
	wire [4-1:0] node5949;
	wire [4-1:0] node5950;
	wire [4-1:0] node5952;
	wire [4-1:0] node5955;
	wire [4-1:0] node5957;
	wire [4-1:0] node5960;
	wire [4-1:0] node5961;
	wire [4-1:0] node5963;
	wire [4-1:0] node5965;
	wire [4-1:0] node5968;
	wire [4-1:0] node5969;
	wire [4-1:0] node5970;
	wire [4-1:0] node5973;
	wire [4-1:0] node5974;
	wire [4-1:0] node5978;
	wire [4-1:0] node5979;
	wire [4-1:0] node5980;
	wire [4-1:0] node5985;
	wire [4-1:0] node5986;
	wire [4-1:0] node5987;
	wire [4-1:0] node5988;
	wire [4-1:0] node5989;
	wire [4-1:0] node5993;
	wire [4-1:0] node5994;
	wire [4-1:0] node5995;
	wire [4-1:0] node5998;
	wire [4-1:0] node5999;
	wire [4-1:0] node6002;
	wire [4-1:0] node6005;
	wire [4-1:0] node6006;
	wire [4-1:0] node6009;
	wire [4-1:0] node6010;
	wire [4-1:0] node6014;
	wire [4-1:0] node6015;
	wire [4-1:0] node6017;
	wire [4-1:0] node6019;
	wire [4-1:0] node6021;
	wire [4-1:0] node6024;
	wire [4-1:0] node6025;
	wire [4-1:0] node6027;
	wire [4-1:0] node6030;
	wire [4-1:0] node6033;
	wire [4-1:0] node6034;
	wire [4-1:0] node6035;
	wire [4-1:0] node6036;
	wire [4-1:0] node6038;
	wire [4-1:0] node6041;
	wire [4-1:0] node6042;
	wire [4-1:0] node6044;
	wire [4-1:0] node6047;
	wire [4-1:0] node6050;
	wire [4-1:0] node6052;
	wire [4-1:0] node6054;
	wire [4-1:0] node6057;
	wire [4-1:0] node6058;
	wire [4-1:0] node6059;
	wire [4-1:0] node6061;
	wire [4-1:0] node6064;
	wire [4-1:0] node6067;
	wire [4-1:0] node6068;
	wire [4-1:0] node6069;
	wire [4-1:0] node6070;
	wire [4-1:0] node6075;
	wire [4-1:0] node6078;
	wire [4-1:0] node6079;
	wire [4-1:0] node6080;
	wire [4-1:0] node6081;
	wire [4-1:0] node6082;
	wire [4-1:0] node6083;
	wire [4-1:0] node6084;
	wire [4-1:0] node6085;
	wire [4-1:0] node6086;
	wire [4-1:0] node6087;
	wire [4-1:0] node6088;
	wire [4-1:0] node6090;
	wire [4-1:0] node6091;
	wire [4-1:0] node6095;
	wire [4-1:0] node6096;
	wire [4-1:0] node6100;
	wire [4-1:0] node6101;
	wire [4-1:0] node6102;
	wire [4-1:0] node6103;
	wire [4-1:0] node6106;
	wire [4-1:0] node6110;
	wire [4-1:0] node6112;
	wire [4-1:0] node6115;
	wire [4-1:0] node6116;
	wire [4-1:0] node6117;
	wire [4-1:0] node6118;
	wire [4-1:0] node6120;
	wire [4-1:0] node6125;
	wire [4-1:0] node6126;
	wire [4-1:0] node6128;
	wire [4-1:0] node6129;
	wire [4-1:0] node6134;
	wire [4-1:0] node6135;
	wire [4-1:0] node6136;
	wire [4-1:0] node6137;
	wire [4-1:0] node6139;
	wire [4-1:0] node6141;
	wire [4-1:0] node6144;
	wire [4-1:0] node6145;
	wire [4-1:0] node6146;
	wire [4-1:0] node6151;
	wire [4-1:0] node6152;
	wire [4-1:0] node6153;
	wire [4-1:0] node6154;
	wire [4-1:0] node6158;
	wire [4-1:0] node6161;
	wire [4-1:0] node6162;
	wire [4-1:0] node6163;
	wire [4-1:0] node6168;
	wire [4-1:0] node6169;
	wire [4-1:0] node6170;
	wire [4-1:0] node6171;
	wire [4-1:0] node6172;
	wire [4-1:0] node6177;
	wire [4-1:0] node6178;
	wire [4-1:0] node6182;
	wire [4-1:0] node6183;
	wire [4-1:0] node6184;
	wire [4-1:0] node6185;
	wire [4-1:0] node6188;
	wire [4-1:0] node6191;
	wire [4-1:0] node6193;
	wire [4-1:0] node6196;
	wire [4-1:0] node6198;
	wire [4-1:0] node6201;
	wire [4-1:0] node6202;
	wire [4-1:0] node6203;
	wire [4-1:0] node6204;
	wire [4-1:0] node6205;
	wire [4-1:0] node6207;
	wire [4-1:0] node6211;
	wire [4-1:0] node6212;
	wire [4-1:0] node6214;
	wire [4-1:0] node6215;
	wire [4-1:0] node6218;
	wire [4-1:0] node6221;
	wire [4-1:0] node6222;
	wire [4-1:0] node6224;
	wire [4-1:0] node6227;
	wire [4-1:0] node6228;
	wire [4-1:0] node6232;
	wire [4-1:0] node6233;
	wire [4-1:0] node6234;
	wire [4-1:0] node6235;
	wire [4-1:0] node6238;
	wire [4-1:0] node6241;
	wire [4-1:0] node6242;
	wire [4-1:0] node6243;
	wire [4-1:0] node6247;
	wire [4-1:0] node6249;
	wire [4-1:0] node6252;
	wire [4-1:0] node6253;
	wire [4-1:0] node6254;
	wire [4-1:0] node6258;
	wire [4-1:0] node6260;
	wire [4-1:0] node6262;
	wire [4-1:0] node6265;
	wire [4-1:0] node6266;
	wire [4-1:0] node6268;
	wire [4-1:0] node6270;
	wire [4-1:0] node6271;
	wire [4-1:0] node6274;
	wire [4-1:0] node6277;
	wire [4-1:0] node6278;
	wire [4-1:0] node6279;
	wire [4-1:0] node6283;
	wire [4-1:0] node6286;
	wire [4-1:0] node6287;
	wire [4-1:0] node6288;
	wire [4-1:0] node6289;
	wire [4-1:0] node6290;
	wire [4-1:0] node6291;
	wire [4-1:0] node6294;
	wire [4-1:0] node6295;
	wire [4-1:0] node6296;
	wire [4-1:0] node6299;
	wire [4-1:0] node6302;
	wire [4-1:0] node6303;
	wire [4-1:0] node6307;
	wire [4-1:0] node6308;
	wire [4-1:0] node6309;
	wire [4-1:0] node6312;
	wire [4-1:0] node6315;
	wire [4-1:0] node6316;
	wire [4-1:0] node6320;
	wire [4-1:0] node6321;
	wire [4-1:0] node6322;
	wire [4-1:0] node6325;
	wire [4-1:0] node6327;
	wire [4-1:0] node6330;
	wire [4-1:0] node6331;
	wire [4-1:0] node6333;
	wire [4-1:0] node6335;
	wire [4-1:0] node6338;
	wire [4-1:0] node6340;
	wire [4-1:0] node6343;
	wire [4-1:0] node6344;
	wire [4-1:0] node6345;
	wire [4-1:0] node6346;
	wire [4-1:0] node6350;
	wire [4-1:0] node6351;
	wire [4-1:0] node6352;
	wire [4-1:0] node6353;
	wire [4-1:0] node6356;
	wire [4-1:0] node6360;
	wire [4-1:0] node6362;
	wire [4-1:0] node6363;
	wire [4-1:0] node6366;
	wire [4-1:0] node6369;
	wire [4-1:0] node6370;
	wire [4-1:0] node6373;
	wire [4-1:0] node6374;
	wire [4-1:0] node6377;
	wire [4-1:0] node6378;
	wire [4-1:0] node6380;
	wire [4-1:0] node6384;
	wire [4-1:0] node6385;
	wire [4-1:0] node6386;
	wire [4-1:0] node6387;
	wire [4-1:0] node6388;
	wire [4-1:0] node6389;
	wire [4-1:0] node6393;
	wire [4-1:0] node6394;
	wire [4-1:0] node6397;
	wire [4-1:0] node6400;
	wire [4-1:0] node6401;
	wire [4-1:0] node6402;
	wire [4-1:0] node6405;
	wire [4-1:0] node6408;
	wire [4-1:0] node6411;
	wire [4-1:0] node6412;
	wire [4-1:0] node6413;
	wire [4-1:0] node6414;
	wire [4-1:0] node6417;
	wire [4-1:0] node6418;
	wire [4-1:0] node6422;
	wire [4-1:0] node6425;
	wire [4-1:0] node6427;
	wire [4-1:0] node6430;
	wire [4-1:0] node6431;
	wire [4-1:0] node6432;
	wire [4-1:0] node6434;
	wire [4-1:0] node6435;
	wire [4-1:0] node6438;
	wire [4-1:0] node6441;
	wire [4-1:0] node6443;
	wire [4-1:0] node6445;
	wire [4-1:0] node6446;
	wire [4-1:0] node6450;
	wire [4-1:0] node6451;
	wire [4-1:0] node6452;
	wire [4-1:0] node6453;
	wire [4-1:0] node6456;
	wire [4-1:0] node6458;
	wire [4-1:0] node6461;
	wire [4-1:0] node6462;
	wire [4-1:0] node6466;
	wire [4-1:0] node6467;
	wire [4-1:0] node6469;
	wire [4-1:0] node6472;
	wire [4-1:0] node6474;
	wire [4-1:0] node6477;
	wire [4-1:0] node6478;
	wire [4-1:0] node6479;
	wire [4-1:0] node6480;
	wire [4-1:0] node6481;
	wire [4-1:0] node6482;
	wire [4-1:0] node6483;
	wire [4-1:0] node6484;
	wire [4-1:0] node6489;
	wire [4-1:0] node6490;
	wire [4-1:0] node6491;
	wire [4-1:0] node6493;
	wire [4-1:0] node6498;
	wire [4-1:0] node6499;
	wire [4-1:0] node6500;
	wire [4-1:0] node6503;
	wire [4-1:0] node6506;
	wire [4-1:0] node6507;
	wire [4-1:0] node6508;
	wire [4-1:0] node6512;
	wire [4-1:0] node6513;
	wire [4-1:0] node6517;
	wire [4-1:0] node6518;
	wire [4-1:0] node6519;
	wire [4-1:0] node6520;
	wire [4-1:0] node6523;
	wire [4-1:0] node6525;
	wire [4-1:0] node6527;
	wire [4-1:0] node6530;
	wire [4-1:0] node6532;
	wire [4-1:0] node6534;
	wire [4-1:0] node6537;
	wire [4-1:0] node6538;
	wire [4-1:0] node6539;
	wire [4-1:0] node6542;
	wire [4-1:0] node6543;
	wire [4-1:0] node6546;
	wire [4-1:0] node6547;
	wire [4-1:0] node6551;
	wire [4-1:0] node6552;
	wire [4-1:0] node6554;
	wire [4-1:0] node6555;
	wire [4-1:0] node6558;
	wire [4-1:0] node6561;
	wire [4-1:0] node6562;
	wire [4-1:0] node6566;
	wire [4-1:0] node6567;
	wire [4-1:0] node6568;
	wire [4-1:0] node6569;
	wire [4-1:0] node6570;
	wire [4-1:0] node6573;
	wire [4-1:0] node6576;
	wire [4-1:0] node6577;
	wire [4-1:0] node6578;
	wire [4-1:0] node6580;
	wire [4-1:0] node6584;
	wire [4-1:0] node6587;
	wire [4-1:0] node6588;
	wire [4-1:0] node6589;
	wire [4-1:0] node6590;
	wire [4-1:0] node6593;
	wire [4-1:0] node6595;
	wire [4-1:0] node6598;
	wire [4-1:0] node6601;
	wire [4-1:0] node6602;
	wire [4-1:0] node6603;
	wire [4-1:0] node6606;
	wire [4-1:0] node6607;
	wire [4-1:0] node6611;
	wire [4-1:0] node6612;
	wire [4-1:0] node6616;
	wire [4-1:0] node6617;
	wire [4-1:0] node6618;
	wire [4-1:0] node6619;
	wire [4-1:0] node6620;
	wire [4-1:0] node6621;
	wire [4-1:0] node6625;
	wire [4-1:0] node6629;
	wire [4-1:0] node6630;
	wire [4-1:0] node6631;
	wire [4-1:0] node6635;
	wire [4-1:0] node6638;
	wire [4-1:0] node6639;
	wire [4-1:0] node6640;
	wire [4-1:0] node6641;
	wire [4-1:0] node6642;
	wire [4-1:0] node6645;
	wire [4-1:0] node6649;
	wire [4-1:0] node6650;
	wire [4-1:0] node6653;
	wire [4-1:0] node6656;
	wire [4-1:0] node6657;
	wire [4-1:0] node6658;
	wire [4-1:0] node6662;
	wire [4-1:0] node6663;
	wire [4-1:0] node6666;
	wire [4-1:0] node6669;
	wire [4-1:0] node6670;
	wire [4-1:0] node6671;
	wire [4-1:0] node6672;
	wire [4-1:0] node6673;
	wire [4-1:0] node6674;
	wire [4-1:0] node6675;
	wire [4-1:0] node6679;
	wire [4-1:0] node6680;
	wire [4-1:0] node6681;
	wire [4-1:0] node6684;
	wire [4-1:0] node6687;
	wire [4-1:0] node6688;
	wire [4-1:0] node6691;
	wire [4-1:0] node6694;
	wire [4-1:0] node6695;
	wire [4-1:0] node6696;
	wire [4-1:0] node6697;
	wire [4-1:0] node6701;
	wire [4-1:0] node6705;
	wire [4-1:0] node6706;
	wire [4-1:0] node6708;
	wire [4-1:0] node6709;
	wire [4-1:0] node6711;
	wire [4-1:0] node6715;
	wire [4-1:0] node6716;
	wire [4-1:0] node6717;
	wire [4-1:0] node6721;
	wire [4-1:0] node6722;
	wire [4-1:0] node6723;
	wire [4-1:0] node6726;
	wire [4-1:0] node6729;
	wire [4-1:0] node6732;
	wire [4-1:0] node6733;
	wire [4-1:0] node6734;
	wire [4-1:0] node6735;
	wire [4-1:0] node6736;
	wire [4-1:0] node6737;
	wire [4-1:0] node6741;
	wire [4-1:0] node6744;
	wire [4-1:0] node6745;
	wire [4-1:0] node6747;
	wire [4-1:0] node6751;
	wire [4-1:0] node6752;
	wire [4-1:0] node6753;
	wire [4-1:0] node6754;
	wire [4-1:0] node6758;
	wire [4-1:0] node6760;
	wire [4-1:0] node6763;
	wire [4-1:0] node6764;
	wire [4-1:0] node6768;
	wire [4-1:0] node6769;
	wire [4-1:0] node6770;
	wire [4-1:0] node6771;
	wire [4-1:0] node6772;
	wire [4-1:0] node6776;
	wire [4-1:0] node6779;
	wire [4-1:0] node6780;
	wire [4-1:0] node6782;
	wire [4-1:0] node6786;
	wire [4-1:0] node6787;
	wire [4-1:0] node6789;
	wire [4-1:0] node6791;
	wire [4-1:0] node6794;
	wire [4-1:0] node6795;
	wire [4-1:0] node6799;
	wire [4-1:0] node6800;
	wire [4-1:0] node6801;
	wire [4-1:0] node6802;
	wire [4-1:0] node6803;
	wire [4-1:0] node6805;
	wire [4-1:0] node6808;
	wire [4-1:0] node6809;
	wire [4-1:0] node6813;
	wire [4-1:0] node6814;
	wire [4-1:0] node6815;
	wire [4-1:0] node6816;
	wire [4-1:0] node6820;
	wire [4-1:0] node6823;
	wire [4-1:0] node6824;
	wire [4-1:0] node6828;
	wire [4-1:0] node6829;
	wire [4-1:0] node6832;
	wire [4-1:0] node6833;
	wire [4-1:0] node6834;
	wire [4-1:0] node6835;
	wire [4-1:0] node6840;
	wire [4-1:0] node6841;
	wire [4-1:0] node6842;
	wire [4-1:0] node6845;
	wire [4-1:0] node6849;
	wire [4-1:0] node6850;
	wire [4-1:0] node6851;
	wire [4-1:0] node6852;
	wire [4-1:0] node6854;
	wire [4-1:0] node6855;
	wire [4-1:0] node6859;
	wire [4-1:0] node6862;
	wire [4-1:0] node6863;
	wire [4-1:0] node6865;
	wire [4-1:0] node6868;
	wire [4-1:0] node6869;
	wire [4-1:0] node6872;
	wire [4-1:0] node6875;
	wire [4-1:0] node6876;
	wire [4-1:0] node6877;
	wire [4-1:0] node6878;
	wire [4-1:0] node6881;
	wire [4-1:0] node6882;
	wire [4-1:0] node6885;
	wire [4-1:0] node6888;
	wire [4-1:0] node6889;
	wire [4-1:0] node6891;
	wire [4-1:0] node6895;
	wire [4-1:0] node6896;
	wire [4-1:0] node6898;
	wire [4-1:0] node6899;
	wire [4-1:0] node6903;
	wire [4-1:0] node6905;
	wire [4-1:0] node6906;
	wire [4-1:0] node6910;
	wire [4-1:0] node6911;
	wire [4-1:0] node6912;
	wire [4-1:0] node6913;
	wire [4-1:0] node6914;
	wire [4-1:0] node6915;
	wire [4-1:0] node6916;
	wire [4-1:0] node6917;
	wire [4-1:0] node6919;
	wire [4-1:0] node6922;
	wire [4-1:0] node6924;
	wire [4-1:0] node6927;
	wire [4-1:0] node6928;
	wire [4-1:0] node6930;
	wire [4-1:0] node6932;
	wire [4-1:0] node6935;
	wire [4-1:0] node6937;
	wire [4-1:0] node6940;
	wire [4-1:0] node6941;
	wire [4-1:0] node6942;
	wire [4-1:0] node6943;
	wire [4-1:0] node6946;
	wire [4-1:0] node6949;
	wire [4-1:0] node6950;
	wire [4-1:0] node6954;
	wire [4-1:0] node6955;
	wire [4-1:0] node6957;
	wire [4-1:0] node6958;
	wire [4-1:0] node6961;
	wire [4-1:0] node6964;
	wire [4-1:0] node6966;
	wire [4-1:0] node6969;
	wire [4-1:0] node6970;
	wire [4-1:0] node6971;
	wire [4-1:0] node6972;
	wire [4-1:0] node6974;
	wire [4-1:0] node6978;
	wire [4-1:0] node6979;
	wire [4-1:0] node6981;
	wire [4-1:0] node6984;
	wire [4-1:0] node6985;
	wire [4-1:0] node6987;
	wire [4-1:0] node6990;
	wire [4-1:0] node6991;
	wire [4-1:0] node6995;
	wire [4-1:0] node6996;
	wire [4-1:0] node6997;
	wire [4-1:0] node7000;
	wire [4-1:0] node7003;
	wire [4-1:0] node7004;
	wire [4-1:0] node7007;
	wire [4-1:0] node7009;
	wire [4-1:0] node7010;
	wire [4-1:0] node7013;
	wire [4-1:0] node7016;
	wire [4-1:0] node7017;
	wire [4-1:0] node7018;
	wire [4-1:0] node7019;
	wire [4-1:0] node7020;
	wire [4-1:0] node7021;
	wire [4-1:0] node7025;
	wire [4-1:0] node7028;
	wire [4-1:0] node7029;
	wire [4-1:0] node7031;
	wire [4-1:0] node7034;
	wire [4-1:0] node7037;
	wire [4-1:0] node7038;
	wire [4-1:0] node7039;
	wire [4-1:0] node7040;
	wire [4-1:0] node7045;
	wire [4-1:0] node7046;
	wire [4-1:0] node7047;
	wire [4-1:0] node7048;
	wire [4-1:0] node7052;
	wire [4-1:0] node7054;
	wire [4-1:0] node7057;
	wire [4-1:0] node7060;
	wire [4-1:0] node7061;
	wire [4-1:0] node7062;
	wire [4-1:0] node7063;
	wire [4-1:0] node7064;
	wire [4-1:0] node7066;
	wire [4-1:0] node7070;
	wire [4-1:0] node7071;
	wire [4-1:0] node7072;
	wire [4-1:0] node7075;
	wire [4-1:0] node7078;
	wire [4-1:0] node7079;
	wire [4-1:0] node7083;
	wire [4-1:0] node7084;
	wire [4-1:0] node7086;
	wire [4-1:0] node7088;
	wire [4-1:0] node7091;
	wire [4-1:0] node7092;
	wire [4-1:0] node7095;
	wire [4-1:0] node7098;
	wire [4-1:0] node7099;
	wire [4-1:0] node7100;
	wire [4-1:0] node7102;
	wire [4-1:0] node7105;
	wire [4-1:0] node7107;
	wire [4-1:0] node7110;
	wire [4-1:0] node7112;
	wire [4-1:0] node7114;
	wire [4-1:0] node7117;
	wire [4-1:0] node7118;
	wire [4-1:0] node7119;
	wire [4-1:0] node7120;
	wire [4-1:0] node7121;
	wire [4-1:0] node7122;
	wire [4-1:0] node7125;
	wire [4-1:0] node7127;
	wire [4-1:0] node7130;
	wire [4-1:0] node7132;
	wire [4-1:0] node7133;
	wire [4-1:0] node7136;
	wire [4-1:0] node7139;
	wire [4-1:0] node7140;
	wire [4-1:0] node7141;
	wire [4-1:0] node7143;
	wire [4-1:0] node7145;
	wire [4-1:0] node7148;
	wire [4-1:0] node7149;
	wire [4-1:0] node7151;
	wire [4-1:0] node7154;
	wire [4-1:0] node7157;
	wire [4-1:0] node7158;
	wire [4-1:0] node7161;
	wire [4-1:0] node7162;
	wire [4-1:0] node7166;
	wire [4-1:0] node7167;
	wire [4-1:0] node7168;
	wire [4-1:0] node7169;
	wire [4-1:0] node7170;
	wire [4-1:0] node7174;
	wire [4-1:0] node7175;
	wire [4-1:0] node7178;
	wire [4-1:0] node7179;
	wire [4-1:0] node7182;
	wire [4-1:0] node7185;
	wire [4-1:0] node7186;
	wire [4-1:0] node7188;
	wire [4-1:0] node7191;
	wire [4-1:0] node7194;
	wire [4-1:0] node7195;
	wire [4-1:0] node7197;
	wire [4-1:0] node7198;
	wire [4-1:0] node7200;
	wire [4-1:0] node7204;
	wire [4-1:0] node7205;
	wire [4-1:0] node7206;
	wire [4-1:0] node7210;
	wire [4-1:0] node7212;
	wire [4-1:0] node7215;
	wire [4-1:0] node7216;
	wire [4-1:0] node7217;
	wire [4-1:0] node7218;
	wire [4-1:0] node7219;
	wire [4-1:0] node7220;
	wire [4-1:0] node7223;
	wire [4-1:0] node7226;
	wire [4-1:0] node7227;
	wire [4-1:0] node7231;
	wire [4-1:0] node7232;
	wire [4-1:0] node7236;
	wire [4-1:0] node7237;
	wire [4-1:0] node7238;
	wire [4-1:0] node7239;
	wire [4-1:0] node7240;
	wire [4-1:0] node7243;
	wire [4-1:0] node7247;
	wire [4-1:0] node7249;
	wire [4-1:0] node7252;
	wire [4-1:0] node7254;
	wire [4-1:0] node7256;
	wire [4-1:0] node7259;
	wire [4-1:0] node7260;
	wire [4-1:0] node7261;
	wire [4-1:0] node7262;
	wire [4-1:0] node7264;
	wire [4-1:0] node7267;
	wire [4-1:0] node7269;
	wire [4-1:0] node7272;
	wire [4-1:0] node7273;
	wire [4-1:0] node7275;
	wire [4-1:0] node7276;
	wire [4-1:0] node7279;
	wire [4-1:0] node7282;
	wire [4-1:0] node7283;
	wire [4-1:0] node7286;
	wire [4-1:0] node7289;
	wire [4-1:0] node7290;
	wire [4-1:0] node7292;
	wire [4-1:0] node7295;
	wire [4-1:0] node7298;
	wire [4-1:0] node7299;
	wire [4-1:0] node7300;
	wire [4-1:0] node7301;
	wire [4-1:0] node7302;
	wire [4-1:0] node7303;
	wire [4-1:0] node7304;
	wire [4-1:0] node7306;
	wire [4-1:0] node7309;
	wire [4-1:0] node7310;
	wire [4-1:0] node7314;
	wire [4-1:0] node7315;
	wire [4-1:0] node7317;
	wire [4-1:0] node7318;
	wire [4-1:0] node7321;
	wire [4-1:0] node7324;
	wire [4-1:0] node7327;
	wire [4-1:0] node7328;
	wire [4-1:0] node7329;
	wire [4-1:0] node7330;
	wire [4-1:0] node7334;
	wire [4-1:0] node7335;
	wire [4-1:0] node7337;
	wire [4-1:0] node7341;
	wire [4-1:0] node7342;
	wire [4-1:0] node7344;
	wire [4-1:0] node7345;
	wire [4-1:0] node7349;
	wire [4-1:0] node7351;
	wire [4-1:0] node7354;
	wire [4-1:0] node7355;
	wire [4-1:0] node7356;
	wire [4-1:0] node7358;
	wire [4-1:0] node7359;
	wire [4-1:0] node7363;
	wire [4-1:0] node7364;
	wire [4-1:0] node7367;
	wire [4-1:0] node7368;
	wire [4-1:0] node7369;
	wire [4-1:0] node7374;
	wire [4-1:0] node7375;
	wire [4-1:0] node7376;
	wire [4-1:0] node7378;
	wire [4-1:0] node7380;
	wire [4-1:0] node7383;
	wire [4-1:0] node7384;
	wire [4-1:0] node7385;
	wire [4-1:0] node7388;
	wire [4-1:0] node7391;
	wire [4-1:0] node7392;
	wire [4-1:0] node7396;
	wire [4-1:0] node7397;
	wire [4-1:0] node7398;
	wire [4-1:0] node7402;
	wire [4-1:0] node7403;
	wire [4-1:0] node7407;
	wire [4-1:0] node7408;
	wire [4-1:0] node7409;
	wire [4-1:0] node7410;
	wire [4-1:0] node7412;
	wire [4-1:0] node7413;
	wire [4-1:0] node7416;
	wire [4-1:0] node7419;
	wire [4-1:0] node7420;
	wire [4-1:0] node7421;
	wire [4-1:0] node7426;
	wire [4-1:0] node7427;
	wire [4-1:0] node7428;
	wire [4-1:0] node7430;
	wire [4-1:0] node7433;
	wire [4-1:0] node7434;
	wire [4-1:0] node7437;
	wire [4-1:0] node7440;
	wire [4-1:0] node7442;
	wire [4-1:0] node7443;
	wire [4-1:0] node7447;
	wire [4-1:0] node7448;
	wire [4-1:0] node7449;
	wire [4-1:0] node7450;
	wire [4-1:0] node7451;
	wire [4-1:0] node7454;
	wire [4-1:0] node7457;
	wire [4-1:0] node7459;
	wire [4-1:0] node7462;
	wire [4-1:0] node7463;
	wire [4-1:0] node7464;
	wire [4-1:0] node7469;
	wire [4-1:0] node7470;
	wire [4-1:0] node7471;
	wire [4-1:0] node7474;
	wire [4-1:0] node7477;
	wire [4-1:0] node7479;
	wire [4-1:0] node7480;
	wire [4-1:0] node7483;
	wire [4-1:0] node7486;
	wire [4-1:0] node7487;
	wire [4-1:0] node7488;
	wire [4-1:0] node7489;
	wire [4-1:0] node7490;
	wire [4-1:0] node7491;
	wire [4-1:0] node7492;
	wire [4-1:0] node7493;
	wire [4-1:0] node7496;
	wire [4-1:0] node7500;
	wire [4-1:0] node7502;
	wire [4-1:0] node7504;
	wire [4-1:0] node7507;
	wire [4-1:0] node7508;
	wire [4-1:0] node7509;
	wire [4-1:0] node7511;
	wire [4-1:0] node7514;
	wire [4-1:0] node7515;
	wire [4-1:0] node7518;
	wire [4-1:0] node7522;
	wire [4-1:0] node7523;
	wire [4-1:0] node7524;
	wire [4-1:0] node7525;
	wire [4-1:0] node7529;
	wire [4-1:0] node7531;
	wire [4-1:0] node7534;
	wire [4-1:0] node7536;
	wire [4-1:0] node7537;
	wire [4-1:0] node7540;
	wire [4-1:0] node7543;
	wire [4-1:0] node7544;
	wire [4-1:0] node7545;
	wire [4-1:0] node7546;
	wire [4-1:0] node7547;
	wire [4-1:0] node7550;
	wire [4-1:0] node7553;
	wire [4-1:0] node7555;
	wire [4-1:0] node7556;
	wire [4-1:0] node7559;
	wire [4-1:0] node7562;
	wire [4-1:0] node7563;
	wire [4-1:0] node7564;
	wire [4-1:0] node7565;
	wire [4-1:0] node7569;
	wire [4-1:0] node7570;
	wire [4-1:0] node7574;
	wire [4-1:0] node7576;
	wire [4-1:0] node7579;
	wire [4-1:0] node7580;
	wire [4-1:0] node7581;
	wire [4-1:0] node7582;
	wire [4-1:0] node7583;
	wire [4-1:0] node7588;
	wire [4-1:0] node7591;
	wire [4-1:0] node7592;
	wire [4-1:0] node7593;
	wire [4-1:0] node7594;
	wire [4-1:0] node7598;
	wire [4-1:0] node7599;
	wire [4-1:0] node7602;
	wire [4-1:0] node7606;
	wire [4-1:0] node7607;
	wire [4-1:0] node7608;
	wire [4-1:0] node7609;
	wire [4-1:0] node7610;
	wire [4-1:0] node7611;
	wire [4-1:0] node7614;
	wire [4-1:0] node7617;
	wire [4-1:0] node7618;
	wire [4-1:0] node7622;
	wire [4-1:0] node7623;
	wire [4-1:0] node7625;
	wire [4-1:0] node7629;
	wire [4-1:0] node7630;
	wire [4-1:0] node7631;
	wire [4-1:0] node7635;
	wire [4-1:0] node7637;
	wire [4-1:0] node7640;
	wire [4-1:0] node7641;
	wire [4-1:0] node7642;
	wire [4-1:0] node7643;
	wire [4-1:0] node7644;
	wire [4-1:0] node7648;
	wire [4-1:0] node7649;
	wire [4-1:0] node7650;
	wire [4-1:0] node7654;
	wire [4-1:0] node7657;
	wire [4-1:0] node7658;
	wire [4-1:0] node7659;
	wire [4-1:0] node7663;
	wire [4-1:0] node7664;
	wire [4-1:0] node7665;
	wire [4-1:0] node7669;
	wire [4-1:0] node7670;
	wire [4-1:0] node7673;
	wire [4-1:0] node7676;
	wire [4-1:0] node7677;
	wire [4-1:0] node7679;
	wire [4-1:0] node7680;
	wire [4-1:0] node7681;
	wire [4-1:0] node7686;
	wire [4-1:0] node7687;
	wire [4-1:0] node7689;
	wire [4-1:0] node7690;
	wire [4-1:0] node7694;
	wire [4-1:0] node7695;
	wire [4-1:0] node7698;
	wire [4-1:0] node7701;
	wire [4-1:0] node7702;
	wire [4-1:0] node7703;
	wire [4-1:0] node7704;
	wire [4-1:0] node7705;
	wire [4-1:0] node7706;
	wire [4-1:0] node7707;
	wire [4-1:0] node7708;
	wire [4-1:0] node7709;
	wire [4-1:0] node7710;
	wire [4-1:0] node7712;
	wire [4-1:0] node7716;
	wire [4-1:0] node7718;
	wire [4-1:0] node7720;
	wire [4-1:0] node7723;
	wire [4-1:0] node7724;
	wire [4-1:0] node7726;
	wire [4-1:0] node7729;
	wire [4-1:0] node7731;
	wire [4-1:0] node7734;
	wire [4-1:0] node7735;
	wire [4-1:0] node7736;
	wire [4-1:0] node7739;
	wire [4-1:0] node7740;
	wire [4-1:0] node7743;
	wire [4-1:0] node7745;
	wire [4-1:0] node7748;
	wire [4-1:0] node7749;
	wire [4-1:0] node7751;
	wire [4-1:0] node7753;
	wire [4-1:0] node7756;
	wire [4-1:0] node7758;
	wire [4-1:0] node7759;
	wire [4-1:0] node7762;
	wire [4-1:0] node7765;
	wire [4-1:0] node7766;
	wire [4-1:0] node7767;
	wire [4-1:0] node7769;
	wire [4-1:0] node7770;
	wire [4-1:0] node7773;
	wire [4-1:0] node7776;
	wire [4-1:0] node7777;
	wire [4-1:0] node7778;
	wire [4-1:0] node7782;
	wire [4-1:0] node7785;
	wire [4-1:0] node7786;
	wire [4-1:0] node7787;
	wire [4-1:0] node7790;
	wire [4-1:0] node7791;
	wire [4-1:0] node7795;
	wire [4-1:0] node7796;
	wire [4-1:0] node7797;
	wire [4-1:0] node7800;
	wire [4-1:0] node7804;
	wire [4-1:0] node7805;
	wire [4-1:0] node7806;
	wire [4-1:0] node7807;
	wire [4-1:0] node7808;
	wire [4-1:0] node7810;
	wire [4-1:0] node7813;
	wire [4-1:0] node7814;
	wire [4-1:0] node7817;
	wire [4-1:0] node7820;
	wire [4-1:0] node7821;
	wire [4-1:0] node7822;
	wire [4-1:0] node7826;
	wire [4-1:0] node7829;
	wire [4-1:0] node7830;
	wire [4-1:0] node7832;
	wire [4-1:0] node7833;
	wire [4-1:0] node7837;
	wire [4-1:0] node7838;
	wire [4-1:0] node7841;
	wire [4-1:0] node7843;
	wire [4-1:0] node7844;
	wire [4-1:0] node7847;
	wire [4-1:0] node7850;
	wire [4-1:0] node7851;
	wire [4-1:0] node7852;
	wire [4-1:0] node7853;
	wire [4-1:0] node7855;
	wire [4-1:0] node7858;
	wire [4-1:0] node7861;
	wire [4-1:0] node7862;
	wire [4-1:0] node7864;
	wire [4-1:0] node7866;
	wire [4-1:0] node7870;
	wire [4-1:0] node7871;
	wire [4-1:0] node7873;
	wire [4-1:0] node7874;
	wire [4-1:0] node7875;
	wire [4-1:0] node7879;
	wire [4-1:0] node7881;
	wire [4-1:0] node7884;
	wire [4-1:0] node7885;
	wire [4-1:0] node7886;
	wire [4-1:0] node7889;
	wire [4-1:0] node7892;
	wire [4-1:0] node7893;
	wire [4-1:0] node7897;
	wire [4-1:0] node7898;
	wire [4-1:0] node7899;
	wire [4-1:0] node7900;
	wire [4-1:0] node7901;
	wire [4-1:0] node7902;
	wire [4-1:0] node7904;
	wire [4-1:0] node7907;
	wire [4-1:0] node7908;
	wire [4-1:0] node7911;
	wire [4-1:0] node7914;
	wire [4-1:0] node7915;
	wire [4-1:0] node7917;
	wire [4-1:0] node7918;
	wire [4-1:0] node7922;
	wire [4-1:0] node7923;
	wire [4-1:0] node7926;
	wire [4-1:0] node7929;
	wire [4-1:0] node7930;
	wire [4-1:0] node7931;
	wire [4-1:0] node7932;
	wire [4-1:0] node7934;
	wire [4-1:0] node7937;
	wire [4-1:0] node7938;
	wire [4-1:0] node7942;
	wire [4-1:0] node7943;
	wire [4-1:0] node7947;
	wire [4-1:0] node7948;
	wire [4-1:0] node7949;
	wire [4-1:0] node7953;
	wire [4-1:0] node7955;
	wire [4-1:0] node7958;
	wire [4-1:0] node7959;
	wire [4-1:0] node7960;
	wire [4-1:0] node7961;
	wire [4-1:0] node7964;
	wire [4-1:0] node7965;
	wire [4-1:0] node7966;
	wire [4-1:0] node7969;
	wire [4-1:0] node7972;
	wire [4-1:0] node7974;
	wire [4-1:0] node7977;
	wire [4-1:0] node7978;
	wire [4-1:0] node7979;
	wire [4-1:0] node7984;
	wire [4-1:0] node7985;
	wire [4-1:0] node7986;
	wire [4-1:0] node7987;
	wire [4-1:0] node7989;
	wire [4-1:0] node7992;
	wire [4-1:0] node7995;
	wire [4-1:0] node7996;
	wire [4-1:0] node7998;
	wire [4-1:0] node8001;
	wire [4-1:0] node8002;
	wire [4-1:0] node8006;
	wire [4-1:0] node8007;
	wire [4-1:0] node8008;
	wire [4-1:0] node8010;
	wire [4-1:0] node8014;
	wire [4-1:0] node8017;
	wire [4-1:0] node8018;
	wire [4-1:0] node8019;
	wire [4-1:0] node8020;
	wire [4-1:0] node8022;
	wire [4-1:0] node8023;
	wire [4-1:0] node8026;
	wire [4-1:0] node8029;
	wire [4-1:0] node8030;
	wire [4-1:0] node8031;
	wire [4-1:0] node8033;
	wire [4-1:0] node8037;
	wire [4-1:0] node8038;
	wire [4-1:0] node8039;
	wire [4-1:0] node8042;
	wire [4-1:0] node8046;
	wire [4-1:0] node8047;
	wire [4-1:0] node8048;
	wire [4-1:0] node8049;
	wire [4-1:0] node8050;
	wire [4-1:0] node8053;
	wire [4-1:0] node8056;
	wire [4-1:0] node8057;
	wire [4-1:0] node8060;
	wire [4-1:0] node8063;
	wire [4-1:0] node8065;
	wire [4-1:0] node8068;
	wire [4-1:0] node8069;
	wire [4-1:0] node8073;
	wire [4-1:0] node8074;
	wire [4-1:0] node8075;
	wire [4-1:0] node8076;
	wire [4-1:0] node8077;
	wire [4-1:0] node8081;
	wire [4-1:0] node8082;
	wire [4-1:0] node8084;
	wire [4-1:0] node8088;
	wire [4-1:0] node8089;
	wire [4-1:0] node8090;
	wire [4-1:0] node8093;
	wire [4-1:0] node8096;
	wire [4-1:0] node8099;
	wire [4-1:0] node8100;
	wire [4-1:0] node8103;
	wire [4-1:0] node8105;
	wire [4-1:0] node8106;
	wire [4-1:0] node8107;
	wire [4-1:0] node8110;
	wire [4-1:0] node8114;
	wire [4-1:0] node8115;
	wire [4-1:0] node8116;
	wire [4-1:0] node8117;
	wire [4-1:0] node8118;
	wire [4-1:0] node8119;
	wire [4-1:0] node8120;
	wire [4-1:0] node8121;
	wire [4-1:0] node8123;
	wire [4-1:0] node8126;
	wire [4-1:0] node8127;
	wire [4-1:0] node8130;
	wire [4-1:0] node8133;
	wire [4-1:0] node8136;
	wire [4-1:0] node8137;
	wire [4-1:0] node8139;
	wire [4-1:0] node8142;
	wire [4-1:0] node8145;
	wire [4-1:0] node8146;
	wire [4-1:0] node8147;
	wire [4-1:0] node8149;
	wire [4-1:0] node8150;
	wire [4-1:0] node8154;
	wire [4-1:0] node8156;
	wire [4-1:0] node8157;
	wire [4-1:0] node8161;
	wire [4-1:0] node8162;
	wire [4-1:0] node8164;
	wire [4-1:0] node8167;
	wire [4-1:0] node8168;
	wire [4-1:0] node8170;
	wire [4-1:0] node8174;
	wire [4-1:0] node8175;
	wire [4-1:0] node8176;
	wire [4-1:0] node8179;
	wire [4-1:0] node8180;
	wire [4-1:0] node8181;
	wire [4-1:0] node8186;
	wire [4-1:0] node8187;
	wire [4-1:0] node8188;
	wire [4-1:0] node8189;
	wire [4-1:0] node8192;
	wire [4-1:0] node8195;
	wire [4-1:0] node8196;
	wire [4-1:0] node8199;
	wire [4-1:0] node8200;
	wire [4-1:0] node8204;
	wire [4-1:0] node8205;
	wire [4-1:0] node8207;
	wire [4-1:0] node8209;
	wire [4-1:0] node8212;
	wire [4-1:0] node8214;
	wire [4-1:0] node8217;
	wire [4-1:0] node8218;
	wire [4-1:0] node8219;
	wire [4-1:0] node8220;
	wire [4-1:0] node8221;
	wire [4-1:0] node8224;
	wire [4-1:0] node8227;
	wire [4-1:0] node8228;
	wire [4-1:0] node8229;
	wire [4-1:0] node8232;
	wire [4-1:0] node8235;
	wire [4-1:0] node8238;
	wire [4-1:0] node8239;
	wire [4-1:0] node8240;
	wire [4-1:0] node8241;
	wire [4-1:0] node8244;
	wire [4-1:0] node8247;
	wire [4-1:0] node8248;
	wire [4-1:0] node8252;
	wire [4-1:0] node8254;
	wire [4-1:0] node8255;
	wire [4-1:0] node8256;
	wire [4-1:0] node8260;
	wire [4-1:0] node8263;
	wire [4-1:0] node8264;
	wire [4-1:0] node8265;
	wire [4-1:0] node8266;
	wire [4-1:0] node8267;
	wire [4-1:0] node8270;
	wire [4-1:0] node8273;
	wire [4-1:0] node8274;
	wire [4-1:0] node8278;
	wire [4-1:0] node8279;
	wire [4-1:0] node8280;
	wire [4-1:0] node8283;
	wire [4-1:0] node8286;
	wire [4-1:0] node8288;
	wire [4-1:0] node8290;
	wire [4-1:0] node8293;
	wire [4-1:0] node8294;
	wire [4-1:0] node8295;
	wire [4-1:0] node8296;
	wire [4-1:0] node8300;
	wire [4-1:0] node8303;
	wire [4-1:0] node8304;
	wire [4-1:0] node8306;
	wire [4-1:0] node8307;
	wire [4-1:0] node8311;
	wire [4-1:0] node8312;
	wire [4-1:0] node8315;
	wire [4-1:0] node8316;
	wire [4-1:0] node8320;
	wire [4-1:0] node8321;
	wire [4-1:0] node8322;
	wire [4-1:0] node8323;
	wire [4-1:0] node8324;
	wire [4-1:0] node8325;
	wire [4-1:0] node8327;
	wire [4-1:0] node8330;
	wire [4-1:0] node8331;
	wire [4-1:0] node8334;
	wire [4-1:0] node8335;
	wire [4-1:0] node8338;
	wire [4-1:0] node8341;
	wire [4-1:0] node8342;
	wire [4-1:0] node8343;
	wire [4-1:0] node8344;
	wire [4-1:0] node8348;
	wire [4-1:0] node8349;
	wire [4-1:0] node8353;
	wire [4-1:0] node8356;
	wire [4-1:0] node8357;
	wire [4-1:0] node8359;
	wire [4-1:0] node8360;
	wire [4-1:0] node8364;
	wire [4-1:0] node8365;
	wire [4-1:0] node8368;
	wire [4-1:0] node8369;
	wire [4-1:0] node8371;
	wire [4-1:0] node8375;
	wire [4-1:0] node8376;
	wire [4-1:0] node8377;
	wire [4-1:0] node8379;
	wire [4-1:0] node8382;
	wire [4-1:0] node8384;
	wire [4-1:0] node8387;
	wire [4-1:0] node8388;
	wire [4-1:0] node8389;
	wire [4-1:0] node8391;
	wire [4-1:0] node8394;
	wire [4-1:0] node8396;
	wire [4-1:0] node8398;
	wire [4-1:0] node8401;
	wire [4-1:0] node8402;
	wire [4-1:0] node8403;
	wire [4-1:0] node8404;
	wire [4-1:0] node8409;
	wire [4-1:0] node8410;
	wire [4-1:0] node8414;
	wire [4-1:0] node8415;
	wire [4-1:0] node8416;
	wire [4-1:0] node8417;
	wire [4-1:0] node8418;
	wire [4-1:0] node8420;
	wire [4-1:0] node8422;
	wire [4-1:0] node8425;
	wire [4-1:0] node8428;
	wire [4-1:0] node8429;
	wire [4-1:0] node8430;
	wire [4-1:0] node8433;
	wire [4-1:0] node8436;
	wire [4-1:0] node8437;
	wire [4-1:0] node8440;
	wire [4-1:0] node8443;
	wire [4-1:0] node8444;
	wire [4-1:0] node8445;
	wire [4-1:0] node8448;
	wire [4-1:0] node8450;
	wire [4-1:0] node8453;
	wire [4-1:0] node8454;
	wire [4-1:0] node8456;
	wire [4-1:0] node8459;
	wire [4-1:0] node8461;
	wire [4-1:0] node8462;
	wire [4-1:0] node8466;
	wire [4-1:0] node8467;
	wire [4-1:0] node8468;
	wire [4-1:0] node8469;
	wire [4-1:0] node8470;
	wire [4-1:0] node8473;
	wire [4-1:0] node8476;
	wire [4-1:0] node8479;
	wire [4-1:0] node8480;
	wire [4-1:0] node8482;
	wire [4-1:0] node8483;
	wire [4-1:0] node8486;
	wire [4-1:0] node8489;
	wire [4-1:0] node8490;
	wire [4-1:0] node8491;
	wire [4-1:0] node8495;
	wire [4-1:0] node8497;
	wire [4-1:0] node8500;
	wire [4-1:0] node8501;
	wire [4-1:0] node8502;
	wire [4-1:0] node8503;
	wire [4-1:0] node8505;
	wire [4-1:0] node8509;
	wire [4-1:0] node8510;
	wire [4-1:0] node8511;
	wire [4-1:0] node8515;
	wire [4-1:0] node8517;
	wire [4-1:0] node8520;
	wire [4-1:0] node8521;
	wire [4-1:0] node8523;
	wire [4-1:0] node8526;
	wire [4-1:0] node8529;
	wire [4-1:0] node8530;
	wire [4-1:0] node8531;
	wire [4-1:0] node8532;
	wire [4-1:0] node8533;
	wire [4-1:0] node8534;
	wire [4-1:0] node8535;
	wire [4-1:0] node8536;
	wire [4-1:0] node8538;
	wire [4-1:0] node8541;
	wire [4-1:0] node8543;
	wire [4-1:0] node8546;
	wire [4-1:0] node8547;
	wire [4-1:0] node8548;
	wire [4-1:0] node8550;
	wire [4-1:0] node8554;
	wire [4-1:0] node8556;
	wire [4-1:0] node8559;
	wire [4-1:0] node8560;
	wire [4-1:0] node8561;
	wire [4-1:0] node8563;
	wire [4-1:0] node8564;
	wire [4-1:0] node8568;
	wire [4-1:0] node8569;
	wire [4-1:0] node8570;
	wire [4-1:0] node8574;
	wire [4-1:0] node8575;
	wire [4-1:0] node8578;
	wire [4-1:0] node8581;
	wire [4-1:0] node8582;
	wire [4-1:0] node8583;
	wire [4-1:0] node8584;
	wire [4-1:0] node8587;
	wire [4-1:0] node8591;
	wire [4-1:0] node8592;
	wire [4-1:0] node8595;
	wire [4-1:0] node8598;
	wire [4-1:0] node8599;
	wire [4-1:0] node8600;
	wire [4-1:0] node8601;
	wire [4-1:0] node8603;
	wire [4-1:0] node8605;
	wire [4-1:0] node8608;
	wire [4-1:0] node8609;
	wire [4-1:0] node8610;
	wire [4-1:0] node8613;
	wire [4-1:0] node8616;
	wire [4-1:0] node8617;
	wire [4-1:0] node8621;
	wire [4-1:0] node8622;
	wire [4-1:0] node8624;
	wire [4-1:0] node8625;
	wire [4-1:0] node8628;
	wire [4-1:0] node8631;
	wire [4-1:0] node8633;
	wire [4-1:0] node8636;
	wire [4-1:0] node8637;
	wire [4-1:0] node8638;
	wire [4-1:0] node8641;
	wire [4-1:0] node8644;
	wire [4-1:0] node8646;
	wire [4-1:0] node8647;
	wire [4-1:0] node8650;
	wire [4-1:0] node8653;
	wire [4-1:0] node8654;
	wire [4-1:0] node8655;
	wire [4-1:0] node8656;
	wire [4-1:0] node8658;
	wire [4-1:0] node8659;
	wire [4-1:0] node8663;
	wire [4-1:0] node8664;
	wire [4-1:0] node8665;
	wire [4-1:0] node8669;
	wire [4-1:0] node8672;
	wire [4-1:0] node8673;
	wire [4-1:0] node8674;
	wire [4-1:0] node8677;
	wire [4-1:0] node8678;
	wire [4-1:0] node8681;
	wire [4-1:0] node8684;
	wire [4-1:0] node8685;
	wire [4-1:0] node8687;
	wire [4-1:0] node8689;
	wire [4-1:0] node8692;
	wire [4-1:0] node8693;
	wire [4-1:0] node8697;
	wire [4-1:0] node8698;
	wire [4-1:0] node8699;
	wire [4-1:0] node8700;
	wire [4-1:0] node8703;
	wire [4-1:0] node8705;
	wire [4-1:0] node8706;
	wire [4-1:0] node8709;
	wire [4-1:0] node8712;
	wire [4-1:0] node8713;
	wire [4-1:0] node8715;
	wire [4-1:0] node8718;
	wire [4-1:0] node8720;
	wire [4-1:0] node8721;
	wire [4-1:0] node8724;
	wire [4-1:0] node8727;
	wire [4-1:0] node8728;
	wire [4-1:0] node8729;
	wire [4-1:0] node8730;
	wire [4-1:0] node8733;
	wire [4-1:0] node8735;
	wire [4-1:0] node8738;
	wire [4-1:0] node8741;
	wire [4-1:0] node8743;
	wire [4-1:0] node8744;
	wire [4-1:0] node8748;
	wire [4-1:0] node8749;
	wire [4-1:0] node8750;
	wire [4-1:0] node8751;
	wire [4-1:0] node8752;
	wire [4-1:0] node8754;
	wire [4-1:0] node8755;
	wire [4-1:0] node8759;
	wire [4-1:0] node8760;
	wire [4-1:0] node8761;
	wire [4-1:0] node8765;
	wire [4-1:0] node8768;
	wire [4-1:0] node8769;
	wire [4-1:0] node8770;
	wire [4-1:0] node8772;
	wire [4-1:0] node8773;
	wire [4-1:0] node8776;
	wire [4-1:0] node8780;
	wire [4-1:0] node8781;
	wire [4-1:0] node8784;
	wire [4-1:0] node8787;
	wire [4-1:0] node8788;
	wire [4-1:0] node8789;
	wire [4-1:0] node8790;
	wire [4-1:0] node8793;
	wire [4-1:0] node8795;
	wire [4-1:0] node8798;
	wire [4-1:0] node8799;
	wire [4-1:0] node8800;
	wire [4-1:0] node8801;
	wire [4-1:0] node8804;
	wire [4-1:0] node8808;
	wire [4-1:0] node8809;
	wire [4-1:0] node8811;
	wire [4-1:0] node8815;
	wire [4-1:0] node8816;
	wire [4-1:0] node8817;
	wire [4-1:0] node8818;
	wire [4-1:0] node8820;
	wire [4-1:0] node8823;
	wire [4-1:0] node8824;
	wire [4-1:0] node8827;
	wire [4-1:0] node8830;
	wire [4-1:0] node8831;
	wire [4-1:0] node8834;
	wire [4-1:0] node8837;
	wire [4-1:0] node8838;
	wire [4-1:0] node8840;
	wire [4-1:0] node8842;
	wire [4-1:0] node8845;
	wire [4-1:0] node8848;
	wire [4-1:0] node8849;
	wire [4-1:0] node8850;
	wire [4-1:0] node8851;
	wire [4-1:0] node8852;
	wire [4-1:0] node8854;
	wire [4-1:0] node8857;
	wire [4-1:0] node8858;
	wire [4-1:0] node8862;
	wire [4-1:0] node8863;
	wire [4-1:0] node8864;
	wire [4-1:0] node8868;
	wire [4-1:0] node8870;
	wire [4-1:0] node8871;
	wire [4-1:0] node8874;
	wire [4-1:0] node8877;
	wire [4-1:0] node8878;
	wire [4-1:0] node8879;
	wire [4-1:0] node8882;
	wire [4-1:0] node8885;
	wire [4-1:0] node8887;
	wire [4-1:0] node8888;
	wire [4-1:0] node8891;
	wire [4-1:0] node8894;
	wire [4-1:0] node8895;
	wire [4-1:0] node8896;
	wire [4-1:0] node8897;
	wire [4-1:0] node8900;
	wire [4-1:0] node8903;
	wire [4-1:0] node8904;
	wire [4-1:0] node8907;
	wire [4-1:0] node8908;
	wire [4-1:0] node8912;
	wire [4-1:0] node8913;
	wire [4-1:0] node8914;
	wire [4-1:0] node8915;
	wire [4-1:0] node8918;
	wire [4-1:0] node8922;
	wire [4-1:0] node8923;
	wire [4-1:0] node8924;
	wire [4-1:0] node8928;
	wire [4-1:0] node8931;
	wire [4-1:0] node8932;
	wire [4-1:0] node8933;
	wire [4-1:0] node8934;
	wire [4-1:0] node8935;
	wire [4-1:0] node8936;
	wire [4-1:0] node8937;
	wire [4-1:0] node8940;
	wire [4-1:0] node8941;
	wire [4-1:0] node8945;
	wire [4-1:0] node8946;
	wire [4-1:0] node8947;
	wire [4-1:0] node8952;
	wire [4-1:0] node8953;
	wire [4-1:0] node8954;
	wire [4-1:0] node8955;
	wire [4-1:0] node8959;
	wire [4-1:0] node8961;
	wire [4-1:0] node8964;
	wire [4-1:0] node8966;
	wire [4-1:0] node8968;
	wire [4-1:0] node8971;
	wire [4-1:0] node8972;
	wire [4-1:0] node8973;
	wire [4-1:0] node8974;
	wire [4-1:0] node8975;
	wire [4-1:0] node8979;
	wire [4-1:0] node8980;
	wire [4-1:0] node8984;
	wire [4-1:0] node8985;
	wire [4-1:0] node8986;
	wire [4-1:0] node8990;
	wire [4-1:0] node8991;
	wire [4-1:0] node8992;
	wire [4-1:0] node8995;
	wire [4-1:0] node8999;
	wire [4-1:0] node9000;
	wire [4-1:0] node9002;
	wire [4-1:0] node9005;
	wire [4-1:0] node9006;
	wire [4-1:0] node9007;
	wire [4-1:0] node9011;
	wire [4-1:0] node9013;
	wire [4-1:0] node9014;
	wire [4-1:0] node9018;
	wire [4-1:0] node9019;
	wire [4-1:0] node9020;
	wire [4-1:0] node9021;
	wire [4-1:0] node9022;
	wire [4-1:0] node9023;
	wire [4-1:0] node9024;
	wire [4-1:0] node9028;
	wire [4-1:0] node9029;
	wire [4-1:0] node9035;
	wire [4-1:0] node9036;
	wire [4-1:0] node9037;
	wire [4-1:0] node9038;
	wire [4-1:0] node9039;
	wire [4-1:0] node9044;
	wire [4-1:0] node9045;
	wire [4-1:0] node9048;
	wire [4-1:0] node9051;
	wire [4-1:0] node9053;
	wire [4-1:0] node9054;
	wire [4-1:0] node9055;
	wire [4-1:0] node9060;
	wire [4-1:0] node9061;
	wire [4-1:0] node9062;
	wire [4-1:0] node9064;
	wire [4-1:0] node9067;
	wire [4-1:0] node9069;
	wire [4-1:0] node9072;
	wire [4-1:0] node9073;
	wire [4-1:0] node9074;
	wire [4-1:0] node9076;
	wire [4-1:0] node9079;
	wire [4-1:0] node9082;
	wire [4-1:0] node9083;
	wire [4-1:0] node9084;
	wire [4-1:0] node9085;
	wire [4-1:0] node9088;
	wire [4-1:0] node9092;
	wire [4-1:0] node9094;
	wire [4-1:0] node9097;
	wire [4-1:0] node9098;
	wire [4-1:0] node9099;
	wire [4-1:0] node9100;
	wire [4-1:0] node9101;
	wire [4-1:0] node9102;
	wire [4-1:0] node9105;
	wire [4-1:0] node9106;
	wire [4-1:0] node9108;
	wire [4-1:0] node9112;
	wire [4-1:0] node9114;
	wire [4-1:0] node9117;
	wire [4-1:0] node9118;
	wire [4-1:0] node9119;
	wire [4-1:0] node9120;
	wire [4-1:0] node9125;
	wire [4-1:0] node9126;
	wire [4-1:0] node9128;
	wire [4-1:0] node9131;
	wire [4-1:0] node9134;
	wire [4-1:0] node9135;
	wire [4-1:0] node9136;
	wire [4-1:0] node9137;
	wire [4-1:0] node9141;
	wire [4-1:0] node9143;
	wire [4-1:0] node9145;
	wire [4-1:0] node9148;
	wire [4-1:0] node9149;
	wire [4-1:0] node9152;
	wire [4-1:0] node9154;
	wire [4-1:0] node9157;
	wire [4-1:0] node9158;
	wire [4-1:0] node9159;
	wire [4-1:0] node9160;
	wire [4-1:0] node9161;
	wire [4-1:0] node9162;
	wire [4-1:0] node9164;
	wire [4-1:0] node9168;
	wire [4-1:0] node9171;
	wire [4-1:0] node9173;
	wire [4-1:0] node9175;
	wire [4-1:0] node9178;
	wire [4-1:0] node9179;
	wire [4-1:0] node9181;
	wire [4-1:0] node9182;
	wire [4-1:0] node9183;
	wire [4-1:0] node9186;
	wire [4-1:0] node9189;
	wire [4-1:0] node9191;
	wire [4-1:0] node9194;
	wire [4-1:0] node9195;
	wire [4-1:0] node9196;
	wire [4-1:0] node9199;
	wire [4-1:0] node9203;
	wire [4-1:0] node9204;
	wire [4-1:0] node9205;
	wire [4-1:0] node9206;
	wire [4-1:0] node9207;
	wire [4-1:0] node9208;
	wire [4-1:0] node9213;
	wire [4-1:0] node9214;
	wire [4-1:0] node9219;
	wire [4-1:0] node9220;
	wire [4-1:0] node9223;
	wire [4-1:0] node9224;
	wire [4-1:0] node9225;
	wire [4-1:0] node9226;
	wire [4-1:0] node9232;
	wire [4-1:0] node9233;
	wire [4-1:0] node9234;
	wire [4-1:0] node9235;
	wire [4-1:0] node9236;
	wire [4-1:0] node9237;
	wire [4-1:0] node9238;
	wire [4-1:0] node9239;
	wire [4-1:0] node9240;
	wire [4-1:0] node9241;
	wire [4-1:0] node9244;
	wire [4-1:0] node9246;
	wire [4-1:0] node9249;
	wire [4-1:0] node9251;
	wire [4-1:0] node9253;
	wire [4-1:0] node9256;
	wire [4-1:0] node9257;
	wire [4-1:0] node9258;
	wire [4-1:0] node9259;
	wire [4-1:0] node9261;
	wire [4-1:0] node9265;
	wire [4-1:0] node9268;
	wire [4-1:0] node9269;
	wire [4-1:0] node9270;
	wire [4-1:0] node9273;
	wire [4-1:0] node9276;
	wire [4-1:0] node9277;
	wire [4-1:0] node9279;
	wire [4-1:0] node9283;
	wire [4-1:0] node9284;
	wire [4-1:0] node9285;
	wire [4-1:0] node9286;
	wire [4-1:0] node9289;
	wire [4-1:0] node9292;
	wire [4-1:0] node9294;
	wire [4-1:0] node9295;
	wire [4-1:0] node9296;
	wire [4-1:0] node9299;
	wire [4-1:0] node9303;
	wire [4-1:0] node9304;
	wire [4-1:0] node9305;
	wire [4-1:0] node9307;
	wire [4-1:0] node9309;
	wire [4-1:0] node9312;
	wire [4-1:0] node9313;
	wire [4-1:0] node9315;
	wire [4-1:0] node9319;
	wire [4-1:0] node9320;
	wire [4-1:0] node9321;
	wire [4-1:0] node9324;
	wire [4-1:0] node9327;
	wire [4-1:0] node9329;
	wire [4-1:0] node9330;
	wire [4-1:0] node9333;
	wire [4-1:0] node9336;
	wire [4-1:0] node9337;
	wire [4-1:0] node9338;
	wire [4-1:0] node9339;
	wire [4-1:0] node9340;
	wire [4-1:0] node9341;
	wire [4-1:0] node9345;
	wire [4-1:0] node9347;
	wire [4-1:0] node9350;
	wire [4-1:0] node9351;
	wire [4-1:0] node9353;
	wire [4-1:0] node9355;
	wire [4-1:0] node9358;
	wire [4-1:0] node9360;
	wire [4-1:0] node9362;
	wire [4-1:0] node9365;
	wire [4-1:0] node9366;
	wire [4-1:0] node9367;
	wire [4-1:0] node9368;
	wire [4-1:0] node9370;
	wire [4-1:0] node9374;
	wire [4-1:0] node9377;
	wire [4-1:0] node9378;
	wire [4-1:0] node9380;
	wire [4-1:0] node9383;
	wire [4-1:0] node9384;
	wire [4-1:0] node9385;
	wire [4-1:0] node9388;
	wire [4-1:0] node9392;
	wire [4-1:0] node9393;
	wire [4-1:0] node9394;
	wire [4-1:0] node9395;
	wire [4-1:0] node9397;
	wire [4-1:0] node9400;
	wire [4-1:0] node9401;
	wire [4-1:0] node9404;
	wire [4-1:0] node9407;
	wire [4-1:0] node9408;
	wire [4-1:0] node9409;
	wire [4-1:0] node9411;
	wire [4-1:0] node9414;
	wire [4-1:0] node9417;
	wire [4-1:0] node9420;
	wire [4-1:0] node9421;
	wire [4-1:0] node9422;
	wire [4-1:0] node9425;
	wire [4-1:0] node9426;
	wire [4-1:0] node9428;
	wire [4-1:0] node9431;
	wire [4-1:0] node9433;
	wire [4-1:0] node9436;
	wire [4-1:0] node9437;
	wire [4-1:0] node9440;
	wire [4-1:0] node9441;
	wire [4-1:0] node9443;
	wire [4-1:0] node9447;
	wire [4-1:0] node9448;
	wire [4-1:0] node9449;
	wire [4-1:0] node9450;
	wire [4-1:0] node9451;
	wire [4-1:0] node9452;
	wire [4-1:0] node9453;
	wire [4-1:0] node9456;
	wire [4-1:0] node9459;
	wire [4-1:0] node9460;
	wire [4-1:0] node9463;
	wire [4-1:0] node9466;
	wire [4-1:0] node9467;
	wire [4-1:0] node9471;
	wire [4-1:0] node9472;
	wire [4-1:0] node9474;
	wire [4-1:0] node9476;
	wire [4-1:0] node9477;
	wire [4-1:0] node9481;
	wire [4-1:0] node9483;
	wire [4-1:0] node9485;
	wire [4-1:0] node9488;
	wire [4-1:0] node9489;
	wire [4-1:0] node9490;
	wire [4-1:0] node9491;
	wire [4-1:0] node9493;
	wire [4-1:0] node9496;
	wire [4-1:0] node9497;
	wire [4-1:0] node9498;
	wire [4-1:0] node9501;
	wire [4-1:0] node9505;
	wire [4-1:0] node9506;
	wire [4-1:0] node9508;
	wire [4-1:0] node9510;
	wire [4-1:0] node9513;
	wire [4-1:0] node9514;
	wire [4-1:0] node9517;
	wire [4-1:0] node9520;
	wire [4-1:0] node9521;
	wire [4-1:0] node9522;
	wire [4-1:0] node9523;
	wire [4-1:0] node9526;
	wire [4-1:0] node9527;
	wire [4-1:0] node9531;
	wire [4-1:0] node9532;
	wire [4-1:0] node9533;
	wire [4-1:0] node9537;
	wire [4-1:0] node9539;
	wire [4-1:0] node9542;
	wire [4-1:0] node9545;
	wire [4-1:0] node9546;
	wire [4-1:0] node9547;
	wire [4-1:0] node9548;
	wire [4-1:0] node9549;
	wire [4-1:0] node9550;
	wire [4-1:0] node9554;
	wire [4-1:0] node9555;
	wire [4-1:0] node9558;
	wire [4-1:0] node9561;
	wire [4-1:0] node9562;
	wire [4-1:0] node9563;
	wire [4-1:0] node9567;
	wire [4-1:0] node9568;
	wire [4-1:0] node9570;
	wire [4-1:0] node9573;
	wire [4-1:0] node9575;
	wire [4-1:0] node9578;
	wire [4-1:0] node9579;
	wire [4-1:0] node9580;
	wire [4-1:0] node9582;
	wire [4-1:0] node9583;
	wire [4-1:0] node9587;
	wire [4-1:0] node9589;
	wire [4-1:0] node9590;
	wire [4-1:0] node9593;
	wire [4-1:0] node9597;
	wire [4-1:0] node9598;
	wire [4-1:0] node9599;
	wire [4-1:0] node9600;
	wire [4-1:0] node9601;
	wire [4-1:0] node9602;
	wire [4-1:0] node9605;
	wire [4-1:0] node9608;
	wire [4-1:0] node9611;
	wire [4-1:0] node9612;
	wire [4-1:0] node9614;
	wire [4-1:0] node9618;
	wire [4-1:0] node9619;
	wire [4-1:0] node9620;
	wire [4-1:0] node9621;
	wire [4-1:0] node9626;
	wire [4-1:0] node9627;
	wire [4-1:0] node9631;
	wire [4-1:0] node9632;
	wire [4-1:0] node9634;
	wire [4-1:0] node9636;
	wire [4-1:0] node9639;
	wire [4-1:0] node9640;
	wire [4-1:0] node9641;
	wire [4-1:0] node9642;
	wire [4-1:0] node9647;
	wire [4-1:0] node9648;
	wire [4-1:0] node9650;
	wire [4-1:0] node9654;
	wire [4-1:0] node9655;
	wire [4-1:0] node9656;
	wire [4-1:0] node9657;
	wire [4-1:0] node9658;
	wire [4-1:0] node9659;
	wire [4-1:0] node9661;
	wire [4-1:0] node9663;
	wire [4-1:0] node9665;
	wire [4-1:0] node9668;
	wire [4-1:0] node9669;
	wire [4-1:0] node9672;
	wire [4-1:0] node9673;
	wire [4-1:0] node9675;
	wire [4-1:0] node9678;
	wire [4-1:0] node9680;
	wire [4-1:0] node9683;
	wire [4-1:0] node9684;
	wire [4-1:0] node9685;
	wire [4-1:0] node9686;
	wire [4-1:0] node9689;
	wire [4-1:0] node9692;
	wire [4-1:0] node9693;
	wire [4-1:0] node9694;
	wire [4-1:0] node9697;
	wire [4-1:0] node9701;
	wire [4-1:0] node9702;
	wire [4-1:0] node9704;
	wire [4-1:0] node9705;
	wire [4-1:0] node9709;
	wire [4-1:0] node9712;
	wire [4-1:0] node9713;
	wire [4-1:0] node9714;
	wire [4-1:0] node9715;
	wire [4-1:0] node9717;
	wire [4-1:0] node9721;
	wire [4-1:0] node9722;
	wire [4-1:0] node9725;
	wire [4-1:0] node9726;
	wire [4-1:0] node9727;
	wire [4-1:0] node9732;
	wire [4-1:0] node9733;
	wire [4-1:0] node9735;
	wire [4-1:0] node9737;
	wire [4-1:0] node9740;
	wire [4-1:0] node9741;
	wire [4-1:0] node9743;
	wire [4-1:0] node9746;
	wire [4-1:0] node9747;
	wire [4-1:0] node9748;
	wire [4-1:0] node9751;
	wire [4-1:0] node9755;
	wire [4-1:0] node9756;
	wire [4-1:0] node9757;
	wire [4-1:0] node9758;
	wire [4-1:0] node9759;
	wire [4-1:0] node9760;
	wire [4-1:0] node9763;
	wire [4-1:0] node9766;
	wire [4-1:0] node9767;
	wire [4-1:0] node9770;
	wire [4-1:0] node9773;
	wire [4-1:0] node9775;
	wire [4-1:0] node9776;
	wire [4-1:0] node9780;
	wire [4-1:0] node9781;
	wire [4-1:0] node9782;
	wire [4-1:0] node9783;
	wire [4-1:0] node9785;
	wire [4-1:0] node9789;
	wire [4-1:0] node9790;
	wire [4-1:0] node9791;
	wire [4-1:0] node9796;
	wire [4-1:0] node9797;
	wire [4-1:0] node9800;
	wire [4-1:0] node9803;
	wire [4-1:0] node9804;
	wire [4-1:0] node9805;
	wire [4-1:0] node9807;
	wire [4-1:0] node9808;
	wire [4-1:0] node9810;
	wire [4-1:0] node9813;
	wire [4-1:0] node9814;
	wire [4-1:0] node9817;
	wire [4-1:0] node9820;
	wire [4-1:0] node9821;
	wire [4-1:0] node9822;
	wire [4-1:0] node9824;
	wire [4-1:0] node9827;
	wire [4-1:0] node9828;
	wire [4-1:0] node9832;
	wire [4-1:0] node9833;
	wire [4-1:0] node9834;
	wire [4-1:0] node9839;
	wire [4-1:0] node9840;
	wire [4-1:0] node9841;
	wire [4-1:0] node9843;
	wire [4-1:0] node9844;
	wire [4-1:0] node9847;
	wire [4-1:0] node9850;
	wire [4-1:0] node9853;
	wire [4-1:0] node9854;
	wire [4-1:0] node9856;
	wire [4-1:0] node9860;
	wire [4-1:0] node9861;
	wire [4-1:0] node9862;
	wire [4-1:0] node9863;
	wire [4-1:0] node9864;
	wire [4-1:0] node9865;
	wire [4-1:0] node9866;
	wire [4-1:0] node9870;
	wire [4-1:0] node9872;
	wire [4-1:0] node9873;
	wire [4-1:0] node9877;
	wire [4-1:0] node9878;
	wire [4-1:0] node9879;
	wire [4-1:0] node9884;
	wire [4-1:0] node9885;
	wire [4-1:0] node9886;
	wire [4-1:0] node9890;
	wire [4-1:0] node9891;
	wire [4-1:0] node9894;
	wire [4-1:0] node9895;
	wire [4-1:0] node9898;
	wire [4-1:0] node9900;
	wire [4-1:0] node9903;
	wire [4-1:0] node9904;
	wire [4-1:0] node9905;
	wire [4-1:0] node9906;
	wire [4-1:0] node9907;
	wire [4-1:0] node9911;
	wire [4-1:0] node9913;
	wire [4-1:0] node9914;
	wire [4-1:0] node9917;
	wire [4-1:0] node9920;
	wire [4-1:0] node9921;
	wire [4-1:0] node9922;
	wire [4-1:0] node9925;
	wire [4-1:0] node9928;
	wire [4-1:0] node9929;
	wire [4-1:0] node9931;
	wire [4-1:0] node9935;
	wire [4-1:0] node9936;
	wire [4-1:0] node9937;
	wire [4-1:0] node9940;
	wire [4-1:0] node9941;
	wire [4-1:0] node9945;
	wire [4-1:0] node9946;
	wire [4-1:0] node9947;
	wire [4-1:0] node9950;
	wire [4-1:0] node9952;
	wire [4-1:0] node9955;
	wire [4-1:0] node9957;
	wire [4-1:0] node9960;
	wire [4-1:0] node9961;
	wire [4-1:0] node9962;
	wire [4-1:0] node9963;
	wire [4-1:0] node9964;
	wire [4-1:0] node9965;
	wire [4-1:0] node9968;
	wire [4-1:0] node9971;
	wire [4-1:0] node9972;
	wire [4-1:0] node9976;
	wire [4-1:0] node9978;
	wire [4-1:0] node9980;
	wire [4-1:0] node9981;
	wire [4-1:0] node9984;
	wire [4-1:0] node9987;
	wire [4-1:0] node9988;
	wire [4-1:0] node9990;
	wire [4-1:0] node9992;
	wire [4-1:0] node9995;
	wire [4-1:0] node9996;
	wire [4-1:0] node9997;
	wire [4-1:0] node10001;
	wire [4-1:0] node10003;
	wire [4-1:0] node10006;
	wire [4-1:0] node10007;
	wire [4-1:0] node10008;
	wire [4-1:0] node10009;
	wire [4-1:0] node10011;
	wire [4-1:0] node10014;
	wire [4-1:0] node10015;
	wire [4-1:0] node10017;
	wire [4-1:0] node10020;
	wire [4-1:0] node10021;
	wire [4-1:0] node10024;
	wire [4-1:0] node10027;
	wire [4-1:0] node10028;
	wire [4-1:0] node10030;
	wire [4-1:0] node10033;
	wire [4-1:0] node10034;
	wire [4-1:0] node10038;
	wire [4-1:0] node10039;
	wire [4-1:0] node10040;
	wire [4-1:0] node10043;
	wire [4-1:0] node10045;
	wire [4-1:0] node10048;
	wire [4-1:0] node10049;
	wire [4-1:0] node10050;
	wire [4-1:0] node10054;
	wire [4-1:0] node10055;
	wire [4-1:0] node10059;
	wire [4-1:0] node10060;
	wire [4-1:0] node10061;
	wire [4-1:0] node10062;
	wire [4-1:0] node10063;
	wire [4-1:0] node10064;
	wire [4-1:0] node10065;
	wire [4-1:0] node10066;
	wire [4-1:0] node10067;
	wire [4-1:0] node10068;
	wire [4-1:0] node10071;
	wire [4-1:0] node10075;
	wire [4-1:0] node10078;
	wire [4-1:0] node10079;
	wire [4-1:0] node10080;
	wire [4-1:0] node10083;
	wire [4-1:0] node10086;
	wire [4-1:0] node10087;
	wire [4-1:0] node10091;
	wire [4-1:0] node10092;
	wire [4-1:0] node10094;
	wire [4-1:0] node10095;
	wire [4-1:0] node10098;
	wire [4-1:0] node10099;
	wire [4-1:0] node10103;
	wire [4-1:0] node10104;
	wire [4-1:0] node10105;
	wire [4-1:0] node10108;
	wire [4-1:0] node10112;
	wire [4-1:0] node10113;
	wire [4-1:0] node10114;
	wire [4-1:0] node10115;
	wire [4-1:0] node10118;
	wire [4-1:0] node10121;
	wire [4-1:0] node10122;
	wire [4-1:0] node10123;
	wire [4-1:0] node10124;
	wire [4-1:0] node10128;
	wire [4-1:0] node10131;
	wire [4-1:0] node10132;
	wire [4-1:0] node10133;
	wire [4-1:0] node10138;
	wire [4-1:0] node10139;
	wire [4-1:0] node10140;
	wire [4-1:0] node10142;
	wire [4-1:0] node10145;
	wire [4-1:0] node10147;
	wire [4-1:0] node10149;
	wire [4-1:0] node10152;
	wire [4-1:0] node10153;
	wire [4-1:0] node10156;
	wire [4-1:0] node10157;
	wire [4-1:0] node10158;
	wire [4-1:0] node10162;
	wire [4-1:0] node10164;
	wire [4-1:0] node10167;
	wire [4-1:0] node10168;
	wire [4-1:0] node10169;
	wire [4-1:0] node10170;
	wire [4-1:0] node10171;
	wire [4-1:0] node10172;
	wire [4-1:0] node10177;
	wire [4-1:0] node10178;
	wire [4-1:0] node10179;
	wire [4-1:0] node10182;
	wire [4-1:0] node10186;
	wire [4-1:0] node10187;
	wire [4-1:0] node10188;
	wire [4-1:0] node10189;
	wire [4-1:0] node10193;
	wire [4-1:0] node10195;
	wire [4-1:0] node10198;
	wire [4-1:0] node10199;
	wire [4-1:0] node10203;
	wire [4-1:0] node10204;
	wire [4-1:0] node10205;
	wire [4-1:0] node10206;
	wire [4-1:0] node10209;
	wire [4-1:0] node10211;
	wire [4-1:0] node10212;
	wire [4-1:0] node10216;
	wire [4-1:0] node10218;
	wire [4-1:0] node10220;
	wire [4-1:0] node10221;
	wire [4-1:0] node10224;
	wire [4-1:0] node10227;
	wire [4-1:0] node10228;
	wire [4-1:0] node10229;
	wire [4-1:0] node10230;
	wire [4-1:0] node10233;
	wire [4-1:0] node10237;
	wire [4-1:0] node10238;
	wire [4-1:0] node10240;
	wire [4-1:0] node10243;
	wire [4-1:0] node10246;
	wire [4-1:0] node10247;
	wire [4-1:0] node10248;
	wire [4-1:0] node10249;
	wire [4-1:0] node10250;
	wire [4-1:0] node10252;
	wire [4-1:0] node10254;
	wire [4-1:0] node10256;
	wire [4-1:0] node10259;
	wire [4-1:0] node10260;
	wire [4-1:0] node10261;
	wire [4-1:0] node10264;
	wire [4-1:0] node10268;
	wire [4-1:0] node10269;
	wire [4-1:0] node10270;
	wire [4-1:0] node10271;
	wire [4-1:0] node10275;
	wire [4-1:0] node10277;
	wire [4-1:0] node10280;
	wire [4-1:0] node10281;
	wire [4-1:0] node10283;
	wire [4-1:0] node10284;
	wire [4-1:0] node10288;
	wire [4-1:0] node10289;
	wire [4-1:0] node10290;
	wire [4-1:0] node10293;
	wire [4-1:0] node10296;
	wire [4-1:0] node10298;
	wire [4-1:0] node10301;
	wire [4-1:0] node10302;
	wire [4-1:0] node10303;
	wire [4-1:0] node10304;
	wire [4-1:0] node10306;
	wire [4-1:0] node10307;
	wire [4-1:0] node10310;
	wire [4-1:0] node10313;
	wire [4-1:0] node10316;
	wire [4-1:0] node10317;
	wire [4-1:0] node10320;
	wire [4-1:0] node10321;
	wire [4-1:0] node10322;
	wire [4-1:0] node10326;
	wire [4-1:0] node10327;
	wire [4-1:0] node10331;
	wire [4-1:0] node10332;
	wire [4-1:0] node10333;
	wire [4-1:0] node10335;
	wire [4-1:0] node10336;
	wire [4-1:0] node10340;
	wire [4-1:0] node10343;
	wire [4-1:0] node10344;
	wire [4-1:0] node10345;
	wire [4-1:0] node10348;
	wire [4-1:0] node10351;
	wire [4-1:0] node10354;
	wire [4-1:0] node10355;
	wire [4-1:0] node10356;
	wire [4-1:0] node10357;
	wire [4-1:0] node10359;
	wire [4-1:0] node10362;
	wire [4-1:0] node10363;
	wire [4-1:0] node10364;
	wire [4-1:0] node10367;
	wire [4-1:0] node10370;
	wire [4-1:0] node10371;
	wire [4-1:0] node10375;
	wire [4-1:0] node10376;
	wire [4-1:0] node10377;
	wire [4-1:0] node10379;
	wire [4-1:0] node10382;
	wire [4-1:0] node10383;
	wire [4-1:0] node10387;
	wire [4-1:0] node10388;
	wire [4-1:0] node10389;
	wire [4-1:0] node10392;
	wire [4-1:0] node10395;
	wire [4-1:0] node10397;
	wire [4-1:0] node10400;
	wire [4-1:0] node10401;
	wire [4-1:0] node10402;
	wire [4-1:0] node10404;
	wire [4-1:0] node10406;
	wire [4-1:0] node10409;
	wire [4-1:0] node10410;
	wire [4-1:0] node10413;
	wire [4-1:0] node10414;
	wire [4-1:0] node10418;
	wire [4-1:0] node10419;
	wire [4-1:0] node10420;
	wire [4-1:0] node10422;
	wire [4-1:0] node10423;
	wire [4-1:0] node10426;
	wire [4-1:0] node10429;
	wire [4-1:0] node10430;
	wire [4-1:0] node10434;
	wire [4-1:0] node10435;
	wire [4-1:0] node10436;
	wire [4-1:0] node10439;
	wire [4-1:0] node10442;
	wire [4-1:0] node10443;
	wire [4-1:0] node10444;
	wire [4-1:0] node10449;
	wire [4-1:0] node10450;
	wire [4-1:0] node10451;
	wire [4-1:0] node10452;
	wire [4-1:0] node10453;
	wire [4-1:0] node10454;
	wire [4-1:0] node10455;
	wire [4-1:0] node10456;
	wire [4-1:0] node10457;
	wire [4-1:0] node10460;
	wire [4-1:0] node10464;
	wire [4-1:0] node10466;
	wire [4-1:0] node10469;
	wire [4-1:0] node10470;
	wire [4-1:0] node10471;
	wire [4-1:0] node10474;
	wire [4-1:0] node10477;
	wire [4-1:0] node10479;
	wire [4-1:0] node10482;
	wire [4-1:0] node10483;
	wire [4-1:0] node10485;
	wire [4-1:0] node10486;
	wire [4-1:0] node10487;
	wire [4-1:0] node10493;
	wire [4-1:0] node10494;
	wire [4-1:0] node10495;
	wire [4-1:0] node10496;
	wire [4-1:0] node10498;
	wire [4-1:0] node10500;
	wire [4-1:0] node10503;
	wire [4-1:0] node10504;
	wire [4-1:0] node10507;
	wire [4-1:0] node10510;
	wire [4-1:0] node10511;
	wire [4-1:0] node10513;
	wire [4-1:0] node10514;
	wire [4-1:0] node10518;
	wire [4-1:0] node10519;
	wire [4-1:0] node10522;
	wire [4-1:0] node10525;
	wire [4-1:0] node10526;
	wire [4-1:0] node10527;
	wire [4-1:0] node10530;
	wire [4-1:0] node10531;
	wire [4-1:0] node10532;
	wire [4-1:0] node10535;
	wire [4-1:0] node10538;
	wire [4-1:0] node10541;
	wire [4-1:0] node10543;
	wire [4-1:0] node10544;
	wire [4-1:0] node10545;
	wire [4-1:0] node10548;
	wire [4-1:0] node10552;
	wire [4-1:0] node10553;
	wire [4-1:0] node10554;
	wire [4-1:0] node10555;
	wire [4-1:0] node10556;
	wire [4-1:0] node10557;
	wire [4-1:0] node10559;
	wire [4-1:0] node10562;
	wire [4-1:0] node10563;
	wire [4-1:0] node10567;
	wire [4-1:0] node10568;
	wire [4-1:0] node10571;
	wire [4-1:0] node10574;
	wire [4-1:0] node10575;
	wire [4-1:0] node10578;
	wire [4-1:0] node10579;
	wire [4-1:0] node10583;
	wire [4-1:0] node10584;
	wire [4-1:0] node10585;
	wire [4-1:0] node10588;
	wire [4-1:0] node10590;
	wire [4-1:0] node10593;
	wire [4-1:0] node10594;
	wire [4-1:0] node10595;
	wire [4-1:0] node10596;
	wire [4-1:0] node10600;
	wire [4-1:0] node10601;
	wire [4-1:0] node10606;
	wire [4-1:0] node10607;
	wire [4-1:0] node10608;
	wire [4-1:0] node10609;
	wire [4-1:0] node10611;
	wire [4-1:0] node10614;
	wire [4-1:0] node10615;
	wire [4-1:0] node10616;
	wire [4-1:0] node10619;
	wire [4-1:0] node10623;
	wire [4-1:0] node10624;
	wire [4-1:0] node10628;
	wire [4-1:0] node10629;
	wire [4-1:0] node10630;
	wire [4-1:0] node10631;
	wire [4-1:0] node10634;
	wire [4-1:0] node10637;
	wire [4-1:0] node10640;
	wire [4-1:0] node10641;
	wire [4-1:0] node10642;
	wire [4-1:0] node10645;
	wire [4-1:0] node10648;
	wire [4-1:0] node10650;
	wire [4-1:0] node10653;
	wire [4-1:0] node10654;
	wire [4-1:0] node10655;
	wire [4-1:0] node10656;
	wire [4-1:0] node10657;
	wire [4-1:0] node10658;
	wire [4-1:0] node10659;
	wire [4-1:0] node10661;
	wire [4-1:0] node10665;
	wire [4-1:0] node10666;
	wire [4-1:0] node10669;
	wire [4-1:0] node10670;
	wire [4-1:0] node10674;
	wire [4-1:0] node10675;
	wire [4-1:0] node10676;
	wire [4-1:0] node10678;
	wire [4-1:0] node10681;
	wire [4-1:0] node10682;
	wire [4-1:0] node10686;
	wire [4-1:0] node10688;
	wire [4-1:0] node10691;
	wire [4-1:0] node10692;
	wire [4-1:0] node10693;
	wire [4-1:0] node10694;
	wire [4-1:0] node10697;
	wire [4-1:0] node10700;
	wire [4-1:0] node10703;
	wire [4-1:0] node10704;
	wire [4-1:0] node10706;
	wire [4-1:0] node10709;
	wire [4-1:0] node10711;
	wire [4-1:0] node10714;
	wire [4-1:0] node10715;
	wire [4-1:0] node10716;
	wire [4-1:0] node10717;
	wire [4-1:0] node10718;
	wire [4-1:0] node10723;
	wire [4-1:0] node10724;
	wire [4-1:0] node10725;
	wire [4-1:0] node10728;
	wire [4-1:0] node10731;
	wire [4-1:0] node10733;
	wire [4-1:0] node10736;
	wire [4-1:0] node10737;
	wire [4-1:0] node10738;
	wire [4-1:0] node10741;
	wire [4-1:0] node10742;
	wire [4-1:0] node10744;
	wire [4-1:0] node10747;
	wire [4-1:0] node10750;
	wire [4-1:0] node10751;
	wire [4-1:0] node10753;
	wire [4-1:0] node10754;
	wire [4-1:0] node10757;
	wire [4-1:0] node10760;
	wire [4-1:0] node10763;
	wire [4-1:0] node10764;
	wire [4-1:0] node10765;
	wire [4-1:0] node10766;
	wire [4-1:0] node10767;
	wire [4-1:0] node10769;
	wire [4-1:0] node10772;
	wire [4-1:0] node10773;
	wire [4-1:0] node10776;
	wire [4-1:0] node10779;
	wire [4-1:0] node10781;
	wire [4-1:0] node10782;
	wire [4-1:0] node10785;
	wire [4-1:0] node10788;
	wire [4-1:0] node10789;
	wire [4-1:0] node10790;
	wire [4-1:0] node10791;
	wire [4-1:0] node10795;
	wire [4-1:0] node10797;
	wire [4-1:0] node10800;
	wire [4-1:0] node10801;
	wire [4-1:0] node10803;
	wire [4-1:0] node10804;
	wire [4-1:0] node10807;
	wire [4-1:0] node10810;
	wire [4-1:0] node10811;
	wire [4-1:0] node10815;
	wire [4-1:0] node10816;
	wire [4-1:0] node10817;
	wire [4-1:0] node10818;
	wire [4-1:0] node10819;
	wire [4-1:0] node10820;
	wire [4-1:0] node10825;
	wire [4-1:0] node10826;
	wire [4-1:0] node10830;
	wire [4-1:0] node10831;
	wire [4-1:0] node10833;
	wire [4-1:0] node10836;
	wire [4-1:0] node10838;
	wire [4-1:0] node10841;
	wire [4-1:0] node10842;
	wire [4-1:0] node10843;
	wire [4-1:0] node10846;
	wire [4-1:0] node10849;
	wire [4-1:0] node10851;
	wire [4-1:0] node10852;
	wire [4-1:0] node10855;
	wire [4-1:0] node10858;
	wire [4-1:0] node10859;
	wire [4-1:0] node10860;
	wire [4-1:0] node10861;
	wire [4-1:0] node10862;
	wire [4-1:0] node10863;
	wire [4-1:0] node10864;
	wire [4-1:0] node10865;
	wire [4-1:0] node10866;
	wire [4-1:0] node10869;
	wire [4-1:0] node10872;
	wire [4-1:0] node10874;
	wire [4-1:0] node10875;
	wire [4-1:0] node10876;
	wire [4-1:0] node10879;
	wire [4-1:0] node10883;
	wire [4-1:0] node10884;
	wire [4-1:0] node10885;
	wire [4-1:0] node10889;
	wire [4-1:0] node10891;
	wire [4-1:0] node10892;
	wire [4-1:0] node10896;
	wire [4-1:0] node10897;
	wire [4-1:0] node10898;
	wire [4-1:0] node10899;
	wire [4-1:0] node10900;
	wire [4-1:0] node10904;
	wire [4-1:0] node10906;
	wire [4-1:0] node10909;
	wire [4-1:0] node10910;
	wire [4-1:0] node10912;
	wire [4-1:0] node10915;
	wire [4-1:0] node10916;
	wire [4-1:0] node10920;
	wire [4-1:0] node10921;
	wire [4-1:0] node10922;
	wire [4-1:0] node10924;
	wire [4-1:0] node10927;
	wire [4-1:0] node10928;
	wire [4-1:0] node10929;
	wire [4-1:0] node10933;
	wire [4-1:0] node10935;
	wire [4-1:0] node10938;
	wire [4-1:0] node10939;
	wire [4-1:0] node10941;
	wire [4-1:0] node10944;
	wire [4-1:0] node10946;
	wire [4-1:0] node10948;
	wire [4-1:0] node10951;
	wire [4-1:0] node10952;
	wire [4-1:0] node10953;
	wire [4-1:0] node10954;
	wire [4-1:0] node10955;
	wire [4-1:0] node10958;
	wire [4-1:0] node10959;
	wire [4-1:0] node10962;
	wire [4-1:0] node10964;
	wire [4-1:0] node10967;
	wire [4-1:0] node10968;
	wire [4-1:0] node10970;
	wire [4-1:0] node10972;
	wire [4-1:0] node10975;
	wire [4-1:0] node10978;
	wire [4-1:0] node10979;
	wire [4-1:0] node10980;
	wire [4-1:0] node10981;
	wire [4-1:0] node10985;
	wire [4-1:0] node10986;
	wire [4-1:0] node10988;
	wire [4-1:0] node10991;
	wire [4-1:0] node10993;
	wire [4-1:0] node10996;
	wire [4-1:0] node10997;
	wire [4-1:0] node11000;
	wire [4-1:0] node11001;
	wire [4-1:0] node11005;
	wire [4-1:0] node11006;
	wire [4-1:0] node11007;
	wire [4-1:0] node11008;
	wire [4-1:0] node11011;
	wire [4-1:0] node11012;
	wire [4-1:0] node11015;
	wire [4-1:0] node11018;
	wire [4-1:0] node11019;
	wire [4-1:0] node11021;
	wire [4-1:0] node11024;
	wire [4-1:0] node11025;
	wire [4-1:0] node11026;
	wire [4-1:0] node11029;
	wire [4-1:0] node11032;
	wire [4-1:0] node11033;
	wire [4-1:0] node11036;
	wire [4-1:0] node11039;
	wire [4-1:0] node11040;
	wire [4-1:0] node11041;
	wire [4-1:0] node11044;
	wire [4-1:0] node11045;
	wire [4-1:0] node11047;
	wire [4-1:0] node11050;
	wire [4-1:0] node11053;
	wire [4-1:0] node11054;
	wire [4-1:0] node11055;
	wire [4-1:0] node11058;
	wire [4-1:0] node11061;
	wire [4-1:0] node11062;
	wire [4-1:0] node11066;
	wire [4-1:0] node11067;
	wire [4-1:0] node11068;
	wire [4-1:0] node11069;
	wire [4-1:0] node11070;
	wire [4-1:0] node11071;
	wire [4-1:0] node11072;
	wire [4-1:0] node11077;
	wire [4-1:0] node11078;
	wire [4-1:0] node11081;
	wire [4-1:0] node11083;
	wire [4-1:0] node11084;
	wire [4-1:0] node11087;
	wire [4-1:0] node11090;
	wire [4-1:0] node11091;
	wire [4-1:0] node11092;
	wire [4-1:0] node11093;
	wire [4-1:0] node11096;
	wire [4-1:0] node11099;
	wire [4-1:0] node11100;
	wire [4-1:0] node11104;
	wire [4-1:0] node11105;
	wire [4-1:0] node11106;
	wire [4-1:0] node11108;
	wire [4-1:0] node11112;
	wire [4-1:0] node11114;
	wire [4-1:0] node11117;
	wire [4-1:0] node11118;
	wire [4-1:0] node11119;
	wire [4-1:0] node11120;
	wire [4-1:0] node11124;
	wire [4-1:0] node11126;
	wire [4-1:0] node11127;
	wire [4-1:0] node11128;
	wire [4-1:0] node11132;
	wire [4-1:0] node11133;
	wire [4-1:0] node11137;
	wire [4-1:0] node11138;
	wire [4-1:0] node11139;
	wire [4-1:0] node11140;
	wire [4-1:0] node11143;
	wire [4-1:0] node11146;
	wire [4-1:0] node11147;
	wire [4-1:0] node11148;
	wire [4-1:0] node11151;
	wire [4-1:0] node11155;
	wire [4-1:0] node11156;
	wire [4-1:0] node11159;
	wire [4-1:0] node11160;
	wire [4-1:0] node11164;
	wire [4-1:0] node11165;
	wire [4-1:0] node11166;
	wire [4-1:0] node11167;
	wire [4-1:0] node11168;
	wire [4-1:0] node11169;
	wire [4-1:0] node11170;
	wire [4-1:0] node11174;
	wire [4-1:0] node11176;
	wire [4-1:0] node11179;
	wire [4-1:0] node11181;
	wire [4-1:0] node11183;
	wire [4-1:0] node11186;
	wire [4-1:0] node11187;
	wire [4-1:0] node11188;
	wire [4-1:0] node11192;
	wire [4-1:0] node11194;
	wire [4-1:0] node11197;
	wire [4-1:0] node11198;
	wire [4-1:0] node11199;
	wire [4-1:0] node11200;
	wire [4-1:0] node11204;
	wire [4-1:0] node11207;
	wire [4-1:0] node11210;
	wire [4-1:0] node11211;
	wire [4-1:0] node11212;
	wire [4-1:0] node11213;
	wire [4-1:0] node11217;
	wire [4-1:0] node11218;
	wire [4-1:0] node11220;
	wire [4-1:0] node11223;
	wire [4-1:0] node11224;
	wire [4-1:0] node11227;
	wire [4-1:0] node11230;
	wire [4-1:0] node11231;
	wire [4-1:0] node11232;
	wire [4-1:0] node11234;
	wire [4-1:0] node11237;
	wire [4-1:0] node11238;
	wire [4-1:0] node11242;
	wire [4-1:0] node11243;
	wire [4-1:0] node11244;
	wire [4-1:0] node11248;
	wire [4-1:0] node11249;
	wire [4-1:0] node11252;
	wire [4-1:0] node11255;
	wire [4-1:0] node11256;
	wire [4-1:0] node11257;
	wire [4-1:0] node11258;
	wire [4-1:0] node11259;
	wire [4-1:0] node11260;
	wire [4-1:0] node11261;
	wire [4-1:0] node11264;
	wire [4-1:0] node11265;
	wire [4-1:0] node11269;
	wire [4-1:0] node11270;
	wire [4-1:0] node11272;
	wire [4-1:0] node11276;
	wire [4-1:0] node11277;
	wire [4-1:0] node11279;
	wire [4-1:0] node11282;
	wire [4-1:0] node11283;
	wire [4-1:0] node11287;
	wire [4-1:0] node11288;
	wire [4-1:0] node11289;
	wire [4-1:0] node11290;
	wire [4-1:0] node11292;
	wire [4-1:0] node11295;
	wire [4-1:0] node11297;
	wire [4-1:0] node11298;
	wire [4-1:0] node11301;
	wire [4-1:0] node11304;
	wire [4-1:0] node11305;
	wire [4-1:0] node11306;
	wire [4-1:0] node11310;
	wire [4-1:0] node11311;
	wire [4-1:0] node11312;
	wire [4-1:0] node11315;
	wire [4-1:0] node11319;
	wire [4-1:0] node11320;
	wire [4-1:0] node11321;
	wire [4-1:0] node11322;
	wire [4-1:0] node11325;
	wire [4-1:0] node11328;
	wire [4-1:0] node11331;
	wire [4-1:0] node11332;
	wire [4-1:0] node11335;
	wire [4-1:0] node11336;
	wire [4-1:0] node11338;
	wire [4-1:0] node11342;
	wire [4-1:0] node11343;
	wire [4-1:0] node11344;
	wire [4-1:0] node11345;
	wire [4-1:0] node11346;
	wire [4-1:0] node11349;
	wire [4-1:0] node11350;
	wire [4-1:0] node11354;
	wire [4-1:0] node11355;
	wire [4-1:0] node11356;
	wire [4-1:0] node11357;
	wire [4-1:0] node11360;
	wire [4-1:0] node11363;
	wire [4-1:0] node11364;
	wire [4-1:0] node11368;
	wire [4-1:0] node11371;
	wire [4-1:0] node11372;
	wire [4-1:0] node11373;
	wire [4-1:0] node11374;
	wire [4-1:0] node11376;
	wire [4-1:0] node11380;
	wire [4-1:0] node11381;
	wire [4-1:0] node11385;
	wire [4-1:0] node11386;
	wire [4-1:0] node11388;
	wire [4-1:0] node11390;
	wire [4-1:0] node11394;
	wire [4-1:0] node11395;
	wire [4-1:0] node11396;
	wire [4-1:0] node11399;
	wire [4-1:0] node11401;
	wire [4-1:0] node11403;
	wire [4-1:0] node11406;
	wire [4-1:0] node11407;
	wire [4-1:0] node11408;
	wire [4-1:0] node11409;
	wire [4-1:0] node11410;
	wire [4-1:0] node11415;
	wire [4-1:0] node11416;
	wire [4-1:0] node11417;
	wire [4-1:0] node11421;
	wire [4-1:0] node11424;
	wire [4-1:0] node11425;
	wire [4-1:0] node11427;
	wire [4-1:0] node11430;
	wire [4-1:0] node11431;
	wire [4-1:0] node11433;
	wire [4-1:0] node11436;
	wire [4-1:0] node11439;
	wire [4-1:0] node11440;
	wire [4-1:0] node11441;
	wire [4-1:0] node11442;
	wire [4-1:0] node11443;
	wire [4-1:0] node11444;
	wire [4-1:0] node11445;
	wire [4-1:0] node11449;
	wire [4-1:0] node11451;
	wire [4-1:0] node11454;
	wire [4-1:0] node11455;
	wire [4-1:0] node11456;
	wire [4-1:0] node11459;
	wire [4-1:0] node11462;
	wire [4-1:0] node11463;
	wire [4-1:0] node11467;
	wire [4-1:0] node11468;
	wire [4-1:0] node11470;
	wire [4-1:0] node11471;
	wire [4-1:0] node11475;
	wire [4-1:0] node11477;
	wire [4-1:0] node11478;
	wire [4-1:0] node11482;
	wire [4-1:0] node11483;
	wire [4-1:0] node11484;
	wire [4-1:0] node11485;
	wire [4-1:0] node11487;
	wire [4-1:0] node11491;
	wire [4-1:0] node11493;
	wire [4-1:0] node11495;
	wire [4-1:0] node11498;
	wire [4-1:0] node11499;
	wire [4-1:0] node11501;
	wire [4-1:0] node11502;
	wire [4-1:0] node11503;
	wire [4-1:0] node11507;
	wire [4-1:0] node11510;
	wire [4-1:0] node11511;
	wire [4-1:0] node11512;
	wire [4-1:0] node11517;
	wire [4-1:0] node11518;
	wire [4-1:0] node11519;
	wire [4-1:0] node11520;
	wire [4-1:0] node11521;
	wire [4-1:0] node11522;
	wire [4-1:0] node11524;
	wire [4-1:0] node11527;
	wire [4-1:0] node11528;
	wire [4-1:0] node11531;
	wire [4-1:0] node11535;
	wire [4-1:0] node11536;
	wire [4-1:0] node11538;
	wire [4-1:0] node11541;
	wire [4-1:0] node11542;
	wire [4-1:0] node11544;
	wire [4-1:0] node11548;
	wire [4-1:0] node11549;
	wire [4-1:0] node11551;
	wire [4-1:0] node11552;
	wire [4-1:0] node11553;
	wire [4-1:0] node11557;
	wire [4-1:0] node11560;
	wire [4-1:0] node11561;
	wire [4-1:0] node11562;
	wire [4-1:0] node11563;
	wire [4-1:0] node11567;
	wire [4-1:0] node11570;
	wire [4-1:0] node11571;
	wire [4-1:0] node11575;
	wire [4-1:0] node11576;
	wire [4-1:0] node11577;
	wire [4-1:0] node11578;
	wire [4-1:0] node11579;
	wire [4-1:0] node11582;
	wire [4-1:0] node11585;
	wire [4-1:0] node11586;
	wire [4-1:0] node11589;
	wire [4-1:0] node11592;
	wire [4-1:0] node11593;
	wire [4-1:0] node11595;
	wire [4-1:0] node11598;
	wire [4-1:0] node11599;
	wire [4-1:0] node11602;
	wire [4-1:0] node11605;
	wire [4-1:0] node11606;
	wire [4-1:0] node11607;
	wire [4-1:0] node11608;
	wire [4-1:0] node11612;
	wire [4-1:0] node11614;
	wire [4-1:0] node11617;
	wire [4-1:0] node11618;
	wire [4-1:0] node11621;
	wire [4-1:0] node11624;
	wire [4-1:0] node11625;
	wire [4-1:0] node11626;
	wire [4-1:0] node11627;
	wire [4-1:0] node11628;
	wire [4-1:0] node11629;
	wire [4-1:0] node11630;
	wire [4-1:0] node11631;
	wire [4-1:0] node11632;
	wire [4-1:0] node11634;
	wire [4-1:0] node11637;
	wire [4-1:0] node11638;
	wire [4-1:0] node11641;
	wire [4-1:0] node11644;
	wire [4-1:0] node11646;
	wire [4-1:0] node11649;
	wire [4-1:0] node11650;
	wire [4-1:0] node11652;
	wire [4-1:0] node11653;
	wire [4-1:0] node11656;
	wire [4-1:0] node11659;
	wire [4-1:0] node11662;
	wire [4-1:0] node11663;
	wire [4-1:0] node11664;
	wire [4-1:0] node11667;
	wire [4-1:0] node11668;
	wire [4-1:0] node11669;
	wire [4-1:0] node11672;
	wire [4-1:0] node11675;
	wire [4-1:0] node11678;
	wire [4-1:0] node11679;
	wire [4-1:0] node11682;
	wire [4-1:0] node11684;
	wire [4-1:0] node11685;
	wire [4-1:0] node11689;
	wire [4-1:0] node11690;
	wire [4-1:0] node11691;
	wire [4-1:0] node11692;
	wire [4-1:0] node11693;
	wire [4-1:0] node11695;
	wire [4-1:0] node11698;
	wire [4-1:0] node11702;
	wire [4-1:0] node11703;
	wire [4-1:0] node11705;
	wire [4-1:0] node11708;
	wire [4-1:0] node11709;
	wire [4-1:0] node11711;
	wire [4-1:0] node11714;
	wire [4-1:0] node11715;
	wire [4-1:0] node11719;
	wire [4-1:0] node11720;
	wire [4-1:0] node11721;
	wire [4-1:0] node11722;
	wire [4-1:0] node11725;
	wire [4-1:0] node11728;
	wire [4-1:0] node11729;
	wire [4-1:0] node11733;
	wire [4-1:0] node11734;
	wire [4-1:0] node11735;
	wire [4-1:0] node11736;
	wire [4-1:0] node11740;
	wire [4-1:0] node11741;
	wire [4-1:0] node11745;
	wire [4-1:0] node11746;
	wire [4-1:0] node11749;
	wire [4-1:0] node11752;
	wire [4-1:0] node11753;
	wire [4-1:0] node11754;
	wire [4-1:0] node11755;
	wire [4-1:0] node11756;
	wire [4-1:0] node11757;
	wire [4-1:0] node11758;
	wire [4-1:0] node11763;
	wire [4-1:0] node11764;
	wire [4-1:0] node11766;
	wire [4-1:0] node11769;
	wire [4-1:0] node11771;
	wire [4-1:0] node11774;
	wire [4-1:0] node11775;
	wire [4-1:0] node11778;
	wire [4-1:0] node11779;
	wire [4-1:0] node11780;
	wire [4-1:0] node11783;
	wire [4-1:0] node11786;
	wire [4-1:0] node11789;
	wire [4-1:0] node11790;
	wire [4-1:0] node11791;
	wire [4-1:0] node11792;
	wire [4-1:0] node11795;
	wire [4-1:0] node11796;
	wire [4-1:0] node11799;
	wire [4-1:0] node11802;
	wire [4-1:0] node11805;
	wire [4-1:0] node11806;
	wire [4-1:0] node11807;
	wire [4-1:0] node11808;
	wire [4-1:0] node11812;
	wire [4-1:0] node11815;
	wire [4-1:0] node11817;
	wire [4-1:0] node11820;
	wire [4-1:0] node11821;
	wire [4-1:0] node11822;
	wire [4-1:0] node11823;
	wire [4-1:0] node11824;
	wire [4-1:0] node11825;
	wire [4-1:0] node11830;
	wire [4-1:0] node11831;
	wire [4-1:0] node11832;
	wire [4-1:0] node11835;
	wire [4-1:0] node11839;
	wire [4-1:0] node11840;
	wire [4-1:0] node11843;
	wire [4-1:0] node11844;
	wire [4-1:0] node11845;
	wire [4-1:0] node11848;
	wire [4-1:0] node11851;
	wire [4-1:0] node11852;
	wire [4-1:0] node11855;
	wire [4-1:0] node11858;
	wire [4-1:0] node11859;
	wire [4-1:0] node11860;
	wire [4-1:0] node11862;
	wire [4-1:0] node11863;
	wire [4-1:0] node11866;
	wire [4-1:0] node11869;
	wire [4-1:0] node11870;
	wire [4-1:0] node11871;
	wire [4-1:0] node11875;
	wire [4-1:0] node11877;
	wire [4-1:0] node11880;
	wire [4-1:0] node11881;
	wire [4-1:0] node11884;
	wire [4-1:0] node11887;
	wire [4-1:0] node11888;
	wire [4-1:0] node11889;
	wire [4-1:0] node11890;
	wire [4-1:0] node11891;
	wire [4-1:0] node11893;
	wire [4-1:0] node11894;
	wire [4-1:0] node11896;
	wire [4-1:0] node11900;
	wire [4-1:0] node11901;
	wire [4-1:0] node11904;
	wire [4-1:0] node11907;
	wire [4-1:0] node11908;
	wire [4-1:0] node11909;
	wire [4-1:0] node11910;
	wire [4-1:0] node11911;
	wire [4-1:0] node11914;
	wire [4-1:0] node11918;
	wire [4-1:0] node11920;
	wire [4-1:0] node11923;
	wire [4-1:0] node11924;
	wire [4-1:0] node11925;
	wire [4-1:0] node11926;
	wire [4-1:0] node11929;
	wire [4-1:0] node11932;
	wire [4-1:0] node11934;
	wire [4-1:0] node11937;
	wire [4-1:0] node11940;
	wire [4-1:0] node11941;
	wire [4-1:0] node11942;
	wire [4-1:0] node11943;
	wire [4-1:0] node11945;
	wire [4-1:0] node11948;
	wire [4-1:0] node11951;
	wire [4-1:0] node11952;
	wire [4-1:0] node11953;
	wire [4-1:0] node11956;
	wire [4-1:0] node11960;
	wire [4-1:0] node11961;
	wire [4-1:0] node11962;
	wire [4-1:0] node11964;
	wire [4-1:0] node11968;
	wire [4-1:0] node11969;
	wire [4-1:0] node11971;
	wire [4-1:0] node11974;
	wire [4-1:0] node11975;
	wire [4-1:0] node11978;
	wire [4-1:0] node11981;
	wire [4-1:0] node11982;
	wire [4-1:0] node11983;
	wire [4-1:0] node11984;
	wire [4-1:0] node11985;
	wire [4-1:0] node11988;
	wire [4-1:0] node11989;
	wire [4-1:0] node11990;
	wire [4-1:0] node11995;
	wire [4-1:0] node11996;
	wire [4-1:0] node11998;
	wire [4-1:0] node12001;
	wire [4-1:0] node12002;
	wire [4-1:0] node12004;
	wire [4-1:0] node12008;
	wire [4-1:0] node12009;
	wire [4-1:0] node12010;
	wire [4-1:0] node12011;
	wire [4-1:0] node12015;
	wire [4-1:0] node12018;
	wire [4-1:0] node12019;
	wire [4-1:0] node12020;
	wire [4-1:0] node12022;
	wire [4-1:0] node12026;
	wire [4-1:0] node12028;
	wire [4-1:0] node12029;
	wire [4-1:0] node12032;
	wire [4-1:0] node12035;
	wire [4-1:0] node12036;
	wire [4-1:0] node12037;
	wire [4-1:0] node12039;
	wire [4-1:0] node12040;
	wire [4-1:0] node12044;
	wire [4-1:0] node12045;
	wire [4-1:0] node12046;
	wire [4-1:0] node12049;
	wire [4-1:0] node12053;
	wire [4-1:0] node12054;
	wire [4-1:0] node12055;
	wire [4-1:0] node12057;
	wire [4-1:0] node12060;
	wire [4-1:0] node12061;
	wire [4-1:0] node12064;
	wire [4-1:0] node12067;
	wire [4-1:0] node12069;
	wire [4-1:0] node12070;
	wire [4-1:0] node12073;
	wire [4-1:0] node12076;
	wire [4-1:0] node12077;
	wire [4-1:0] node12078;
	wire [4-1:0] node12079;
	wire [4-1:0] node12080;
	wire [4-1:0] node12081;
	wire [4-1:0] node12082;
	wire [4-1:0] node12084;
	wire [4-1:0] node12087;
	wire [4-1:0] node12088;
	wire [4-1:0] node12089;
	wire [4-1:0] node12092;
	wire [4-1:0] node12095;
	wire [4-1:0] node12097;
	wire [4-1:0] node12100;
	wire [4-1:0] node12101;
	wire [4-1:0] node12102;
	wire [4-1:0] node12107;
	wire [4-1:0] node12108;
	wire [4-1:0] node12109;
	wire [4-1:0] node12111;
	wire [4-1:0] node12113;
	wire [4-1:0] node12116;
	wire [4-1:0] node12117;
	wire [4-1:0] node12118;
	wire [4-1:0] node12121;
	wire [4-1:0] node12125;
	wire [4-1:0] node12126;
	wire [4-1:0] node12129;
	wire [4-1:0] node12132;
	wire [4-1:0] node12133;
	wire [4-1:0] node12134;
	wire [4-1:0] node12137;
	wire [4-1:0] node12138;
	wire [4-1:0] node12141;
	wire [4-1:0] node12142;
	wire [4-1:0] node12146;
	wire [4-1:0] node12147;
	wire [4-1:0] node12148;
	wire [4-1:0] node12149;
	wire [4-1:0] node12152;
	wire [4-1:0] node12155;
	wire [4-1:0] node12157;
	wire [4-1:0] node12159;
	wire [4-1:0] node12162;
	wire [4-1:0] node12163;
	wire [4-1:0] node12164;
	wire [4-1:0] node12167;
	wire [4-1:0] node12168;
	wire [4-1:0] node12172;
	wire [4-1:0] node12175;
	wire [4-1:0] node12176;
	wire [4-1:0] node12177;
	wire [4-1:0] node12178;
	wire [4-1:0] node12179;
	wire [4-1:0] node12180;
	wire [4-1:0] node12181;
	wire [4-1:0] node12184;
	wire [4-1:0] node12188;
	wire [4-1:0] node12189;
	wire [4-1:0] node12193;
	wire [4-1:0] node12194;
	wire [4-1:0] node12195;
	wire [4-1:0] node12196;
	wire [4-1:0] node12199;
	wire [4-1:0] node12204;
	wire [4-1:0] node12205;
	wire [4-1:0] node12206;
	wire [4-1:0] node12209;
	wire [4-1:0] node12212;
	wire [4-1:0] node12213;
	wire [4-1:0] node12214;
	wire [4-1:0] node12215;
	wire [4-1:0] node12218;
	wire [4-1:0] node12222;
	wire [4-1:0] node12223;
	wire [4-1:0] node12224;
	wire [4-1:0] node12228;
	wire [4-1:0] node12229;
	wire [4-1:0] node12232;
	wire [4-1:0] node12235;
	wire [4-1:0] node12236;
	wire [4-1:0] node12237;
	wire [4-1:0] node12238;
	wire [4-1:0] node12241;
	wire [4-1:0] node12243;
	wire [4-1:0] node12244;
	wire [4-1:0] node12248;
	wire [4-1:0] node12249;
	wire [4-1:0] node12252;
	wire [4-1:0] node12253;
	wire [4-1:0] node12256;
	wire [4-1:0] node12259;
	wire [4-1:0] node12260;
	wire [4-1:0] node12261;
	wire [4-1:0] node12263;
	wire [4-1:0] node12267;
	wire [4-1:0] node12268;
	wire [4-1:0] node12271;
	wire [4-1:0] node12272;
	wire [4-1:0] node12275;
	wire [4-1:0] node12278;
	wire [4-1:0] node12279;
	wire [4-1:0] node12280;
	wire [4-1:0] node12281;
	wire [4-1:0] node12282;
	wire [4-1:0] node12283;
	wire [4-1:0] node12287;
	wire [4-1:0] node12288;
	wire [4-1:0] node12289;
	wire [4-1:0] node12291;
	wire [4-1:0] node12294;
	wire [4-1:0] node12296;
	wire [4-1:0] node12299;
	wire [4-1:0] node12300;
	wire [4-1:0] node12304;
	wire [4-1:0] node12305;
	wire [4-1:0] node12307;
	wire [4-1:0] node12308;
	wire [4-1:0] node12311;
	wire [4-1:0] node12314;
	wire [4-1:0] node12315;
	wire [4-1:0] node12316;
	wire [4-1:0] node12317;
	wire [4-1:0] node12320;
	wire [4-1:0] node12324;
	wire [4-1:0] node12325;
	wire [4-1:0] node12329;
	wire [4-1:0] node12330;
	wire [4-1:0] node12331;
	wire [4-1:0] node12333;
	wire [4-1:0] node12336;
	wire [4-1:0] node12338;
	wire [4-1:0] node12339;
	wire [4-1:0] node12342;
	wire [4-1:0] node12345;
	wire [4-1:0] node12346;
	wire [4-1:0] node12347;
	wire [4-1:0] node12349;
	wire [4-1:0] node12350;
	wire [4-1:0] node12353;
	wire [4-1:0] node12356;
	wire [4-1:0] node12357;
	wire [4-1:0] node12359;
	wire [4-1:0] node12363;
	wire [4-1:0] node12364;
	wire [4-1:0] node12365;
	wire [4-1:0] node12369;
	wire [4-1:0] node12370;
	wire [4-1:0] node12373;
	wire [4-1:0] node12376;
	wire [4-1:0] node12377;
	wire [4-1:0] node12378;
	wire [4-1:0] node12379;
	wire [4-1:0] node12380;
	wire [4-1:0] node12381;
	wire [4-1:0] node12385;
	wire [4-1:0] node12386;
	wire [4-1:0] node12388;
	wire [4-1:0] node12391;
	wire [4-1:0] node12394;
	wire [4-1:0] node12395;
	wire [4-1:0] node12397;
	wire [4-1:0] node12399;
	wire [4-1:0] node12402;
	wire [4-1:0] node12403;
	wire [4-1:0] node12404;
	wire [4-1:0] node12407;
	wire [4-1:0] node12411;
	wire [4-1:0] node12412;
	wire [4-1:0] node12413;
	wire [4-1:0] node12415;
	wire [4-1:0] node12418;
	wire [4-1:0] node12419;
	wire [4-1:0] node12423;
	wire [4-1:0] node12424;
	wire [4-1:0] node12425;
	wire [4-1:0] node12426;
	wire [4-1:0] node12430;
	wire [4-1:0] node12431;
	wire [4-1:0] node12435;
	wire [4-1:0] node12436;
	wire [4-1:0] node12440;
	wire [4-1:0] node12441;
	wire [4-1:0] node12442;
	wire [4-1:0] node12443;
	wire [4-1:0] node12444;
	wire [4-1:0] node12445;
	wire [4-1:0] node12449;
	wire [4-1:0] node12451;
	wire [4-1:0] node12454;
	wire [4-1:0] node12455;
	wire [4-1:0] node12459;
	wire [4-1:0] node12460;
	wire [4-1:0] node12461;
	wire [4-1:0] node12464;
	wire [4-1:0] node12467;
	wire [4-1:0] node12469;
	wire [4-1:0] node12472;
	wire [4-1:0] node12473;
	wire [4-1:0] node12474;
	wire [4-1:0] node12476;
	wire [4-1:0] node12479;
	wire [4-1:0] node12481;
	wire [4-1:0] node12483;
	wire [4-1:0] node12486;
	wire [4-1:0] node12488;
	wire [4-1:0] node12490;
	wire [4-1:0] node12493;
	wire [4-1:0] node12494;
	wire [4-1:0] node12495;
	wire [4-1:0] node12496;
	wire [4-1:0] node12497;
	wire [4-1:0] node12498;
	wire [4-1:0] node12499;
	wire [4-1:0] node12500;
	wire [4-1:0] node12501;
	wire [4-1:0] node12502;
	wire [4-1:0] node12503;
	wire [4-1:0] node12504;
	wire [4-1:0] node12506;
	wire [4-1:0] node12509;
	wire [4-1:0] node12512;
	wire [4-1:0] node12513;
	wire [4-1:0] node12514;
	wire [4-1:0] node12517;
	wire [4-1:0] node12521;
	wire [4-1:0] node12522;
	wire [4-1:0] node12523;
	wire [4-1:0] node12524;
	wire [4-1:0] node12527;
	wire [4-1:0] node12530;
	wire [4-1:0] node12532;
	wire [4-1:0] node12534;
	wire [4-1:0] node12537;
	wire [4-1:0] node12538;
	wire [4-1:0] node12539;
	wire [4-1:0] node12541;
	wire [4-1:0] node12544;
	wire [4-1:0] node12545;
	wire [4-1:0] node12548;
	wire [4-1:0] node12551;
	wire [4-1:0] node12554;
	wire [4-1:0] node12555;
	wire [4-1:0] node12556;
	wire [4-1:0] node12557;
	wire [4-1:0] node12559;
	wire [4-1:0] node12560;
	wire [4-1:0] node12563;
	wire [4-1:0] node12566;
	wire [4-1:0] node12569;
	wire [4-1:0] node12570;
	wire [4-1:0] node12571;
	wire [4-1:0] node12572;
	wire [4-1:0] node12575;
	wire [4-1:0] node12579;
	wire [4-1:0] node12582;
	wire [4-1:0] node12583;
	wire [4-1:0] node12584;
	wire [4-1:0] node12587;
	wire [4-1:0] node12588;
	wire [4-1:0] node12591;
	wire [4-1:0] node12592;
	wire [4-1:0] node12596;
	wire [4-1:0] node12597;
	wire [4-1:0] node12598;
	wire [4-1:0] node12602;
	wire [4-1:0] node12605;
	wire [4-1:0] node12606;
	wire [4-1:0] node12607;
	wire [4-1:0] node12608;
	wire [4-1:0] node12609;
	wire [4-1:0] node12610;
	wire [4-1:0] node12611;
	wire [4-1:0] node12614;
	wire [4-1:0] node12618;
	wire [4-1:0] node12619;
	wire [4-1:0] node12622;
	wire [4-1:0] node12625;
	wire [4-1:0] node12627;
	wire [4-1:0] node12628;
	wire [4-1:0] node12631;
	wire [4-1:0] node12634;
	wire [4-1:0] node12635;
	wire [4-1:0] node12636;
	wire [4-1:0] node12638;
	wire [4-1:0] node12639;
	wire [4-1:0] node12643;
	wire [4-1:0] node12645;
	wire [4-1:0] node12647;
	wire [4-1:0] node12651;
	wire [4-1:0] node12652;
	wire [4-1:0] node12653;
	wire [4-1:0] node12655;
	wire [4-1:0] node12656;
	wire [4-1:0] node12657;
	wire [4-1:0] node12661;
	wire [4-1:0] node12664;
	wire [4-1:0] node12665;
	wire [4-1:0] node12666;
	wire [4-1:0] node12668;
	wire [4-1:0] node12671;
	wire [4-1:0] node12672;
	wire [4-1:0] node12676;
	wire [4-1:0] node12677;
	wire [4-1:0] node12680;
	wire [4-1:0] node12681;
	wire [4-1:0] node12685;
	wire [4-1:0] node12686;
	wire [4-1:0] node12687;
	wire [4-1:0] node12691;
	wire [4-1:0] node12692;
	wire [4-1:0] node12694;
	wire [4-1:0] node12697;
	wire [4-1:0] node12698;
	wire [4-1:0] node12701;
	wire [4-1:0] node12704;
	wire [4-1:0] node12705;
	wire [4-1:0] node12706;
	wire [4-1:0] node12707;
	wire [4-1:0] node12708;
	wire [4-1:0] node12709;
	wire [4-1:0] node12711;
	wire [4-1:0] node12714;
	wire [4-1:0] node12717;
	wire [4-1:0] node12718;
	wire [4-1:0] node12720;
	wire [4-1:0] node12722;
	wire [4-1:0] node12725;
	wire [4-1:0] node12728;
	wire [4-1:0] node12729;
	wire [4-1:0] node12730;
	wire [4-1:0] node12731;
	wire [4-1:0] node12735;
	wire [4-1:0] node12736;
	wire [4-1:0] node12738;
	wire [4-1:0] node12742;
	wire [4-1:0] node12743;
	wire [4-1:0] node12745;
	wire [4-1:0] node12746;
	wire [4-1:0] node12750;
	wire [4-1:0] node12751;
	wire [4-1:0] node12755;
	wire [4-1:0] node12756;
	wire [4-1:0] node12757;
	wire [4-1:0] node12758;
	wire [4-1:0] node12760;
	wire [4-1:0] node12761;
	wire [4-1:0] node12764;
	wire [4-1:0] node12767;
	wire [4-1:0] node12768;
	wire [4-1:0] node12772;
	wire [4-1:0] node12773;
	wire [4-1:0] node12774;
	wire [4-1:0] node12777;
	wire [4-1:0] node12779;
	wire [4-1:0] node12782;
	wire [4-1:0] node12785;
	wire [4-1:0] node12786;
	wire [4-1:0] node12787;
	wire [4-1:0] node12788;
	wire [4-1:0] node12791;
	wire [4-1:0] node12794;
	wire [4-1:0] node12796;
	wire [4-1:0] node12798;
	wire [4-1:0] node12801;
	wire [4-1:0] node12802;
	wire [4-1:0] node12803;
	wire [4-1:0] node12807;
	wire [4-1:0] node12808;
	wire [4-1:0] node12810;
	wire [4-1:0] node12813;
	wire [4-1:0] node12816;
	wire [4-1:0] node12817;
	wire [4-1:0] node12818;
	wire [4-1:0] node12819;
	wire [4-1:0] node12820;
	wire [4-1:0] node12821;
	wire [4-1:0] node12823;
	wire [4-1:0] node12827;
	wire [4-1:0] node12830;
	wire [4-1:0] node12831;
	wire [4-1:0] node12832;
	wire [4-1:0] node12835;
	wire [4-1:0] node12838;
	wire [4-1:0] node12839;
	wire [4-1:0] node12843;
	wire [4-1:0] node12844;
	wire [4-1:0] node12845;
	wire [4-1:0] node12846;
	wire [4-1:0] node12851;
	wire [4-1:0] node12852;
	wire [4-1:0] node12853;
	wire [4-1:0] node12857;
	wire [4-1:0] node12859;
	wire [4-1:0] node12862;
	wire [4-1:0] node12863;
	wire [4-1:0] node12864;
	wire [4-1:0] node12865;
	wire [4-1:0] node12866;
	wire [4-1:0] node12870;
	wire [4-1:0] node12872;
	wire [4-1:0] node12874;
	wire [4-1:0] node12877;
	wire [4-1:0] node12878;
	wire [4-1:0] node12879;
	wire [4-1:0] node12883;
	wire [4-1:0] node12884;
	wire [4-1:0] node12887;
	wire [4-1:0] node12889;
	wire [4-1:0] node12892;
	wire [4-1:0] node12893;
	wire [4-1:0] node12895;
	wire [4-1:0] node12897;
	wire [4-1:0] node12898;
	wire [4-1:0] node12901;
	wire [4-1:0] node12904;
	wire [4-1:0] node12905;
	wire [4-1:0] node12907;
	wire [4-1:0] node12910;
	wire [4-1:0] node12911;
	wire [4-1:0] node12914;
	wire [4-1:0] node12917;
	wire [4-1:0] node12918;
	wire [4-1:0] node12919;
	wire [4-1:0] node12920;
	wire [4-1:0] node12921;
	wire [4-1:0] node12922;
	wire [4-1:0] node12923;
	wire [4-1:0] node12924;
	wire [4-1:0] node12926;
	wire [4-1:0] node12929;
	wire [4-1:0] node12930;
	wire [4-1:0] node12934;
	wire [4-1:0] node12937;
	wire [4-1:0] node12938;
	wire [4-1:0] node12940;
	wire [4-1:0] node12944;
	wire [4-1:0] node12945;
	wire [4-1:0] node12946;
	wire [4-1:0] node12950;
	wire [4-1:0] node12951;
	wire [4-1:0] node12953;
	wire [4-1:0] node12955;
	wire [4-1:0] node12958;
	wire [4-1:0] node12960;
	wire [4-1:0] node12963;
	wire [4-1:0] node12964;
	wire [4-1:0] node12965;
	wire [4-1:0] node12966;
	wire [4-1:0] node12968;
	wire [4-1:0] node12969;
	wire [4-1:0] node12973;
	wire [4-1:0] node12976;
	wire [4-1:0] node12977;
	wire [4-1:0] node12980;
	wire [4-1:0] node12982;
	wire [4-1:0] node12983;
	wire [4-1:0] node12986;
	wire [4-1:0] node12989;
	wire [4-1:0] node12990;
	wire [4-1:0] node12991;
	wire [4-1:0] node12992;
	wire [4-1:0] node12997;
	wire [4-1:0] node12998;
	wire [4-1:0] node12999;
	wire [4-1:0] node13002;
	wire [4-1:0] node13005;
	wire [4-1:0] node13007;
	wire [4-1:0] node13009;
	wire [4-1:0] node13012;
	wire [4-1:0] node13013;
	wire [4-1:0] node13014;
	wire [4-1:0] node13015;
	wire [4-1:0] node13017;
	wire [4-1:0] node13019;
	wire [4-1:0] node13020;
	wire [4-1:0] node13023;
	wire [4-1:0] node13026;
	wire [4-1:0] node13027;
	wire [4-1:0] node13028;
	wire [4-1:0] node13030;
	wire [4-1:0] node13033;
	wire [4-1:0] node13036;
	wire [4-1:0] node13037;
	wire [4-1:0] node13041;
	wire [4-1:0] node13042;
	wire [4-1:0] node13043;
	wire [4-1:0] node13044;
	wire [4-1:0] node13045;
	wire [4-1:0] node13050;
	wire [4-1:0] node13051;
	wire [4-1:0] node13052;
	wire [4-1:0] node13055;
	wire [4-1:0] node13059;
	wire [4-1:0] node13060;
	wire [4-1:0] node13062;
	wire [4-1:0] node13063;
	wire [4-1:0] node13067;
	wire [4-1:0] node13068;
	wire [4-1:0] node13071;
	wire [4-1:0] node13073;
	wire [4-1:0] node13076;
	wire [4-1:0] node13077;
	wire [4-1:0] node13078;
	wire [4-1:0] node13079;
	wire [4-1:0] node13082;
	wire [4-1:0] node13085;
	wire [4-1:0] node13086;
	wire [4-1:0] node13087;
	wire [4-1:0] node13089;
	wire [4-1:0] node13092;
	wire [4-1:0] node13093;
	wire [4-1:0] node13096;
	wire [4-1:0] node13099;
	wire [4-1:0] node13100;
	wire [4-1:0] node13101;
	wire [4-1:0] node13106;
	wire [4-1:0] node13107;
	wire [4-1:0] node13108;
	wire [4-1:0] node13110;
	wire [4-1:0] node13113;
	wire [4-1:0] node13114;
	wire [4-1:0] node13117;
	wire [4-1:0] node13118;
	wire [4-1:0] node13121;
	wire [4-1:0] node13124;
	wire [4-1:0] node13125;
	wire [4-1:0] node13126;
	wire [4-1:0] node13127;
	wire [4-1:0] node13132;
	wire [4-1:0] node13133;
	wire [4-1:0] node13137;
	wire [4-1:0] node13138;
	wire [4-1:0] node13139;
	wire [4-1:0] node13140;
	wire [4-1:0] node13141;
	wire [4-1:0] node13142;
	wire [4-1:0] node13143;
	wire [4-1:0] node13144;
	wire [4-1:0] node13147;
	wire [4-1:0] node13150;
	wire [4-1:0] node13151;
	wire [4-1:0] node13155;
	wire [4-1:0] node13158;
	wire [4-1:0] node13159;
	wire [4-1:0] node13160;
	wire [4-1:0] node13163;
	wire [4-1:0] node13165;
	wire [4-1:0] node13168;
	wire [4-1:0] node13171;
	wire [4-1:0] node13172;
	wire [4-1:0] node13173;
	wire [4-1:0] node13176;
	wire [4-1:0] node13177;
	wire [4-1:0] node13178;
	wire [4-1:0] node13183;
	wire [4-1:0] node13184;
	wire [4-1:0] node13187;
	wire [4-1:0] node13189;
	wire [4-1:0] node13190;
	wire [4-1:0] node13193;
	wire [4-1:0] node13196;
	wire [4-1:0] node13197;
	wire [4-1:0] node13198;
	wire [4-1:0] node13199;
	wire [4-1:0] node13201;
	wire [4-1:0] node13204;
	wire [4-1:0] node13205;
	wire [4-1:0] node13209;
	wire [4-1:0] node13210;
	wire [4-1:0] node13212;
	wire [4-1:0] node13216;
	wire [4-1:0] node13217;
	wire [4-1:0] node13218;
	wire [4-1:0] node13221;
	wire [4-1:0] node13222;
	wire [4-1:0] node13226;
	wire [4-1:0] node13227;
	wire [4-1:0] node13228;
	wire [4-1:0] node13229;
	wire [4-1:0] node13233;
	wire [4-1:0] node13236;
	wire [4-1:0] node13237;
	wire [4-1:0] node13240;
	wire [4-1:0] node13243;
	wire [4-1:0] node13244;
	wire [4-1:0] node13245;
	wire [4-1:0] node13246;
	wire [4-1:0] node13247;
	wire [4-1:0] node13248;
	wire [4-1:0] node13251;
	wire [4-1:0] node13254;
	wire [4-1:0] node13255;
	wire [4-1:0] node13256;
	wire [4-1:0] node13261;
	wire [4-1:0] node13262;
	wire [4-1:0] node13263;
	wire [4-1:0] node13266;
	wire [4-1:0] node13267;
	wire [4-1:0] node13271;
	wire [4-1:0] node13273;
	wire [4-1:0] node13276;
	wire [4-1:0] node13277;
	wire [4-1:0] node13279;
	wire [4-1:0] node13280;
	wire [4-1:0] node13282;
	wire [4-1:0] node13286;
	wire [4-1:0] node13288;
	wire [4-1:0] node13289;
	wire [4-1:0] node13291;
	wire [4-1:0] node13294;
	wire [4-1:0] node13297;
	wire [4-1:0] node13298;
	wire [4-1:0] node13299;
	wire [4-1:0] node13300;
	wire [4-1:0] node13302;
	wire [4-1:0] node13303;
	wire [4-1:0] node13306;
	wire [4-1:0] node13309;
	wire [4-1:0] node13310;
	wire [4-1:0] node13311;
	wire [4-1:0] node13315;
	wire [4-1:0] node13316;
	wire [4-1:0] node13320;
	wire [4-1:0] node13321;
	wire [4-1:0] node13323;
	wire [4-1:0] node13324;
	wire [4-1:0] node13328;
	wire [4-1:0] node13329;
	wire [4-1:0] node13333;
	wire [4-1:0] node13334;
	wire [4-1:0] node13335;
	wire [4-1:0] node13338;
	wire [4-1:0] node13339;
	wire [4-1:0] node13342;
	wire [4-1:0] node13344;
	wire [4-1:0] node13347;
	wire [4-1:0] node13348;
	wire [4-1:0] node13349;
	wire [4-1:0] node13351;
	wire [4-1:0] node13354;
	wire [4-1:0] node13355;
	wire [4-1:0] node13358;
	wire [4-1:0] node13361;
	wire [4-1:0] node13363;
	wire [4-1:0] node13364;
	wire [4-1:0] node13367;
	wire [4-1:0] node13370;
	wire [4-1:0] node13371;
	wire [4-1:0] node13372;
	wire [4-1:0] node13373;
	wire [4-1:0] node13374;
	wire [4-1:0] node13375;
	wire [4-1:0] node13376;
	wire [4-1:0] node13377;
	wire [4-1:0] node13378;
	wire [4-1:0] node13381;
	wire [4-1:0] node13383;
	wire [4-1:0] node13387;
	wire [4-1:0] node13388;
	wire [4-1:0] node13390;
	wire [4-1:0] node13393;
	wire [4-1:0] node13395;
	wire [4-1:0] node13396;
	wire [4-1:0] node13400;
	wire [4-1:0] node13401;
	wire [4-1:0] node13403;
	wire [4-1:0] node13404;
	wire [4-1:0] node13408;
	wire [4-1:0] node13409;
	wire [4-1:0] node13410;
	wire [4-1:0] node13412;
	wire [4-1:0] node13415;
	wire [4-1:0] node13417;
	wire [4-1:0] node13421;
	wire [4-1:0] node13422;
	wire [4-1:0] node13423;
	wire [4-1:0] node13424;
	wire [4-1:0] node13426;
	wire [4-1:0] node13429;
	wire [4-1:0] node13430;
	wire [4-1:0] node13432;
	wire [4-1:0] node13436;
	wire [4-1:0] node13437;
	wire [4-1:0] node13439;
	wire [4-1:0] node13441;
	wire [4-1:0] node13445;
	wire [4-1:0] node13446;
	wire [4-1:0] node13447;
	wire [4-1:0] node13448;
	wire [4-1:0] node13451;
	wire [4-1:0] node13454;
	wire [4-1:0] node13457;
	wire [4-1:0] node13458;
	wire [4-1:0] node13460;
	wire [4-1:0] node13462;
	wire [4-1:0] node13465;
	wire [4-1:0] node13467;
	wire [4-1:0] node13470;
	wire [4-1:0] node13471;
	wire [4-1:0] node13472;
	wire [4-1:0] node13473;
	wire [4-1:0] node13474;
	wire [4-1:0] node13477;
	wire [4-1:0] node13478;
	wire [4-1:0] node13482;
	wire [4-1:0] node13483;
	wire [4-1:0] node13484;
	wire [4-1:0] node13486;
	wire [4-1:0] node13491;
	wire [4-1:0] node13492;
	wire [4-1:0] node13493;
	wire [4-1:0] node13494;
	wire [4-1:0] node13498;
	wire [4-1:0] node13499;
	wire [4-1:0] node13502;
	wire [4-1:0] node13503;
	wire [4-1:0] node13507;
	wire [4-1:0] node13508;
	wire [4-1:0] node13509;
	wire [4-1:0] node13512;
	wire [4-1:0] node13515;
	wire [4-1:0] node13517;
	wire [4-1:0] node13520;
	wire [4-1:0] node13521;
	wire [4-1:0] node13522;
	wire [4-1:0] node13523;
	wire [4-1:0] node13526;
	wire [4-1:0] node13529;
	wire [4-1:0] node13531;
	wire [4-1:0] node13532;
	wire [4-1:0] node13535;
	wire [4-1:0] node13538;
	wire [4-1:0] node13539;
	wire [4-1:0] node13540;
	wire [4-1:0] node13542;
	wire [4-1:0] node13543;
	wire [4-1:0] node13547;
	wire [4-1:0] node13550;
	wire [4-1:0] node13551;
	wire [4-1:0] node13553;
	wire [4-1:0] node13556;
	wire [4-1:0] node13557;
	wire [4-1:0] node13558;
	wire [4-1:0] node13563;
	wire [4-1:0] node13564;
	wire [4-1:0] node13565;
	wire [4-1:0] node13566;
	wire [4-1:0] node13567;
	wire [4-1:0] node13568;
	wire [4-1:0] node13570;
	wire [4-1:0] node13573;
	wire [4-1:0] node13574;
	wire [4-1:0] node13576;
	wire [4-1:0] node13579;
	wire [4-1:0] node13582;
	wire [4-1:0] node13583;
	wire [4-1:0] node13585;
	wire [4-1:0] node13588;
	wire [4-1:0] node13590;
	wire [4-1:0] node13592;
	wire [4-1:0] node13595;
	wire [4-1:0] node13596;
	wire [4-1:0] node13599;
	wire [4-1:0] node13600;
	wire [4-1:0] node13601;
	wire [4-1:0] node13603;
	wire [4-1:0] node13606;
	wire [4-1:0] node13608;
	wire [4-1:0] node13611;
	wire [4-1:0] node13613;
	wire [4-1:0] node13616;
	wire [4-1:0] node13617;
	wire [4-1:0] node13618;
	wire [4-1:0] node13619;
	wire [4-1:0] node13620;
	wire [4-1:0] node13621;
	wire [4-1:0] node13624;
	wire [4-1:0] node13627;
	wire [4-1:0] node13629;
	wire [4-1:0] node13632;
	wire [4-1:0] node13634;
	wire [4-1:0] node13636;
	wire [4-1:0] node13639;
	wire [4-1:0] node13640;
	wire [4-1:0] node13642;
	wire [4-1:0] node13645;
	wire [4-1:0] node13647;
	wire [4-1:0] node13650;
	wire [4-1:0] node13651;
	wire [4-1:0] node13652;
	wire [4-1:0] node13655;
	wire [4-1:0] node13657;
	wire [4-1:0] node13660;
	wire [4-1:0] node13661;
	wire [4-1:0] node13662;
	wire [4-1:0] node13665;
	wire [4-1:0] node13668;
	wire [4-1:0] node13669;
	wire [4-1:0] node13670;
	wire [4-1:0] node13675;
	wire [4-1:0] node13676;
	wire [4-1:0] node13677;
	wire [4-1:0] node13678;
	wire [4-1:0] node13679;
	wire [4-1:0] node13680;
	wire [4-1:0] node13684;
	wire [4-1:0] node13687;
	wire [4-1:0] node13688;
	wire [4-1:0] node13689;
	wire [4-1:0] node13692;
	wire [4-1:0] node13695;
	wire [4-1:0] node13697;
	wire [4-1:0] node13700;
	wire [4-1:0] node13701;
	wire [4-1:0] node13702;
	wire [4-1:0] node13703;
	wire [4-1:0] node13706;
	wire [4-1:0] node13709;
	wire [4-1:0] node13710;
	wire [4-1:0] node13713;
	wire [4-1:0] node13715;
	wire [4-1:0] node13718;
	wire [4-1:0] node13719;
	wire [4-1:0] node13720;
	wire [4-1:0] node13724;
	wire [4-1:0] node13725;
	wire [4-1:0] node13726;
	wire [4-1:0] node13730;
	wire [4-1:0] node13732;
	wire [4-1:0] node13735;
	wire [4-1:0] node13736;
	wire [4-1:0] node13737;
	wire [4-1:0] node13739;
	wire [4-1:0] node13740;
	wire [4-1:0] node13742;
	wire [4-1:0] node13746;
	wire [4-1:0] node13747;
	wire [4-1:0] node13751;
	wire [4-1:0] node13752;
	wire [4-1:0] node13753;
	wire [4-1:0] node13755;
	wire [4-1:0] node13758;
	wire [4-1:0] node13761;
	wire [4-1:0] node13763;
	wire [4-1:0] node13764;
	wire [4-1:0] node13765;
	wire [4-1:0] node13768;
	wire [4-1:0] node13772;
	wire [4-1:0] node13773;
	wire [4-1:0] node13774;
	wire [4-1:0] node13775;
	wire [4-1:0] node13776;
	wire [4-1:0] node13777;
	wire [4-1:0] node13780;
	wire [4-1:0] node13781;
	wire [4-1:0] node13782;
	wire [4-1:0] node13786;
	wire [4-1:0] node13787;
	wire [4-1:0] node13788;
	wire [4-1:0] node13793;
	wire [4-1:0] node13794;
	wire [4-1:0] node13795;
	wire [4-1:0] node13797;
	wire [4-1:0] node13799;
	wire [4-1:0] node13802;
	wire [4-1:0] node13805;
	wire [4-1:0] node13806;
	wire [4-1:0] node13808;
	wire [4-1:0] node13811;
	wire [4-1:0] node13812;
	wire [4-1:0] node13814;
	wire [4-1:0] node13818;
	wire [4-1:0] node13819;
	wire [4-1:0] node13820;
	wire [4-1:0] node13821;
	wire [4-1:0] node13822;
	wire [4-1:0] node13826;
	wire [4-1:0] node13827;
	wire [4-1:0] node13830;
	wire [4-1:0] node13831;
	wire [4-1:0] node13835;
	wire [4-1:0] node13836;
	wire [4-1:0] node13838;
	wire [4-1:0] node13839;
	wire [4-1:0] node13842;
	wire [4-1:0] node13845;
	wire [4-1:0] node13846;
	wire [4-1:0] node13847;
	wire [4-1:0] node13851;
	wire [4-1:0] node13853;
	wire [4-1:0] node13856;
	wire [4-1:0] node13857;
	wire [4-1:0] node13858;
	wire [4-1:0] node13859;
	wire [4-1:0] node13862;
	wire [4-1:0] node13865;
	wire [4-1:0] node13866;
	wire [4-1:0] node13870;
	wire [4-1:0] node13871;
	wire [4-1:0] node13875;
	wire [4-1:0] node13876;
	wire [4-1:0] node13877;
	wire [4-1:0] node13878;
	wire [4-1:0] node13879;
	wire [4-1:0] node13880;
	wire [4-1:0] node13883;
	wire [4-1:0] node13886;
	wire [4-1:0] node13889;
	wire [4-1:0] node13890;
	wire [4-1:0] node13891;
	wire [4-1:0] node13894;
	wire [4-1:0] node13897;
	wire [4-1:0] node13898;
	wire [4-1:0] node13901;
	wire [4-1:0] node13904;
	wire [4-1:0] node13905;
	wire [4-1:0] node13906;
	wire [4-1:0] node13908;
	wire [4-1:0] node13911;
	wire [4-1:0] node13913;
	wire [4-1:0] node13915;
	wire [4-1:0] node13918;
	wire [4-1:0] node13919;
	wire [4-1:0] node13920;
	wire [4-1:0] node13921;
	wire [4-1:0] node13924;
	wire [4-1:0] node13927;
	wire [4-1:0] node13929;
	wire [4-1:0] node13932;
	wire [4-1:0] node13935;
	wire [4-1:0] node13936;
	wire [4-1:0] node13937;
	wire [4-1:0] node13938;
	wire [4-1:0] node13939;
	wire [4-1:0] node13943;
	wire [4-1:0] node13946;
	wire [4-1:0] node13947;
	wire [4-1:0] node13949;
	wire [4-1:0] node13952;
	wire [4-1:0] node13953;
	wire [4-1:0] node13954;
	wire [4-1:0] node13957;
	wire [4-1:0] node13960;
	wire [4-1:0] node13963;
	wire [4-1:0] node13964;
	wire [4-1:0] node13965;
	wire [4-1:0] node13966;
	wire [4-1:0] node13967;
	wire [4-1:0] node13970;
	wire [4-1:0] node13973;
	wire [4-1:0] node13976;
	wire [4-1:0] node13978;
	wire [4-1:0] node13980;
	wire [4-1:0] node13983;
	wire [4-1:0] node13984;
	wire [4-1:0] node13987;
	wire [4-1:0] node13988;
	wire [4-1:0] node13990;
	wire [4-1:0] node13994;
	wire [4-1:0] node13995;
	wire [4-1:0] node13996;
	wire [4-1:0] node13997;
	wire [4-1:0] node13998;
	wire [4-1:0] node14000;
	wire [4-1:0] node14001;
	wire [4-1:0] node14002;
	wire [4-1:0] node14005;
	wire [4-1:0] node14009;
	wire [4-1:0] node14010;
	wire [4-1:0] node14011;
	wire [4-1:0] node14013;
	wire [4-1:0] node14016;
	wire [4-1:0] node14018;
	wire [4-1:0] node14021;
	wire [4-1:0] node14023;
	wire [4-1:0] node14024;
	wire [4-1:0] node14028;
	wire [4-1:0] node14029;
	wire [4-1:0] node14030;
	wire [4-1:0] node14032;
	wire [4-1:0] node14035;
	wire [4-1:0] node14036;
	wire [4-1:0] node14038;
	wire [4-1:0] node14041;
	wire [4-1:0] node14042;
	wire [4-1:0] node14046;
	wire [4-1:0] node14047;
	wire [4-1:0] node14049;
	wire [4-1:0] node14051;
	wire [4-1:0] node14054;
	wire [4-1:0] node14055;
	wire [4-1:0] node14056;
	wire [4-1:0] node14060;
	wire [4-1:0] node14063;
	wire [4-1:0] node14064;
	wire [4-1:0] node14065;
	wire [4-1:0] node14066;
	wire [4-1:0] node14067;
	wire [4-1:0] node14070;
	wire [4-1:0] node14073;
	wire [4-1:0] node14076;
	wire [4-1:0] node14077;
	wire [4-1:0] node14079;
	wire [4-1:0] node14080;
	wire [4-1:0] node14083;
	wire [4-1:0] node14086;
	wire [4-1:0] node14087;
	wire [4-1:0] node14088;
	wire [4-1:0] node14092;
	wire [4-1:0] node14095;
	wire [4-1:0] node14096;
	wire [4-1:0] node14097;
	wire [4-1:0] node14098;
	wire [4-1:0] node14102;
	wire [4-1:0] node14105;
	wire [4-1:0] node14106;
	wire [4-1:0] node14107;
	wire [4-1:0] node14110;
	wire [4-1:0] node14113;
	wire [4-1:0] node14114;
	wire [4-1:0] node14117;
	wire [4-1:0] node14119;
	wire [4-1:0] node14122;
	wire [4-1:0] node14123;
	wire [4-1:0] node14124;
	wire [4-1:0] node14125;
	wire [4-1:0] node14127;
	wire [4-1:0] node14129;
	wire [4-1:0] node14132;
	wire [4-1:0] node14133;
	wire [4-1:0] node14134;
	wire [4-1:0] node14137;
	wire [4-1:0] node14140;
	wire [4-1:0] node14141;
	wire [4-1:0] node14143;
	wire [4-1:0] node14147;
	wire [4-1:0] node14148;
	wire [4-1:0] node14149;
	wire [4-1:0] node14153;
	wire [4-1:0] node14155;
	wire [4-1:0] node14156;
	wire [4-1:0] node14158;
	wire [4-1:0] node14162;
	wire [4-1:0] node14163;
	wire [4-1:0] node14164;
	wire [4-1:0] node14166;
	wire [4-1:0] node14167;
	wire [4-1:0] node14171;
	wire [4-1:0] node14172;
	wire [4-1:0] node14174;
	wire [4-1:0] node14178;
	wire [4-1:0] node14179;
	wire [4-1:0] node14181;
	wire [4-1:0] node14182;
	wire [4-1:0] node14183;
	wire [4-1:0] node14186;
	wire [4-1:0] node14189;
	wire [4-1:0] node14191;
	wire [4-1:0] node14194;
	wire [4-1:0] node14195;
	wire [4-1:0] node14198;
	wire [4-1:0] node14201;
	wire [4-1:0] node14202;
	wire [4-1:0] node14203;
	wire [4-1:0] node14204;
	wire [4-1:0] node14205;
	wire [4-1:0] node14206;
	wire [4-1:0] node14207;
	wire [4-1:0] node14208;
	wire [4-1:0] node14209;
	wire [4-1:0] node14212;
	wire [4-1:0] node14215;
	wire [4-1:0] node14216;
	wire [4-1:0] node14217;
	wire [4-1:0] node14219;
	wire [4-1:0] node14222;
	wire [4-1:0] node14224;
	wire [4-1:0] node14227;
	wire [4-1:0] node14228;
	wire [4-1:0] node14232;
	wire [4-1:0] node14233;
	wire [4-1:0] node14235;
	wire [4-1:0] node14236;
	wire [4-1:0] node14240;
	wire [4-1:0] node14241;
	wire [4-1:0] node14244;
	wire [4-1:0] node14246;
	wire [4-1:0] node14249;
	wire [4-1:0] node14250;
	wire [4-1:0] node14251;
	wire [4-1:0] node14252;
	wire [4-1:0] node14253;
	wire [4-1:0] node14254;
	wire [4-1:0] node14257;
	wire [4-1:0] node14260;
	wire [4-1:0] node14261;
	wire [4-1:0] node14265;
	wire [4-1:0] node14267;
	wire [4-1:0] node14269;
	wire [4-1:0] node14272;
	wire [4-1:0] node14273;
	wire [4-1:0] node14274;
	wire [4-1:0] node14277;
	wire [4-1:0] node14280;
	wire [4-1:0] node14281;
	wire [4-1:0] node14283;
	wire [4-1:0] node14287;
	wire [4-1:0] node14288;
	wire [4-1:0] node14289;
	wire [4-1:0] node14290;
	wire [4-1:0] node14291;
	wire [4-1:0] node14294;
	wire [4-1:0] node14297;
	wire [4-1:0] node14300;
	wire [4-1:0] node14303;
	wire [4-1:0] node14304;
	wire [4-1:0] node14305;
	wire [4-1:0] node14306;
	wire [4-1:0] node14310;
	wire [4-1:0] node14312;
	wire [4-1:0] node14315;
	wire [4-1:0] node14316;
	wire [4-1:0] node14318;
	wire [4-1:0] node14322;
	wire [4-1:0] node14323;
	wire [4-1:0] node14324;
	wire [4-1:0] node14325;
	wire [4-1:0] node14327;
	wire [4-1:0] node14330;
	wire [4-1:0] node14331;
	wire [4-1:0] node14332;
	wire [4-1:0] node14336;
	wire [4-1:0] node14339;
	wire [4-1:0] node14340;
	wire [4-1:0] node14341;
	wire [4-1:0] node14342;
	wire [4-1:0] node14346;
	wire [4-1:0] node14348;
	wire [4-1:0] node14351;
	wire [4-1:0] node14353;
	wire [4-1:0] node14355;
	wire [4-1:0] node14358;
	wire [4-1:0] node14359;
	wire [4-1:0] node14360;
	wire [4-1:0] node14361;
	wire [4-1:0] node14365;
	wire [4-1:0] node14368;
	wire [4-1:0] node14369;
	wire [4-1:0] node14370;
	wire [4-1:0] node14373;
	wire [4-1:0] node14376;
	wire [4-1:0] node14377;
	wire [4-1:0] node14378;
	wire [4-1:0] node14382;
	wire [4-1:0] node14383;
	wire [4-1:0] node14387;
	wire [4-1:0] node14388;
	wire [4-1:0] node14389;
	wire [4-1:0] node14390;
	wire [4-1:0] node14391;
	wire [4-1:0] node14393;
	wire [4-1:0] node14396;
	wire [4-1:0] node14397;
	wire [4-1:0] node14398;
	wire [4-1:0] node14402;
	wire [4-1:0] node14404;
	wire [4-1:0] node14406;
	wire [4-1:0] node14409;
	wire [4-1:0] node14410;
	wire [4-1:0] node14412;
	wire [4-1:0] node14414;
	wire [4-1:0] node14417;
	wire [4-1:0] node14418;
	wire [4-1:0] node14419;
	wire [4-1:0] node14424;
	wire [4-1:0] node14425;
	wire [4-1:0] node14426;
	wire [4-1:0] node14428;
	wire [4-1:0] node14430;
	wire [4-1:0] node14431;
	wire [4-1:0] node14434;
	wire [4-1:0] node14437;
	wire [4-1:0] node14438;
	wire [4-1:0] node14439;
	wire [4-1:0] node14443;
	wire [4-1:0] node14445;
	wire [4-1:0] node14446;
	wire [4-1:0] node14449;
	wire [4-1:0] node14452;
	wire [4-1:0] node14453;
	wire [4-1:0] node14454;
	wire [4-1:0] node14456;
	wire [4-1:0] node14459;
	wire [4-1:0] node14461;
	wire [4-1:0] node14462;
	wire [4-1:0] node14466;
	wire [4-1:0] node14467;
	wire [4-1:0] node14468;
	wire [4-1:0] node14472;
	wire [4-1:0] node14473;
	wire [4-1:0] node14474;
	wire [4-1:0] node14479;
	wire [4-1:0] node14480;
	wire [4-1:0] node14481;
	wire [4-1:0] node14482;
	wire [4-1:0] node14483;
	wire [4-1:0] node14485;
	wire [4-1:0] node14488;
	wire [4-1:0] node14491;
	wire [4-1:0] node14492;
	wire [4-1:0] node14494;
	wire [4-1:0] node14497;
	wire [4-1:0] node14499;
	wire [4-1:0] node14502;
	wire [4-1:0] node14503;
	wire [4-1:0] node14504;
	wire [4-1:0] node14505;
	wire [4-1:0] node14509;
	wire [4-1:0] node14512;
	wire [4-1:0] node14513;
	wire [4-1:0] node14514;
	wire [4-1:0] node14515;
	wire [4-1:0] node14520;
	wire [4-1:0] node14521;
	wire [4-1:0] node14522;
	wire [4-1:0] node14527;
	wire [4-1:0] node14528;
	wire [4-1:0] node14529;
	wire [4-1:0] node14530;
	wire [4-1:0] node14534;
	wire [4-1:0] node14535;
	wire [4-1:0] node14536;
	wire [4-1:0] node14541;
	wire [4-1:0] node14542;
	wire [4-1:0] node14543;
	wire [4-1:0] node14544;
	wire [4-1:0] node14545;
	wire [4-1:0] node14549;
	wire [4-1:0] node14550;
	wire [4-1:0] node14554;
	wire [4-1:0] node14555;
	wire [4-1:0] node14559;
	wire [4-1:0] node14560;
	wire [4-1:0] node14561;
	wire [4-1:0] node14562;
	wire [4-1:0] node14567;
	wire [4-1:0] node14569;
	wire [4-1:0] node14572;
	wire [4-1:0] node14573;
	wire [4-1:0] node14574;
	wire [4-1:0] node14575;
	wire [4-1:0] node14576;
	wire [4-1:0] node14577;
	wire [4-1:0] node14579;
	wire [4-1:0] node14580;
	wire [4-1:0] node14584;
	wire [4-1:0] node14586;
	wire [4-1:0] node14588;
	wire [4-1:0] node14591;
	wire [4-1:0] node14592;
	wire [4-1:0] node14594;
	wire [4-1:0] node14595;
	wire [4-1:0] node14599;
	wire [4-1:0] node14600;
	wire [4-1:0] node14601;
	wire [4-1:0] node14604;
	wire [4-1:0] node14606;
	wire [4-1:0] node14610;
	wire [4-1:0] node14611;
	wire [4-1:0] node14612;
	wire [4-1:0] node14613;
	wire [4-1:0] node14617;
	wire [4-1:0] node14618;
	wire [4-1:0] node14620;
	wire [4-1:0] node14621;
	wire [4-1:0] node14624;
	wire [4-1:0] node14627;
	wire [4-1:0] node14628;
	wire [4-1:0] node14629;
	wire [4-1:0] node14633;
	wire [4-1:0] node14636;
	wire [4-1:0] node14637;
	wire [4-1:0] node14638;
	wire [4-1:0] node14639;
	wire [4-1:0] node14641;
	wire [4-1:0] node14645;
	wire [4-1:0] node14646;
	wire [4-1:0] node14650;
	wire [4-1:0] node14651;
	wire [4-1:0] node14653;
	wire [4-1:0] node14656;
	wire [4-1:0] node14658;
	wire [4-1:0] node14661;
	wire [4-1:0] node14662;
	wire [4-1:0] node14663;
	wire [4-1:0] node14664;
	wire [4-1:0] node14665;
	wire [4-1:0] node14667;
	wire [4-1:0] node14670;
	wire [4-1:0] node14671;
	wire [4-1:0] node14672;
	wire [4-1:0] node14676;
	wire [4-1:0] node14677;
	wire [4-1:0] node14681;
	wire [4-1:0] node14682;
	wire [4-1:0] node14684;
	wire [4-1:0] node14687;
	wire [4-1:0] node14690;
	wire [4-1:0] node14691;
	wire [4-1:0] node14692;
	wire [4-1:0] node14693;
	wire [4-1:0] node14696;
	wire [4-1:0] node14698;
	wire [4-1:0] node14701;
	wire [4-1:0] node14703;
	wire [4-1:0] node14705;
	wire [4-1:0] node14708;
	wire [4-1:0] node14710;
	wire [4-1:0] node14712;
	wire [4-1:0] node14714;
	wire [4-1:0] node14717;
	wire [4-1:0] node14718;
	wire [4-1:0] node14719;
	wire [4-1:0] node14720;
	wire [4-1:0] node14721;
	wire [4-1:0] node14723;
	wire [4-1:0] node14727;
	wire [4-1:0] node14730;
	wire [4-1:0] node14731;
	wire [4-1:0] node14732;
	wire [4-1:0] node14734;
	wire [4-1:0] node14738;
	wire [4-1:0] node14739;
	wire [4-1:0] node14743;
	wire [4-1:0] node14744;
	wire [4-1:0] node14745;
	wire [4-1:0] node14748;
	wire [4-1:0] node14749;
	wire [4-1:0] node14751;
	wire [4-1:0] node14755;
	wire [4-1:0] node14756;
	wire [4-1:0] node14759;
	wire [4-1:0] node14760;
	wire [4-1:0] node14762;
	wire [4-1:0] node14765;
	wire [4-1:0] node14767;
	wire [4-1:0] node14770;
	wire [4-1:0] node14771;
	wire [4-1:0] node14772;
	wire [4-1:0] node14773;
	wire [4-1:0] node14774;
	wire [4-1:0] node14775;
	wire [4-1:0] node14776;
	wire [4-1:0] node14779;
	wire [4-1:0] node14782;
	wire [4-1:0] node14783;
	wire [4-1:0] node14787;
	wire [4-1:0] node14788;
	wire [4-1:0] node14789;
	wire [4-1:0] node14792;
	wire [4-1:0] node14796;
	wire [4-1:0] node14797;
	wire [4-1:0] node14798;
	wire [4-1:0] node14799;
	wire [4-1:0] node14802;
	wire [4-1:0] node14805;
	wire [4-1:0] node14807;
	wire [4-1:0] node14810;
	wire [4-1:0] node14811;
	wire [4-1:0] node14812;
	wire [4-1:0] node14814;
	wire [4-1:0] node14818;
	wire [4-1:0] node14820;
	wire [4-1:0] node14822;
	wire [4-1:0] node14825;
	wire [4-1:0] node14826;
	wire [4-1:0] node14827;
	wire [4-1:0] node14828;
	wire [4-1:0] node14832;
	wire [4-1:0] node14834;
	wire [4-1:0] node14835;
	wire [4-1:0] node14838;
	wire [4-1:0] node14841;
	wire [4-1:0] node14842;
	wire [4-1:0] node14843;
	wire [4-1:0] node14846;
	wire [4-1:0] node14849;
	wire [4-1:0] node14850;
	wire [4-1:0] node14853;
	wire [4-1:0] node14855;
	wire [4-1:0] node14858;
	wire [4-1:0] node14859;
	wire [4-1:0] node14860;
	wire [4-1:0] node14861;
	wire [4-1:0] node14862;
	wire [4-1:0] node14863;
	wire [4-1:0] node14867;
	wire [4-1:0] node14871;
	wire [4-1:0] node14872;
	wire [4-1:0] node14873;
	wire [4-1:0] node14874;
	wire [4-1:0] node14875;
	wire [4-1:0] node14878;
	wire [4-1:0] node14881;
	wire [4-1:0] node14883;
	wire [4-1:0] node14886;
	wire [4-1:0] node14887;
	wire [4-1:0] node14891;
	wire [4-1:0] node14892;
	wire [4-1:0] node14893;
	wire [4-1:0] node14894;
	wire [4-1:0] node14899;
	wire [4-1:0] node14900;
	wire [4-1:0] node14901;
	wire [4-1:0] node14904;
	wire [4-1:0] node14908;
	wire [4-1:0] node14909;
	wire [4-1:0] node14910;
	wire [4-1:0] node14911;
	wire [4-1:0] node14912;
	wire [4-1:0] node14916;
	wire [4-1:0] node14919;
	wire [4-1:0] node14920;
	wire [4-1:0] node14923;
	wire [4-1:0] node14926;
	wire [4-1:0] node14927;
	wire [4-1:0] node14928;
	wire [4-1:0] node14931;
	wire [4-1:0] node14932;
	wire [4-1:0] node14934;
	wire [4-1:0] node14938;
	wire [4-1:0] node14939;
	wire [4-1:0] node14940;
	wire [4-1:0] node14944;
	wire [4-1:0] node14947;
	wire [4-1:0] node14948;
	wire [4-1:0] node14949;
	wire [4-1:0] node14950;
	wire [4-1:0] node14951;
	wire [4-1:0] node14952;
	wire [4-1:0] node14953;
	wire [4-1:0] node14954;
	wire [4-1:0] node14955;
	wire [4-1:0] node14959;
	wire [4-1:0] node14960;
	wire [4-1:0] node14963;
	wire [4-1:0] node14966;
	wire [4-1:0] node14967;
	wire [4-1:0] node14968;
	wire [4-1:0] node14969;
	wire [4-1:0] node14973;
	wire [4-1:0] node14977;
	wire [4-1:0] node14978;
	wire [4-1:0] node14979;
	wire [4-1:0] node14981;
	wire [4-1:0] node14984;
	wire [4-1:0] node14986;
	wire [4-1:0] node14989;
	wire [4-1:0] node14990;
	wire [4-1:0] node14991;
	wire [4-1:0] node14994;
	wire [4-1:0] node14997;
	wire [4-1:0] node15000;
	wire [4-1:0] node15001;
	wire [4-1:0] node15002;
	wire [4-1:0] node15003;
	wire [4-1:0] node15004;
	wire [4-1:0] node15007;
	wire [4-1:0] node15010;
	wire [4-1:0] node15011;
	wire [4-1:0] node15015;
	wire [4-1:0] node15016;
	wire [4-1:0] node15017;
	wire [4-1:0] node15020;
	wire [4-1:0] node15022;
	wire [4-1:0] node15025;
	wire [4-1:0] node15026;
	wire [4-1:0] node15030;
	wire [4-1:0] node15031;
	wire [4-1:0] node15032;
	wire [4-1:0] node15033;
	wire [4-1:0] node15035;
	wire [4-1:0] node15040;
	wire [4-1:0] node15042;
	wire [4-1:0] node15043;
	wire [4-1:0] node15046;
	wire [4-1:0] node15049;
	wire [4-1:0] node15050;
	wire [4-1:0] node15051;
	wire [4-1:0] node15052;
	wire [4-1:0] node15053;
	wire [4-1:0] node15054;
	wire [4-1:0] node15059;
	wire [4-1:0] node15061;
	wire [4-1:0] node15062;
	wire [4-1:0] node15063;
	wire [4-1:0] node15066;
	wire [4-1:0] node15069;
	wire [4-1:0] node15070;
	wire [4-1:0] node15073;
	wire [4-1:0] node15076;
	wire [4-1:0] node15077;
	wire [4-1:0] node15078;
	wire [4-1:0] node15079;
	wire [4-1:0] node15082;
	wire [4-1:0] node15085;
	wire [4-1:0] node15087;
	wire [4-1:0] node15090;
	wire [4-1:0] node15091;
	wire [4-1:0] node15093;
	wire [4-1:0] node15096;
	wire [4-1:0] node15097;
	wire [4-1:0] node15098;
	wire [4-1:0] node15102;
	wire [4-1:0] node15105;
	wire [4-1:0] node15106;
	wire [4-1:0] node15107;
	wire [4-1:0] node15108;
	wire [4-1:0] node15109;
	wire [4-1:0] node15113;
	wire [4-1:0] node15116;
	wire [4-1:0] node15118;
	wire [4-1:0] node15119;
	wire [4-1:0] node15123;
	wire [4-1:0] node15124;
	wire [4-1:0] node15125;
	wire [4-1:0] node15126;
	wire [4-1:0] node15131;
	wire [4-1:0] node15134;
	wire [4-1:0] node15135;
	wire [4-1:0] node15136;
	wire [4-1:0] node15137;
	wire [4-1:0] node15138;
	wire [4-1:0] node15139;
	wire [4-1:0] node15140;
	wire [4-1:0] node15142;
	wire [4-1:0] node15146;
	wire [4-1:0] node15147;
	wire [4-1:0] node15148;
	wire [4-1:0] node15151;
	wire [4-1:0] node15155;
	wire [4-1:0] node15156;
	wire [4-1:0] node15160;
	wire [4-1:0] node15161;
	wire [4-1:0] node15162;
	wire [4-1:0] node15164;
	wire [4-1:0] node15167;
	wire [4-1:0] node15169;
	wire [4-1:0] node15172;
	wire [4-1:0] node15174;
	wire [4-1:0] node15177;
	wire [4-1:0] node15178;
	wire [4-1:0] node15179;
	wire [4-1:0] node15181;
	wire [4-1:0] node15183;
	wire [4-1:0] node15184;
	wire [4-1:0] node15187;
	wire [4-1:0] node15190;
	wire [4-1:0] node15191;
	wire [4-1:0] node15193;
	wire [4-1:0] node15196;
	wire [4-1:0] node15198;
	wire [4-1:0] node15201;
	wire [4-1:0] node15202;
	wire [4-1:0] node15203;
	wire [4-1:0] node15207;
	wire [4-1:0] node15208;
	wire [4-1:0] node15209;
	wire [4-1:0] node15211;
	wire [4-1:0] node15214;
	wire [4-1:0] node15215;
	wire [4-1:0] node15218;
	wire [4-1:0] node15222;
	wire [4-1:0] node15223;
	wire [4-1:0] node15224;
	wire [4-1:0] node15225;
	wire [4-1:0] node15226;
	wire [4-1:0] node15227;
	wire [4-1:0] node15230;
	wire [4-1:0] node15233;
	wire [4-1:0] node15234;
	wire [4-1:0] node15235;
	wire [4-1:0] node15238;
	wire [4-1:0] node15242;
	wire [4-1:0] node15243;
	wire [4-1:0] node15245;
	wire [4-1:0] node15248;
	wire [4-1:0] node15251;
	wire [4-1:0] node15252;
	wire [4-1:0] node15253;
	wire [4-1:0] node15254;
	wire [4-1:0] node15258;
	wire [4-1:0] node15260;
	wire [4-1:0] node15263;
	wire [4-1:0] node15264;
	wire [4-1:0] node15268;
	wire [4-1:0] node15269;
	wire [4-1:0] node15270;
	wire [4-1:0] node15271;
	wire [4-1:0] node15273;
	wire [4-1:0] node15274;
	wire [4-1:0] node15277;
	wire [4-1:0] node15281;
	wire [4-1:0] node15283;
	wire [4-1:0] node15284;
	wire [4-1:0] node15288;
	wire [4-1:0] node15289;
	wire [4-1:0] node15291;
	wire [4-1:0] node15293;
	wire [4-1:0] node15296;
	wire [4-1:0] node15297;
	wire [4-1:0] node15299;
	wire [4-1:0] node15302;
	wire [4-1:0] node15303;
	wire [4-1:0] node15307;
	wire [4-1:0] node15308;
	wire [4-1:0] node15309;
	wire [4-1:0] node15310;
	wire [4-1:0] node15311;
	wire [4-1:0] node15312;
	wire [4-1:0] node15314;
	wire [4-1:0] node15317;
	wire [4-1:0] node15319;
	wire [4-1:0] node15321;
	wire [4-1:0] node15324;
	wire [4-1:0] node15325;
	wire [4-1:0] node15327;
	wire [4-1:0] node15329;
	wire [4-1:0] node15332;
	wire [4-1:0] node15333;
	wire [4-1:0] node15335;
	wire [4-1:0] node15338;
	wire [4-1:0] node15340;
	wire [4-1:0] node15343;
	wire [4-1:0] node15344;
	wire [4-1:0] node15345;
	wire [4-1:0] node15346;
	wire [4-1:0] node15347;
	wire [4-1:0] node15350;
	wire [4-1:0] node15353;
	wire [4-1:0] node15355;
	wire [4-1:0] node15358;
	wire [4-1:0] node15359;
	wire [4-1:0] node15360;
	wire [4-1:0] node15361;
	wire [4-1:0] node15364;
	wire [4-1:0] node15368;
	wire [4-1:0] node15370;
	wire [4-1:0] node15373;
	wire [4-1:0] node15374;
	wire [4-1:0] node15375;
	wire [4-1:0] node15377;
	wire [4-1:0] node15380;
	wire [4-1:0] node15381;
	wire [4-1:0] node15382;
	wire [4-1:0] node15387;
	wire [4-1:0] node15389;
	wire [4-1:0] node15390;
	wire [4-1:0] node15393;
	wire [4-1:0] node15396;
	wire [4-1:0] node15397;
	wire [4-1:0] node15398;
	wire [4-1:0] node15399;
	wire [4-1:0] node15400;
	wire [4-1:0] node15401;
	wire [4-1:0] node15406;
	wire [4-1:0] node15407;
	wire [4-1:0] node15408;
	wire [4-1:0] node15410;
	wire [4-1:0] node15415;
	wire [4-1:0] node15416;
	wire [4-1:0] node15417;
	wire [4-1:0] node15419;
	wire [4-1:0] node15422;
	wire [4-1:0] node15424;
	wire [4-1:0] node15427;
	wire [4-1:0] node15429;
	wire [4-1:0] node15430;
	wire [4-1:0] node15433;
	wire [4-1:0] node15436;
	wire [4-1:0] node15437;
	wire [4-1:0] node15438;
	wire [4-1:0] node15439;
	wire [4-1:0] node15440;
	wire [4-1:0] node15441;
	wire [4-1:0] node15444;
	wire [4-1:0] node15447;
	wire [4-1:0] node15449;
	wire [4-1:0] node15452;
	wire [4-1:0] node15454;
	wire [4-1:0] node15456;
	wire [4-1:0] node15459;
	wire [4-1:0] node15461;
	wire [4-1:0] node15462;
	wire [4-1:0] node15466;
	wire [4-1:0] node15468;
	wire [4-1:0] node15469;
	wire [4-1:0] node15470;
	wire [4-1:0] node15474;
	wire [4-1:0] node15475;
	wire [4-1:0] node15479;
	wire [4-1:0] node15480;
	wire [4-1:0] node15481;
	wire [4-1:0] node15482;
	wire [4-1:0] node15483;
	wire [4-1:0] node15484;
	wire [4-1:0] node15485;
	wire [4-1:0] node15489;
	wire [4-1:0] node15490;
	wire [4-1:0] node15491;
	wire [4-1:0] node15494;
	wire [4-1:0] node15497;
	wire [4-1:0] node15499;
	wire [4-1:0] node15502;
	wire [4-1:0] node15504;
	wire [4-1:0] node15505;
	wire [4-1:0] node15506;
	wire [4-1:0] node15509;
	wire [4-1:0] node15513;
	wire [4-1:0] node15514;
	wire [4-1:0] node15516;
	wire [4-1:0] node15517;
	wire [4-1:0] node15518;
	wire [4-1:0] node15521;
	wire [4-1:0] node15524;
	wire [4-1:0] node15526;
	wire [4-1:0] node15529;
	wire [4-1:0] node15530;
	wire [4-1:0] node15532;
	wire [4-1:0] node15533;
	wire [4-1:0] node15536;
	wire [4-1:0] node15539;
	wire [4-1:0] node15541;
	wire [4-1:0] node15542;
	wire [4-1:0] node15546;
	wire [4-1:0] node15547;
	wire [4-1:0] node15548;
	wire [4-1:0] node15549;
	wire [4-1:0] node15551;
	wire [4-1:0] node15552;
	wire [4-1:0] node15556;
	wire [4-1:0] node15558;
	wire [4-1:0] node15561;
	wire [4-1:0] node15562;
	wire [4-1:0] node15563;
	wire [4-1:0] node15567;
	wire [4-1:0] node15568;
	wire [4-1:0] node15572;
	wire [4-1:0] node15573;
	wire [4-1:0] node15574;
	wire [4-1:0] node15576;
	wire [4-1:0] node15577;
	wire [4-1:0] node15580;
	wire [4-1:0] node15584;
	wire [4-1:0] node15585;
	wire [4-1:0] node15586;
	wire [4-1:0] node15590;
	wire [4-1:0] node15591;
	wire [4-1:0] node15594;
	wire [4-1:0] node15597;
	wire [4-1:0] node15598;
	wire [4-1:0] node15599;
	wire [4-1:0] node15600;
	wire [4-1:0] node15601;
	wire [4-1:0] node15602;
	wire [4-1:0] node15605;
	wire [4-1:0] node15609;
	wire [4-1:0] node15610;
	wire [4-1:0] node15611;
	wire [4-1:0] node15613;
	wire [4-1:0] node15616;
	wire [4-1:0] node15619;
	wire [4-1:0] node15621;
	wire [4-1:0] node15622;
	wire [4-1:0] node15625;
	wire [4-1:0] node15628;
	wire [4-1:0] node15629;
	wire [4-1:0] node15630;
	wire [4-1:0] node15632;
	wire [4-1:0] node15634;
	wire [4-1:0] node15638;
	wire [4-1:0] node15640;
	wire [4-1:0] node15641;
	wire [4-1:0] node15644;
	wire [4-1:0] node15645;
	wire [4-1:0] node15649;
	wire [4-1:0] node15650;
	wire [4-1:0] node15651;
	wire [4-1:0] node15652;
	wire [4-1:0] node15654;
	wire [4-1:0] node15658;
	wire [4-1:0] node15659;
	wire [4-1:0] node15660;
	wire [4-1:0] node15661;
	wire [4-1:0] node15665;
	wire [4-1:0] node15668;
	wire [4-1:0] node15671;
	wire [4-1:0] node15672;
	wire [4-1:0] node15673;
	wire [4-1:0] node15676;
	wire [4-1:0] node15677;
	wire [4-1:0] node15679;
	wire [4-1:0] node15683;
	wire [4-1:0] node15684;
	wire [4-1:0] node15687;
	wire [4-1:0] node15689;
	wire [4-1:0] node15692;
	wire [4-1:0] node15693;
	wire [4-1:0] node15694;
	wire [4-1:0] node15695;
	wire [4-1:0] node15696;
	wire [4-1:0] node15697;
	wire [4-1:0] node15698;
	wire [4-1:0] node15699;
	wire [4-1:0] node15700;
	wire [4-1:0] node15701;
	wire [4-1:0] node15703;
	wire [4-1:0] node15707;
	wire [4-1:0] node15708;
	wire [4-1:0] node15711;
	wire [4-1:0] node15713;
	wire [4-1:0] node15716;
	wire [4-1:0] node15717;
	wire [4-1:0] node15719;
	wire [4-1:0] node15721;
	wire [4-1:0] node15722;
	wire [4-1:0] node15725;
	wire [4-1:0] node15728;
	wire [4-1:0] node15730;
	wire [4-1:0] node15731;
	wire [4-1:0] node15735;
	wire [4-1:0] node15736;
	wire [4-1:0] node15737;
	wire [4-1:0] node15739;
	wire [4-1:0] node15742;
	wire [4-1:0] node15743;
	wire [4-1:0] node15745;
	wire [4-1:0] node15748;
	wire [4-1:0] node15749;
	wire [4-1:0] node15752;
	wire [4-1:0] node15754;
	wire [4-1:0] node15757;
	wire [4-1:0] node15758;
	wire [4-1:0] node15759;
	wire [4-1:0] node15760;
	wire [4-1:0] node15763;
	wire [4-1:0] node15767;
	wire [4-1:0] node15769;
	wire [4-1:0] node15770;
	wire [4-1:0] node15773;
	wire [4-1:0] node15774;
	wire [4-1:0] node15778;
	wire [4-1:0] node15779;
	wire [4-1:0] node15780;
	wire [4-1:0] node15781;
	wire [4-1:0] node15783;
	wire [4-1:0] node15784;
	wire [4-1:0] node15788;
	wire [4-1:0] node15789;
	wire [4-1:0] node15790;
	wire [4-1:0] node15794;
	wire [4-1:0] node15796;
	wire [4-1:0] node15797;
	wire [4-1:0] node15800;
	wire [4-1:0] node15803;
	wire [4-1:0] node15804;
	wire [4-1:0] node15805;
	wire [4-1:0] node15806;
	wire [4-1:0] node15809;
	wire [4-1:0] node15812;
	wire [4-1:0] node15814;
	wire [4-1:0] node15817;
	wire [4-1:0] node15818;
	wire [4-1:0] node15819;
	wire [4-1:0] node15824;
	wire [4-1:0] node15825;
	wire [4-1:0] node15826;
	wire [4-1:0] node15827;
	wire [4-1:0] node15828;
	wire [4-1:0] node15832;
	wire [4-1:0] node15833;
	wire [4-1:0] node15835;
	wire [4-1:0] node15838;
	wire [4-1:0] node15839;
	wire [4-1:0] node15843;
	wire [4-1:0] node15844;
	wire [4-1:0] node15846;
	wire [4-1:0] node15850;
	wire [4-1:0] node15851;
	wire [4-1:0] node15852;
	wire [4-1:0] node15856;
	wire [4-1:0] node15857;
	wire [4-1:0] node15859;
	wire [4-1:0] node15862;
	wire [4-1:0] node15863;
	wire [4-1:0] node15867;
	wire [4-1:0] node15868;
	wire [4-1:0] node15869;
	wire [4-1:0] node15870;
	wire [4-1:0] node15871;
	wire [4-1:0] node15872;
	wire [4-1:0] node15873;
	wire [4-1:0] node15878;
	wire [4-1:0] node15880;
	wire [4-1:0] node15883;
	wire [4-1:0] node15884;
	wire [4-1:0] node15885;
	wire [4-1:0] node15887;
	wire [4-1:0] node15891;
	wire [4-1:0] node15892;
	wire [4-1:0] node15893;
	wire [4-1:0] node15897;
	wire [4-1:0] node15899;
	wire [4-1:0] node15902;
	wire [4-1:0] node15903;
	wire [4-1:0] node15904;
	wire [4-1:0] node15905;
	wire [4-1:0] node15906;
	wire [4-1:0] node15910;
	wire [4-1:0] node15913;
	wire [4-1:0] node15914;
	wire [4-1:0] node15917;
	wire [4-1:0] node15918;
	wire [4-1:0] node15921;
	wire [4-1:0] node15924;
	wire [4-1:0] node15925;
	wire [4-1:0] node15926;
	wire [4-1:0] node15928;
	wire [4-1:0] node15930;
	wire [4-1:0] node15933;
	wire [4-1:0] node15935;
	wire [4-1:0] node15936;
	wire [4-1:0] node15939;
	wire [4-1:0] node15942;
	wire [4-1:0] node15943;
	wire [4-1:0] node15945;
	wire [4-1:0] node15948;
	wire [4-1:0] node15951;
	wire [4-1:0] node15952;
	wire [4-1:0] node15953;
	wire [4-1:0] node15954;
	wire [4-1:0] node15955;
	wire [4-1:0] node15956;
	wire [4-1:0] node15960;
	wire [4-1:0] node15961;
	wire [4-1:0] node15965;
	wire [4-1:0] node15966;
	wire [4-1:0] node15968;
	wire [4-1:0] node15969;
	wire [4-1:0] node15973;
	wire [4-1:0] node15974;
	wire [4-1:0] node15975;
	wire [4-1:0] node15978;
	wire [4-1:0] node15982;
	wire [4-1:0] node15983;
	wire [4-1:0] node15984;
	wire [4-1:0] node15985;
	wire [4-1:0] node15989;
	wire [4-1:0] node15990;
	wire [4-1:0] node15993;
	wire [4-1:0] node15996;
	wire [4-1:0] node15997;
	wire [4-1:0] node15998;
	wire [4-1:0] node16002;
	wire [4-1:0] node16005;
	wire [4-1:0] node16006;
	wire [4-1:0] node16007;
	wire [4-1:0] node16009;
	wire [4-1:0] node16010;
	wire [4-1:0] node16013;
	wire [4-1:0] node16016;
	wire [4-1:0] node16017;
	wire [4-1:0] node16019;
	wire [4-1:0] node16021;
	wire [4-1:0] node16024;
	wire [4-1:0] node16025;
	wire [4-1:0] node16029;
	wire [4-1:0] node16030;
	wire [4-1:0] node16031;
	wire [4-1:0] node16033;
	wire [4-1:0] node16034;
	wire [4-1:0] node16037;
	wire [4-1:0] node16040;
	wire [4-1:0] node16041;
	wire [4-1:0] node16045;
	wire [4-1:0] node16046;
	wire [4-1:0] node16047;
	wire [4-1:0] node16050;
	wire [4-1:0] node16053;
	wire [4-1:0] node16055;
	wire [4-1:0] node16058;
	wire [4-1:0] node16059;
	wire [4-1:0] node16060;
	wire [4-1:0] node16061;
	wire [4-1:0] node16062;
	wire [4-1:0] node16063;
	wire [4-1:0] node16064;
	wire [4-1:0] node16065;
	wire [4-1:0] node16069;
	wire [4-1:0] node16072;
	wire [4-1:0] node16073;
	wire [4-1:0] node16074;
	wire [4-1:0] node16077;
	wire [4-1:0] node16081;
	wire [4-1:0] node16082;
	wire [4-1:0] node16083;
	wire [4-1:0] node16084;
	wire [4-1:0] node16087;
	wire [4-1:0] node16088;
	wire [4-1:0] node16092;
	wire [4-1:0] node16093;
	wire [4-1:0] node16095;
	wire [4-1:0] node16098;
	wire [4-1:0] node16100;
	wire [4-1:0] node16103;
	wire [4-1:0] node16104;
	wire [4-1:0] node16106;
	wire [4-1:0] node16109;
	wire [4-1:0] node16110;
	wire [4-1:0] node16114;
	wire [4-1:0] node16115;
	wire [4-1:0] node16116;
	wire [4-1:0] node16117;
	wire [4-1:0] node16119;
	wire [4-1:0] node16122;
	wire [4-1:0] node16124;
	wire [4-1:0] node16127;
	wire [4-1:0] node16128;
	wire [4-1:0] node16129;
	wire [4-1:0] node16133;
	wire [4-1:0] node16134;
	wire [4-1:0] node16137;
	wire [4-1:0] node16140;
	wire [4-1:0] node16141;
	wire [4-1:0] node16143;
	wire [4-1:0] node16146;
	wire [4-1:0] node16147;
	wire [4-1:0] node16148;
	wire [4-1:0] node16149;
	wire [4-1:0] node16154;
	wire [4-1:0] node16155;
	wire [4-1:0] node16156;
	wire [4-1:0] node16159;
	wire [4-1:0] node16163;
	wire [4-1:0] node16164;
	wire [4-1:0] node16165;
	wire [4-1:0] node16166;
	wire [4-1:0] node16167;
	wire [4-1:0] node16169;
	wire [4-1:0] node16172;
	wire [4-1:0] node16174;
	wire [4-1:0] node16176;
	wire [4-1:0] node16179;
	wire [4-1:0] node16180;
	wire [4-1:0] node16181;
	wire [4-1:0] node16185;
	wire [4-1:0] node16186;
	wire [4-1:0] node16190;
	wire [4-1:0] node16191;
	wire [4-1:0] node16192;
	wire [4-1:0] node16194;
	wire [4-1:0] node16196;
	wire [4-1:0] node16199;
	wire [4-1:0] node16200;
	wire [4-1:0] node16203;
	wire [4-1:0] node16206;
	wire [4-1:0] node16207;
	wire [4-1:0] node16208;
	wire [4-1:0] node16212;
	wire [4-1:0] node16214;
	wire [4-1:0] node16217;
	wire [4-1:0] node16218;
	wire [4-1:0] node16219;
	wire [4-1:0] node16220;
	wire [4-1:0] node16223;
	wire [4-1:0] node16225;
	wire [4-1:0] node16228;
	wire [4-1:0] node16230;
	wire [4-1:0] node16233;
	wire [4-1:0] node16234;
	wire [4-1:0] node16235;
	wire [4-1:0] node16236;
	wire [4-1:0] node16238;
	wire [4-1:0] node16242;
	wire [4-1:0] node16243;
	wire [4-1:0] node16247;
	wire [4-1:0] node16249;
	wire [4-1:0] node16251;
	wire [4-1:0] node16254;
	wire [4-1:0] node16255;
	wire [4-1:0] node16256;
	wire [4-1:0] node16257;
	wire [4-1:0] node16258;
	wire [4-1:0] node16259;
	wire [4-1:0] node16260;
	wire [4-1:0] node16263;
	wire [4-1:0] node16267;
	wire [4-1:0] node16268;
	wire [4-1:0] node16270;
	wire [4-1:0] node16271;
	wire [4-1:0] node16274;
	wire [4-1:0] node16277;
	wire [4-1:0] node16279;
	wire [4-1:0] node16282;
	wire [4-1:0] node16283;
	wire [4-1:0] node16284;
	wire [4-1:0] node16286;
	wire [4-1:0] node16289;
	wire [4-1:0] node16291;
	wire [4-1:0] node16292;
	wire [4-1:0] node16295;
	wire [4-1:0] node16298;
	wire [4-1:0] node16299;
	wire [4-1:0] node16300;
	wire [4-1:0] node16301;
	wire [4-1:0] node16305;
	wire [4-1:0] node16306;
	wire [4-1:0] node16309;
	wire [4-1:0] node16312;
	wire [4-1:0] node16314;
	wire [4-1:0] node16316;
	wire [4-1:0] node16319;
	wire [4-1:0] node16320;
	wire [4-1:0] node16321;
	wire [4-1:0] node16323;
	wire [4-1:0] node16325;
	wire [4-1:0] node16326;
	wire [4-1:0] node16330;
	wire [4-1:0] node16331;
	wire [4-1:0] node16332;
	wire [4-1:0] node16336;
	wire [4-1:0] node16337;
	wire [4-1:0] node16341;
	wire [4-1:0] node16342;
	wire [4-1:0] node16343;
	wire [4-1:0] node16344;
	wire [4-1:0] node16345;
	wire [4-1:0] node16350;
	wire [4-1:0] node16351;
	wire [4-1:0] node16354;
	wire [4-1:0] node16357;
	wire [4-1:0] node16358;
	wire [4-1:0] node16359;
	wire [4-1:0] node16362;
	wire [4-1:0] node16365;
	wire [4-1:0] node16368;
	wire [4-1:0] node16369;
	wire [4-1:0] node16370;
	wire [4-1:0] node16371;
	wire [4-1:0] node16372;
	wire [4-1:0] node16374;
	wire [4-1:0] node16378;
	wire [4-1:0] node16379;
	wire [4-1:0] node16382;
	wire [4-1:0] node16384;
	wire [4-1:0] node16387;
	wire [4-1:0] node16388;
	wire [4-1:0] node16389;
	wire [4-1:0] node16393;
	wire [4-1:0] node16394;
	wire [4-1:0] node16398;
	wire [4-1:0] node16399;
	wire [4-1:0] node16400;
	wire [4-1:0] node16401;
	wire [4-1:0] node16403;
	wire [4-1:0] node16406;
	wire [4-1:0] node16407;
	wire [4-1:0] node16411;
	wire [4-1:0] node16413;
	wire [4-1:0] node16414;
	wire [4-1:0] node16415;
	wire [4-1:0] node16418;
	wire [4-1:0] node16422;
	wire [4-1:0] node16423;
	wire [4-1:0] node16424;
	wire [4-1:0] node16426;
	wire [4-1:0] node16427;
	wire [4-1:0] node16431;
	wire [4-1:0] node16434;
	wire [4-1:0] node16435;
	wire [4-1:0] node16439;
	wire [4-1:0] node16440;
	wire [4-1:0] node16441;
	wire [4-1:0] node16442;
	wire [4-1:0] node16443;
	wire [4-1:0] node16444;
	wire [4-1:0] node16445;
	wire [4-1:0] node16446;
	wire [4-1:0] node16448;
	wire [4-1:0] node16451;
	wire [4-1:0] node16454;
	wire [4-1:0] node16455;
	wire [4-1:0] node16459;
	wire [4-1:0] node16460;
	wire [4-1:0] node16462;
	wire [4-1:0] node16465;
	wire [4-1:0] node16468;
	wire [4-1:0] node16469;
	wire [4-1:0] node16470;
	wire [4-1:0] node16472;
	wire [4-1:0] node16475;
	wire [4-1:0] node16477;
	wire [4-1:0] node16478;
	wire [4-1:0] node16482;
	wire [4-1:0] node16483;
	wire [4-1:0] node16484;
	wire [4-1:0] node16487;
	wire [4-1:0] node16491;
	wire [4-1:0] node16492;
	wire [4-1:0] node16493;
	wire [4-1:0] node16494;
	wire [4-1:0] node16495;
	wire [4-1:0] node16497;
	wire [4-1:0] node16500;
	wire [4-1:0] node16501;
	wire [4-1:0] node16505;
	wire [4-1:0] node16507;
	wire [4-1:0] node16509;
	wire [4-1:0] node16512;
	wire [4-1:0] node16513;
	wire [4-1:0] node16514;
	wire [4-1:0] node16515;
	wire [4-1:0] node16516;
	wire [4-1:0] node16519;
	wire [4-1:0] node16523;
	wire [4-1:0] node16524;
	wire [4-1:0] node16526;
	wire [4-1:0] node16530;
	wire [4-1:0] node16531;
	wire [4-1:0] node16532;
	wire [4-1:0] node16534;
	wire [4-1:0] node16537;
	wire [4-1:0] node16538;
	wire [4-1:0] node16542;
	wire [4-1:0] node16545;
	wire [4-1:0] node16546;
	wire [4-1:0] node16547;
	wire [4-1:0] node16548;
	wire [4-1:0] node16549;
	wire [4-1:0] node16552;
	wire [4-1:0] node16555;
	wire [4-1:0] node16556;
	wire [4-1:0] node16559;
	wire [4-1:0] node16560;
	wire [4-1:0] node16563;
	wire [4-1:0] node16566;
	wire [4-1:0] node16567;
	wire [4-1:0] node16568;
	wire [4-1:0] node16572;
	wire [4-1:0] node16575;
	wire [4-1:0] node16576;
	wire [4-1:0] node16577;
	wire [4-1:0] node16578;
	wire [4-1:0] node16579;
	wire [4-1:0] node16584;
	wire [4-1:0] node16585;
	wire [4-1:0] node16588;
	wire [4-1:0] node16591;
	wire [4-1:0] node16593;
	wire [4-1:0] node16596;
	wire [4-1:0] node16597;
	wire [4-1:0] node16598;
	wire [4-1:0] node16599;
	wire [4-1:0] node16600;
	wire [4-1:0] node16601;
	wire [4-1:0] node16603;
	wire [4-1:0] node16606;
	wire [4-1:0] node16607;
	wire [4-1:0] node16611;
	wire [4-1:0] node16612;
	wire [4-1:0] node16613;
	wire [4-1:0] node16614;
	wire [4-1:0] node16617;
	wire [4-1:0] node16622;
	wire [4-1:0] node16623;
	wire [4-1:0] node16624;
	wire [4-1:0] node16625;
	wire [4-1:0] node16629;
	wire [4-1:0] node16631;
	wire [4-1:0] node16634;
	wire [4-1:0] node16635;
	wire [4-1:0] node16636;
	wire [4-1:0] node16638;
	wire [4-1:0] node16641;
	wire [4-1:0] node16644;
	wire [4-1:0] node16646;
	wire [4-1:0] node16647;
	wire [4-1:0] node16650;
	wire [4-1:0] node16653;
	wire [4-1:0] node16654;
	wire [4-1:0] node16655;
	wire [4-1:0] node16656;
	wire [4-1:0] node16658;
	wire [4-1:0] node16661;
	wire [4-1:0] node16664;
	wire [4-1:0] node16665;
	wire [4-1:0] node16667;
	wire [4-1:0] node16671;
	wire [4-1:0] node16672;
	wire [4-1:0] node16673;
	wire [4-1:0] node16674;
	wire [4-1:0] node16676;
	wire [4-1:0] node16680;
	wire [4-1:0] node16681;
	wire [4-1:0] node16682;
	wire [4-1:0] node16685;
	wire [4-1:0] node16689;
	wire [4-1:0] node16690;
	wire [4-1:0] node16694;
	wire [4-1:0] node16695;
	wire [4-1:0] node16696;
	wire [4-1:0] node16697;
	wire [4-1:0] node16698;
	wire [4-1:0] node16699;
	wire [4-1:0] node16700;
	wire [4-1:0] node16704;
	wire [4-1:0] node16707;
	wire [4-1:0] node16709;
	wire [4-1:0] node16711;
	wire [4-1:0] node16714;
	wire [4-1:0] node16715;
	wire [4-1:0] node16716;
	wire [4-1:0] node16719;
	wire [4-1:0] node16720;
	wire [4-1:0] node16724;
	wire [4-1:0] node16727;
	wire [4-1:0] node16728;
	wire [4-1:0] node16729;
	wire [4-1:0] node16730;
	wire [4-1:0] node16732;
	wire [4-1:0] node16735;
	wire [4-1:0] node16737;
	wire [4-1:0] node16740;
	wire [4-1:0] node16741;
	wire [4-1:0] node16742;
	wire [4-1:0] node16747;
	wire [4-1:0] node16748;
	wire [4-1:0] node16749;
	wire [4-1:0] node16752;
	wire [4-1:0] node16755;
	wire [4-1:0] node16758;
	wire [4-1:0] node16759;
	wire [4-1:0] node16760;
	wire [4-1:0] node16761;
	wire [4-1:0] node16764;
	wire [4-1:0] node16765;
	wire [4-1:0] node16769;
	wire [4-1:0] node16770;
	wire [4-1:0] node16773;
	wire [4-1:0] node16776;
	wire [4-1:0] node16778;
	wire [4-1:0] node16779;
	wire [4-1:0] node16782;
	wire [4-1:0] node16785;
	wire [4-1:0] node16786;
	wire [4-1:0] node16787;
	wire [4-1:0] node16788;
	wire [4-1:0] node16789;
	wire [4-1:0] node16790;
	wire [4-1:0] node16791;
	wire [4-1:0] node16793;
	wire [4-1:0] node16796;
	wire [4-1:0] node16799;
	wire [4-1:0] node16800;
	wire [4-1:0] node16802;
	wire [4-1:0] node16805;
	wire [4-1:0] node16806;
	wire [4-1:0] node16809;
	wire [4-1:0] node16811;
	wire [4-1:0] node16814;
	wire [4-1:0] node16815;
	wire [4-1:0] node16816;
	wire [4-1:0] node16819;
	wire [4-1:0] node16820;
	wire [4-1:0] node16823;
	wire [4-1:0] node16824;
	wire [4-1:0] node16827;
	wire [4-1:0] node16830;
	wire [4-1:0] node16831;
	wire [4-1:0] node16832;
	wire [4-1:0] node16836;
	wire [4-1:0] node16837;
	wire [4-1:0] node16841;
	wire [4-1:0] node16842;
	wire [4-1:0] node16843;
	wire [4-1:0] node16846;
	wire [4-1:0] node16847;
	wire [4-1:0] node16850;
	wire [4-1:0] node16851;
	wire [4-1:0] node16855;
	wire [4-1:0] node16856;
	wire [4-1:0] node16857;
	wire [4-1:0] node16860;
	wire [4-1:0] node16861;
	wire [4-1:0] node16865;
	wire [4-1:0] node16868;
	wire [4-1:0] node16869;
	wire [4-1:0] node16870;
	wire [4-1:0] node16871;
	wire [4-1:0] node16872;
	wire [4-1:0] node16874;
	wire [4-1:0] node16877;
	wire [4-1:0] node16878;
	wire [4-1:0] node16880;
	wire [4-1:0] node16883;
	wire [4-1:0] node16884;
	wire [4-1:0] node16888;
	wire [4-1:0] node16889;
	wire [4-1:0] node16890;
	wire [4-1:0] node16894;
	wire [4-1:0] node16895;
	wire [4-1:0] node16897;
	wire [4-1:0] node16900;
	wire [4-1:0] node16901;
	wire [4-1:0] node16904;
	wire [4-1:0] node16907;
	wire [4-1:0] node16908;
	wire [4-1:0] node16909;
	wire [4-1:0] node16910;
	wire [4-1:0] node16913;
	wire [4-1:0] node16916;
	wire [4-1:0] node16917;
	wire [4-1:0] node16919;
	wire [4-1:0] node16922;
	wire [4-1:0] node16923;
	wire [4-1:0] node16926;
	wire [4-1:0] node16929;
	wire [4-1:0] node16932;
	wire [4-1:0] node16933;
	wire [4-1:0] node16934;
	wire [4-1:0] node16935;
	wire [4-1:0] node16936;
	wire [4-1:0] node16941;
	wire [4-1:0] node16942;
	wire [4-1:0] node16943;
	wire [4-1:0] node16948;
	wire [4-1:0] node16949;
	wire [4-1:0] node16951;
	wire [4-1:0] node16954;
	wire [4-1:0] node16956;
	wire [4-1:0] node16957;
	wire [4-1:0] node16961;
	wire [4-1:0] node16962;
	wire [4-1:0] node16963;
	wire [4-1:0] node16964;
	wire [4-1:0] node16965;
	wire [4-1:0] node16967;
	wire [4-1:0] node16969;
	wire [4-1:0] node16971;
	wire [4-1:0] node16974;
	wire [4-1:0] node16975;
	wire [4-1:0] node16976;
	wire [4-1:0] node16980;
	wire [4-1:0] node16981;
	wire [4-1:0] node16982;
	wire [4-1:0] node16987;
	wire [4-1:0] node16988;
	wire [4-1:0] node16989;
	wire [4-1:0] node16991;
	wire [4-1:0] node16994;
	wire [4-1:0] node16996;
	wire [4-1:0] node16997;
	wire [4-1:0] node17000;
	wire [4-1:0] node17003;
	wire [4-1:0] node17005;
	wire [4-1:0] node17007;
	wire [4-1:0] node17010;
	wire [4-1:0] node17011;
	wire [4-1:0] node17012;
	wire [4-1:0] node17013;
	wire [4-1:0] node17014;
	wire [4-1:0] node17017;
	wire [4-1:0] node17020;
	wire [4-1:0] node17022;
	wire [4-1:0] node17024;
	wire [4-1:0] node17027;
	wire [4-1:0] node17028;
	wire [4-1:0] node17030;
	wire [4-1:0] node17032;
	wire [4-1:0] node17035;
	wire [4-1:0] node17036;
	wire [4-1:0] node17038;
	wire [4-1:0] node17041;
	wire [4-1:0] node17042;
	wire [4-1:0] node17046;
	wire [4-1:0] node17047;
	wire [4-1:0] node17048;
	wire [4-1:0] node17049;
	wire [4-1:0] node17050;
	wire [4-1:0] node17053;
	wire [4-1:0] node17057;
	wire [4-1:0] node17059;
	wire [4-1:0] node17062;
	wire [4-1:0] node17063;
	wire [4-1:0] node17066;
	wire [4-1:0] node17067;
	wire [4-1:0] node17071;
	wire [4-1:0] node17072;
	wire [4-1:0] node17073;
	wire [4-1:0] node17074;
	wire [4-1:0] node17075;
	wire [4-1:0] node17077;
	wire [4-1:0] node17080;
	wire [4-1:0] node17081;
	wire [4-1:0] node17083;
	wire [4-1:0] node17087;
	wire [4-1:0] node17089;
	wire [4-1:0] node17090;
	wire [4-1:0] node17093;
	wire [4-1:0] node17096;
	wire [4-1:0] node17097;
	wire [4-1:0] node17098;
	wire [4-1:0] node17099;
	wire [4-1:0] node17102;
	wire [4-1:0] node17103;
	wire [4-1:0] node17107;
	wire [4-1:0] node17109;
	wire [4-1:0] node17112;
	wire [4-1:0] node17113;
	wire [4-1:0] node17114;
	wire [4-1:0] node17115;
	wire [4-1:0] node17119;
	wire [4-1:0] node17120;
	wire [4-1:0] node17125;
	wire [4-1:0] node17126;
	wire [4-1:0] node17127;
	wire [4-1:0] node17128;
	wire [4-1:0] node17129;
	wire [4-1:0] node17132;
	wire [4-1:0] node17134;
	wire [4-1:0] node17137;
	wire [4-1:0] node17138;
	wire [4-1:0] node17141;
	wire [4-1:0] node17144;
	wire [4-1:0] node17147;
	wire [4-1:0] node17148;
	wire [4-1:0] node17149;
	wire [4-1:0] node17150;
	wire [4-1:0] node17151;
	wire [4-1:0] node17156;
	wire [4-1:0] node17157;
	wire [4-1:0] node17161;
	wire [4-1:0] node17162;
	wire [4-1:0] node17164;
	wire [4-1:0] node17167;
	wire [4-1:0] node17168;
	wire [4-1:0] node17171;
	wire [4-1:0] node17174;
	wire [4-1:0] node17175;
	wire [4-1:0] node17176;
	wire [4-1:0] node17177;
	wire [4-1:0] node17178;
	wire [4-1:0] node17179;
	wire [4-1:0] node17180;
	wire [4-1:0] node17181;
	wire [4-1:0] node17182;
	wire [4-1:0] node17183;
	wire [4-1:0] node17188;
	wire [4-1:0] node17190;
	wire [4-1:0] node17192;
	wire [4-1:0] node17195;
	wire [4-1:0] node17196;
	wire [4-1:0] node17197;
	wire [4-1:0] node17199;
	wire [4-1:0] node17201;
	wire [4-1:0] node17204;
	wire [4-1:0] node17205;
	wire [4-1:0] node17208;
	wire [4-1:0] node17211;
	wire [4-1:0] node17212;
	wire [4-1:0] node17213;
	wire [4-1:0] node17214;
	wire [4-1:0] node17218;
	wire [4-1:0] node17219;
	wire [4-1:0] node17223;
	wire [4-1:0] node17225;
	wire [4-1:0] node17228;
	wire [4-1:0] node17229;
	wire [4-1:0] node17230;
	wire [4-1:0] node17231;
	wire [4-1:0] node17233;
	wire [4-1:0] node17236;
	wire [4-1:0] node17237;
	wire [4-1:0] node17238;
	wire [4-1:0] node17243;
	wire [4-1:0] node17244;
	wire [4-1:0] node17247;
	wire [4-1:0] node17248;
	wire [4-1:0] node17250;
	wire [4-1:0] node17253;
	wire [4-1:0] node17256;
	wire [4-1:0] node17257;
	wire [4-1:0] node17258;
	wire [4-1:0] node17259;
	wire [4-1:0] node17260;
	wire [4-1:0] node17264;
	wire [4-1:0] node17267;
	wire [4-1:0] node17268;
	wire [4-1:0] node17272;
	wire [4-1:0] node17274;
	wire [4-1:0] node17275;
	wire [4-1:0] node17276;
	wire [4-1:0] node17280;
	wire [4-1:0] node17283;
	wire [4-1:0] node17284;
	wire [4-1:0] node17285;
	wire [4-1:0] node17286;
	wire [4-1:0] node17289;
	wire [4-1:0] node17290;
	wire [4-1:0] node17292;
	wire [4-1:0] node17294;
	wire [4-1:0] node17298;
	wire [4-1:0] node17299;
	wire [4-1:0] node17300;
	wire [4-1:0] node17301;
	wire [4-1:0] node17303;
	wire [4-1:0] node17307;
	wire [4-1:0] node17308;
	wire [4-1:0] node17309;
	wire [4-1:0] node17312;
	wire [4-1:0] node17315;
	wire [4-1:0] node17318;
	wire [4-1:0] node17319;
	wire [4-1:0] node17320;
	wire [4-1:0] node17323;
	wire [4-1:0] node17326;
	wire [4-1:0] node17329;
	wire [4-1:0] node17330;
	wire [4-1:0] node17331;
	wire [4-1:0] node17333;
	wire [4-1:0] node17334;
	wire [4-1:0] node17335;
	wire [4-1:0] node17338;
	wire [4-1:0] node17342;
	wire [4-1:0] node17343;
	wire [4-1:0] node17346;
	wire [4-1:0] node17348;
	wire [4-1:0] node17351;
	wire [4-1:0] node17352;
	wire [4-1:0] node17354;
	wire [4-1:0] node17355;
	wire [4-1:0] node17358;
	wire [4-1:0] node17359;
	wire [4-1:0] node17363;
	wire [4-1:0] node17364;
	wire [4-1:0] node17365;
	wire [4-1:0] node17368;
	wire [4-1:0] node17369;
	wire [4-1:0] node17372;
	wire [4-1:0] node17375;
	wire [4-1:0] node17376;
	wire [4-1:0] node17378;
	wire [4-1:0] node17382;
	wire [4-1:0] node17383;
	wire [4-1:0] node17384;
	wire [4-1:0] node17385;
	wire [4-1:0] node17386;
	wire [4-1:0] node17387;
	wire [4-1:0] node17388;
	wire [4-1:0] node17389;
	wire [4-1:0] node17392;
	wire [4-1:0] node17395;
	wire [4-1:0] node17397;
	wire [4-1:0] node17400;
	wire [4-1:0] node17401;
	wire [4-1:0] node17405;
	wire [4-1:0] node17406;
	wire [4-1:0] node17409;
	wire [4-1:0] node17412;
	wire [4-1:0] node17413;
	wire [4-1:0] node17414;
	wire [4-1:0] node17417;
	wire [4-1:0] node17419;
	wire [4-1:0] node17421;
	wire [4-1:0] node17424;
	wire [4-1:0] node17425;
	wire [4-1:0] node17427;
	wire [4-1:0] node17428;
	wire [4-1:0] node17431;
	wire [4-1:0] node17434;
	wire [4-1:0] node17435;
	wire [4-1:0] node17438;
	wire [4-1:0] node17441;
	wire [4-1:0] node17442;
	wire [4-1:0] node17443;
	wire [4-1:0] node17444;
	wire [4-1:0] node17447;
	wire [4-1:0] node17450;
	wire [4-1:0] node17451;
	wire [4-1:0] node17453;
	wire [4-1:0] node17456;
	wire [4-1:0] node17457;
	wire [4-1:0] node17458;
	wire [4-1:0] node17461;
	wire [4-1:0] node17464;
	wire [4-1:0] node17466;
	wire [4-1:0] node17469;
	wire [4-1:0] node17470;
	wire [4-1:0] node17471;
	wire [4-1:0] node17474;
	wire [4-1:0] node17475;
	wire [4-1:0] node17477;
	wire [4-1:0] node17481;
	wire [4-1:0] node17482;
	wire [4-1:0] node17484;
	wire [4-1:0] node17485;
	wire [4-1:0] node17488;
	wire [4-1:0] node17491;
	wire [4-1:0] node17492;
	wire [4-1:0] node17493;
	wire [4-1:0] node17498;
	wire [4-1:0] node17499;
	wire [4-1:0] node17500;
	wire [4-1:0] node17501;
	wire [4-1:0] node17502;
	wire [4-1:0] node17503;
	wire [4-1:0] node17504;
	wire [4-1:0] node17507;
	wire [4-1:0] node17510;
	wire [4-1:0] node17512;
	wire [4-1:0] node17516;
	wire [4-1:0] node17518;
	wire [4-1:0] node17519;
	wire [4-1:0] node17522;
	wire [4-1:0] node17525;
	wire [4-1:0] node17526;
	wire [4-1:0] node17527;
	wire [4-1:0] node17528;
	wire [4-1:0] node17529;
	wire [4-1:0] node17533;
	wire [4-1:0] node17534;
	wire [4-1:0] node17537;
	wire [4-1:0] node17540;
	wire [4-1:0] node17541;
	wire [4-1:0] node17542;
	wire [4-1:0] node17546;
	wire [4-1:0] node17547;
	wire [4-1:0] node17551;
	wire [4-1:0] node17552;
	wire [4-1:0] node17553;
	wire [4-1:0] node17554;
	wire [4-1:0] node17557;
	wire [4-1:0] node17561;
	wire [4-1:0] node17563;
	wire [4-1:0] node17564;
	wire [4-1:0] node17567;
	wire [4-1:0] node17570;
	wire [4-1:0] node17571;
	wire [4-1:0] node17572;
	wire [4-1:0] node17573;
	wire [4-1:0] node17576;
	wire [4-1:0] node17578;
	wire [4-1:0] node17581;
	wire [4-1:0] node17582;
	wire [4-1:0] node17583;
	wire [4-1:0] node17584;
	wire [4-1:0] node17588;
	wire [4-1:0] node17590;
	wire [4-1:0] node17593;
	wire [4-1:0] node17596;
	wire [4-1:0] node17597;
	wire [4-1:0] node17599;
	wire [4-1:0] node17602;
	wire [4-1:0] node17605;
	wire [4-1:0] node17606;
	wire [4-1:0] node17607;
	wire [4-1:0] node17608;
	wire [4-1:0] node17609;
	wire [4-1:0] node17610;
	wire [4-1:0] node17611;
	wire [4-1:0] node17614;
	wire [4-1:0] node17615;
	wire [4-1:0] node17616;
	wire [4-1:0] node17621;
	wire [4-1:0] node17622;
	wire [4-1:0] node17624;
	wire [4-1:0] node17627;
	wire [4-1:0] node17628;
	wire [4-1:0] node17632;
	wire [4-1:0] node17633;
	wire [4-1:0] node17634;
	wire [4-1:0] node17635;
	wire [4-1:0] node17636;
	wire [4-1:0] node17639;
	wire [4-1:0] node17642;
	wire [4-1:0] node17643;
	wire [4-1:0] node17648;
	wire [4-1:0] node17649;
	wire [4-1:0] node17651;
	wire [4-1:0] node17652;
	wire [4-1:0] node17655;
	wire [4-1:0] node17658;
	wire [4-1:0] node17661;
	wire [4-1:0] node17662;
	wire [4-1:0] node17663;
	wire [4-1:0] node17665;
	wire [4-1:0] node17666;
	wire [4-1:0] node17669;
	wire [4-1:0] node17672;
	wire [4-1:0] node17674;
	wire [4-1:0] node17675;
	wire [4-1:0] node17677;
	wire [4-1:0] node17680;
	wire [4-1:0] node17683;
	wire [4-1:0] node17684;
	wire [4-1:0] node17685;
	wire [4-1:0] node17688;
	wire [4-1:0] node17691;
	wire [4-1:0] node17692;
	wire [4-1:0] node17694;
	wire [4-1:0] node17697;
	wire [4-1:0] node17698;
	wire [4-1:0] node17699;
	wire [4-1:0] node17703;
	wire [4-1:0] node17706;
	wire [4-1:0] node17707;
	wire [4-1:0] node17708;
	wire [4-1:0] node17709;
	wire [4-1:0] node17710;
	wire [4-1:0] node17711;
	wire [4-1:0] node17715;
	wire [4-1:0] node17717;
	wire [4-1:0] node17720;
	wire [4-1:0] node17722;
	wire [4-1:0] node17723;
	wire [4-1:0] node17727;
	wire [4-1:0] node17728;
	wire [4-1:0] node17729;
	wire [4-1:0] node17730;
	wire [4-1:0] node17732;
	wire [4-1:0] node17736;
	wire [4-1:0] node17737;
	wire [4-1:0] node17741;
	wire [4-1:0] node17742;
	wire [4-1:0] node17745;
	wire [4-1:0] node17748;
	wire [4-1:0] node17749;
	wire [4-1:0] node17750;
	wire [4-1:0] node17751;
	wire [4-1:0] node17753;
	wire [4-1:0] node17756;
	wire [4-1:0] node17758;
	wire [4-1:0] node17761;
	wire [4-1:0] node17762;
	wire [4-1:0] node17763;
	wire [4-1:0] node17766;
	wire [4-1:0] node17770;
	wire [4-1:0] node17771;
	wire [4-1:0] node17772;
	wire [4-1:0] node17775;
	wire [4-1:0] node17777;
	wire [4-1:0] node17780;
	wire [4-1:0] node17781;
	wire [4-1:0] node17784;
	wire [4-1:0] node17787;
	wire [4-1:0] node17788;
	wire [4-1:0] node17789;
	wire [4-1:0] node17790;
	wire [4-1:0] node17791;
	wire [4-1:0] node17792;
	wire [4-1:0] node17794;
	wire [4-1:0] node17796;
	wire [4-1:0] node17799;
	wire [4-1:0] node17800;
	wire [4-1:0] node17804;
	wire [4-1:0] node17805;
	wire [4-1:0] node17806;
	wire [4-1:0] node17810;
	wire [4-1:0] node17811;
	wire [4-1:0] node17813;
	wire [4-1:0] node17817;
	wire [4-1:0] node17818;
	wire [4-1:0] node17819;
	wire [4-1:0] node17820;
	wire [4-1:0] node17824;
	wire [4-1:0] node17826;
	wire [4-1:0] node17829;
	wire [4-1:0] node17830;
	wire [4-1:0] node17833;
	wire [4-1:0] node17836;
	wire [4-1:0] node17837;
	wire [4-1:0] node17838;
	wire [4-1:0] node17839;
	wire [4-1:0] node17840;
	wire [4-1:0] node17842;
	wire [4-1:0] node17846;
	wire [4-1:0] node17847;
	wire [4-1:0] node17848;
	wire [4-1:0] node17852;
	wire [4-1:0] node17854;
	wire [4-1:0] node17857;
	wire [4-1:0] node17858;
	wire [4-1:0] node17860;
	wire [4-1:0] node17863;
	wire [4-1:0] node17865;
	wire [4-1:0] node17868;
	wire [4-1:0] node17869;
	wire [4-1:0] node17870;
	wire [4-1:0] node17872;
	wire [4-1:0] node17873;
	wire [4-1:0] node17878;
	wire [4-1:0] node17879;
	wire [4-1:0] node17881;
	wire [4-1:0] node17884;
	wire [4-1:0] node17886;
	wire [4-1:0] node17889;
	wire [4-1:0] node17890;
	wire [4-1:0] node17891;
	wire [4-1:0] node17892;
	wire [4-1:0] node17894;
	wire [4-1:0] node17895;
	wire [4-1:0] node17896;
	wire [4-1:0] node17899;
	wire [4-1:0] node17903;
	wire [4-1:0] node17906;
	wire [4-1:0] node17907;
	wire [4-1:0] node17908;
	wire [4-1:0] node17909;
	wire [4-1:0] node17910;
	wire [4-1:0] node17914;
	wire [4-1:0] node17918;
	wire [4-1:0] node17920;
	wire [4-1:0] node17923;
	wire [4-1:0] node17924;
	wire [4-1:0] node17925;
	wire [4-1:0] node17926;
	wire [4-1:0] node17928;
	wire [4-1:0] node17931;
	wire [4-1:0] node17934;
	wire [4-1:0] node17935;
	wire [4-1:0] node17937;
	wire [4-1:0] node17941;
	wire [4-1:0] node17942;
	wire [4-1:0] node17943;
	wire [4-1:0] node17945;
	wire [4-1:0] node17948;
	wire [4-1:0] node17951;
	wire [4-1:0] node17952;
	wire [4-1:0] node17953;
	wire [4-1:0] node17954;
	wire [4-1:0] node17957;
	wire [4-1:0] node17962;
	wire [4-1:0] node17963;
	wire [4-1:0] node17964;
	wire [4-1:0] node17965;
	wire [4-1:0] node17966;
	wire [4-1:0] node17967;
	wire [4-1:0] node17968;
	wire [4-1:0] node17970;
	wire [4-1:0] node17973;
	wire [4-1:0] node17974;
	wire [4-1:0] node17976;
	wire [4-1:0] node17979;
	wire [4-1:0] node17980;
	wire [4-1:0] node17981;
	wire [4-1:0] node17984;
	wire [4-1:0] node17987;
	wire [4-1:0] node17988;
	wire [4-1:0] node17992;
	wire [4-1:0] node17993;
	wire [4-1:0] node17994;
	wire [4-1:0] node17995;
	wire [4-1:0] node17999;
	wire [4-1:0] node18002;
	wire [4-1:0] node18004;
	wire [4-1:0] node18006;
	wire [4-1:0] node18008;
	wire [4-1:0] node18011;
	wire [4-1:0] node18012;
	wire [4-1:0] node18013;
	wire [4-1:0] node18014;
	wire [4-1:0] node18015;
	wire [4-1:0] node18019;
	wire [4-1:0] node18022;
	wire [4-1:0] node18023;
	wire [4-1:0] node18024;
	wire [4-1:0] node18026;
	wire [4-1:0] node18031;
	wire [4-1:0] node18032;
	wire [4-1:0] node18033;
	wire [4-1:0] node18034;
	wire [4-1:0] node18038;
	wire [4-1:0] node18039;
	wire [4-1:0] node18042;
	wire [4-1:0] node18045;
	wire [4-1:0] node18047;
	wire [4-1:0] node18049;
	wire [4-1:0] node18050;
	wire [4-1:0] node18053;
	wire [4-1:0] node18056;
	wire [4-1:0] node18057;
	wire [4-1:0] node18058;
	wire [4-1:0] node18059;
	wire [4-1:0] node18061;
	wire [4-1:0] node18063;
	wire [4-1:0] node18066;
	wire [4-1:0] node18067;
	wire [4-1:0] node18068;
	wire [4-1:0] node18072;
	wire [4-1:0] node18075;
	wire [4-1:0] node18076;
	wire [4-1:0] node18077;
	wire [4-1:0] node18079;
	wire [4-1:0] node18083;
	wire [4-1:0] node18084;
	wire [4-1:0] node18087;
	wire [4-1:0] node18090;
	wire [4-1:0] node18091;
	wire [4-1:0] node18092;
	wire [4-1:0] node18093;
	wire [4-1:0] node18096;
	wire [4-1:0] node18099;
	wire [4-1:0] node18100;
	wire [4-1:0] node18102;
	wire [4-1:0] node18103;
	wire [4-1:0] node18107;
	wire [4-1:0] node18108;
	wire [4-1:0] node18109;
	wire [4-1:0] node18112;
	wire [4-1:0] node18116;
	wire [4-1:0] node18117;
	wire [4-1:0] node18118;
	wire [4-1:0] node18119;
	wire [4-1:0] node18122;
	wire [4-1:0] node18124;
	wire [4-1:0] node18127;
	wire [4-1:0] node18130;
	wire [4-1:0] node18131;
	wire [4-1:0] node18134;
	wire [4-1:0] node18135;
	wire [4-1:0] node18137;
	wire [4-1:0] node18141;
	wire [4-1:0] node18142;
	wire [4-1:0] node18143;
	wire [4-1:0] node18144;
	wire [4-1:0] node18145;
	wire [4-1:0] node18146;
	wire [4-1:0] node18147;
	wire [4-1:0] node18150;
	wire [4-1:0] node18153;
	wire [4-1:0] node18156;
	wire [4-1:0] node18157;
	wire [4-1:0] node18158;
	wire [4-1:0] node18162;
	wire [4-1:0] node18164;
	wire [4-1:0] node18167;
	wire [4-1:0] node18168;
	wire [4-1:0] node18169;
	wire [4-1:0] node18173;
	wire [4-1:0] node18175;
	wire [4-1:0] node18176;
	wire [4-1:0] node18177;
	wire [4-1:0] node18180;
	wire [4-1:0] node18183;
	wire [4-1:0] node18184;
	wire [4-1:0] node18188;
	wire [4-1:0] node18189;
	wire [4-1:0] node18190;
	wire [4-1:0] node18191;
	wire [4-1:0] node18193;
	wire [4-1:0] node18196;
	wire [4-1:0] node18198;
	wire [4-1:0] node18201;
	wire [4-1:0] node18202;
	wire [4-1:0] node18203;
	wire [4-1:0] node18204;
	wire [4-1:0] node18207;
	wire [4-1:0] node18211;
	wire [4-1:0] node18212;
	wire [4-1:0] node18214;
	wire [4-1:0] node18217;
	wire [4-1:0] node18219;
	wire [4-1:0] node18222;
	wire [4-1:0] node18223;
	wire [4-1:0] node18224;
	wire [4-1:0] node18225;
	wire [4-1:0] node18228;
	wire [4-1:0] node18232;
	wire [4-1:0] node18233;
	wire [4-1:0] node18234;
	wire [4-1:0] node18237;
	wire [4-1:0] node18239;
	wire [4-1:0] node18242;
	wire [4-1:0] node18244;
	wire [4-1:0] node18247;
	wire [4-1:0] node18248;
	wire [4-1:0] node18249;
	wire [4-1:0] node18250;
	wire [4-1:0] node18251;
	wire [4-1:0] node18253;
	wire [4-1:0] node18256;
	wire [4-1:0] node18258;
	wire [4-1:0] node18261;
	wire [4-1:0] node18263;
	wire [4-1:0] node18264;
	wire [4-1:0] node18265;
	wire [4-1:0] node18268;
	wire [4-1:0] node18271;
	wire [4-1:0] node18273;
	wire [4-1:0] node18276;
	wire [4-1:0] node18277;
	wire [4-1:0] node18278;
	wire [4-1:0] node18279;
	wire [4-1:0] node18282;
	wire [4-1:0] node18285;
	wire [4-1:0] node18288;
	wire [4-1:0] node18289;
	wire [4-1:0] node18290;
	wire [4-1:0] node18292;
	wire [4-1:0] node18295;
	wire [4-1:0] node18297;
	wire [4-1:0] node18300;
	wire [4-1:0] node18301;
	wire [4-1:0] node18304;
	wire [4-1:0] node18307;
	wire [4-1:0] node18308;
	wire [4-1:0] node18309;
	wire [4-1:0] node18310;
	wire [4-1:0] node18313;
	wire [4-1:0] node18316;
	wire [4-1:0] node18317;
	wire [4-1:0] node18320;
	wire [4-1:0] node18323;
	wire [4-1:0] node18324;
	wire [4-1:0] node18325;
	wire [4-1:0] node18328;
	wire [4-1:0] node18331;
	wire [4-1:0] node18332;
	wire [4-1:0] node18335;
	wire [4-1:0] node18338;
	wire [4-1:0] node18339;
	wire [4-1:0] node18340;
	wire [4-1:0] node18341;
	wire [4-1:0] node18342;
	wire [4-1:0] node18343;
	wire [4-1:0] node18344;
	wire [4-1:0] node18345;
	wire [4-1:0] node18347;
	wire [4-1:0] node18350;
	wire [4-1:0] node18351;
	wire [4-1:0] node18355;
	wire [4-1:0] node18357;
	wire [4-1:0] node18358;
	wire [4-1:0] node18361;
	wire [4-1:0] node18364;
	wire [4-1:0] node18367;
	wire [4-1:0] node18368;
	wire [4-1:0] node18369;
	wire [4-1:0] node18371;
	wire [4-1:0] node18375;
	wire [4-1:0] node18376;
	wire [4-1:0] node18378;
	wire [4-1:0] node18381;
	wire [4-1:0] node18384;
	wire [4-1:0] node18385;
	wire [4-1:0] node18386;
	wire [4-1:0] node18388;
	wire [4-1:0] node18389;
	wire [4-1:0] node18390;
	wire [4-1:0] node18393;
	wire [4-1:0] node18396;
	wire [4-1:0] node18397;
	wire [4-1:0] node18401;
	wire [4-1:0] node18403;
	wire [4-1:0] node18404;
	wire [4-1:0] node18408;
	wire [4-1:0] node18409;
	wire [4-1:0] node18410;
	wire [4-1:0] node18411;
	wire [4-1:0] node18413;
	wire [4-1:0] node18416;
	wire [4-1:0] node18417;
	wire [4-1:0] node18422;
	wire [4-1:0] node18423;
	wire [4-1:0] node18424;
	wire [4-1:0] node18425;
	wire [4-1:0] node18429;
	wire [4-1:0] node18430;
	wire [4-1:0] node18435;
	wire [4-1:0] node18436;
	wire [4-1:0] node18437;
	wire [4-1:0] node18438;
	wire [4-1:0] node18439;
	wire [4-1:0] node18440;
	wire [4-1:0] node18445;
	wire [4-1:0] node18446;
	wire [4-1:0] node18447;
	wire [4-1:0] node18451;
	wire [4-1:0] node18452;
	wire [4-1:0] node18455;
	wire [4-1:0] node18458;
	wire [4-1:0] node18459;
	wire [4-1:0] node18460;
	wire [4-1:0] node18461;
	wire [4-1:0] node18464;
	wire [4-1:0] node18467;
	wire [4-1:0] node18470;
	wire [4-1:0] node18471;
	wire [4-1:0] node18473;
	wire [4-1:0] node18476;
	wire [4-1:0] node18479;
	wire [4-1:0] node18480;
	wire [4-1:0] node18481;
	wire [4-1:0] node18482;
	wire [4-1:0] node18484;
	wire [4-1:0] node18485;
	wire [4-1:0] node18489;
	wire [4-1:0] node18490;
	wire [4-1:0] node18492;
	wire [4-1:0] node18495;
	wire [4-1:0] node18498;
	wire [4-1:0] node18499;
	wire [4-1:0] node18500;
	wire [4-1:0] node18501;
	wire [4-1:0] node18505;
	wire [4-1:0] node18507;
	wire [4-1:0] node18510;
	wire [4-1:0] node18511;
	wire [4-1:0] node18514;
	wire [4-1:0] node18516;
	wire [4-1:0] node18519;
	wire [4-1:0] node18520;
	wire [4-1:0] node18521;
	wire [4-1:0] node18522;
	wire [4-1:0] node18525;
	wire [4-1:0] node18528;
	wire [4-1:0] node18530;
	wire [4-1:0] node18533;
	wire [4-1:0] node18535;
	wire [4-1:0] node18536;
	wire [4-1:0] node18539;
	wire [4-1:0] node18542;
	wire [4-1:0] node18543;
	wire [4-1:0] node18544;
	wire [4-1:0] node18545;
	wire [4-1:0] node18546;
	wire [4-1:0] node18547;
	wire [4-1:0] node18548;
	wire [4-1:0] node18550;
	wire [4-1:0] node18553;
	wire [4-1:0] node18556;
	wire [4-1:0] node18557;
	wire [4-1:0] node18560;
	wire [4-1:0] node18563;
	wire [4-1:0] node18564;
	wire [4-1:0] node18567;
	wire [4-1:0] node18568;
	wire [4-1:0] node18571;
	wire [4-1:0] node18574;
	wire [4-1:0] node18575;
	wire [4-1:0] node18576;
	wire [4-1:0] node18577;
	wire [4-1:0] node18578;
	wire [4-1:0] node18581;
	wire [4-1:0] node18586;
	wire [4-1:0] node18587;
	wire [4-1:0] node18588;
	wire [4-1:0] node18591;
	wire [4-1:0] node18594;
	wire [4-1:0] node18595;
	wire [4-1:0] node18597;
	wire [4-1:0] node18600;
	wire [4-1:0] node18601;
	wire [4-1:0] node18605;
	wire [4-1:0] node18606;
	wire [4-1:0] node18607;
	wire [4-1:0] node18608;
	wire [4-1:0] node18610;
	wire [4-1:0] node18613;
	wire [4-1:0] node18616;
	wire [4-1:0] node18618;
	wire [4-1:0] node18621;
	wire [4-1:0] node18622;
	wire [4-1:0] node18623;
	wire [4-1:0] node18624;
	wire [4-1:0] node18628;
	wire [4-1:0] node18629;
	wire [4-1:0] node18630;
	wire [4-1:0] node18633;
	wire [4-1:0] node18637;
	wire [4-1:0] node18639;
	wire [4-1:0] node18640;
	wire [4-1:0] node18641;
	wire [4-1:0] node18646;
	wire [4-1:0] node18647;
	wire [4-1:0] node18648;
	wire [4-1:0] node18649;
	wire [4-1:0] node18650;
	wire [4-1:0] node18651;
	wire [4-1:0] node18655;
	wire [4-1:0] node18656;
	wire [4-1:0] node18660;
	wire [4-1:0] node18661;
	wire [4-1:0] node18662;
	wire [4-1:0] node18664;
	wire [4-1:0] node18667;
	wire [4-1:0] node18670;
	wire [4-1:0] node18671;
	wire [4-1:0] node18675;
	wire [4-1:0] node18676;
	wire [4-1:0] node18677;
	wire [4-1:0] node18678;
	wire [4-1:0] node18681;
	wire [4-1:0] node18685;
	wire [4-1:0] node18686;
	wire [4-1:0] node18687;
	wire [4-1:0] node18688;
	wire [4-1:0] node18692;
	wire [4-1:0] node18694;
	wire [4-1:0] node18697;
	wire [4-1:0] node18698;
	wire [4-1:0] node18701;
	wire [4-1:0] node18704;
	wire [4-1:0] node18705;
	wire [4-1:0] node18706;
	wire [4-1:0] node18707;
	wire [4-1:0] node18710;
	wire [4-1:0] node18713;
	wire [4-1:0] node18714;
	wire [4-1:0] node18717;
	wire [4-1:0] node18720;
	wire [4-1:0] node18721;
	wire [4-1:0] node18722;
	wire [4-1:0] node18724;
	wire [4-1:0] node18727;
	wire [4-1:0] node18728;
	wire [4-1:0] node18732;
	wire [4-1:0] node18733;
	wire [4-1:0] node18734;
	wire [4-1:0] node18738;
	wire [4-1:0] node18740;
	wire [4-1:0] node18743;
	wire [4-1:0] node18744;
	wire [4-1:0] node18745;
	wire [4-1:0] node18746;
	wire [4-1:0] node18747;
	wire [4-1:0] node18748;
	wire [4-1:0] node18749;
	wire [4-1:0] node18750;
	wire [4-1:0] node18751;
	wire [4-1:0] node18752;
	wire [4-1:0] node18753;
	wire [4-1:0] node18754;
	wire [4-1:0] node18758;
	wire [4-1:0] node18759;
	wire [4-1:0] node18763;
	wire [4-1:0] node18764;
	wire [4-1:0] node18765;
	wire [4-1:0] node18767;
	wire [4-1:0] node18770;
	wire [4-1:0] node18772;
	wire [4-1:0] node18775;
	wire [4-1:0] node18777;
	wire [4-1:0] node18778;
	wire [4-1:0] node18782;
	wire [4-1:0] node18783;
	wire [4-1:0] node18784;
	wire [4-1:0] node18786;
	wire [4-1:0] node18789;
	wire [4-1:0] node18791;
	wire [4-1:0] node18793;
	wire [4-1:0] node18796;
	wire [4-1:0] node18797;
	wire [4-1:0] node18799;
	wire [4-1:0] node18801;
	wire [4-1:0] node18804;
	wire [4-1:0] node18805;
	wire [4-1:0] node18807;
	wire [4-1:0] node18811;
	wire [4-1:0] node18812;
	wire [4-1:0] node18813;
	wire [4-1:0] node18814;
	wire [4-1:0] node18817;
	wire [4-1:0] node18818;
	wire [4-1:0] node18821;
	wire [4-1:0] node18824;
	wire [4-1:0] node18826;
	wire [4-1:0] node18829;
	wire [4-1:0] node18830;
	wire [4-1:0] node18831;
	wire [4-1:0] node18834;
	wire [4-1:0] node18835;
	wire [4-1:0] node18836;
	wire [4-1:0] node18840;
	wire [4-1:0] node18842;
	wire [4-1:0] node18845;
	wire [4-1:0] node18847;
	wire [4-1:0] node18848;
	wire [4-1:0] node18851;
	wire [4-1:0] node18854;
	wire [4-1:0] node18855;
	wire [4-1:0] node18856;
	wire [4-1:0] node18857;
	wire [4-1:0] node18858;
	wire [4-1:0] node18859;
	wire [4-1:0] node18861;
	wire [4-1:0] node18864;
	wire [4-1:0] node18866;
	wire [4-1:0] node18869;
	wire [4-1:0] node18870;
	wire [4-1:0] node18874;
	wire [4-1:0] node18875;
	wire [4-1:0] node18877;
	wire [4-1:0] node18880;
	wire [4-1:0] node18882;
	wire [4-1:0] node18884;
	wire [4-1:0] node18887;
	wire [4-1:0] node18888;
	wire [4-1:0] node18889;
	wire [4-1:0] node18890;
	wire [4-1:0] node18891;
	wire [4-1:0] node18895;
	wire [4-1:0] node18897;
	wire [4-1:0] node18900;
	wire [4-1:0] node18903;
	wire [4-1:0] node18904;
	wire [4-1:0] node18906;
	wire [4-1:0] node18909;
	wire [4-1:0] node18911;
	wire [4-1:0] node18913;
	wire [4-1:0] node18916;
	wire [4-1:0] node18917;
	wire [4-1:0] node18918;
	wire [4-1:0] node18919;
	wire [4-1:0] node18920;
	wire [4-1:0] node18921;
	wire [4-1:0] node18924;
	wire [4-1:0] node18927;
	wire [4-1:0] node18929;
	wire [4-1:0] node18932;
	wire [4-1:0] node18933;
	wire [4-1:0] node18937;
	wire [4-1:0] node18938;
	wire [4-1:0] node18939;
	wire [4-1:0] node18943;
	wire [4-1:0] node18944;
	wire [4-1:0] node18945;
	wire [4-1:0] node18948;
	wire [4-1:0] node18951;
	wire [4-1:0] node18952;
	wire [4-1:0] node18956;
	wire [4-1:0] node18957;
	wire [4-1:0] node18959;
	wire [4-1:0] node18960;
	wire [4-1:0] node18961;
	wire [4-1:0] node18964;
	wire [4-1:0] node18968;
	wire [4-1:0] node18970;
	wire [4-1:0] node18971;
	wire [4-1:0] node18974;
	wire [4-1:0] node18977;
	wire [4-1:0] node18978;
	wire [4-1:0] node18979;
	wire [4-1:0] node18980;
	wire [4-1:0] node18981;
	wire [4-1:0] node18983;
	wire [4-1:0] node18984;
	wire [4-1:0] node18988;
	wire [4-1:0] node18989;
	wire [4-1:0] node18990;
	wire [4-1:0] node18995;
	wire [4-1:0] node18996;
	wire [4-1:0] node18997;
	wire [4-1:0] node18998;
	wire [4-1:0] node18999;
	wire [4-1:0] node19004;
	wire [4-1:0] node19005;
	wire [4-1:0] node19006;
	wire [4-1:0] node19011;
	wire [4-1:0] node19012;
	wire [4-1:0] node19013;
	wire [4-1:0] node19016;
	wire [4-1:0] node19019;
	wire [4-1:0] node19021;
	wire [4-1:0] node19024;
	wire [4-1:0] node19025;
	wire [4-1:0] node19026;
	wire [4-1:0] node19027;
	wire [4-1:0] node19030;
	wire [4-1:0] node19032;
	wire [4-1:0] node19035;
	wire [4-1:0] node19037;
	wire [4-1:0] node19038;
	wire [4-1:0] node19039;
	wire [4-1:0] node19042;
	wire [4-1:0] node19046;
	wire [4-1:0] node19047;
	wire [4-1:0] node19048;
	wire [4-1:0] node19050;
	wire [4-1:0] node19053;
	wire [4-1:0] node19054;
	wire [4-1:0] node19055;
	wire [4-1:0] node19060;
	wire [4-1:0] node19062;
	wire [4-1:0] node19063;
	wire [4-1:0] node19067;
	wire [4-1:0] node19068;
	wire [4-1:0] node19069;
	wire [4-1:0] node19070;
	wire [4-1:0] node19071;
	wire [4-1:0] node19072;
	wire [4-1:0] node19073;
	wire [4-1:0] node19076;
	wire [4-1:0] node19080;
	wire [4-1:0] node19081;
	wire [4-1:0] node19085;
	wire [4-1:0] node19086;
	wire [4-1:0] node19087;
	wire [4-1:0] node19088;
	wire [4-1:0] node19092;
	wire [4-1:0] node19093;
	wire [4-1:0] node19097;
	wire [4-1:0] node19098;
	wire [4-1:0] node19101;
	wire [4-1:0] node19104;
	wire [4-1:0] node19105;
	wire [4-1:0] node19106;
	wire [4-1:0] node19110;
	wire [4-1:0] node19111;
	wire [4-1:0] node19112;
	wire [4-1:0] node19116;
	wire [4-1:0] node19119;
	wire [4-1:0] node19120;
	wire [4-1:0] node19121;
	wire [4-1:0] node19122;
	wire [4-1:0] node19123;
	wire [4-1:0] node19125;
	wire [4-1:0] node19129;
	wire [4-1:0] node19130;
	wire [4-1:0] node19133;
	wire [4-1:0] node19136;
	wire [4-1:0] node19137;
	wire [4-1:0] node19138;
	wire [4-1:0] node19142;
	wire [4-1:0] node19143;
	wire [4-1:0] node19147;
	wire [4-1:0] node19148;
	wire [4-1:0] node19149;
	wire [4-1:0] node19151;
	wire [4-1:0] node19154;
	wire [4-1:0] node19155;
	wire [4-1:0] node19158;
	wire [4-1:0] node19161;
	wire [4-1:0] node19162;
	wire [4-1:0] node19166;
	wire [4-1:0] node19167;
	wire [4-1:0] node19168;
	wire [4-1:0] node19169;
	wire [4-1:0] node19170;
	wire [4-1:0] node19171;
	wire [4-1:0] node19174;
	wire [4-1:0] node19175;
	wire [4-1:0] node19177;
	wire [4-1:0] node19181;
	wire [4-1:0] node19182;
	wire [4-1:0] node19183;
	wire [4-1:0] node19185;
	wire [4-1:0] node19186;
	wire [4-1:0] node19189;
	wire [4-1:0] node19192;
	wire [4-1:0] node19193;
	wire [4-1:0] node19196;
	wire [4-1:0] node19198;
	wire [4-1:0] node19201;
	wire [4-1:0] node19202;
	wire [4-1:0] node19205;
	wire [4-1:0] node19206;
	wire [4-1:0] node19209;
	wire [4-1:0] node19212;
	wire [4-1:0] node19213;
	wire [4-1:0] node19214;
	wire [4-1:0] node19215;
	wire [4-1:0] node19219;
	wire [4-1:0] node19220;
	wire [4-1:0] node19221;
	wire [4-1:0] node19225;
	wire [4-1:0] node19226;
	wire [4-1:0] node19229;
	wire [4-1:0] node19232;
	wire [4-1:0] node19233;
	wire [4-1:0] node19234;
	wire [4-1:0] node19235;
	wire [4-1:0] node19236;
	wire [4-1:0] node19241;
	wire [4-1:0] node19242;
	wire [4-1:0] node19245;
	wire [4-1:0] node19247;
	wire [4-1:0] node19250;
	wire [4-1:0] node19251;
	wire [4-1:0] node19252;
	wire [4-1:0] node19255;
	wire [4-1:0] node19258;
	wire [4-1:0] node19261;
	wire [4-1:0] node19262;
	wire [4-1:0] node19263;
	wire [4-1:0] node19264;
	wire [4-1:0] node19267;
	wire [4-1:0] node19268;
	wire [4-1:0] node19270;
	wire [4-1:0] node19273;
	wire [4-1:0] node19275;
	wire [4-1:0] node19278;
	wire [4-1:0] node19279;
	wire [4-1:0] node19280;
	wire [4-1:0] node19281;
	wire [4-1:0] node19282;
	wire [4-1:0] node19285;
	wire [4-1:0] node19289;
	wire [4-1:0] node19290;
	wire [4-1:0] node19291;
	wire [4-1:0] node19296;
	wire [4-1:0] node19298;
	wire [4-1:0] node19299;
	wire [4-1:0] node19302;
	wire [4-1:0] node19305;
	wire [4-1:0] node19306;
	wire [4-1:0] node19307;
	wire [4-1:0] node19308;
	wire [4-1:0] node19309;
	wire [4-1:0] node19310;
	wire [4-1:0] node19313;
	wire [4-1:0] node19317;
	wire [4-1:0] node19318;
	wire [4-1:0] node19320;
	wire [4-1:0] node19324;
	wire [4-1:0] node19325;
	wire [4-1:0] node19326;
	wire [4-1:0] node19328;
	wire [4-1:0] node19332;
	wire [4-1:0] node19333;
	wire [4-1:0] node19335;
	wire [4-1:0] node19339;
	wire [4-1:0] node19340;
	wire [4-1:0] node19341;
	wire [4-1:0] node19345;
	wire [4-1:0] node19346;
	wire [4-1:0] node19349;
	wire [4-1:0] node19351;
	wire [4-1:0] node19354;
	wire [4-1:0] node19355;
	wire [4-1:0] node19356;
	wire [4-1:0] node19357;
	wire [4-1:0] node19358;
	wire [4-1:0] node19359;
	wire [4-1:0] node19361;
	wire [4-1:0] node19363;
	wire [4-1:0] node19367;
	wire [4-1:0] node19368;
	wire [4-1:0] node19369;
	wire [4-1:0] node19370;
	wire [4-1:0] node19376;
	wire [4-1:0] node19377;
	wire [4-1:0] node19378;
	wire [4-1:0] node19380;
	wire [4-1:0] node19381;
	wire [4-1:0] node19384;
	wire [4-1:0] node19388;
	wire [4-1:0] node19390;
	wire [4-1:0] node19391;
	wire [4-1:0] node19394;
	wire [4-1:0] node19397;
	wire [4-1:0] node19398;
	wire [4-1:0] node19399;
	wire [4-1:0] node19400;
	wire [4-1:0] node19401;
	wire [4-1:0] node19403;
	wire [4-1:0] node19407;
	wire [4-1:0] node19408;
	wire [4-1:0] node19412;
	wire [4-1:0] node19413;
	wire [4-1:0] node19414;
	wire [4-1:0] node19415;
	wire [4-1:0] node19419;
	wire [4-1:0] node19421;
	wire [4-1:0] node19424;
	wire [4-1:0] node19425;
	wire [4-1:0] node19426;
	wire [4-1:0] node19429;
	wire [4-1:0] node19433;
	wire [4-1:0] node19434;
	wire [4-1:0] node19435;
	wire [4-1:0] node19438;
	wire [4-1:0] node19439;
	wire [4-1:0] node19440;
	wire [4-1:0] node19445;
	wire [4-1:0] node19446;
	wire [4-1:0] node19447;
	wire [4-1:0] node19450;
	wire [4-1:0] node19453;
	wire [4-1:0] node19455;
	wire [4-1:0] node19458;
	wire [4-1:0] node19459;
	wire [4-1:0] node19460;
	wire [4-1:0] node19461;
	wire [4-1:0] node19462;
	wire [4-1:0] node19466;
	wire [4-1:0] node19469;
	wire [4-1:0] node19470;
	wire [4-1:0] node19471;
	wire [4-1:0] node19473;
	wire [4-1:0] node19475;
	wire [4-1:0] node19478;
	wire [4-1:0] node19479;
	wire [4-1:0] node19483;
	wire [4-1:0] node19484;
	wire [4-1:0] node19487;
	wire [4-1:0] node19488;
	wire [4-1:0] node19489;
	wire [4-1:0] node19493;
	wire [4-1:0] node19494;
	wire [4-1:0] node19498;
	wire [4-1:0] node19499;
	wire [4-1:0] node19500;
	wire [4-1:0] node19501;
	wire [4-1:0] node19502;
	wire [4-1:0] node19504;
	wire [4-1:0] node19509;
	wire [4-1:0] node19511;
	wire [4-1:0] node19513;
	wire [4-1:0] node19516;
	wire [4-1:0] node19517;
	wire [4-1:0] node19518;
	wire [4-1:0] node19519;
	wire [4-1:0] node19522;
	wire [4-1:0] node19525;
	wire [4-1:0] node19526;
	wire [4-1:0] node19530;
	wire [4-1:0] node19531;
	wire [4-1:0] node19532;
	wire [4-1:0] node19533;
	wire [4-1:0] node19538;
	wire [4-1:0] node19539;
	wire [4-1:0] node19540;
	wire [4-1:0] node19543;
	wire [4-1:0] node19547;
	wire [4-1:0] node19548;
	wire [4-1:0] node19549;
	wire [4-1:0] node19550;
	wire [4-1:0] node19551;
	wire [4-1:0] node19552;
	wire [4-1:0] node19553;
	wire [4-1:0] node19554;
	wire [4-1:0] node19555;
	wire [4-1:0] node19556;
	wire [4-1:0] node19559;
	wire [4-1:0] node19563;
	wire [4-1:0] node19565;
	wire [4-1:0] node19568;
	wire [4-1:0] node19569;
	wire [4-1:0] node19571;
	wire [4-1:0] node19574;
	wire [4-1:0] node19576;
	wire [4-1:0] node19577;
	wire [4-1:0] node19581;
	wire [4-1:0] node19582;
	wire [4-1:0] node19583;
	wire [4-1:0] node19584;
	wire [4-1:0] node19585;
	wire [4-1:0] node19588;
	wire [4-1:0] node19591;
	wire [4-1:0] node19592;
	wire [4-1:0] node19595;
	wire [4-1:0] node19598;
	wire [4-1:0] node19599;
	wire [4-1:0] node19602;
	wire [4-1:0] node19605;
	wire [4-1:0] node19606;
	wire [4-1:0] node19608;
	wire [4-1:0] node19611;
	wire [4-1:0] node19614;
	wire [4-1:0] node19615;
	wire [4-1:0] node19616;
	wire [4-1:0] node19617;
	wire [4-1:0] node19618;
	wire [4-1:0] node19619;
	wire [4-1:0] node19624;
	wire [4-1:0] node19625;
	wire [4-1:0] node19626;
	wire [4-1:0] node19631;
	wire [4-1:0] node19633;
	wire [4-1:0] node19635;
	wire [4-1:0] node19636;
	wire [4-1:0] node19639;
	wire [4-1:0] node19642;
	wire [4-1:0] node19643;
	wire [4-1:0] node19645;
	wire [4-1:0] node19646;
	wire [4-1:0] node19648;
	wire [4-1:0] node19652;
	wire [4-1:0] node19653;
	wire [4-1:0] node19655;
	wire [4-1:0] node19656;
	wire [4-1:0] node19659;
	wire [4-1:0] node19662;
	wire [4-1:0] node19663;
	wire [4-1:0] node19664;
	wire [4-1:0] node19667;
	wire [4-1:0] node19671;
	wire [4-1:0] node19672;
	wire [4-1:0] node19673;
	wire [4-1:0] node19674;
	wire [4-1:0] node19675;
	wire [4-1:0] node19677;
	wire [4-1:0] node19679;
	wire [4-1:0] node19683;
	wire [4-1:0] node19684;
	wire [4-1:0] node19685;
	wire [4-1:0] node19690;
	wire [4-1:0] node19691;
	wire [4-1:0] node19692;
	wire [4-1:0] node19693;
	wire [4-1:0] node19694;
	wire [4-1:0] node19697;
	wire [4-1:0] node19700;
	wire [4-1:0] node19701;
	wire [4-1:0] node19705;
	wire [4-1:0] node19706;
	wire [4-1:0] node19710;
	wire [4-1:0] node19712;
	wire [4-1:0] node19714;
	wire [4-1:0] node19715;
	wire [4-1:0] node19718;
	wire [4-1:0] node19721;
	wire [4-1:0] node19722;
	wire [4-1:0] node19723;
	wire [4-1:0] node19724;
	wire [4-1:0] node19725;
	wire [4-1:0] node19726;
	wire [4-1:0] node19729;
	wire [4-1:0] node19733;
	wire [4-1:0] node19734;
	wire [4-1:0] node19735;
	wire [4-1:0] node19740;
	wire [4-1:0] node19741;
	wire [4-1:0] node19744;
	wire [4-1:0] node19745;
	wire [4-1:0] node19746;
	wire [4-1:0] node19751;
	wire [4-1:0] node19752;
	wire [4-1:0] node19754;
	wire [4-1:0] node19755;
	wire [4-1:0] node19756;
	wire [4-1:0] node19759;
	wire [4-1:0] node19763;
	wire [4-1:0] node19764;
	wire [4-1:0] node19765;
	wire [4-1:0] node19767;
	wire [4-1:0] node19771;
	wire [4-1:0] node19774;
	wire [4-1:0] node19775;
	wire [4-1:0] node19776;
	wire [4-1:0] node19777;
	wire [4-1:0] node19778;
	wire [4-1:0] node19779;
	wire [4-1:0] node19780;
	wire [4-1:0] node19781;
	wire [4-1:0] node19786;
	wire [4-1:0] node19787;
	wire [4-1:0] node19788;
	wire [4-1:0] node19791;
	wire [4-1:0] node19794;
	wire [4-1:0] node19796;
	wire [4-1:0] node19799;
	wire [4-1:0] node19800;
	wire [4-1:0] node19801;
	wire [4-1:0] node19802;
	wire [4-1:0] node19807;
	wire [4-1:0] node19808;
	wire [4-1:0] node19811;
	wire [4-1:0] node19814;
	wire [4-1:0] node19815;
	wire [4-1:0] node19816;
	wire [4-1:0] node19817;
	wire [4-1:0] node19818;
	wire [4-1:0] node19823;
	wire [4-1:0] node19826;
	wire [4-1:0] node19827;
	wire [4-1:0] node19829;
	wire [4-1:0] node19831;
	wire [4-1:0] node19834;
	wire [4-1:0] node19835;
	wire [4-1:0] node19838;
	wire [4-1:0] node19839;
	wire [4-1:0] node19842;
	wire [4-1:0] node19845;
	wire [4-1:0] node19846;
	wire [4-1:0] node19847;
	wire [4-1:0] node19849;
	wire [4-1:0] node19850;
	wire [4-1:0] node19854;
	wire [4-1:0] node19855;
	wire [4-1:0] node19859;
	wire [4-1:0] node19860;
	wire [4-1:0] node19861;
	wire [4-1:0] node19862;
	wire [4-1:0] node19865;
	wire [4-1:0] node19868;
	wire [4-1:0] node19871;
	wire [4-1:0] node19872;
	wire [4-1:0] node19876;
	wire [4-1:0] node19877;
	wire [4-1:0] node19878;
	wire [4-1:0] node19879;
	wire [4-1:0] node19881;
	wire [4-1:0] node19883;
	wire [4-1:0] node19886;
	wire [4-1:0] node19887;
	wire [4-1:0] node19888;
	wire [4-1:0] node19892;
	wire [4-1:0] node19893;
	wire [4-1:0] node19897;
	wire [4-1:0] node19898;
	wire [4-1:0] node19899;
	wire [4-1:0] node19900;
	wire [4-1:0] node19902;
	wire [4-1:0] node19905;
	wire [4-1:0] node19906;
	wire [4-1:0] node19909;
	wire [4-1:0] node19912;
	wire [4-1:0] node19913;
	wire [4-1:0] node19916;
	wire [4-1:0] node19919;
	wire [4-1:0] node19920;
	wire [4-1:0] node19921;
	wire [4-1:0] node19924;
	wire [4-1:0] node19927;
	wire [4-1:0] node19929;
	wire [4-1:0] node19930;
	wire [4-1:0] node19934;
	wire [4-1:0] node19935;
	wire [4-1:0] node19936;
	wire [4-1:0] node19937;
	wire [4-1:0] node19938;
	wire [4-1:0] node19941;
	wire [4-1:0] node19944;
	wire [4-1:0] node19945;
	wire [4-1:0] node19948;
	wire [4-1:0] node19951;
	wire [4-1:0] node19952;
	wire [4-1:0] node19953;
	wire [4-1:0] node19954;
	wire [4-1:0] node19959;
	wire [4-1:0] node19960;
	wire [4-1:0] node19961;
	wire [4-1:0] node19965;
	wire [4-1:0] node19968;
	wire [4-1:0] node19969;
	wire [4-1:0] node19970;
	wire [4-1:0] node19971;
	wire [4-1:0] node19972;
	wire [4-1:0] node19977;
	wire [4-1:0] node19978;
	wire [4-1:0] node19980;
	wire [4-1:0] node19983;
	wire [4-1:0] node19986;
	wire [4-1:0] node19988;
	wire [4-1:0] node19991;
	wire [4-1:0] node19992;
	wire [4-1:0] node19993;
	wire [4-1:0] node19994;
	wire [4-1:0] node19995;
	wire [4-1:0] node19996;
	wire [4-1:0] node19997;
	wire [4-1:0] node19998;
	wire [4-1:0] node19999;
	wire [4-1:0] node20002;
	wire [4-1:0] node20005;
	wire [4-1:0] node20007;
	wire [4-1:0] node20010;
	wire [4-1:0] node20013;
	wire [4-1:0] node20014;
	wire [4-1:0] node20018;
	wire [4-1:0] node20019;
	wire [4-1:0] node20020;
	wire [4-1:0] node20021;
	wire [4-1:0] node20024;
	wire [4-1:0] node20027;
	wire [4-1:0] node20028;
	wire [4-1:0] node20029;
	wire [4-1:0] node20033;
	wire [4-1:0] node20036;
	wire [4-1:0] node20037;
	wire [4-1:0] node20038;
	wire [4-1:0] node20039;
	wire [4-1:0] node20044;
	wire [4-1:0] node20046;
	wire [4-1:0] node20049;
	wire [4-1:0] node20050;
	wire [4-1:0] node20051;
	wire [4-1:0] node20052;
	wire [4-1:0] node20054;
	wire [4-1:0] node20055;
	wire [4-1:0] node20058;
	wire [4-1:0] node20061;
	wire [4-1:0] node20062;
	wire [4-1:0] node20064;
	wire [4-1:0] node20068;
	wire [4-1:0] node20069;
	wire [4-1:0] node20070;
	wire [4-1:0] node20074;
	wire [4-1:0] node20076;
	wire [4-1:0] node20077;
	wire [4-1:0] node20080;
	wire [4-1:0] node20083;
	wire [4-1:0] node20084;
	wire [4-1:0] node20085;
	wire [4-1:0] node20086;
	wire [4-1:0] node20089;
	wire [4-1:0] node20092;
	wire [4-1:0] node20093;
	wire [4-1:0] node20096;
	wire [4-1:0] node20099;
	wire [4-1:0] node20100;
	wire [4-1:0] node20102;
	wire [4-1:0] node20105;
	wire [4-1:0] node20106;
	wire [4-1:0] node20109;
	wire [4-1:0] node20112;
	wire [4-1:0] node20113;
	wire [4-1:0] node20114;
	wire [4-1:0] node20115;
	wire [4-1:0] node20116;
	wire [4-1:0] node20117;
	wire [4-1:0] node20121;
	wire [4-1:0] node20122;
	wire [4-1:0] node20125;
	wire [4-1:0] node20128;
	wire [4-1:0] node20129;
	wire [4-1:0] node20131;
	wire [4-1:0] node20132;
	wire [4-1:0] node20135;
	wire [4-1:0] node20138;
	wire [4-1:0] node20139;
	wire [4-1:0] node20143;
	wire [4-1:0] node20144;
	wire [4-1:0] node20146;
	wire [4-1:0] node20148;
	wire [4-1:0] node20149;
	wire [4-1:0] node20152;
	wire [4-1:0] node20155;
	wire [4-1:0] node20156;
	wire [4-1:0] node20157;
	wire [4-1:0] node20158;
	wire [4-1:0] node20164;
	wire [4-1:0] node20165;
	wire [4-1:0] node20166;
	wire [4-1:0] node20167;
	wire [4-1:0] node20169;
	wire [4-1:0] node20172;
	wire [4-1:0] node20173;
	wire [4-1:0] node20174;
	wire [4-1:0] node20178;
	wire [4-1:0] node20179;
	wire [4-1:0] node20182;
	wire [4-1:0] node20185;
	wire [4-1:0] node20186;
	wire [4-1:0] node20188;
	wire [4-1:0] node20191;
	wire [4-1:0] node20192;
	wire [4-1:0] node20195;
	wire [4-1:0] node20198;
	wire [4-1:0] node20199;
	wire [4-1:0] node20201;
	wire [4-1:0] node20204;
	wire [4-1:0] node20205;
	wire [4-1:0] node20206;
	wire [4-1:0] node20209;
	wire [4-1:0] node20213;
	wire [4-1:0] node20214;
	wire [4-1:0] node20215;
	wire [4-1:0] node20216;
	wire [4-1:0] node20217;
	wire [4-1:0] node20218;
	wire [4-1:0] node20219;
	wire [4-1:0] node20222;
	wire [4-1:0] node20225;
	wire [4-1:0] node20226;
	wire [4-1:0] node20230;
	wire [4-1:0] node20232;
	wire [4-1:0] node20235;
	wire [4-1:0] node20236;
	wire [4-1:0] node20237;
	wire [4-1:0] node20239;
	wire [4-1:0] node20242;
	wire [4-1:0] node20243;
	wire [4-1:0] node20247;
	wire [4-1:0] node20248;
	wire [4-1:0] node20250;
	wire [4-1:0] node20253;
	wire [4-1:0] node20255;
	wire [4-1:0] node20258;
	wire [4-1:0] node20259;
	wire [4-1:0] node20260;
	wire [4-1:0] node20261;
	wire [4-1:0] node20262;
	wire [4-1:0] node20266;
	wire [4-1:0] node20267;
	wire [4-1:0] node20269;
	wire [4-1:0] node20272;
	wire [4-1:0] node20274;
	wire [4-1:0] node20277;
	wire [4-1:0] node20278;
	wire [4-1:0] node20280;
	wire [4-1:0] node20282;
	wire [4-1:0] node20286;
	wire [4-1:0] node20287;
	wire [4-1:0] node20289;
	wire [4-1:0] node20291;
	wire [4-1:0] node20292;
	wire [4-1:0] node20296;
	wire [4-1:0] node20298;
	wire [4-1:0] node20299;
	wire [4-1:0] node20300;
	wire [4-1:0] node20304;
	wire [4-1:0] node20305;
	wire [4-1:0] node20308;
	wire [4-1:0] node20311;
	wire [4-1:0] node20312;
	wire [4-1:0] node20313;
	wire [4-1:0] node20314;
	wire [4-1:0] node20315;
	wire [4-1:0] node20317;
	wire [4-1:0] node20320;
	wire [4-1:0] node20321;
	wire [4-1:0] node20322;
	wire [4-1:0] node20327;
	wire [4-1:0] node20330;
	wire [4-1:0] node20331;
	wire [4-1:0] node20332;
	wire [4-1:0] node20336;
	wire [4-1:0] node20337;
	wire [4-1:0] node20339;
	wire [4-1:0] node20342;
	wire [4-1:0] node20344;
	wire [4-1:0] node20347;
	wire [4-1:0] node20348;
	wire [4-1:0] node20349;
	wire [4-1:0] node20350;
	wire [4-1:0] node20351;
	wire [4-1:0] node20354;
	wire [4-1:0] node20357;
	wire [4-1:0] node20358;
	wire [4-1:0] node20362;
	wire [4-1:0] node20363;
	wire [4-1:0] node20364;
	wire [4-1:0] node20366;
	wire [4-1:0] node20369;
	wire [4-1:0] node20370;
	wire [4-1:0] node20373;
	wire [4-1:0] node20377;
	wire [4-1:0] node20378;
	wire [4-1:0] node20379;
	wire [4-1:0] node20383;
	wire [4-1:0] node20384;
	wire [4-1:0] node20387;
	wire [4-1:0] node20388;
	wire [4-1:0] node20392;
	wire [4-1:0] node20393;
	wire [4-1:0] node20394;
	wire [4-1:0] node20395;
	wire [4-1:0] node20396;
	wire [4-1:0] node20397;
	wire [4-1:0] node20398;
	wire [4-1:0] node20399;
	wire [4-1:0] node20400;
	wire [4-1:0] node20403;
	wire [4-1:0] node20404;
	wire [4-1:0] node20408;
	wire [4-1:0] node20409;
	wire [4-1:0] node20410;
	wire [4-1:0] node20414;
	wire [4-1:0] node20416;
	wire [4-1:0] node20417;
	wire [4-1:0] node20420;
	wire [4-1:0] node20423;
	wire [4-1:0] node20424;
	wire [4-1:0] node20427;
	wire [4-1:0] node20428;
	wire [4-1:0] node20430;
	wire [4-1:0] node20434;
	wire [4-1:0] node20435;
	wire [4-1:0] node20436;
	wire [4-1:0] node20437;
	wire [4-1:0] node20438;
	wire [4-1:0] node20441;
	wire [4-1:0] node20443;
	wire [4-1:0] node20446;
	wire [4-1:0] node20448;
	wire [4-1:0] node20450;
	wire [4-1:0] node20453;
	wire [4-1:0] node20455;
	wire [4-1:0] node20456;
	wire [4-1:0] node20457;
	wire [4-1:0] node20461;
	wire [4-1:0] node20463;
	wire [4-1:0] node20466;
	wire [4-1:0] node20467;
	wire [4-1:0] node20468;
	wire [4-1:0] node20472;
	wire [4-1:0] node20473;
	wire [4-1:0] node20474;
	wire [4-1:0] node20476;
	wire [4-1:0] node20480;
	wire [4-1:0] node20481;
	wire [4-1:0] node20482;
	wire [4-1:0] node20486;
	wire [4-1:0] node20487;
	wire [4-1:0] node20491;
	wire [4-1:0] node20492;
	wire [4-1:0] node20493;
	wire [4-1:0] node20494;
	wire [4-1:0] node20495;
	wire [4-1:0] node20496;
	wire [4-1:0] node20499;
	wire [4-1:0] node20501;
	wire [4-1:0] node20505;
	wire [4-1:0] node20506;
	wire [4-1:0] node20507;
	wire [4-1:0] node20508;
	wire [4-1:0] node20513;
	wire [4-1:0] node20514;
	wire [4-1:0] node20515;
	wire [4-1:0] node20520;
	wire [4-1:0] node20521;
	wire [4-1:0] node20522;
	wire [4-1:0] node20523;
	wire [4-1:0] node20526;
	wire [4-1:0] node20528;
	wire [4-1:0] node20531;
	wire [4-1:0] node20532;
	wire [4-1:0] node20536;
	wire [4-1:0] node20538;
	wire [4-1:0] node20539;
	wire [4-1:0] node20542;
	wire [4-1:0] node20545;
	wire [4-1:0] node20546;
	wire [4-1:0] node20547;
	wire [4-1:0] node20548;
	wire [4-1:0] node20551;
	wire [4-1:0] node20554;
	wire [4-1:0] node20555;
	wire [4-1:0] node20557;
	wire [4-1:0] node20558;
	wire [4-1:0] node20562;
	wire [4-1:0] node20563;
	wire [4-1:0] node20566;
	wire [4-1:0] node20567;
	wire [4-1:0] node20570;
	wire [4-1:0] node20573;
	wire [4-1:0] node20574;
	wire [4-1:0] node20575;
	wire [4-1:0] node20576;
	wire [4-1:0] node20580;
	wire [4-1:0] node20583;
	wire [4-1:0] node20584;
	wire [4-1:0] node20587;
	wire [4-1:0] node20588;
	wire [4-1:0] node20592;
	wire [4-1:0] node20593;
	wire [4-1:0] node20594;
	wire [4-1:0] node20595;
	wire [4-1:0] node20596;
	wire [4-1:0] node20599;
	wire [4-1:0] node20600;
	wire [4-1:0] node20602;
	wire [4-1:0] node20605;
	wire [4-1:0] node20608;
	wire [4-1:0] node20609;
	wire [4-1:0] node20611;
	wire [4-1:0] node20612;
	wire [4-1:0] node20614;
	wire [4-1:0] node20617;
	wire [4-1:0] node20620;
	wire [4-1:0] node20621;
	wire [4-1:0] node20622;
	wire [4-1:0] node20625;
	wire [4-1:0] node20628;
	wire [4-1:0] node20631;
	wire [4-1:0] node20632;
	wire [4-1:0] node20633;
	wire [4-1:0] node20634;
	wire [4-1:0] node20635;
	wire [4-1:0] node20639;
	wire [4-1:0] node20640;
	wire [4-1:0] node20644;
	wire [4-1:0] node20645;
	wire [4-1:0] node20648;
	wire [4-1:0] node20651;
	wire [4-1:0] node20652;
	wire [4-1:0] node20653;
	wire [4-1:0] node20654;
	wire [4-1:0] node20655;
	wire [4-1:0] node20659;
	wire [4-1:0] node20660;
	wire [4-1:0] node20664;
	wire [4-1:0] node20667;
	wire [4-1:0] node20668;
	wire [4-1:0] node20670;
	wire [4-1:0] node20673;
	wire [4-1:0] node20674;
	wire [4-1:0] node20677;
	wire [4-1:0] node20678;
	wire [4-1:0] node20682;
	wire [4-1:0] node20683;
	wire [4-1:0] node20684;
	wire [4-1:0] node20685;
	wire [4-1:0] node20686;
	wire [4-1:0] node20687;
	wire [4-1:0] node20692;
	wire [4-1:0] node20693;
	wire [4-1:0] node20696;
	wire [4-1:0] node20699;
	wire [4-1:0] node20700;
	wire [4-1:0] node20701;
	wire [4-1:0] node20704;
	wire [4-1:0] node20707;
	wire [4-1:0] node20709;
	wire [4-1:0] node20710;
	wire [4-1:0] node20714;
	wire [4-1:0] node20715;
	wire [4-1:0] node20716;
	wire [4-1:0] node20717;
	wire [4-1:0] node20719;
	wire [4-1:0] node20722;
	wire [4-1:0] node20723;
	wire [4-1:0] node20727;
	wire [4-1:0] node20728;
	wire [4-1:0] node20729;
	wire [4-1:0] node20731;
	wire [4-1:0] node20735;
	wire [4-1:0] node20738;
	wire [4-1:0] node20739;
	wire [4-1:0] node20740;
	wire [4-1:0] node20741;
	wire [4-1:0] node20742;
	wire [4-1:0] node20746;
	wire [4-1:0] node20749;
	wire [4-1:0] node20752;
	wire [4-1:0] node20753;
	wire [4-1:0] node20754;
	wire [4-1:0] node20758;
	wire [4-1:0] node20759;
	wire [4-1:0] node20763;
	wire [4-1:0] node20764;
	wire [4-1:0] node20765;
	wire [4-1:0] node20766;
	wire [4-1:0] node20767;
	wire [4-1:0] node20768;
	wire [4-1:0] node20769;
	wire [4-1:0] node20770;
	wire [4-1:0] node20773;
	wire [4-1:0] node20776;
	wire [4-1:0] node20778;
	wire [4-1:0] node20781;
	wire [4-1:0] node20782;
	wire [4-1:0] node20786;
	wire [4-1:0] node20787;
	wire [4-1:0] node20788;
	wire [4-1:0] node20790;
	wire [4-1:0] node20794;
	wire [4-1:0] node20795;
	wire [4-1:0] node20799;
	wire [4-1:0] node20800;
	wire [4-1:0] node20801;
	wire [4-1:0] node20803;
	wire [4-1:0] node20804;
	wire [4-1:0] node20808;
	wire [4-1:0] node20809;
	wire [4-1:0] node20812;
	wire [4-1:0] node20813;
	wire [4-1:0] node20817;
	wire [4-1:0] node20818;
	wire [4-1:0] node20819;
	wire [4-1:0] node20820;
	wire [4-1:0] node20825;
	wire [4-1:0] node20826;
	wire [4-1:0] node20828;
	wire [4-1:0] node20831;
	wire [4-1:0] node20834;
	wire [4-1:0] node20835;
	wire [4-1:0] node20836;
	wire [4-1:0] node20837;
	wire [4-1:0] node20838;
	wire [4-1:0] node20839;
	wire [4-1:0] node20842;
	wire [4-1:0] node20844;
	wire [4-1:0] node20847;
	wire [4-1:0] node20848;
	wire [4-1:0] node20852;
	wire [4-1:0] node20854;
	wire [4-1:0] node20857;
	wire [4-1:0] node20858;
	wire [4-1:0] node20859;
	wire [4-1:0] node20860;
	wire [4-1:0] node20863;
	wire [4-1:0] node20866;
	wire [4-1:0] node20869;
	wire [4-1:0] node20871;
	wire [4-1:0] node20874;
	wire [4-1:0] node20875;
	wire [4-1:0] node20876;
	wire [4-1:0] node20877;
	wire [4-1:0] node20879;
	wire [4-1:0] node20882;
	wire [4-1:0] node20885;
	wire [4-1:0] node20886;
	wire [4-1:0] node20888;
	wire [4-1:0] node20891;
	wire [4-1:0] node20893;
	wire [4-1:0] node20896;
	wire [4-1:0] node20897;
	wire [4-1:0] node20898;
	wire [4-1:0] node20900;
	wire [4-1:0] node20903;
	wire [4-1:0] node20905;
	wire [4-1:0] node20908;
	wire [4-1:0] node20909;
	wire [4-1:0] node20911;
	wire [4-1:0] node20914;
	wire [4-1:0] node20915;
	wire [4-1:0] node20918;
	wire [4-1:0] node20921;
	wire [4-1:0] node20922;
	wire [4-1:0] node20923;
	wire [4-1:0] node20924;
	wire [4-1:0] node20925;
	wire [4-1:0] node20926;
	wire [4-1:0] node20929;
	wire [4-1:0] node20930;
	wire [4-1:0] node20935;
	wire [4-1:0] node20936;
	wire [4-1:0] node20937;
	wire [4-1:0] node20938;
	wire [4-1:0] node20942;
	wire [4-1:0] node20944;
	wire [4-1:0] node20947;
	wire [4-1:0] node20948;
	wire [4-1:0] node20949;
	wire [4-1:0] node20953;
	wire [4-1:0] node20956;
	wire [4-1:0] node20957;
	wire [4-1:0] node20958;
	wire [4-1:0] node20959;
	wire [4-1:0] node20961;
	wire [4-1:0] node20964;
	wire [4-1:0] node20966;
	wire [4-1:0] node20969;
	wire [4-1:0] node20970;
	wire [4-1:0] node20971;
	wire [4-1:0] node20975;
	wire [4-1:0] node20976;
	wire [4-1:0] node20980;
	wire [4-1:0] node20981;
	wire [4-1:0] node20982;
	wire [4-1:0] node20986;
	wire [4-1:0] node20987;
	wire [4-1:0] node20991;
	wire [4-1:0] node20992;
	wire [4-1:0] node20993;
	wire [4-1:0] node20994;
	wire [4-1:0] node20997;
	wire [4-1:0] node20999;
	wire [4-1:0] node21000;
	wire [4-1:0] node21001;
	wire [4-1:0] node21005;
	wire [4-1:0] node21008;
	wire [4-1:0] node21009;
	wire [4-1:0] node21011;
	wire [4-1:0] node21012;
	wire [4-1:0] node21013;
	wire [4-1:0] node21017;
	wire [4-1:0] node21020;
	wire [4-1:0] node21022;
	wire [4-1:0] node21024;
	wire [4-1:0] node21025;
	wire [4-1:0] node21029;
	wire [4-1:0] node21030;
	wire [4-1:0] node21031;
	wire [4-1:0] node21032;
	wire [4-1:0] node21034;
	wire [4-1:0] node21038;
	wire [4-1:0] node21039;
	wire [4-1:0] node21040;
	wire [4-1:0] node21044;
	wire [4-1:0] node21047;
	wire [4-1:0] node21048;
	wire [4-1:0] node21050;
	wire [4-1:0] node21051;
	wire [4-1:0] node21054;
	wire [4-1:0] node21055;
	wire [4-1:0] node21059;
	wire [4-1:0] node21060;
	wire [4-1:0] node21062;
	wire [4-1:0] node21065;
	wire [4-1:0] node21067;
	wire [4-1:0] node21070;
	wire [4-1:0] node21071;
	wire [4-1:0] node21072;
	wire [4-1:0] node21073;
	wire [4-1:0] node21074;
	wire [4-1:0] node21075;
	wire [4-1:0] node21076;
	wire [4-1:0] node21077;
	wire [4-1:0] node21079;
	wire [4-1:0] node21082;
	wire [4-1:0] node21084;
	wire [4-1:0] node21086;
	wire [4-1:0] node21089;
	wire [4-1:0] node21090;
	wire [4-1:0] node21091;
	wire [4-1:0] node21096;
	wire [4-1:0] node21097;
	wire [4-1:0] node21098;
	wire [4-1:0] node21102;
	wire [4-1:0] node21103;
	wire [4-1:0] node21105;
	wire [4-1:0] node21106;
	wire [4-1:0] node21109;
	wire [4-1:0] node21113;
	wire [4-1:0] node21114;
	wire [4-1:0] node21115;
	wire [4-1:0] node21116;
	wire [4-1:0] node21118;
	wire [4-1:0] node21120;
	wire [4-1:0] node21124;
	wire [4-1:0] node21125;
	wire [4-1:0] node21127;
	wire [4-1:0] node21130;
	wire [4-1:0] node21132;
	wire [4-1:0] node21135;
	wire [4-1:0] node21136;
	wire [4-1:0] node21137;
	wire [4-1:0] node21138;
	wire [4-1:0] node21140;
	wire [4-1:0] node21144;
	wire [4-1:0] node21145;
	wire [4-1:0] node21147;
	wire [4-1:0] node21151;
	wire [4-1:0] node21152;
	wire [4-1:0] node21154;
	wire [4-1:0] node21157;
	wire [4-1:0] node21160;
	wire [4-1:0] node21161;
	wire [4-1:0] node21162;
	wire [4-1:0] node21163;
	wire [4-1:0] node21164;
	wire [4-1:0] node21166;
	wire [4-1:0] node21167;
	wire [4-1:0] node21170;
	wire [4-1:0] node21173;
	wire [4-1:0] node21174;
	wire [4-1:0] node21176;
	wire [4-1:0] node21180;
	wire [4-1:0] node21182;
	wire [4-1:0] node21183;
	wire [4-1:0] node21187;
	wire [4-1:0] node21188;
	wire [4-1:0] node21191;
	wire [4-1:0] node21192;
	wire [4-1:0] node21193;
	wire [4-1:0] node21194;
	wire [4-1:0] node21199;
	wire [4-1:0] node21200;
	wire [4-1:0] node21204;
	wire [4-1:0] node21205;
	wire [4-1:0] node21206;
	wire [4-1:0] node21207;
	wire [4-1:0] node21211;
	wire [4-1:0] node21212;
	wire [4-1:0] node21213;
	wire [4-1:0] node21214;
	wire [4-1:0] node21219;
	wire [4-1:0] node21222;
	wire [4-1:0] node21223;
	wire [4-1:0] node21224;
	wire [4-1:0] node21225;
	wire [4-1:0] node21230;
	wire [4-1:0] node21231;
	wire [4-1:0] node21232;
	wire [4-1:0] node21236;
	wire [4-1:0] node21237;
	wire [4-1:0] node21241;
	wire [4-1:0] node21242;
	wire [4-1:0] node21243;
	wire [4-1:0] node21244;
	wire [4-1:0] node21245;
	wire [4-1:0] node21246;
	wire [4-1:0] node21249;
	wire [4-1:0] node21251;
	wire [4-1:0] node21252;
	wire [4-1:0] node21256;
	wire [4-1:0] node21257;
	wire [4-1:0] node21258;
	wire [4-1:0] node21260;
	wire [4-1:0] node21264;
	wire [4-1:0] node21265;
	wire [4-1:0] node21268;
	wire [4-1:0] node21270;
	wire [4-1:0] node21273;
	wire [4-1:0] node21274;
	wire [4-1:0] node21275;
	wire [4-1:0] node21278;
	wire [4-1:0] node21279;
	wire [4-1:0] node21283;
	wire [4-1:0] node21284;
	wire [4-1:0] node21285;
	wire [4-1:0] node21287;
	wire [4-1:0] node21291;
	wire [4-1:0] node21294;
	wire [4-1:0] node21295;
	wire [4-1:0] node21296;
	wire [4-1:0] node21297;
	wire [4-1:0] node21298;
	wire [4-1:0] node21299;
	wire [4-1:0] node21304;
	wire [4-1:0] node21307;
	wire [4-1:0] node21308;
	wire [4-1:0] node21310;
	wire [4-1:0] node21313;
	wire [4-1:0] node21314;
	wire [4-1:0] node21318;
	wire [4-1:0] node21319;
	wire [4-1:0] node21320;
	wire [4-1:0] node21321;
	wire [4-1:0] node21323;
	wire [4-1:0] node21327;
	wire [4-1:0] node21328;
	wire [4-1:0] node21329;
	wire [4-1:0] node21332;
	wire [4-1:0] node21336;
	wire [4-1:0] node21338;
	wire [4-1:0] node21341;
	wire [4-1:0] node21342;
	wire [4-1:0] node21343;
	wire [4-1:0] node21344;
	wire [4-1:0] node21345;
	wire [4-1:0] node21346;
	wire [4-1:0] node21347;
	wire [4-1:0] node21350;
	wire [4-1:0] node21354;
	wire [4-1:0] node21356;
	wire [4-1:0] node21358;
	wire [4-1:0] node21361;
	wire [4-1:0] node21362;
	wire [4-1:0] node21363;
	wire [4-1:0] node21366;
	wire [4-1:0] node21370;
	wire [4-1:0] node21371;
	wire [4-1:0] node21372;
	wire [4-1:0] node21373;
	wire [4-1:0] node21374;
	wire [4-1:0] node21378;
	wire [4-1:0] node21381;
	wire [4-1:0] node21382;
	wire [4-1:0] node21386;
	wire [4-1:0] node21387;
	wire [4-1:0] node21390;
	wire [4-1:0] node21393;
	wire [4-1:0] node21394;
	wire [4-1:0] node21395;
	wire [4-1:0] node21396;
	wire [4-1:0] node21397;
	wire [4-1:0] node21398;
	wire [4-1:0] node21402;
	wire [4-1:0] node21405;
	wire [4-1:0] node21408;
	wire [4-1:0] node21410;
	wire [4-1:0] node21411;
	wire [4-1:0] node21415;
	wire [4-1:0] node21416;
	wire [4-1:0] node21417;
	wire [4-1:0] node21419;
	wire [4-1:0] node21420;
	wire [4-1:0] node21424;
	wire [4-1:0] node21425;
	wire [4-1:0] node21429;
	wire [4-1:0] node21430;
	wire [4-1:0] node21434;
	wire [4-1:0] node21435;
	wire [4-1:0] node21436;
	wire [4-1:0] node21437;
	wire [4-1:0] node21438;
	wire [4-1:0] node21439;
	wire [4-1:0] node21440;
	wire [4-1:0] node21442;
	wire [4-1:0] node21445;
	wire [4-1:0] node21446;
	wire [4-1:0] node21449;
	wire [4-1:0] node21451;
	wire [4-1:0] node21454;
	wire [4-1:0] node21455;
	wire [4-1:0] node21456;
	wire [4-1:0] node21459;
	wire [4-1:0] node21463;
	wire [4-1:0] node21464;
	wire [4-1:0] node21466;
	wire [4-1:0] node21467;
	wire [4-1:0] node21470;
	wire [4-1:0] node21473;
	wire [4-1:0] node21474;
	wire [4-1:0] node21476;
	wire [4-1:0] node21479;
	wire [4-1:0] node21480;
	wire [4-1:0] node21484;
	wire [4-1:0] node21485;
	wire [4-1:0] node21486;
	wire [4-1:0] node21487;
	wire [4-1:0] node21491;
	wire [4-1:0] node21492;
	wire [4-1:0] node21493;
	wire [4-1:0] node21497;
	wire [4-1:0] node21500;
	wire [4-1:0] node21501;
	wire [4-1:0] node21502;
	wire [4-1:0] node21503;
	wire [4-1:0] node21504;
	wire [4-1:0] node21508;
	wire [4-1:0] node21509;
	wire [4-1:0] node21513;
	wire [4-1:0] node21515;
	wire [4-1:0] node21518;
	wire [4-1:0] node21519;
	wire [4-1:0] node21520;
	wire [4-1:0] node21521;
	wire [4-1:0] node21524;
	wire [4-1:0] node21528;
	wire [4-1:0] node21531;
	wire [4-1:0] node21532;
	wire [4-1:0] node21533;
	wire [4-1:0] node21534;
	wire [4-1:0] node21535;
	wire [4-1:0] node21536;
	wire [4-1:0] node21540;
	wire [4-1:0] node21542;
	wire [4-1:0] node21544;
	wire [4-1:0] node21547;
	wire [4-1:0] node21548;
	wire [4-1:0] node21550;
	wire [4-1:0] node21551;
	wire [4-1:0] node21554;
	wire [4-1:0] node21557;
	wire [4-1:0] node21558;
	wire [4-1:0] node21560;
	wire [4-1:0] node21563;
	wire [4-1:0] node21564;
	wire [4-1:0] node21568;
	wire [4-1:0] node21569;
	wire [4-1:0] node21570;
	wire [4-1:0] node21571;
	wire [4-1:0] node21572;
	wire [4-1:0] node21575;
	wire [4-1:0] node21578;
	wire [4-1:0] node21580;
	wire [4-1:0] node21583;
	wire [4-1:0] node21586;
	wire [4-1:0] node21587;
	wire [4-1:0] node21590;
	wire [4-1:0] node21591;
	wire [4-1:0] node21594;
	wire [4-1:0] node21597;
	wire [4-1:0] node21598;
	wire [4-1:0] node21599;
	wire [4-1:0] node21600;
	wire [4-1:0] node21603;
	wire [4-1:0] node21606;
	wire [4-1:0] node21607;
	wire [4-1:0] node21610;
	wire [4-1:0] node21613;
	wire [4-1:0] node21614;
	wire [4-1:0] node21615;
	wire [4-1:0] node21618;
	wire [4-1:0] node21619;
	wire [4-1:0] node21623;
	wire [4-1:0] node21625;
	wire [4-1:0] node21626;
	wire [4-1:0] node21629;
	wire [4-1:0] node21632;
	wire [4-1:0] node21633;
	wire [4-1:0] node21634;
	wire [4-1:0] node21635;
	wire [4-1:0] node21636;
	wire [4-1:0] node21638;
	wire [4-1:0] node21639;
	wire [4-1:0] node21641;
	wire [4-1:0] node21645;
	wire [4-1:0] node21647;
	wire [4-1:0] node21648;
	wire [4-1:0] node21649;
	wire [4-1:0] node21654;
	wire [4-1:0] node21655;
	wire [4-1:0] node21656;
	wire [4-1:0] node21657;
	wire [4-1:0] node21660;
	wire [4-1:0] node21663;
	wire [4-1:0] node21664;
	wire [4-1:0] node21665;
	wire [4-1:0] node21669;
	wire [4-1:0] node21671;
	wire [4-1:0] node21674;
	wire [4-1:0] node21675;
	wire [4-1:0] node21676;
	wire [4-1:0] node21680;
	wire [4-1:0] node21682;
	wire [4-1:0] node21685;
	wire [4-1:0] node21686;
	wire [4-1:0] node21687;
	wire [4-1:0] node21688;
	wire [4-1:0] node21689;
	wire [4-1:0] node21692;
	wire [4-1:0] node21695;
	wire [4-1:0] node21697;
	wire [4-1:0] node21698;
	wire [4-1:0] node21701;
	wire [4-1:0] node21704;
	wire [4-1:0] node21706;
	wire [4-1:0] node21707;
	wire [4-1:0] node21709;
	wire [4-1:0] node21713;
	wire [4-1:0] node21714;
	wire [4-1:0] node21717;
	wire [4-1:0] node21718;
	wire [4-1:0] node21719;
	wire [4-1:0] node21722;
	wire [4-1:0] node21726;
	wire [4-1:0] node21727;
	wire [4-1:0] node21728;
	wire [4-1:0] node21729;
	wire [4-1:0] node21730;
	wire [4-1:0] node21732;
	wire [4-1:0] node21735;
	wire [4-1:0] node21737;
	wire [4-1:0] node21740;
	wire [4-1:0] node21741;
	wire [4-1:0] node21742;
	wire [4-1:0] node21746;
	wire [4-1:0] node21747;
	wire [4-1:0] node21751;
	wire [4-1:0] node21752;
	wire [4-1:0] node21753;
	wire [4-1:0] node21756;
	wire [4-1:0] node21759;
	wire [4-1:0] node21760;
	wire [4-1:0] node21761;
	wire [4-1:0] node21765;
	wire [4-1:0] node21767;
	wire [4-1:0] node21768;
	wire [4-1:0] node21772;
	wire [4-1:0] node21773;
	wire [4-1:0] node21774;
	wire [4-1:0] node21776;
	wire [4-1:0] node21777;
	wire [4-1:0] node21778;
	wire [4-1:0] node21781;
	wire [4-1:0] node21785;
	wire [4-1:0] node21786;
	wire [4-1:0] node21787;
	wire [4-1:0] node21791;
	wire [4-1:0] node21792;
	wire [4-1:0] node21796;
	wire [4-1:0] node21797;
	wire [4-1:0] node21798;
	wire [4-1:0] node21801;
	wire [4-1:0] node21803;
	wire [4-1:0] node21804;
	wire [4-1:0] node21808;
	wire [4-1:0] node21809;
	wire [4-1:0] node21813;
	wire [4-1:0] node21814;
	wire [4-1:0] node21815;
	wire [4-1:0] node21816;
	wire [4-1:0] node21817;
	wire [4-1:0] node21818;
	wire [4-1:0] node21819;
	wire [4-1:0] node21820;
	wire [4-1:0] node21821;
	wire [4-1:0] node21822;
	wire [4-1:0] node21824;
	wire [4-1:0] node21827;
	wire [4-1:0] node21830;
	wire [4-1:0] node21831;
	wire [4-1:0] node21832;
	wire [4-1:0] node21836;
	wire [4-1:0] node21838;
	wire [4-1:0] node21841;
	wire [4-1:0] node21842;
	wire [4-1:0] node21843;
	wire [4-1:0] node21844;
	wire [4-1:0] node21848;
	wire [4-1:0] node21851;
	wire [4-1:0] node21853;
	wire [4-1:0] node21856;
	wire [4-1:0] node21857;
	wire [4-1:0] node21858;
	wire [4-1:0] node21860;
	wire [4-1:0] node21861;
	wire [4-1:0] node21865;
	wire [4-1:0] node21866;
	wire [4-1:0] node21868;
	wire [4-1:0] node21869;
	wire [4-1:0] node21874;
	wire [4-1:0] node21875;
	wire [4-1:0] node21876;
	wire [4-1:0] node21879;
	wire [4-1:0] node21880;
	wire [4-1:0] node21884;
	wire [4-1:0] node21885;
	wire [4-1:0] node21888;
	wire [4-1:0] node21891;
	wire [4-1:0] node21892;
	wire [4-1:0] node21893;
	wire [4-1:0] node21894;
	wire [4-1:0] node21895;
	wire [4-1:0] node21897;
	wire [4-1:0] node21901;
	wire [4-1:0] node21902;
	wire [4-1:0] node21906;
	wire [4-1:0] node21907;
	wire [4-1:0] node21909;
	wire [4-1:0] node21912;
	wire [4-1:0] node21914;
	wire [4-1:0] node21917;
	wire [4-1:0] node21918;
	wire [4-1:0] node21919;
	wire [4-1:0] node21920;
	wire [4-1:0] node21924;
	wire [4-1:0] node21925;
	wire [4-1:0] node21926;
	wire [4-1:0] node21927;
	wire [4-1:0] node21930;
	wire [4-1:0] node21935;
	wire [4-1:0] node21936;
	wire [4-1:0] node21937;
	wire [4-1:0] node21939;
	wire [4-1:0] node21942;
	wire [4-1:0] node21943;
	wire [4-1:0] node21946;
	wire [4-1:0] node21949;
	wire [4-1:0] node21950;
	wire [4-1:0] node21952;
	wire [4-1:0] node21953;
	wire [4-1:0] node21957;
	wire [4-1:0] node21959;
	wire [4-1:0] node21962;
	wire [4-1:0] node21963;
	wire [4-1:0] node21964;
	wire [4-1:0] node21965;
	wire [4-1:0] node21966;
	wire [4-1:0] node21967;
	wire [4-1:0] node21968;
	wire [4-1:0] node21971;
	wire [4-1:0] node21975;
	wire [4-1:0] node21976;
	wire [4-1:0] node21978;
	wire [4-1:0] node21981;
	wire [4-1:0] node21984;
	wire [4-1:0] node21985;
	wire [4-1:0] node21986;
	wire [4-1:0] node21988;
	wire [4-1:0] node21991;
	wire [4-1:0] node21993;
	wire [4-1:0] node21996;
	wire [4-1:0] node21997;
	wire [4-1:0] node21998;
	wire [4-1:0] node21999;
	wire [4-1:0] node22003;
	wire [4-1:0] node22007;
	wire [4-1:0] node22008;
	wire [4-1:0] node22009;
	wire [4-1:0] node22011;
	wire [4-1:0] node22012;
	wire [4-1:0] node22015;
	wire [4-1:0] node22018;
	wire [4-1:0] node22019;
	wire [4-1:0] node22020;
	wire [4-1:0] node22021;
	wire [4-1:0] node22027;
	wire [4-1:0] node22028;
	wire [4-1:0] node22029;
	wire [4-1:0] node22030;
	wire [4-1:0] node22031;
	wire [4-1:0] node22036;
	wire [4-1:0] node22039;
	wire [4-1:0] node22040;
	wire [4-1:0] node22043;
	wire [4-1:0] node22045;
	wire [4-1:0] node22046;
	wire [4-1:0] node22050;
	wire [4-1:0] node22051;
	wire [4-1:0] node22052;
	wire [4-1:0] node22053;
	wire [4-1:0] node22054;
	wire [4-1:0] node22055;
	wire [4-1:0] node22058;
	wire [4-1:0] node22063;
	wire [4-1:0] node22064;
	wire [4-1:0] node22066;
	wire [4-1:0] node22067;
	wire [4-1:0] node22071;
	wire [4-1:0] node22072;
	wire [4-1:0] node22074;
	wire [4-1:0] node22075;
	wire [4-1:0] node22079;
	wire [4-1:0] node22081;
	wire [4-1:0] node22084;
	wire [4-1:0] node22085;
	wire [4-1:0] node22086;
	wire [4-1:0] node22087;
	wire [4-1:0] node22088;
	wire [4-1:0] node22091;
	wire [4-1:0] node22095;
	wire [4-1:0] node22096;
	wire [4-1:0] node22097;
	wire [4-1:0] node22101;
	wire [4-1:0] node22102;
	wire [4-1:0] node22106;
	wire [4-1:0] node22107;
	wire [4-1:0] node22108;
	wire [4-1:0] node22109;
	wire [4-1:0] node22110;
	wire [4-1:0] node22115;
	wire [4-1:0] node22116;
	wire [4-1:0] node22119;
	wire [4-1:0] node22120;
	wire [4-1:0] node22124;
	wire [4-1:0] node22125;
	wire [4-1:0] node22127;
	wire [4-1:0] node22128;
	wire [4-1:0] node22131;
	wire [4-1:0] node22134;
	wire [4-1:0] node22135;
	wire [4-1:0] node22137;
	wire [4-1:0] node22140;
	wire [4-1:0] node22141;
	wire [4-1:0] node22144;
	wire [4-1:0] node22147;
	wire [4-1:0] node22148;
	wire [4-1:0] node22149;
	wire [4-1:0] node22150;
	wire [4-1:0] node22151;
	wire [4-1:0] node22152;
	wire [4-1:0] node22153;
	wire [4-1:0] node22154;
	wire [4-1:0] node22158;
	wire [4-1:0] node22159;
	wire [4-1:0] node22163;
	wire [4-1:0] node22164;
	wire [4-1:0] node22167;
	wire [4-1:0] node22168;
	wire [4-1:0] node22170;
	wire [4-1:0] node22174;
	wire [4-1:0] node22175;
	wire [4-1:0] node22176;
	wire [4-1:0] node22177;
	wire [4-1:0] node22178;
	wire [4-1:0] node22183;
	wire [4-1:0] node22186;
	wire [4-1:0] node22188;
	wire [4-1:0] node22189;
	wire [4-1:0] node22190;
	wire [4-1:0] node22193;
	wire [4-1:0] node22197;
	wire [4-1:0] node22198;
	wire [4-1:0] node22199;
	wire [4-1:0] node22200;
	wire [4-1:0] node22201;
	wire [4-1:0] node22202;
	wire [4-1:0] node22206;
	wire [4-1:0] node22207;
	wire [4-1:0] node22211;
	wire [4-1:0] node22213;
	wire [4-1:0] node22216;
	wire [4-1:0] node22217;
	wire [4-1:0] node22220;
	wire [4-1:0] node22222;
	wire [4-1:0] node22225;
	wire [4-1:0] node22226;
	wire [4-1:0] node22227;
	wire [4-1:0] node22228;
	wire [4-1:0] node22232;
	wire [4-1:0] node22233;
	wire [4-1:0] node22235;
	wire [4-1:0] node22239;
	wire [4-1:0] node22240;
	wire [4-1:0] node22242;
	wire [4-1:0] node22243;
	wire [4-1:0] node22248;
	wire [4-1:0] node22249;
	wire [4-1:0] node22250;
	wire [4-1:0] node22251;
	wire [4-1:0] node22252;
	wire [4-1:0] node22255;
	wire [4-1:0] node22257;
	wire [4-1:0] node22260;
	wire [4-1:0] node22261;
	wire [4-1:0] node22262;
	wire [4-1:0] node22267;
	wire [4-1:0] node22268;
	wire [4-1:0] node22269;
	wire [4-1:0] node22270;
	wire [4-1:0] node22271;
	wire [4-1:0] node22275;
	wire [4-1:0] node22277;
	wire [4-1:0] node22280;
	wire [4-1:0] node22282;
	wire [4-1:0] node22285;
	wire [4-1:0] node22286;
	wire [4-1:0] node22289;
	wire [4-1:0] node22292;
	wire [4-1:0] node22293;
	wire [4-1:0] node22294;
	wire [4-1:0] node22295;
	wire [4-1:0] node22297;
	wire [4-1:0] node22300;
	wire [4-1:0] node22302;
	wire [4-1:0] node22305;
	wire [4-1:0] node22306;
	wire [4-1:0] node22309;
	wire [4-1:0] node22312;
	wire [4-1:0] node22313;
	wire [4-1:0] node22315;
	wire [4-1:0] node22316;
	wire [4-1:0] node22320;
	wire [4-1:0] node22323;
	wire [4-1:0] node22324;
	wire [4-1:0] node22325;
	wire [4-1:0] node22326;
	wire [4-1:0] node22327;
	wire [4-1:0] node22329;
	wire [4-1:0] node22331;
	wire [4-1:0] node22332;
	wire [4-1:0] node22336;
	wire [4-1:0] node22337;
	wire [4-1:0] node22339;
	wire [4-1:0] node22343;
	wire [4-1:0] node22344;
	wire [4-1:0] node22345;
	wire [4-1:0] node22348;
	wire [4-1:0] node22351;
	wire [4-1:0] node22352;
	wire [4-1:0] node22353;
	wire [4-1:0] node22357;
	wire [4-1:0] node22358;
	wire [4-1:0] node22362;
	wire [4-1:0] node22363;
	wire [4-1:0] node22364;
	wire [4-1:0] node22365;
	wire [4-1:0] node22367;
	wire [4-1:0] node22368;
	wire [4-1:0] node22371;
	wire [4-1:0] node22375;
	wire [4-1:0] node22376;
	wire [4-1:0] node22377;
	wire [4-1:0] node22378;
	wire [4-1:0] node22382;
	wire [4-1:0] node22383;
	wire [4-1:0] node22386;
	wire [4-1:0] node22390;
	wire [4-1:0] node22391;
	wire [4-1:0] node22392;
	wire [4-1:0] node22393;
	wire [4-1:0] node22395;
	wire [4-1:0] node22400;
	wire [4-1:0] node22401;
	wire [4-1:0] node22402;
	wire [4-1:0] node22403;
	wire [4-1:0] node22406;
	wire [4-1:0] node22410;
	wire [4-1:0] node22412;
	wire [4-1:0] node22415;
	wire [4-1:0] node22416;
	wire [4-1:0] node22417;
	wire [4-1:0] node22418;
	wire [4-1:0] node22419;
	wire [4-1:0] node22420;
	wire [4-1:0] node22422;
	wire [4-1:0] node22425;
	wire [4-1:0] node22429;
	wire [4-1:0] node22430;
	wire [4-1:0] node22432;
	wire [4-1:0] node22435;
	wire [4-1:0] node22436;
	wire [4-1:0] node22439;
	wire [4-1:0] node22442;
	wire [4-1:0] node22443;
	wire [4-1:0] node22444;
	wire [4-1:0] node22446;
	wire [4-1:0] node22449;
	wire [4-1:0] node22450;
	wire [4-1:0] node22451;
	wire [4-1:0] node22455;
	wire [4-1:0] node22456;
	wire [4-1:0] node22460;
	wire [4-1:0] node22461;
	wire [4-1:0] node22462;
	wire [4-1:0] node22463;
	wire [4-1:0] node22467;
	wire [4-1:0] node22470;
	wire [4-1:0] node22472;
	wire [4-1:0] node22475;
	wire [4-1:0] node22476;
	wire [4-1:0] node22477;
	wire [4-1:0] node22478;
	wire [4-1:0] node22479;
	wire [4-1:0] node22482;
	wire [4-1:0] node22486;
	wire [4-1:0] node22488;
	wire [4-1:0] node22489;
	wire [4-1:0] node22490;
	wire [4-1:0] node22494;
	wire [4-1:0] node22495;
	wire [4-1:0] node22499;
	wire [4-1:0] node22500;
	wire [4-1:0] node22501;
	wire [4-1:0] node22502;
	wire [4-1:0] node22503;
	wire [4-1:0] node22507;
	wire [4-1:0] node22509;
	wire [4-1:0] node22513;
	wire [4-1:0] node22514;
	wire [4-1:0] node22515;
	wire [4-1:0] node22516;
	wire [4-1:0] node22519;
	wire [4-1:0] node22523;
	wire [4-1:0] node22524;
	wire [4-1:0] node22528;
	wire [4-1:0] node22529;
	wire [4-1:0] node22530;
	wire [4-1:0] node22531;
	wire [4-1:0] node22532;
	wire [4-1:0] node22533;
	wire [4-1:0] node22534;
	wire [4-1:0] node22536;
	wire [4-1:0] node22538;
	wire [4-1:0] node22541;
	wire [4-1:0] node22542;
	wire [4-1:0] node22544;
	wire [4-1:0] node22547;
	wire [4-1:0] node22549;
	wire [4-1:0] node22550;
	wire [4-1:0] node22554;
	wire [4-1:0] node22555;
	wire [4-1:0] node22556;
	wire [4-1:0] node22559;
	wire [4-1:0] node22561;
	wire [4-1:0] node22564;
	wire [4-1:0] node22565;
	wire [4-1:0] node22566;
	wire [4-1:0] node22571;
	wire [4-1:0] node22572;
	wire [4-1:0] node22573;
	wire [4-1:0] node22574;
	wire [4-1:0] node22577;
	wire [4-1:0] node22579;
	wire [4-1:0] node22582;
	wire [4-1:0] node22583;
	wire [4-1:0] node22584;
	wire [4-1:0] node22587;
	wire [4-1:0] node22590;
	wire [4-1:0] node22592;
	wire [4-1:0] node22595;
	wire [4-1:0] node22596;
	wire [4-1:0] node22598;
	wire [4-1:0] node22599;
	wire [4-1:0] node22602;
	wire [4-1:0] node22605;
	wire [4-1:0] node22606;
	wire [4-1:0] node22609;
	wire [4-1:0] node22612;
	wire [4-1:0] node22613;
	wire [4-1:0] node22614;
	wire [4-1:0] node22615;
	wire [4-1:0] node22617;
	wire [4-1:0] node22618;
	wire [4-1:0] node22621;
	wire [4-1:0] node22623;
	wire [4-1:0] node22626;
	wire [4-1:0] node22627;
	wire [4-1:0] node22631;
	wire [4-1:0] node22632;
	wire [4-1:0] node22633;
	wire [4-1:0] node22635;
	wire [4-1:0] node22638;
	wire [4-1:0] node22639;
	wire [4-1:0] node22643;
	wire [4-1:0] node22644;
	wire [4-1:0] node22648;
	wire [4-1:0] node22649;
	wire [4-1:0] node22650;
	wire [4-1:0] node22652;
	wire [4-1:0] node22653;
	wire [4-1:0] node22656;
	wire [4-1:0] node22659;
	wire [4-1:0] node22660;
	wire [4-1:0] node22663;
	wire [4-1:0] node22665;
	wire [4-1:0] node22668;
	wire [4-1:0] node22669;
	wire [4-1:0] node22670;
	wire [4-1:0] node22672;
	wire [4-1:0] node22674;
	wire [4-1:0] node22677;
	wire [4-1:0] node22678;
	wire [4-1:0] node22680;
	wire [4-1:0] node22684;
	wire [4-1:0] node22685;
	wire [4-1:0] node22688;
	wire [4-1:0] node22691;
	wire [4-1:0] node22692;
	wire [4-1:0] node22693;
	wire [4-1:0] node22694;
	wire [4-1:0] node22695;
	wire [4-1:0] node22696;
	wire [4-1:0] node22697;
	wire [4-1:0] node22699;
	wire [4-1:0] node22702;
	wire [4-1:0] node22705;
	wire [4-1:0] node22706;
	wire [4-1:0] node22710;
	wire [4-1:0] node22712;
	wire [4-1:0] node22713;
	wire [4-1:0] node22714;
	wire [4-1:0] node22718;
	wire [4-1:0] node22719;
	wire [4-1:0] node22723;
	wire [4-1:0] node22724;
	wire [4-1:0] node22725;
	wire [4-1:0] node22729;
	wire [4-1:0] node22731;
	wire [4-1:0] node22732;
	wire [4-1:0] node22736;
	wire [4-1:0] node22737;
	wire [4-1:0] node22738;
	wire [4-1:0] node22739;
	wire [4-1:0] node22740;
	wire [4-1:0] node22744;
	wire [4-1:0] node22746;
	wire [4-1:0] node22747;
	wire [4-1:0] node22750;
	wire [4-1:0] node22753;
	wire [4-1:0] node22754;
	wire [4-1:0] node22755;
	wire [4-1:0] node22758;
	wire [4-1:0] node22761;
	wire [4-1:0] node22763;
	wire [4-1:0] node22766;
	wire [4-1:0] node22767;
	wire [4-1:0] node22768;
	wire [4-1:0] node22769;
	wire [4-1:0] node22770;
	wire [4-1:0] node22775;
	wire [4-1:0] node22776;
	wire [4-1:0] node22777;
	wire [4-1:0] node22782;
	wire [4-1:0] node22783;
	wire [4-1:0] node22785;
	wire [4-1:0] node22788;
	wire [4-1:0] node22789;
	wire [4-1:0] node22790;
	wire [4-1:0] node22795;
	wire [4-1:0] node22796;
	wire [4-1:0] node22797;
	wire [4-1:0] node22798;
	wire [4-1:0] node22799;
	wire [4-1:0] node22800;
	wire [4-1:0] node22803;
	wire [4-1:0] node22806;
	wire [4-1:0] node22809;
	wire [4-1:0] node22810;
	wire [4-1:0] node22811;
	wire [4-1:0] node22813;
	wire [4-1:0] node22817;
	wire [4-1:0] node22819;
	wire [4-1:0] node22821;
	wire [4-1:0] node22824;
	wire [4-1:0] node22825;
	wire [4-1:0] node22826;
	wire [4-1:0] node22828;
	wire [4-1:0] node22831;
	wire [4-1:0] node22832;
	wire [4-1:0] node22836;
	wire [4-1:0] node22837;
	wire [4-1:0] node22840;
	wire [4-1:0] node22843;
	wire [4-1:0] node22844;
	wire [4-1:0] node22845;
	wire [4-1:0] node22846;
	wire [4-1:0] node22847;
	wire [4-1:0] node22850;
	wire [4-1:0] node22853;
	wire [4-1:0] node22854;
	wire [4-1:0] node22857;
	wire [4-1:0] node22860;
	wire [4-1:0] node22861;
	wire [4-1:0] node22862;
	wire [4-1:0] node22864;
	wire [4-1:0] node22868;
	wire [4-1:0] node22870;
	wire [4-1:0] node22873;
	wire [4-1:0] node22874;
	wire [4-1:0] node22875;
	wire [4-1:0] node22876;
	wire [4-1:0] node22880;
	wire [4-1:0] node22883;
	wire [4-1:0] node22884;
	wire [4-1:0] node22888;
	wire [4-1:0] node22889;
	wire [4-1:0] node22890;
	wire [4-1:0] node22891;
	wire [4-1:0] node22892;
	wire [4-1:0] node22893;
	wire [4-1:0] node22894;
	wire [4-1:0] node22895;
	wire [4-1:0] node22897;
	wire [4-1:0] node22900;
	wire [4-1:0] node22903;
	wire [4-1:0] node22905;
	wire [4-1:0] node22908;
	wire [4-1:0] node22909;
	wire [4-1:0] node22910;
	wire [4-1:0] node22911;
	wire [4-1:0] node22916;
	wire [4-1:0] node22918;
	wire [4-1:0] node22921;
	wire [4-1:0] node22922;
	wire [4-1:0] node22923;
	wire [4-1:0] node22924;
	wire [4-1:0] node22925;
	wire [4-1:0] node22928;
	wire [4-1:0] node22931;
	wire [4-1:0] node22932;
	wire [4-1:0] node22935;
	wire [4-1:0] node22938;
	wire [4-1:0] node22939;
	wire [4-1:0] node22941;
	wire [4-1:0] node22944;
	wire [4-1:0] node22946;
	wire [4-1:0] node22949;
	wire [4-1:0] node22950;
	wire [4-1:0] node22952;
	wire [4-1:0] node22955;
	wire [4-1:0] node22957;
	wire [4-1:0] node22958;
	wire [4-1:0] node22962;
	wire [4-1:0] node22963;
	wire [4-1:0] node22964;
	wire [4-1:0] node22965;
	wire [4-1:0] node22966;
	wire [4-1:0] node22970;
	wire [4-1:0] node22973;
	wire [4-1:0] node22974;
	wire [4-1:0] node22975;
	wire [4-1:0] node22979;
	wire [4-1:0] node22982;
	wire [4-1:0] node22983;
	wire [4-1:0] node22984;
	wire [4-1:0] node22985;
	wire [4-1:0] node22987;
	wire [4-1:0] node22990;
	wire [4-1:0] node22993;
	wire [4-1:0] node22996;
	wire [4-1:0] node22997;
	wire [4-1:0] node22999;
	wire [4-1:0] node23000;
	wire [4-1:0] node23004;
	wire [4-1:0] node23005;
	wire [4-1:0] node23006;
	wire [4-1:0] node23009;
	wire [4-1:0] node23013;
	wire [4-1:0] node23014;
	wire [4-1:0] node23015;
	wire [4-1:0] node23016;
	wire [4-1:0] node23017;
	wire [4-1:0] node23019;
	wire [4-1:0] node23022;
	wire [4-1:0] node23023;
	wire [4-1:0] node23026;
	wire [4-1:0] node23029;
	wire [4-1:0] node23031;
	wire [4-1:0] node23032;
	wire [4-1:0] node23035;
	wire [4-1:0] node23038;
	wire [4-1:0] node23039;
	wire [4-1:0] node23040;
	wire [4-1:0] node23043;
	wire [4-1:0] node23044;
	wire [4-1:0] node23048;
	wire [4-1:0] node23049;
	wire [4-1:0] node23050;
	wire [4-1:0] node23053;
	wire [4-1:0] node23056;
	wire [4-1:0] node23058;
	wire [4-1:0] node23061;
	wire [4-1:0] node23062;
	wire [4-1:0] node23063;
	wire [4-1:0] node23065;
	wire [4-1:0] node23066;
	wire [4-1:0] node23068;
	wire [4-1:0] node23072;
	wire [4-1:0] node23074;
	wire [4-1:0] node23075;
	wire [4-1:0] node23078;
	wire [4-1:0] node23081;
	wire [4-1:0] node23082;
	wire [4-1:0] node23083;
	wire [4-1:0] node23084;
	wire [4-1:0] node23088;
	wire [4-1:0] node23089;
	wire [4-1:0] node23093;
	wire [4-1:0] node23094;
	wire [4-1:0] node23097;
	wire [4-1:0] node23098;
	wire [4-1:0] node23102;
	wire [4-1:0] node23103;
	wire [4-1:0] node23104;
	wire [4-1:0] node23105;
	wire [4-1:0] node23106;
	wire [4-1:0] node23107;
	wire [4-1:0] node23108;
	wire [4-1:0] node23111;
	wire [4-1:0] node23115;
	wire [4-1:0] node23117;
	wire [4-1:0] node23118;
	wire [4-1:0] node23119;
	wire [4-1:0] node23124;
	wire [4-1:0] node23125;
	wire [4-1:0] node23126;
	wire [4-1:0] node23129;
	wire [4-1:0] node23131;
	wire [4-1:0] node23134;
	wire [4-1:0] node23135;
	wire [4-1:0] node23136;
	wire [4-1:0] node23137;
	wire [4-1:0] node23140;
	wire [4-1:0] node23143;
	wire [4-1:0] node23146;
	wire [4-1:0] node23147;
	wire [4-1:0] node23150;
	wire [4-1:0] node23153;
	wire [4-1:0] node23154;
	wire [4-1:0] node23155;
	wire [4-1:0] node23156;
	wire [4-1:0] node23157;
	wire [4-1:0] node23158;
	wire [4-1:0] node23162;
	wire [4-1:0] node23165;
	wire [4-1:0] node23168;
	wire [4-1:0] node23170;
	wire [4-1:0] node23172;
	wire [4-1:0] node23175;
	wire [4-1:0] node23176;
	wire [4-1:0] node23178;
	wire [4-1:0] node23180;
	wire [4-1:0] node23183;
	wire [4-1:0] node23185;
	wire [4-1:0] node23186;
	wire [4-1:0] node23189;
	wire [4-1:0] node23192;
	wire [4-1:0] node23193;
	wire [4-1:0] node23194;
	wire [4-1:0] node23195;
	wire [4-1:0] node23198;
	wire [4-1:0] node23200;
	wire [4-1:0] node23201;
	wire [4-1:0] node23205;
	wire [4-1:0] node23206;
	wire [4-1:0] node23207;
	wire [4-1:0] node23208;
	wire [4-1:0] node23211;
	wire [4-1:0] node23215;
	wire [4-1:0] node23217;
	wire [4-1:0] node23218;
	wire [4-1:0] node23222;
	wire [4-1:0] node23223;
	wire [4-1:0] node23224;
	wire [4-1:0] node23225;
	wire [4-1:0] node23226;
	wire [4-1:0] node23229;
	wire [4-1:0] node23230;
	wire [4-1:0] node23235;
	wire [4-1:0] node23236;
	wire [4-1:0] node23237;
	wire [4-1:0] node23241;
	wire [4-1:0] node23242;
	wire [4-1:0] node23246;
	wire [4-1:0] node23247;
	wire [4-1:0] node23248;
	wire [4-1:0] node23249;
	wire [4-1:0] node23250;
	wire [4-1:0] node23255;
	wire [4-1:0] node23256;
	wire [4-1:0] node23260;
	wire [4-1:0] node23262;
	wire [4-1:0] node23263;
	wire [4-1:0] node23267;
	wire [4-1:0] node23268;
	wire [4-1:0] node23269;
	wire [4-1:0] node23270;
	wire [4-1:0] node23271;
	wire [4-1:0] node23272;
	wire [4-1:0] node23273;
	wire [4-1:0] node23274;
	wire [4-1:0] node23275;
	wire [4-1:0] node23276;
	wire [4-1:0] node23277;
	wire [4-1:0] node23282;
	wire [4-1:0] node23283;
	wire [4-1:0] node23287;
	wire [4-1:0] node23288;
	wire [4-1:0] node23291;
	wire [4-1:0] node23292;
	wire [4-1:0] node23293;
	wire [4-1:0] node23298;
	wire [4-1:0] node23299;
	wire [4-1:0] node23300;
	wire [4-1:0] node23302;
	wire [4-1:0] node23303;
	wire [4-1:0] node23306;
	wire [4-1:0] node23309;
	wire [4-1:0] node23310;
	wire [4-1:0] node23314;
	wire [4-1:0] node23315;
	wire [4-1:0] node23318;
	wire [4-1:0] node23320;
	wire [4-1:0] node23321;
	wire [4-1:0] node23325;
	wire [4-1:0] node23326;
	wire [4-1:0] node23327;
	wire [4-1:0] node23328;
	wire [4-1:0] node23330;
	wire [4-1:0] node23333;
	wire [4-1:0] node23334;
	wire [4-1:0] node23337;
	wire [4-1:0] node23340;
	wire [4-1:0] node23341;
	wire [4-1:0] node23344;
	wire [4-1:0] node23347;
	wire [4-1:0] node23348;
	wire [4-1:0] node23350;
	wire [4-1:0] node23352;
	wire [4-1:0] node23353;
	wire [4-1:0] node23356;
	wire [4-1:0] node23359;
	wire [4-1:0] node23362;
	wire [4-1:0] node23363;
	wire [4-1:0] node23364;
	wire [4-1:0] node23365;
	wire [4-1:0] node23366;
	wire [4-1:0] node23368;
	wire [4-1:0] node23371;
	wire [4-1:0] node23374;
	wire [4-1:0] node23376;
	wire [4-1:0] node23377;
	wire [4-1:0] node23380;
	wire [4-1:0] node23383;
	wire [4-1:0] node23384;
	wire [4-1:0] node23385;
	wire [4-1:0] node23388;
	wire [4-1:0] node23389;
	wire [4-1:0] node23393;
	wire [4-1:0] node23394;
	wire [4-1:0] node23395;
	wire [4-1:0] node23398;
	wire [4-1:0] node23401;
	wire [4-1:0] node23402;
	wire [4-1:0] node23404;
	wire [4-1:0] node23407;
	wire [4-1:0] node23408;
	wire [4-1:0] node23412;
	wire [4-1:0] node23413;
	wire [4-1:0] node23414;
	wire [4-1:0] node23415;
	wire [4-1:0] node23416;
	wire [4-1:0] node23417;
	wire [4-1:0] node23420;
	wire [4-1:0] node23424;
	wire [4-1:0] node23426;
	wire [4-1:0] node23427;
	wire [4-1:0] node23430;
	wire [4-1:0] node23433;
	wire [4-1:0] node23434;
	wire [4-1:0] node23435;
	wire [4-1:0] node23436;
	wire [4-1:0] node23440;
	wire [4-1:0] node23441;
	wire [4-1:0] node23445;
	wire [4-1:0] node23448;
	wire [4-1:0] node23449;
	wire [4-1:0] node23450;
	wire [4-1:0] node23451;
	wire [4-1:0] node23452;
	wire [4-1:0] node23455;
	wire [4-1:0] node23458;
	wire [4-1:0] node23460;
	wire [4-1:0] node23464;
	wire [4-1:0] node23465;
	wire [4-1:0] node23467;
	wire [4-1:0] node23470;
	wire [4-1:0] node23473;
	wire [4-1:0] node23474;
	wire [4-1:0] node23475;
	wire [4-1:0] node23476;
	wire [4-1:0] node23477;
	wire [4-1:0] node23478;
	wire [4-1:0] node23480;
	wire [4-1:0] node23484;
	wire [4-1:0] node23485;
	wire [4-1:0] node23487;
	wire [4-1:0] node23490;
	wire [4-1:0] node23492;
	wire [4-1:0] node23495;
	wire [4-1:0] node23496;
	wire [4-1:0] node23498;
	wire [4-1:0] node23500;
	wire [4-1:0] node23504;
	wire [4-1:0] node23505;
	wire [4-1:0] node23506;
	wire [4-1:0] node23507;
	wire [4-1:0] node23509;
	wire [4-1:0] node23510;
	wire [4-1:0] node23514;
	wire [4-1:0] node23517;
	wire [4-1:0] node23518;
	wire [4-1:0] node23519;
	wire [4-1:0] node23521;
	wire [4-1:0] node23524;
	wire [4-1:0] node23527;
	wire [4-1:0] node23528;
	wire [4-1:0] node23529;
	wire [4-1:0] node23532;
	wire [4-1:0] node23536;
	wire [4-1:0] node23537;
	wire [4-1:0] node23538;
	wire [4-1:0] node23541;
	wire [4-1:0] node23544;
	wire [4-1:0] node23545;
	wire [4-1:0] node23547;
	wire [4-1:0] node23550;
	wire [4-1:0] node23552;
	wire [4-1:0] node23555;
	wire [4-1:0] node23556;
	wire [4-1:0] node23557;
	wire [4-1:0] node23558;
	wire [4-1:0] node23559;
	wire [4-1:0] node23561;
	wire [4-1:0] node23564;
	wire [4-1:0] node23566;
	wire [4-1:0] node23569;
	wire [4-1:0] node23570;
	wire [4-1:0] node23571;
	wire [4-1:0] node23573;
	wire [4-1:0] node23577;
	wire [4-1:0] node23579;
	wire [4-1:0] node23582;
	wire [4-1:0] node23583;
	wire [4-1:0] node23584;
	wire [4-1:0] node23586;
	wire [4-1:0] node23587;
	wire [4-1:0] node23591;
	wire [4-1:0] node23592;
	wire [4-1:0] node23595;
	wire [4-1:0] node23598;
	wire [4-1:0] node23599;
	wire [4-1:0] node23602;
	wire [4-1:0] node23603;
	wire [4-1:0] node23607;
	wire [4-1:0] node23608;
	wire [4-1:0] node23609;
	wire [4-1:0] node23610;
	wire [4-1:0] node23611;
	wire [4-1:0] node23612;
	wire [4-1:0] node23615;
	wire [4-1:0] node23619;
	wire [4-1:0] node23620;
	wire [4-1:0] node23621;
	wire [4-1:0] node23626;
	wire [4-1:0] node23627;
	wire [4-1:0] node23628;
	wire [4-1:0] node23631;
	wire [4-1:0] node23635;
	wire [4-1:0] node23636;
	wire [4-1:0] node23637;
	wire [4-1:0] node23639;
	wire [4-1:0] node23642;
	wire [4-1:0] node23643;
	wire [4-1:0] node23647;
	wire [4-1:0] node23649;
	wire [4-1:0] node23652;
	wire [4-1:0] node23653;
	wire [4-1:0] node23654;
	wire [4-1:0] node23655;
	wire [4-1:0] node23656;
	wire [4-1:0] node23657;
	wire [4-1:0] node23658;
	wire [4-1:0] node23659;
	wire [4-1:0] node23663;
	wire [4-1:0] node23664;
	wire [4-1:0] node23668;
	wire [4-1:0] node23669;
	wire [4-1:0] node23672;
	wire [4-1:0] node23673;
	wire [4-1:0] node23674;
	wire [4-1:0] node23678;
	wire [4-1:0] node23679;
	wire [4-1:0] node23683;
	wire [4-1:0] node23684;
	wire [4-1:0] node23685;
	wire [4-1:0] node23686;
	wire [4-1:0] node23690;
	wire [4-1:0] node23692;
	wire [4-1:0] node23695;
	wire [4-1:0] node23696;
	wire [4-1:0] node23697;
	wire [4-1:0] node23699;
	wire [4-1:0] node23702;
	wire [4-1:0] node23705;
	wire [4-1:0] node23706;
	wire [4-1:0] node23710;
	wire [4-1:0] node23711;
	wire [4-1:0] node23712;
	wire [4-1:0] node23713;
	wire [4-1:0] node23714;
	wire [4-1:0] node23715;
	wire [4-1:0] node23718;
	wire [4-1:0] node23722;
	wire [4-1:0] node23723;
	wire [4-1:0] node23726;
	wire [4-1:0] node23729;
	wire [4-1:0] node23730;
	wire [4-1:0] node23731;
	wire [4-1:0] node23732;
	wire [4-1:0] node23737;
	wire [4-1:0] node23738;
	wire [4-1:0] node23741;
	wire [4-1:0] node23743;
	wire [4-1:0] node23746;
	wire [4-1:0] node23747;
	wire [4-1:0] node23748;
	wire [4-1:0] node23752;
	wire [4-1:0] node23754;
	wire [4-1:0] node23756;
	wire [4-1:0] node23759;
	wire [4-1:0] node23760;
	wire [4-1:0] node23761;
	wire [4-1:0] node23762;
	wire [4-1:0] node23763;
	wire [4-1:0] node23766;
	wire [4-1:0] node23768;
	wire [4-1:0] node23771;
	wire [4-1:0] node23772;
	wire [4-1:0] node23773;
	wire [4-1:0] node23774;
	wire [4-1:0] node23779;
	wire [4-1:0] node23780;
	wire [4-1:0] node23783;
	wire [4-1:0] node23786;
	wire [4-1:0] node23787;
	wire [4-1:0] node23788;
	wire [4-1:0] node23789;
	wire [4-1:0] node23792;
	wire [4-1:0] node23795;
	wire [4-1:0] node23797;
	wire [4-1:0] node23800;
	wire [4-1:0] node23801;
	wire [4-1:0] node23802;
	wire [4-1:0] node23803;
	wire [4-1:0] node23806;
	wire [4-1:0] node23809;
	wire [4-1:0] node23811;
	wire [4-1:0] node23815;
	wire [4-1:0] node23816;
	wire [4-1:0] node23817;
	wire [4-1:0] node23818;
	wire [4-1:0] node23819;
	wire [4-1:0] node23822;
	wire [4-1:0] node23823;
	wire [4-1:0] node23828;
	wire [4-1:0] node23829;
	wire [4-1:0] node23830;
	wire [4-1:0] node23831;
	wire [4-1:0] node23834;
	wire [4-1:0] node23839;
	wire [4-1:0] node23840;
	wire [4-1:0] node23841;
	wire [4-1:0] node23843;
	wire [4-1:0] node23844;
	wire [4-1:0] node23847;
	wire [4-1:0] node23850;
	wire [4-1:0] node23851;
	wire [4-1:0] node23853;
	wire [4-1:0] node23856;
	wire [4-1:0] node23859;
	wire [4-1:0] node23861;
	wire [4-1:0] node23862;
	wire [4-1:0] node23865;
	wire [4-1:0] node23867;
	wire [4-1:0] node23870;
	wire [4-1:0] node23871;
	wire [4-1:0] node23872;
	wire [4-1:0] node23873;
	wire [4-1:0] node23874;
	wire [4-1:0] node23875;
	wire [4-1:0] node23878;
	wire [4-1:0] node23879;
	wire [4-1:0] node23883;
	wire [4-1:0] node23884;
	wire [4-1:0] node23886;
	wire [4-1:0] node23887;
	wire [4-1:0] node23891;
	wire [4-1:0] node23893;
	wire [4-1:0] node23896;
	wire [4-1:0] node23897;
	wire [4-1:0] node23898;
	wire [4-1:0] node23900;
	wire [4-1:0] node23902;
	wire [4-1:0] node23905;
	wire [4-1:0] node23906;
	wire [4-1:0] node23909;
	wire [4-1:0] node23912;
	wire [4-1:0] node23913;
	wire [4-1:0] node23914;
	wire [4-1:0] node23915;
	wire [4-1:0] node23920;
	wire [4-1:0] node23921;
	wire [4-1:0] node23924;
	wire [4-1:0] node23927;
	wire [4-1:0] node23928;
	wire [4-1:0] node23929;
	wire [4-1:0] node23930;
	wire [4-1:0] node23931;
	wire [4-1:0] node23933;
	wire [4-1:0] node23937;
	wire [4-1:0] node23938;
	wire [4-1:0] node23942;
	wire [4-1:0] node23943;
	wire [4-1:0] node23944;
	wire [4-1:0] node23946;
	wire [4-1:0] node23950;
	wire [4-1:0] node23951;
	wire [4-1:0] node23955;
	wire [4-1:0] node23956;
	wire [4-1:0] node23959;
	wire [4-1:0] node23960;
	wire [4-1:0] node23961;
	wire [4-1:0] node23965;
	wire [4-1:0] node23966;
	wire [4-1:0] node23969;
	wire [4-1:0] node23972;
	wire [4-1:0] node23973;
	wire [4-1:0] node23974;
	wire [4-1:0] node23975;
	wire [4-1:0] node23976;
	wire [4-1:0] node23978;
	wire [4-1:0] node23981;
	wire [4-1:0] node23982;
	wire [4-1:0] node23983;
	wire [4-1:0] node23988;
	wire [4-1:0] node23989;
	wire [4-1:0] node23990;
	wire [4-1:0] node23992;
	wire [4-1:0] node23996;
	wire [4-1:0] node23999;
	wire [4-1:0] node24000;
	wire [4-1:0] node24001;
	wire [4-1:0] node24002;
	wire [4-1:0] node24006;
	wire [4-1:0] node24008;
	wire [4-1:0] node24011;
	wire [4-1:0] node24012;
	wire [4-1:0] node24013;
	wire [4-1:0] node24017;
	wire [4-1:0] node24018;
	wire [4-1:0] node24019;
	wire [4-1:0] node24022;
	wire [4-1:0] node24026;
	wire [4-1:0] node24027;
	wire [4-1:0] node24028;
	wire [4-1:0] node24029;
	wire [4-1:0] node24031;
	wire [4-1:0] node24032;
	wire [4-1:0] node24036;
	wire [4-1:0] node24037;
	wire [4-1:0] node24038;
	wire [4-1:0] node24041;
	wire [4-1:0] node24045;
	wire [4-1:0] node24046;
	wire [4-1:0] node24047;
	wire [4-1:0] node24051;
	wire [4-1:0] node24053;
	wire [4-1:0] node24056;
	wire [4-1:0] node24057;
	wire [4-1:0] node24058;
	wire [4-1:0] node24059;
	wire [4-1:0] node24063;
	wire [4-1:0] node24066;
	wire [4-1:0] node24067;
	wire [4-1:0] node24068;
	wire [4-1:0] node24069;
	wire [4-1:0] node24074;
	wire [4-1:0] node24076;
	wire [4-1:0] node24079;
	wire [4-1:0] node24080;
	wire [4-1:0] node24081;
	wire [4-1:0] node24082;
	wire [4-1:0] node24083;
	wire [4-1:0] node24084;
	wire [4-1:0] node24085;
	wire [4-1:0] node24086;
	wire [4-1:0] node24087;
	wire [4-1:0] node24090;
	wire [4-1:0] node24092;
	wire [4-1:0] node24095;
	wire [4-1:0] node24097;
	wire [4-1:0] node24100;
	wire [4-1:0] node24101;
	wire [4-1:0] node24102;
	wire [4-1:0] node24105;
	wire [4-1:0] node24108;
	wire [4-1:0] node24109;
	wire [4-1:0] node24113;
	wire [4-1:0] node24114;
	wire [4-1:0] node24115;
	wire [4-1:0] node24117;
	wire [4-1:0] node24121;
	wire [4-1:0] node24122;
	wire [4-1:0] node24124;
	wire [4-1:0] node24127;
	wire [4-1:0] node24129;
	wire [4-1:0] node24132;
	wire [4-1:0] node24133;
	wire [4-1:0] node24134;
	wire [4-1:0] node24135;
	wire [4-1:0] node24136;
	wire [4-1:0] node24139;
	wire [4-1:0] node24143;
	wire [4-1:0] node24145;
	wire [4-1:0] node24146;
	wire [4-1:0] node24149;
	wire [4-1:0] node24152;
	wire [4-1:0] node24153;
	wire [4-1:0] node24155;
	wire [4-1:0] node24158;
	wire [4-1:0] node24159;
	wire [4-1:0] node24163;
	wire [4-1:0] node24164;
	wire [4-1:0] node24165;
	wire [4-1:0] node24166;
	wire [4-1:0] node24167;
	wire [4-1:0] node24169;
	wire [4-1:0] node24172;
	wire [4-1:0] node24173;
	wire [4-1:0] node24174;
	wire [4-1:0] node24179;
	wire [4-1:0] node24180;
	wire [4-1:0] node24183;
	wire [4-1:0] node24184;
	wire [4-1:0] node24188;
	wire [4-1:0] node24189;
	wire [4-1:0] node24190;
	wire [4-1:0] node24191;
	wire [4-1:0] node24192;
	wire [4-1:0] node24195;
	wire [4-1:0] node24199;
	wire [4-1:0] node24202;
	wire [4-1:0] node24203;
	wire [4-1:0] node24204;
	wire [4-1:0] node24208;
	wire [4-1:0] node24209;
	wire [4-1:0] node24211;
	wire [4-1:0] node24214;
	wire [4-1:0] node24217;
	wire [4-1:0] node24218;
	wire [4-1:0] node24219;
	wire [4-1:0] node24220;
	wire [4-1:0] node24223;
	wire [4-1:0] node24225;
	wire [4-1:0] node24228;
	wire [4-1:0] node24229;
	wire [4-1:0] node24233;
	wire [4-1:0] node24234;
	wire [4-1:0] node24235;
	wire [4-1:0] node24236;
	wire [4-1:0] node24239;
	wire [4-1:0] node24242;
	wire [4-1:0] node24244;
	wire [4-1:0] node24247;
	wire [4-1:0] node24248;
	wire [4-1:0] node24249;
	wire [4-1:0] node24251;
	wire [4-1:0] node24256;
	wire [4-1:0] node24257;
	wire [4-1:0] node24258;
	wire [4-1:0] node24259;
	wire [4-1:0] node24260;
	wire [4-1:0] node24262;
	wire [4-1:0] node24263;
	wire [4-1:0] node24266;
	wire [4-1:0] node24269;
	wire [4-1:0] node24270;
	wire [4-1:0] node24271;
	wire [4-1:0] node24275;
	wire [4-1:0] node24278;
	wire [4-1:0] node24279;
	wire [4-1:0] node24281;
	wire [4-1:0] node24282;
	wire [4-1:0] node24283;
	wire [4-1:0] node24287;
	wire [4-1:0] node24288;
	wire [4-1:0] node24292;
	wire [4-1:0] node24293;
	wire [4-1:0] node24296;
	wire [4-1:0] node24297;
	wire [4-1:0] node24299;
	wire [4-1:0] node24303;
	wire [4-1:0] node24304;
	wire [4-1:0] node24305;
	wire [4-1:0] node24306;
	wire [4-1:0] node24308;
	wire [4-1:0] node24312;
	wire [4-1:0] node24313;
	wire [4-1:0] node24314;
	wire [4-1:0] node24317;
	wire [4-1:0] node24320;
	wire [4-1:0] node24323;
	wire [4-1:0] node24324;
	wire [4-1:0] node24325;
	wire [4-1:0] node24326;
	wire [4-1:0] node24327;
	wire [4-1:0] node24331;
	wire [4-1:0] node24333;
	wire [4-1:0] node24336;
	wire [4-1:0] node24338;
	wire [4-1:0] node24341;
	wire [4-1:0] node24342;
	wire [4-1:0] node24343;
	wire [4-1:0] node24345;
	wire [4-1:0] node24349;
	wire [4-1:0] node24352;
	wire [4-1:0] node24353;
	wire [4-1:0] node24354;
	wire [4-1:0] node24355;
	wire [4-1:0] node24356;
	wire [4-1:0] node24358;
	wire [4-1:0] node24360;
	wire [4-1:0] node24363;
	wire [4-1:0] node24366;
	wire [4-1:0] node24367;
	wire [4-1:0] node24368;
	wire [4-1:0] node24371;
	wire [4-1:0] node24374;
	wire [4-1:0] node24376;
	wire [4-1:0] node24379;
	wire [4-1:0] node24380;
	wire [4-1:0] node24381;
	wire [4-1:0] node24383;
	wire [4-1:0] node24386;
	wire [4-1:0] node24387;
	wire [4-1:0] node24388;
	wire [4-1:0] node24393;
	wire [4-1:0] node24395;
	wire [4-1:0] node24396;
	wire [4-1:0] node24397;
	wire [4-1:0] node24400;
	wire [4-1:0] node24404;
	wire [4-1:0] node24405;
	wire [4-1:0] node24406;
	wire [4-1:0] node24407;
	wire [4-1:0] node24409;
	wire [4-1:0] node24412;
	wire [4-1:0] node24415;
	wire [4-1:0] node24416;
	wire [4-1:0] node24417;
	wire [4-1:0] node24420;
	wire [4-1:0] node24423;
	wire [4-1:0] node24426;
	wire [4-1:0] node24427;
	wire [4-1:0] node24428;
	wire [4-1:0] node24429;
	wire [4-1:0] node24432;
	wire [4-1:0] node24436;
	wire [4-1:0] node24437;
	wire [4-1:0] node24440;
	wire [4-1:0] node24441;
	wire [4-1:0] node24444;
	wire [4-1:0] node24447;
	wire [4-1:0] node24448;
	wire [4-1:0] node24449;
	wire [4-1:0] node24450;
	wire [4-1:0] node24451;
	wire [4-1:0] node24452;
	wire [4-1:0] node24453;
	wire [4-1:0] node24454;
	wire [4-1:0] node24457;
	wire [4-1:0] node24460;
	wire [4-1:0] node24461;
	wire [4-1:0] node24464;
	wire [4-1:0] node24466;
	wire [4-1:0] node24469;
	wire [4-1:0] node24471;
	wire [4-1:0] node24472;
	wire [4-1:0] node24475;
	wire [4-1:0] node24478;
	wire [4-1:0] node24479;
	wire [4-1:0] node24480;
	wire [4-1:0] node24481;
	wire [4-1:0] node24484;
	wire [4-1:0] node24487;
	wire [4-1:0] node24488;
	wire [4-1:0] node24491;
	wire [4-1:0] node24493;
	wire [4-1:0] node24496;
	wire [4-1:0] node24498;
	wire [4-1:0] node24499;
	wire [4-1:0] node24502;
	wire [4-1:0] node24505;
	wire [4-1:0] node24506;
	wire [4-1:0] node24507;
	wire [4-1:0] node24508;
	wire [4-1:0] node24509;
	wire [4-1:0] node24510;
	wire [4-1:0] node24513;
	wire [4-1:0] node24516;
	wire [4-1:0] node24518;
	wire [4-1:0] node24521;
	wire [4-1:0] node24522;
	wire [4-1:0] node24526;
	wire [4-1:0] node24527;
	wire [4-1:0] node24529;
	wire [4-1:0] node24532;
	wire [4-1:0] node24533;
	wire [4-1:0] node24534;
	wire [4-1:0] node24538;
	wire [4-1:0] node24541;
	wire [4-1:0] node24542;
	wire [4-1:0] node24543;
	wire [4-1:0] node24544;
	wire [4-1:0] node24547;
	wire [4-1:0] node24550;
	wire [4-1:0] node24551;
	wire [4-1:0] node24555;
	wire [4-1:0] node24556;
	wire [4-1:0] node24558;
	wire [4-1:0] node24560;
	wire [4-1:0] node24563;
	wire [4-1:0] node24564;
	wire [4-1:0] node24568;
	wire [4-1:0] node24569;
	wire [4-1:0] node24570;
	wire [4-1:0] node24571;
	wire [4-1:0] node24572;
	wire [4-1:0] node24573;
	wire [4-1:0] node24574;
	wire [4-1:0] node24577;
	wire [4-1:0] node24580;
	wire [4-1:0] node24583;
	wire [4-1:0] node24584;
	wire [4-1:0] node24585;
	wire [4-1:0] node24588;
	wire [4-1:0] node24592;
	wire [4-1:0] node24593;
	wire [4-1:0] node24595;
	wire [4-1:0] node24598;
	wire [4-1:0] node24599;
	wire [4-1:0] node24601;
	wire [4-1:0] node24604;
	wire [4-1:0] node24606;
	wire [4-1:0] node24609;
	wire [4-1:0] node24610;
	wire [4-1:0] node24611;
	wire [4-1:0] node24612;
	wire [4-1:0] node24615;
	wire [4-1:0] node24616;
	wire [4-1:0] node24619;
	wire [4-1:0] node24622;
	wire [4-1:0] node24625;
	wire [4-1:0] node24626;
	wire [4-1:0] node24627;
	wire [4-1:0] node24630;
	wire [4-1:0] node24631;
	wire [4-1:0] node24634;
	wire [4-1:0] node24637;
	wire [4-1:0] node24639;
	wire [4-1:0] node24640;
	wire [4-1:0] node24643;
	wire [4-1:0] node24646;
	wire [4-1:0] node24647;
	wire [4-1:0] node24648;
	wire [4-1:0] node24649;
	wire [4-1:0] node24651;
	wire [4-1:0] node24653;
	wire [4-1:0] node24656;
	wire [4-1:0] node24659;
	wire [4-1:0] node24660;
	wire [4-1:0] node24663;
	wire [4-1:0] node24665;
	wire [4-1:0] node24666;
	wire [4-1:0] node24670;
	wire [4-1:0] node24671;
	wire [4-1:0] node24672;
	wire [4-1:0] node24673;
	wire [4-1:0] node24675;
	wire [4-1:0] node24678;
	wire [4-1:0] node24679;
	wire [4-1:0] node24683;
	wire [4-1:0] node24686;
	wire [4-1:0] node24687;
	wire [4-1:0] node24691;
	wire [4-1:0] node24692;
	wire [4-1:0] node24693;
	wire [4-1:0] node24694;
	wire [4-1:0] node24695;
	wire [4-1:0] node24696;
	wire [4-1:0] node24697;
	wire [4-1:0] node24698;
	wire [4-1:0] node24702;
	wire [4-1:0] node24705;
	wire [4-1:0] node24706;
	wire [4-1:0] node24708;
	wire [4-1:0] node24711;
	wire [4-1:0] node24712;
	wire [4-1:0] node24716;
	wire [4-1:0] node24717;
	wire [4-1:0] node24718;
	wire [4-1:0] node24719;
	wire [4-1:0] node24722;
	wire [4-1:0] node24725;
	wire [4-1:0] node24728;
	wire [4-1:0] node24729;
	wire [4-1:0] node24732;
	wire [4-1:0] node24733;
	wire [4-1:0] node24736;
	wire [4-1:0] node24739;
	wire [4-1:0] node24740;
	wire [4-1:0] node24741;
	wire [4-1:0] node24742;
	wire [4-1:0] node24744;
	wire [4-1:0] node24747;
	wire [4-1:0] node24749;
	wire [4-1:0] node24753;
	wire [4-1:0] node24754;
	wire [4-1:0] node24756;
	wire [4-1:0] node24759;
	wire [4-1:0] node24761;
	wire [4-1:0] node24764;
	wire [4-1:0] node24765;
	wire [4-1:0] node24766;
	wire [4-1:0] node24767;
	wire [4-1:0] node24768;
	wire [4-1:0] node24769;
	wire [4-1:0] node24772;
	wire [4-1:0] node24776;
	wire [4-1:0] node24777;
	wire [4-1:0] node24781;
	wire [4-1:0] node24782;
	wire [4-1:0] node24783;
	wire [4-1:0] node24788;
	wire [4-1:0] node24789;
	wire [4-1:0] node24790;
	wire [4-1:0] node24792;
	wire [4-1:0] node24795;
	wire [4-1:0] node24796;
	wire [4-1:0] node24799;
	wire [4-1:0] node24802;
	wire [4-1:0] node24805;
	wire [4-1:0] node24806;
	wire [4-1:0] node24807;
	wire [4-1:0] node24808;
	wire [4-1:0] node24809;
	wire [4-1:0] node24811;
	wire [4-1:0] node24814;
	wire [4-1:0] node24817;
	wire [4-1:0] node24818;
	wire [4-1:0] node24821;
	wire [4-1:0] node24824;
	wire [4-1:0] node24825;
	wire [4-1:0] node24826;
	wire [4-1:0] node24827;
	wire [4-1:0] node24832;
	wire [4-1:0] node24833;
	wire [4-1:0] node24836;
	wire [4-1:0] node24839;
	wire [4-1:0] node24840;
	wire [4-1:0] node24841;
	wire [4-1:0] node24843;
	wire [4-1:0] node24846;
	wire [4-1:0] node24848;
	wire [4-1:0] node24851;
	wire [4-1:0] node24852;
	wire [4-1:0] node24853;
	wire [4-1:0] node24856;
	wire [4-1:0] node24859;
	wire [4-1:0] node24861;
	wire [4-1:0] node24864;
	wire [4-1:0] node24865;
	wire [4-1:0] node24866;
	wire [4-1:0] node24867;
	wire [4-1:0] node24868;
	wire [4-1:0] node24869;
	wire [4-1:0] node24870;
	wire [4-1:0] node24871;
	wire [4-1:0] node24872;
	wire [4-1:0] node24873;
	wire [4-1:0] node24874;
	wire [4-1:0] node24877;
	wire [4-1:0] node24880;
	wire [4-1:0] node24881;
	wire [4-1:0] node24882;
	wire [4-1:0] node24883;
	wire [4-1:0] node24887;
	wire [4-1:0] node24889;
	wire [4-1:0] node24890;
	wire [4-1:0] node24893;
	wire [4-1:0] node24896;
	wire [4-1:0] node24897;
	wire [4-1:0] node24899;
	wire [4-1:0] node24902;
	wire [4-1:0] node24904;
	wire [4-1:0] node24905;
	wire [4-1:0] node24908;
	wire [4-1:0] node24911;
	wire [4-1:0] node24912;
	wire [4-1:0] node24913;
	wire [4-1:0] node24916;
	wire [4-1:0] node24919;
	wire [4-1:0] node24920;
	wire [4-1:0] node24921;
	wire [4-1:0] node24924;
	wire [4-1:0] node24927;
	wire [4-1:0] node24929;
	wire [4-1:0] node24930;
	wire [4-1:0] node24934;
	wire [4-1:0] node24935;
	wire [4-1:0] node24936;
	wire [4-1:0] node24937;
	wire [4-1:0] node24940;
	wire [4-1:0] node24943;
	wire [4-1:0] node24944;
	wire [4-1:0] node24945;
	wire [4-1:0] node24946;
	wire [4-1:0] node24949;
	wire [4-1:0] node24952;
	wire [4-1:0] node24953;
	wire [4-1:0] node24954;
	wire [4-1:0] node24956;
	wire [4-1:0] node24959;
	wire [4-1:0] node24963;
	wire [4-1:0] node24964;
	wire [4-1:0] node24966;
	wire [4-1:0] node24968;
	wire [4-1:0] node24971;
	wire [4-1:0] node24973;
	wire [4-1:0] node24975;
	wire [4-1:0] node24978;
	wire [4-1:0] node24979;
	wire [4-1:0] node24980;
	wire [4-1:0] node24981;
	wire [4-1:0] node24982;
	wire [4-1:0] node24985;
	wire [4-1:0] node24987;
	wire [4-1:0] node24991;
	wire [4-1:0] node24992;
	wire [4-1:0] node24993;
	wire [4-1:0] node24996;
	wire [4-1:0] node24999;
	wire [4-1:0] node25000;
	wire [4-1:0] node25003;
	wire [4-1:0] node25006;
	wire [4-1:0] node25007;
	wire [4-1:0] node25008;
	wire [4-1:0] node25009;
	wire [4-1:0] node25012;
	wire [4-1:0] node25015;
	wire [4-1:0] node25017;
	wire [4-1:0] node25019;
	wire [4-1:0] node25021;
	wire [4-1:0] node25024;
	wire [4-1:0] node25025;
	wire [4-1:0] node25026;
	wire [4-1:0] node25027;
	wire [4-1:0] node25032;
	wire [4-1:0] node25034;
	wire [4-1:0] node25036;
	wire [4-1:0] node25038;
	wire [4-1:0] node25041;
	wire [4-1:0] node25042;
	wire [4-1:0] node25043;
	wire [4-1:0] node25044;
	wire [4-1:0] node25045;
	wire [4-1:0] node25046;
	wire [4-1:0] node25047;
	wire [4-1:0] node25050;
	wire [4-1:0] node25053;
	wire [4-1:0] node25054;
	wire [4-1:0] node25056;
	wire [4-1:0] node25059;
	wire [4-1:0] node25062;
	wire [4-1:0] node25063;
	wire [4-1:0] node25065;
	wire [4-1:0] node25066;
	wire [4-1:0] node25070;
	wire [4-1:0] node25071;
	wire [4-1:0] node25074;
	wire [4-1:0] node25075;
	wire [4-1:0] node25079;
	wire [4-1:0] node25080;
	wire [4-1:0] node25081;
	wire [4-1:0] node25082;
	wire [4-1:0] node25083;
	wire [4-1:0] node25086;
	wire [4-1:0] node25089;
	wire [4-1:0] node25091;
	wire [4-1:0] node25094;
	wire [4-1:0] node25096;
	wire [4-1:0] node25099;
	wire [4-1:0] node25100;
	wire [4-1:0] node25101;
	wire [4-1:0] node25103;
	wire [4-1:0] node25106;
	wire [4-1:0] node25108;
	wire [4-1:0] node25111;
	wire [4-1:0] node25112;
	wire [4-1:0] node25114;
	wire [4-1:0] node25117;
	wire [4-1:0] node25118;
	wire [4-1:0] node25121;
	wire [4-1:0] node25124;
	wire [4-1:0] node25125;
	wire [4-1:0] node25126;
	wire [4-1:0] node25127;
	wire [4-1:0] node25128;
	wire [4-1:0] node25131;
	wire [4-1:0] node25133;
	wire [4-1:0] node25135;
	wire [4-1:0] node25138;
	wire [4-1:0] node25139;
	wire [4-1:0] node25140;
	wire [4-1:0] node25141;
	wire [4-1:0] node25147;
	wire [4-1:0] node25148;
	wire [4-1:0] node25151;
	wire [4-1:0] node25152;
	wire [4-1:0] node25155;
	wire [4-1:0] node25157;
	wire [4-1:0] node25160;
	wire [4-1:0] node25161;
	wire [4-1:0] node25162;
	wire [4-1:0] node25163;
	wire [4-1:0] node25164;
	wire [4-1:0] node25165;
	wire [4-1:0] node25169;
	wire [4-1:0] node25170;
	wire [4-1:0] node25174;
	wire [4-1:0] node25175;
	wire [4-1:0] node25178;
	wire [4-1:0] node25181;
	wire [4-1:0] node25182;
	wire [4-1:0] node25183;
	wire [4-1:0] node25184;
	wire [4-1:0] node25187;
	wire [4-1:0] node25190;
	wire [4-1:0] node25191;
	wire [4-1:0] node25194;
	wire [4-1:0] node25198;
	wire [4-1:0] node25199;
	wire [4-1:0] node25200;
	wire [4-1:0] node25201;
	wire [4-1:0] node25204;
	wire [4-1:0] node25205;
	wire [4-1:0] node25208;
	wire [4-1:0] node25211;
	wire [4-1:0] node25214;
	wire [4-1:0] node25215;
	wire [4-1:0] node25217;
	wire [4-1:0] node25218;
	wire [4-1:0] node25221;
	wire [4-1:0] node25224;
	wire [4-1:0] node25225;
	wire [4-1:0] node25227;
	wire [4-1:0] node25231;
	wire [4-1:0] node25232;
	wire [4-1:0] node25233;
	wire [4-1:0] node25234;
	wire [4-1:0] node25235;
	wire [4-1:0] node25238;
	wire [4-1:0] node25240;
	wire [4-1:0] node25242;
	wire [4-1:0] node25245;
	wire [4-1:0] node25246;
	wire [4-1:0] node25248;
	wire [4-1:0] node25250;
	wire [4-1:0] node25253;
	wire [4-1:0] node25254;
	wire [4-1:0] node25255;
	wire [4-1:0] node25257;
	wire [4-1:0] node25260;
	wire [4-1:0] node25263;
	wire [4-1:0] node25265;
	wire [4-1:0] node25268;
	wire [4-1:0] node25269;
	wire [4-1:0] node25270;
	wire [4-1:0] node25271;
	wire [4-1:0] node25275;
	wire [4-1:0] node25276;
	wire [4-1:0] node25277;
	wire [4-1:0] node25281;
	wire [4-1:0] node25282;
	wire [4-1:0] node25283;
	wire [4-1:0] node25288;
	wire [4-1:0] node25289;
	wire [4-1:0] node25290;
	wire [4-1:0] node25292;
	wire [4-1:0] node25295;
	wire [4-1:0] node25296;
	wire [4-1:0] node25298;
	wire [4-1:0] node25301;
	wire [4-1:0] node25302;
	wire [4-1:0] node25306;
	wire [4-1:0] node25307;
	wire [4-1:0] node25308;
	wire [4-1:0] node25311;
	wire [4-1:0] node25314;
	wire [4-1:0] node25317;
	wire [4-1:0] node25318;
	wire [4-1:0] node25319;
	wire [4-1:0] node25320;
	wire [4-1:0] node25321;
	wire [4-1:0] node25325;
	wire [4-1:0] node25327;
	wire [4-1:0] node25328;
	wire [4-1:0] node25331;
	wire [4-1:0] node25334;
	wire [4-1:0] node25336;
	wire [4-1:0] node25337;
	wire [4-1:0] node25338;
	wire [4-1:0] node25343;
	wire [4-1:0] node25344;
	wire [4-1:0] node25345;
	wire [4-1:0] node25346;
	wire [4-1:0] node25348;
	wire [4-1:0] node25351;
	wire [4-1:0] node25354;
	wire [4-1:0] node25355;
	wire [4-1:0] node25358;
	wire [4-1:0] node25359;
	wire [4-1:0] node25362;
	wire [4-1:0] node25365;
	wire [4-1:0] node25366;
	wire [4-1:0] node25367;
	wire [4-1:0] node25368;
	wire [4-1:0] node25369;
	wire [4-1:0] node25372;
	wire [4-1:0] node25375;
	wire [4-1:0] node25378;
	wire [4-1:0] node25381;
	wire [4-1:0] node25382;
	wire [4-1:0] node25385;
	wire [4-1:0] node25386;
	wire [4-1:0] node25389;
	wire [4-1:0] node25392;
	wire [4-1:0] node25393;
	wire [4-1:0] node25394;
	wire [4-1:0] node25395;
	wire [4-1:0] node25396;
	wire [4-1:0] node25397;
	wire [4-1:0] node25398;
	wire [4-1:0] node25400;
	wire [4-1:0] node25403;
	wire [4-1:0] node25405;
	wire [4-1:0] node25408;
	wire [4-1:0] node25409;
	wire [4-1:0] node25411;
	wire [4-1:0] node25414;
	wire [4-1:0] node25416;
	wire [4-1:0] node25419;
	wire [4-1:0] node25420;
	wire [4-1:0] node25421;
	wire [4-1:0] node25423;
	wire [4-1:0] node25424;
	wire [4-1:0] node25427;
	wire [4-1:0] node25430;
	wire [4-1:0] node25432;
	wire [4-1:0] node25433;
	wire [4-1:0] node25436;
	wire [4-1:0] node25439;
	wire [4-1:0] node25440;
	wire [4-1:0] node25441;
	wire [4-1:0] node25442;
	wire [4-1:0] node25447;
	wire [4-1:0] node25448;
	wire [4-1:0] node25450;
	wire [4-1:0] node25454;
	wire [4-1:0] node25455;
	wire [4-1:0] node25456;
	wire [4-1:0] node25457;
	wire [4-1:0] node25458;
	wire [4-1:0] node25460;
	wire [4-1:0] node25462;
	wire [4-1:0] node25465;
	wire [4-1:0] node25466;
	wire [4-1:0] node25470;
	wire [4-1:0] node25471;
	wire [4-1:0] node25475;
	wire [4-1:0] node25476;
	wire [4-1:0] node25478;
	wire [4-1:0] node25480;
	wire [4-1:0] node25483;
	wire [4-1:0] node25484;
	wire [4-1:0] node25487;
	wire [4-1:0] node25490;
	wire [4-1:0] node25491;
	wire [4-1:0] node25493;
	wire [4-1:0] node25494;
	wire [4-1:0] node25495;
	wire [4-1:0] node25498;
	wire [4-1:0] node25500;
	wire [4-1:0] node25503;
	wire [4-1:0] node25504;
	wire [4-1:0] node25505;
	wire [4-1:0] node25508;
	wire [4-1:0] node25512;
	wire [4-1:0] node25513;
	wire [4-1:0] node25514;
	wire [4-1:0] node25516;
	wire [4-1:0] node25519;
	wire [4-1:0] node25520;
	wire [4-1:0] node25523;
	wire [4-1:0] node25526;
	wire [4-1:0] node25527;
	wire [4-1:0] node25529;
	wire [4-1:0] node25532;
	wire [4-1:0] node25534;
	wire [4-1:0] node25535;
	wire [4-1:0] node25538;
	wire [4-1:0] node25541;
	wire [4-1:0] node25542;
	wire [4-1:0] node25543;
	wire [4-1:0] node25544;
	wire [4-1:0] node25545;
	wire [4-1:0] node25547;
	wire [4-1:0] node25550;
	wire [4-1:0] node25552;
	wire [4-1:0] node25555;
	wire [4-1:0] node25556;
	wire [4-1:0] node25558;
	wire [4-1:0] node25561;
	wire [4-1:0] node25563;
	wire [4-1:0] node25566;
	wire [4-1:0] node25567;
	wire [4-1:0] node25568;
	wire [4-1:0] node25569;
	wire [4-1:0] node25573;
	wire [4-1:0] node25574;
	wire [4-1:0] node25576;
	wire [4-1:0] node25580;
	wire [4-1:0] node25581;
	wire [4-1:0] node25582;
	wire [4-1:0] node25583;
	wire [4-1:0] node25584;
	wire [4-1:0] node25587;
	wire [4-1:0] node25591;
	wire [4-1:0] node25592;
	wire [4-1:0] node25593;
	wire [4-1:0] node25598;
	wire [4-1:0] node25600;
	wire [4-1:0] node25602;
	wire [4-1:0] node25605;
	wire [4-1:0] node25606;
	wire [4-1:0] node25607;
	wire [4-1:0] node25608;
	wire [4-1:0] node25609;
	wire [4-1:0] node25612;
	wire [4-1:0] node25615;
	wire [4-1:0] node25616;
	wire [4-1:0] node25620;
	wire [4-1:0] node25621;
	wire [4-1:0] node25622;
	wire [4-1:0] node25624;
	wire [4-1:0] node25627;
	wire [4-1:0] node25628;
	wire [4-1:0] node25631;
	wire [4-1:0] node25634;
	wire [4-1:0] node25636;
	wire [4-1:0] node25637;
	wire [4-1:0] node25638;
	wire [4-1:0] node25641;
	wire [4-1:0] node25645;
	wire [4-1:0] node25646;
	wire [4-1:0] node25647;
	wire [4-1:0] node25648;
	wire [4-1:0] node25650;
	wire [4-1:0] node25653;
	wire [4-1:0] node25655;
	wire [4-1:0] node25658;
	wire [4-1:0] node25660;
	wire [4-1:0] node25663;
	wire [4-1:0] node25664;
	wire [4-1:0] node25665;
	wire [4-1:0] node25668;
	wire [4-1:0] node25671;
	wire [4-1:0] node25673;
	wire [4-1:0] node25674;
	wire [4-1:0] node25677;
	wire [4-1:0] node25680;
	wire [4-1:0] node25681;
	wire [4-1:0] node25682;
	wire [4-1:0] node25683;
	wire [4-1:0] node25684;
	wire [4-1:0] node25685;
	wire [4-1:0] node25687;
	wire [4-1:0] node25688;
	wire [4-1:0] node25691;
	wire [4-1:0] node25693;
	wire [4-1:0] node25696;
	wire [4-1:0] node25697;
	wire [4-1:0] node25699;
	wire [4-1:0] node25702;
	wire [4-1:0] node25705;
	wire [4-1:0] node25706;
	wire [4-1:0] node25709;
	wire [4-1:0] node25710;
	wire [4-1:0] node25711;
	wire [4-1:0] node25714;
	wire [4-1:0] node25717;
	wire [4-1:0] node25718;
	wire [4-1:0] node25722;
	wire [4-1:0] node25723;
	wire [4-1:0] node25724;
	wire [4-1:0] node25725;
	wire [4-1:0] node25726;
	wire [4-1:0] node25727;
	wire [4-1:0] node25730;
	wire [4-1:0] node25734;
	wire [4-1:0] node25735;
	wire [4-1:0] node25736;
	wire [4-1:0] node25741;
	wire [4-1:0] node25742;
	wire [4-1:0] node25743;
	wire [4-1:0] node25745;
	wire [4-1:0] node25748;
	wire [4-1:0] node25750;
	wire [4-1:0] node25753;
	wire [4-1:0] node25754;
	wire [4-1:0] node25758;
	wire [4-1:0] node25759;
	wire [4-1:0] node25761;
	wire [4-1:0] node25762;
	wire [4-1:0] node25765;
	wire [4-1:0] node25768;
	wire [4-1:0] node25769;
	wire [4-1:0] node25772;
	wire [4-1:0] node25775;
	wire [4-1:0] node25776;
	wire [4-1:0] node25777;
	wire [4-1:0] node25778;
	wire [4-1:0] node25779;
	wire [4-1:0] node25781;
	wire [4-1:0] node25785;
	wire [4-1:0] node25786;
	wire [4-1:0] node25789;
	wire [4-1:0] node25790;
	wire [4-1:0] node25794;
	wire [4-1:0] node25795;
	wire [4-1:0] node25797;
	wire [4-1:0] node25800;
	wire [4-1:0] node25801;
	wire [4-1:0] node25803;
	wire [4-1:0] node25806;
	wire [4-1:0] node25809;
	wire [4-1:0] node25810;
	wire [4-1:0] node25811;
	wire [4-1:0] node25812;
	wire [4-1:0] node25816;
	wire [4-1:0] node25817;
	wire [4-1:0] node25820;
	wire [4-1:0] node25823;
	wire [4-1:0] node25824;
	wire [4-1:0] node25825;
	wire [4-1:0] node25826;
	wire [4-1:0] node25830;
	wire [4-1:0] node25831;
	wire [4-1:0] node25835;
	wire [4-1:0] node25836;
	wire [4-1:0] node25837;
	wire [4-1:0] node25841;
	wire [4-1:0] node25842;
	wire [4-1:0] node25846;
	wire [4-1:0] node25847;
	wire [4-1:0] node25848;
	wire [4-1:0] node25849;
	wire [4-1:0] node25850;
	wire [4-1:0] node25852;
	wire [4-1:0] node25853;
	wire [4-1:0] node25854;
	wire [4-1:0] node25859;
	wire [4-1:0] node25860;
	wire [4-1:0] node25861;
	wire [4-1:0] node25866;
	wire [4-1:0] node25867;
	wire [4-1:0] node25868;
	wire [4-1:0] node25869;
	wire [4-1:0] node25873;
	wire [4-1:0] node25875;
	wire [4-1:0] node25878;
	wire [4-1:0] node25879;
	wire [4-1:0] node25880;
	wire [4-1:0] node25883;
	wire [4-1:0] node25886;
	wire [4-1:0] node25887;
	wire [4-1:0] node25890;
	wire [4-1:0] node25893;
	wire [4-1:0] node25894;
	wire [4-1:0] node25895;
	wire [4-1:0] node25896;
	wire [4-1:0] node25898;
	wire [4-1:0] node25901;
	wire [4-1:0] node25902;
	wire [4-1:0] node25903;
	wire [4-1:0] node25908;
	wire [4-1:0] node25909;
	wire [4-1:0] node25910;
	wire [4-1:0] node25911;
	wire [4-1:0] node25916;
	wire [4-1:0] node25917;
	wire [4-1:0] node25920;
	wire [4-1:0] node25923;
	wire [4-1:0] node25924;
	wire [4-1:0] node25925;
	wire [4-1:0] node25926;
	wire [4-1:0] node25929;
	wire [4-1:0] node25932;
	wire [4-1:0] node25933;
	wire [4-1:0] node25934;
	wire [4-1:0] node25938;
	wire [4-1:0] node25940;
	wire [4-1:0] node25943;
	wire [4-1:0] node25945;
	wire [4-1:0] node25947;
	wire [4-1:0] node25950;
	wire [4-1:0] node25951;
	wire [4-1:0] node25952;
	wire [4-1:0] node25953;
	wire [4-1:0] node25954;
	wire [4-1:0] node25956;
	wire [4-1:0] node25959;
	wire [4-1:0] node25960;
	wire [4-1:0] node25964;
	wire [4-1:0] node25965;
	wire [4-1:0] node25966;
	wire [4-1:0] node25969;
	wire [4-1:0] node25972;
	wire [4-1:0] node25973;
	wire [4-1:0] node25976;
	wire [4-1:0] node25979;
	wire [4-1:0] node25980;
	wire [4-1:0] node25981;
	wire [4-1:0] node25982;
	wire [4-1:0] node25986;
	wire [4-1:0] node25988;
	wire [4-1:0] node25991;
	wire [4-1:0] node25992;
	wire [4-1:0] node25993;
	wire [4-1:0] node25996;
	wire [4-1:0] node26000;
	wire [4-1:0] node26001;
	wire [4-1:0] node26002;
	wire [4-1:0] node26004;
	wire [4-1:0] node26005;
	wire [4-1:0] node26008;
	wire [4-1:0] node26011;
	wire [4-1:0] node26012;
	wire [4-1:0] node26013;
	wire [4-1:0] node26017;
	wire [4-1:0] node26019;
	wire [4-1:0] node26022;
	wire [4-1:0] node26023;
	wire [4-1:0] node26024;
	wire [4-1:0] node26025;
	wire [4-1:0] node26028;
	wire [4-1:0] node26029;
	wire [4-1:0] node26033;
	wire [4-1:0] node26035;
	wire [4-1:0] node26038;
	wire [4-1:0] node26039;
	wire [4-1:0] node26040;
	wire [4-1:0] node26043;
	wire [4-1:0] node26046;
	wire [4-1:0] node26047;
	wire [4-1:0] node26051;
	wire [4-1:0] node26052;
	wire [4-1:0] node26053;
	wire [4-1:0] node26054;
	wire [4-1:0] node26055;
	wire [4-1:0] node26056;
	wire [4-1:0] node26057;
	wire [4-1:0] node26058;
	wire [4-1:0] node26060;
	wire [4-1:0] node26063;
	wire [4-1:0] node26065;
	wire [4-1:0] node26068;
	wire [4-1:0] node26069;
	wire [4-1:0] node26072;
	wire [4-1:0] node26075;
	wire [4-1:0] node26076;
	wire [4-1:0] node26077;
	wire [4-1:0] node26080;
	wire [4-1:0] node26083;
	wire [4-1:0] node26084;
	wire [4-1:0] node26085;
	wire [4-1:0] node26088;
	wire [4-1:0] node26091;
	wire [4-1:0] node26092;
	wire [4-1:0] node26093;
	wire [4-1:0] node26097;
	wire [4-1:0] node26099;
	wire [4-1:0] node26101;
	wire [4-1:0] node26104;
	wire [4-1:0] node26105;
	wire [4-1:0] node26106;
	wire [4-1:0] node26107;
	wire [4-1:0] node26108;
	wire [4-1:0] node26111;
	wire [4-1:0] node26114;
	wire [4-1:0] node26116;
	wire [4-1:0] node26119;
	wire [4-1:0] node26120;
	wire [4-1:0] node26121;
	wire [4-1:0] node26123;
	wire [4-1:0] node26124;
	wire [4-1:0] node26127;
	wire [4-1:0] node26130;
	wire [4-1:0] node26131;
	wire [4-1:0] node26132;
	wire [4-1:0] node26135;
	wire [4-1:0] node26139;
	wire [4-1:0] node26141;
	wire [4-1:0] node26144;
	wire [4-1:0] node26145;
	wire [4-1:0] node26146;
	wire [4-1:0] node26147;
	wire [4-1:0] node26148;
	wire [4-1:0] node26152;
	wire [4-1:0] node26153;
	wire [4-1:0] node26154;
	wire [4-1:0] node26157;
	wire [4-1:0] node26161;
	wire [4-1:0] node26162;
	wire [4-1:0] node26164;
	wire [4-1:0] node26167;
	wire [4-1:0] node26170;
	wire [4-1:0] node26171;
	wire [4-1:0] node26174;
	wire [4-1:0] node26177;
	wire [4-1:0] node26178;
	wire [4-1:0] node26179;
	wire [4-1:0] node26180;
	wire [4-1:0] node26181;
	wire [4-1:0] node26184;
	wire [4-1:0] node26186;
	wire [4-1:0] node26189;
	wire [4-1:0] node26190;
	wire [4-1:0] node26191;
	wire [4-1:0] node26192;
	wire [4-1:0] node26195;
	wire [4-1:0] node26199;
	wire [4-1:0] node26200;
	wire [4-1:0] node26203;
	wire [4-1:0] node26206;
	wire [4-1:0] node26207;
	wire [4-1:0] node26208;
	wire [4-1:0] node26209;
	wire [4-1:0] node26211;
	wire [4-1:0] node26212;
	wire [4-1:0] node26216;
	wire [4-1:0] node26218;
	wire [4-1:0] node26221;
	wire [4-1:0] node26222;
	wire [4-1:0] node26225;
	wire [4-1:0] node26228;
	wire [4-1:0] node26229;
	wire [4-1:0] node26230;
	wire [4-1:0] node26234;
	wire [4-1:0] node26236;
	wire [4-1:0] node26239;
	wire [4-1:0] node26240;
	wire [4-1:0] node26241;
	wire [4-1:0] node26242;
	wire [4-1:0] node26243;
	wire [4-1:0] node26244;
	wire [4-1:0] node26248;
	wire [4-1:0] node26250;
	wire [4-1:0] node26253;
	wire [4-1:0] node26254;
	wire [4-1:0] node26255;
	wire [4-1:0] node26256;
	wire [4-1:0] node26260;
	wire [4-1:0] node26261;
	wire [4-1:0] node26264;
	wire [4-1:0] node26267;
	wire [4-1:0] node26270;
	wire [4-1:0] node26271;
	wire [4-1:0] node26272;
	wire [4-1:0] node26275;
	wire [4-1:0] node26276;
	wire [4-1:0] node26279;
	wire [4-1:0] node26282;
	wire [4-1:0] node26283;
	wire [4-1:0] node26284;
	wire [4-1:0] node26286;
	wire [4-1:0] node26290;
	wire [4-1:0] node26291;
	wire [4-1:0] node26293;
	wire [4-1:0] node26296;
	wire [4-1:0] node26299;
	wire [4-1:0] node26300;
	wire [4-1:0] node26301;
	wire [4-1:0] node26302;
	wire [4-1:0] node26303;
	wire [4-1:0] node26306;
	wire [4-1:0] node26309;
	wire [4-1:0] node26311;
	wire [4-1:0] node26314;
	wire [4-1:0] node26316;
	wire [4-1:0] node26318;
	wire [4-1:0] node26321;
	wire [4-1:0] node26322;
	wire [4-1:0] node26323;
	wire [4-1:0] node26324;
	wire [4-1:0] node26327;
	wire [4-1:0] node26328;
	wire [4-1:0] node26333;
	wire [4-1:0] node26334;
	wire [4-1:0] node26336;
	wire [4-1:0] node26337;
	wire [4-1:0] node26341;
	wire [4-1:0] node26342;
	wire [4-1:0] node26345;
	wire [4-1:0] node26348;
	wire [4-1:0] node26349;
	wire [4-1:0] node26350;
	wire [4-1:0] node26351;
	wire [4-1:0] node26352;
	wire [4-1:0] node26353;
	wire [4-1:0] node26354;
	wire [4-1:0] node26356;
	wire [4-1:0] node26359;
	wire [4-1:0] node26360;
	wire [4-1:0] node26361;
	wire [4-1:0] node26365;
	wire [4-1:0] node26366;
	wire [4-1:0] node26369;
	wire [4-1:0] node26372;
	wire [4-1:0] node26373;
	wire [4-1:0] node26377;
	wire [4-1:0] node26378;
	wire [4-1:0] node26379;
	wire [4-1:0] node26380;
	wire [4-1:0] node26381;
	wire [4-1:0] node26384;
	wire [4-1:0] node26388;
	wire [4-1:0] node26390;
	wire [4-1:0] node26391;
	wire [4-1:0] node26394;
	wire [4-1:0] node26397;
	wire [4-1:0] node26398;
	wire [4-1:0] node26400;
	wire [4-1:0] node26403;
	wire [4-1:0] node26404;
	wire [4-1:0] node26407;
	wire [4-1:0] node26410;
	wire [4-1:0] node26411;
	wire [4-1:0] node26412;
	wire [4-1:0] node26413;
	wire [4-1:0] node26414;
	wire [4-1:0] node26415;
	wire [4-1:0] node26419;
	wire [4-1:0] node26423;
	wire [4-1:0] node26425;
	wire [4-1:0] node26428;
	wire [4-1:0] node26429;
	wire [4-1:0] node26430;
	wire [4-1:0] node26433;
	wire [4-1:0] node26436;
	wire [4-1:0] node26438;
	wire [4-1:0] node26441;
	wire [4-1:0] node26442;
	wire [4-1:0] node26443;
	wire [4-1:0] node26444;
	wire [4-1:0] node26445;
	wire [4-1:0] node26448;
	wire [4-1:0] node26451;
	wire [4-1:0] node26453;
	wire [4-1:0] node26454;
	wire [4-1:0] node26457;
	wire [4-1:0] node26460;
	wire [4-1:0] node26461;
	wire [4-1:0] node26462;
	wire [4-1:0] node26463;
	wire [4-1:0] node26467;
	wire [4-1:0] node26468;
	wire [4-1:0] node26472;
	wire [4-1:0] node26473;
	wire [4-1:0] node26477;
	wire [4-1:0] node26478;
	wire [4-1:0] node26479;
	wire [4-1:0] node26481;
	wire [4-1:0] node26482;
	wire [4-1:0] node26485;
	wire [4-1:0] node26488;
	wire [4-1:0] node26490;
	wire [4-1:0] node26492;
	wire [4-1:0] node26495;
	wire [4-1:0] node26496;
	wire [4-1:0] node26497;
	wire [4-1:0] node26498;
	wire [4-1:0] node26501;
	wire [4-1:0] node26504;
	wire [4-1:0] node26505;
	wire [4-1:0] node26509;
	wire [4-1:0] node26510;
	wire [4-1:0] node26511;
	wire [4-1:0] node26512;
	wire [4-1:0] node26516;
	wire [4-1:0] node26517;
	wire [4-1:0] node26521;
	wire [4-1:0] node26523;
	wire [4-1:0] node26524;
	wire [4-1:0] node26527;
	wire [4-1:0] node26530;
	wire [4-1:0] node26531;
	wire [4-1:0] node26532;
	wire [4-1:0] node26533;
	wire [4-1:0] node26534;
	wire [4-1:0] node26535;
	wire [4-1:0] node26536;
	wire [4-1:0] node26540;
	wire [4-1:0] node26541;
	wire [4-1:0] node26545;
	wire [4-1:0] node26546;
	wire [4-1:0] node26547;
	wire [4-1:0] node26548;
	wire [4-1:0] node26554;
	wire [4-1:0] node26555;
	wire [4-1:0] node26556;
	wire [4-1:0] node26560;
	wire [4-1:0] node26561;
	wire [4-1:0] node26562;
	wire [4-1:0] node26565;
	wire [4-1:0] node26568;
	wire [4-1:0] node26570;
	wire [4-1:0] node26573;
	wire [4-1:0] node26574;
	wire [4-1:0] node26575;
	wire [4-1:0] node26577;
	wire [4-1:0] node26580;
	wire [4-1:0] node26582;
	wire [4-1:0] node26585;
	wire [4-1:0] node26587;
	wire [4-1:0] node26590;
	wire [4-1:0] node26591;
	wire [4-1:0] node26592;
	wire [4-1:0] node26595;
	wire [4-1:0] node26598;
	wire [4-1:0] node26599;
	wire [4-1:0] node26600;
	wire [4-1:0] node26601;
	wire [4-1:0] node26604;
	wire [4-1:0] node26608;
	wire [4-1:0] node26610;
	wire [4-1:0] node26611;
	wire [4-1:0] node26612;
	wire [4-1:0] node26615;
	wire [4-1:0] node26618;
	wire [4-1:0] node26621;
	wire [4-1:0] node26622;
	wire [4-1:0] node26623;
	wire [4-1:0] node26624;
	wire [4-1:0] node26625;
	wire [4-1:0] node26626;
	wire [4-1:0] node26627;
	wire [4-1:0] node26628;
	wire [4-1:0] node26630;
	wire [4-1:0] node26631;
	wire [4-1:0] node26634;
	wire [4-1:0] node26637;
	wire [4-1:0] node26638;
	wire [4-1:0] node26640;
	wire [4-1:0] node26643;
	wire [4-1:0] node26645;
	wire [4-1:0] node26648;
	wire [4-1:0] node26649;
	wire [4-1:0] node26650;
	wire [4-1:0] node26652;
	wire [4-1:0] node26657;
	wire [4-1:0] node26658;
	wire [4-1:0] node26659;
	wire [4-1:0] node26660;
	wire [4-1:0] node26662;
	wire [4-1:0] node26665;
	wire [4-1:0] node26668;
	wire [4-1:0] node26670;
	wire [4-1:0] node26673;
	wire [4-1:0] node26675;
	wire [4-1:0] node26676;
	wire [4-1:0] node26680;
	wire [4-1:0] node26681;
	wire [4-1:0] node26682;
	wire [4-1:0] node26684;
	wire [4-1:0] node26686;
	wire [4-1:0] node26687;
	wire [4-1:0] node26691;
	wire [4-1:0] node26692;
	wire [4-1:0] node26693;
	wire [4-1:0] node26696;
	wire [4-1:0] node26699;
	wire [4-1:0] node26701;
	wire [4-1:0] node26704;
	wire [4-1:0] node26705;
	wire [4-1:0] node26706;
	wire [4-1:0] node26707;
	wire [4-1:0] node26710;
	wire [4-1:0] node26714;
	wire [4-1:0] node26715;
	wire [4-1:0] node26717;
	wire [4-1:0] node26718;
	wire [4-1:0] node26721;
	wire [4-1:0] node26724;
	wire [4-1:0] node26725;
	wire [4-1:0] node26726;
	wire [4-1:0] node26731;
	wire [4-1:0] node26732;
	wire [4-1:0] node26733;
	wire [4-1:0] node26734;
	wire [4-1:0] node26735;
	wire [4-1:0] node26738;
	wire [4-1:0] node26739;
	wire [4-1:0] node26741;
	wire [4-1:0] node26745;
	wire [4-1:0] node26746;
	wire [4-1:0] node26748;
	wire [4-1:0] node26751;
	wire [4-1:0] node26754;
	wire [4-1:0] node26755;
	wire [4-1:0] node26757;
	wire [4-1:0] node26759;
	wire [4-1:0] node26762;
	wire [4-1:0] node26763;
	wire [4-1:0] node26766;
	wire [4-1:0] node26767;
	wire [4-1:0] node26771;
	wire [4-1:0] node26772;
	wire [4-1:0] node26773;
	wire [4-1:0] node26775;
	wire [4-1:0] node26777;
	wire [4-1:0] node26780;
	wire [4-1:0] node26781;
	wire [4-1:0] node26783;
	wire [4-1:0] node26787;
	wire [4-1:0] node26788;
	wire [4-1:0] node26789;
	wire [4-1:0] node26790;
	wire [4-1:0] node26793;
	wire [4-1:0] node26797;
	wire [4-1:0] node26798;
	wire [4-1:0] node26800;
	wire [4-1:0] node26801;
	wire [4-1:0] node26804;
	wire [4-1:0] node26808;
	wire [4-1:0] node26809;
	wire [4-1:0] node26810;
	wire [4-1:0] node26811;
	wire [4-1:0] node26812;
	wire [4-1:0] node26814;
	wire [4-1:0] node26817;
	wire [4-1:0] node26819;
	wire [4-1:0] node26822;
	wire [4-1:0] node26823;
	wire [4-1:0] node26825;
	wire [4-1:0] node26828;
	wire [4-1:0] node26830;
	wire [4-1:0] node26833;
	wire [4-1:0] node26834;
	wire [4-1:0] node26835;
	wire [4-1:0] node26837;
	wire [4-1:0] node26840;
	wire [4-1:0] node26841;
	wire [4-1:0] node26843;
	wire [4-1:0] node26846;
	wire [4-1:0] node26848;
	wire [4-1:0] node26851;
	wire [4-1:0] node26852;
	wire [4-1:0] node26853;
	wire [4-1:0] node26854;
	wire [4-1:0] node26859;
	wire [4-1:0] node26860;
	wire [4-1:0] node26861;
	wire [4-1:0] node26866;
	wire [4-1:0] node26867;
	wire [4-1:0] node26868;
	wire [4-1:0] node26869;
	wire [4-1:0] node26871;
	wire [4-1:0] node26872;
	wire [4-1:0] node26873;
	wire [4-1:0] node26876;
	wire [4-1:0] node26880;
	wire [4-1:0] node26881;
	wire [4-1:0] node26884;
	wire [4-1:0] node26887;
	wire [4-1:0] node26888;
	wire [4-1:0] node26889;
	wire [4-1:0] node26892;
	wire [4-1:0] node26895;
	wire [4-1:0] node26897;
	wire [4-1:0] node26900;
	wire [4-1:0] node26901;
	wire [4-1:0] node26902;
	wire [4-1:0] node26903;
	wire [4-1:0] node26907;
	wire [4-1:0] node26908;
	wire [4-1:0] node26910;
	wire [4-1:0] node26913;
	wire [4-1:0] node26915;
	wire [4-1:0] node26916;
	wire [4-1:0] node26919;
	wire [4-1:0] node26922;
	wire [4-1:0] node26923;
	wire [4-1:0] node26924;
	wire [4-1:0] node26925;
	wire [4-1:0] node26927;
	wire [4-1:0] node26931;
	wire [4-1:0] node26932;
	wire [4-1:0] node26936;
	wire [4-1:0] node26937;
	wire [4-1:0] node26938;
	wire [4-1:0] node26939;
	wire [4-1:0] node26942;
	wire [4-1:0] node26947;
	wire [4-1:0] node26948;
	wire [4-1:0] node26949;
	wire [4-1:0] node26950;
	wire [4-1:0] node26951;
	wire [4-1:0] node26952;
	wire [4-1:0] node26953;
	wire [4-1:0] node26954;
	wire [4-1:0] node26959;
	wire [4-1:0] node26960;
	wire [4-1:0] node26961;
	wire [4-1:0] node26965;
	wire [4-1:0] node26968;
	wire [4-1:0] node26969;
	wire [4-1:0] node26970;
	wire [4-1:0] node26971;
	wire [4-1:0] node26975;
	wire [4-1:0] node26978;
	wire [4-1:0] node26980;
	wire [4-1:0] node26983;
	wire [4-1:0] node26984;
	wire [4-1:0] node26985;
	wire [4-1:0] node26988;
	wire [4-1:0] node26991;
	wire [4-1:0] node26992;
	wire [4-1:0] node26993;
	wire [4-1:0] node26997;
	wire [4-1:0] node26998;
	wire [4-1:0] node27002;
	wire [4-1:0] node27003;
	wire [4-1:0] node27004;
	wire [4-1:0] node27005;
	wire [4-1:0] node27006;
	wire [4-1:0] node27008;
	wire [4-1:0] node27012;
	wire [4-1:0] node27013;
	wire [4-1:0] node27017;
	wire [4-1:0] node27018;
	wire [4-1:0] node27019;
	wire [4-1:0] node27020;
	wire [4-1:0] node27024;
	wire [4-1:0] node27027;
	wire [4-1:0] node27028;
	wire [4-1:0] node27029;
	wire [4-1:0] node27034;
	wire [4-1:0] node27035;
	wire [4-1:0] node27036;
	wire [4-1:0] node27037;
	wire [4-1:0] node27038;
	wire [4-1:0] node27043;
	wire [4-1:0] node27044;
	wire [4-1:0] node27046;
	wire [4-1:0] node27049;
	wire [4-1:0] node27050;
	wire [4-1:0] node27053;
	wire [4-1:0] node27056;
	wire [4-1:0] node27057;
	wire [4-1:0] node27059;
	wire [4-1:0] node27060;
	wire [4-1:0] node27061;
	wire [4-1:0] node27066;
	wire [4-1:0] node27067;
	wire [4-1:0] node27068;
	wire [4-1:0] node27071;
	wire [4-1:0] node27072;
	wire [4-1:0] node27076;
	wire [4-1:0] node27077;
	wire [4-1:0] node27080;
	wire [4-1:0] node27081;
	wire [4-1:0] node27085;
	wire [4-1:0] node27086;
	wire [4-1:0] node27087;
	wire [4-1:0] node27088;
	wire [4-1:0] node27089;
	wire [4-1:0] node27090;
	wire [4-1:0] node27092;
	wire [4-1:0] node27095;
	wire [4-1:0] node27097;
	wire [4-1:0] node27100;
	wire [4-1:0] node27101;
	wire [4-1:0] node27105;
	wire [4-1:0] node27106;
	wire [4-1:0] node27108;
	wire [4-1:0] node27111;
	wire [4-1:0] node27113;
	wire [4-1:0] node27116;
	wire [4-1:0] node27117;
	wire [4-1:0] node27118;
	wire [4-1:0] node27120;
	wire [4-1:0] node27121;
	wire [4-1:0] node27125;
	wire [4-1:0] node27126;
	wire [4-1:0] node27130;
	wire [4-1:0] node27131;
	wire [4-1:0] node27133;
	wire [4-1:0] node27134;
	wire [4-1:0] node27138;
	wire [4-1:0] node27139;
	wire [4-1:0] node27143;
	wire [4-1:0] node27144;
	wire [4-1:0] node27145;
	wire [4-1:0] node27146;
	wire [4-1:0] node27148;
	wire [4-1:0] node27150;
	wire [4-1:0] node27152;
	wire [4-1:0] node27155;
	wire [4-1:0] node27156;
	wire [4-1:0] node27157;
	wire [4-1:0] node27162;
	wire [4-1:0] node27163;
	wire [4-1:0] node27164;
	wire [4-1:0] node27168;
	wire [4-1:0] node27169;
	wire [4-1:0] node27173;
	wire [4-1:0] node27174;
	wire [4-1:0] node27175;
	wire [4-1:0] node27177;
	wire [4-1:0] node27181;
	wire [4-1:0] node27182;
	wire [4-1:0] node27183;
	wire [4-1:0] node27184;
	wire [4-1:0] node27188;
	wire [4-1:0] node27189;
	wire [4-1:0] node27193;
	wire [4-1:0] node27194;
	wire [4-1:0] node27198;
	wire [4-1:0] node27199;
	wire [4-1:0] node27200;
	wire [4-1:0] node27201;
	wire [4-1:0] node27202;
	wire [4-1:0] node27203;
	wire [4-1:0] node27204;
	wire [4-1:0] node27205;
	wire [4-1:0] node27207;
	wire [4-1:0] node27210;
	wire [4-1:0] node27212;
	wire [4-1:0] node27215;
	wire [4-1:0] node27216;
	wire [4-1:0] node27218;
	wire [4-1:0] node27221;
	wire [4-1:0] node27223;
	wire [4-1:0] node27226;
	wire [4-1:0] node27227;
	wire [4-1:0] node27228;
	wire [4-1:0] node27229;
	wire [4-1:0] node27231;
	wire [4-1:0] node27234;
	wire [4-1:0] node27236;
	wire [4-1:0] node27239;
	wire [4-1:0] node27240;
	wire [4-1:0] node27242;
	wire [4-1:0] node27245;
	wire [4-1:0] node27248;
	wire [4-1:0] node27249;
	wire [4-1:0] node27250;
	wire [4-1:0] node27251;
	wire [4-1:0] node27252;
	wire [4-1:0] node27256;
	wire [4-1:0] node27257;
	wire [4-1:0] node27261;
	wire [4-1:0] node27262;
	wire [4-1:0] node27263;
	wire [4-1:0] node27264;
	wire [4-1:0] node27267;
	wire [4-1:0] node27272;
	wire [4-1:0] node27273;
	wire [4-1:0] node27275;
	wire [4-1:0] node27278;
	wire [4-1:0] node27279;
	wire [4-1:0] node27282;
	wire [4-1:0] node27283;
	wire [4-1:0] node27287;
	wire [4-1:0] node27288;
	wire [4-1:0] node27289;
	wire [4-1:0] node27290;
	wire [4-1:0] node27292;
	wire [4-1:0] node27295;
	wire [4-1:0] node27297;
	wire [4-1:0] node27300;
	wire [4-1:0] node27301;
	wire [4-1:0] node27303;
	wire [4-1:0] node27306;
	wire [4-1:0] node27308;
	wire [4-1:0] node27311;
	wire [4-1:0] node27312;
	wire [4-1:0] node27313;
	wire [4-1:0] node27314;
	wire [4-1:0] node27316;
	wire [4-1:0] node27317;
	wire [4-1:0] node27319;
	wire [4-1:0] node27323;
	wire [4-1:0] node27325;
	wire [4-1:0] node27328;
	wire [4-1:0] node27329;
	wire [4-1:0] node27331;
	wire [4-1:0] node27332;
	wire [4-1:0] node27333;
	wire [4-1:0] node27337;
	wire [4-1:0] node27338;
	wire [4-1:0] node27342;
	wire [4-1:0] node27343;
	wire [4-1:0] node27344;
	wire [4-1:0] node27347;
	wire [4-1:0] node27348;
	wire [4-1:0] node27352;
	wire [4-1:0] node27353;
	wire [4-1:0] node27357;
	wire [4-1:0] node27358;
	wire [4-1:0] node27359;
	wire [4-1:0] node27360;
	wire [4-1:0] node27363;
	wire [4-1:0] node27366;
	wire [4-1:0] node27368;
	wire [4-1:0] node27369;
	wire [4-1:0] node27372;
	wire [4-1:0] node27375;
	wire [4-1:0] node27376;
	wire [4-1:0] node27378;
	wire [4-1:0] node27380;
	wire [4-1:0] node27383;
	wire [4-1:0] node27384;
	wire [4-1:0] node27385;
	wire [4-1:0] node27388;
	wire [4-1:0] node27392;
	wire [4-1:0] node27393;
	wire [4-1:0] node27394;
	wire [4-1:0] node27395;
	wire [4-1:0] node27396;
	wire [4-1:0] node27397;
	wire [4-1:0] node27400;
	wire [4-1:0] node27401;
	wire [4-1:0] node27405;
	wire [4-1:0] node27406;
	wire [4-1:0] node27409;
	wire [4-1:0] node27411;
	wire [4-1:0] node27414;
	wire [4-1:0] node27415;
	wire [4-1:0] node27416;
	wire [4-1:0] node27417;
	wire [4-1:0] node27419;
	wire [4-1:0] node27423;
	wire [4-1:0] node27425;
	wire [4-1:0] node27428;
	wire [4-1:0] node27429;
	wire [4-1:0] node27430;
	wire [4-1:0] node27432;
	wire [4-1:0] node27435;
	wire [4-1:0] node27438;
	wire [4-1:0] node27439;
	wire [4-1:0] node27443;
	wire [4-1:0] node27444;
	wire [4-1:0] node27445;
	wire [4-1:0] node27447;
	wire [4-1:0] node27450;
	wire [4-1:0] node27451;
	wire [4-1:0] node27453;
	wire [4-1:0] node27456;
	wire [4-1:0] node27458;
	wire [4-1:0] node27461;
	wire [4-1:0] node27462;
	wire [4-1:0] node27463;
	wire [4-1:0] node27464;
	wire [4-1:0] node27468;
	wire [4-1:0] node27469;
	wire [4-1:0] node27473;
	wire [4-1:0] node27474;
	wire [4-1:0] node27475;
	wire [4-1:0] node27479;
	wire [4-1:0] node27482;
	wire [4-1:0] node27483;
	wire [4-1:0] node27484;
	wire [4-1:0] node27485;
	wire [4-1:0] node27486;
	wire [4-1:0] node27490;
	wire [4-1:0] node27491;
	wire [4-1:0] node27495;
	wire [4-1:0] node27496;
	wire [4-1:0] node27497;
	wire [4-1:0] node27501;
	wire [4-1:0] node27502;
	wire [4-1:0] node27506;
	wire [4-1:0] node27507;
	wire [4-1:0] node27508;
	wire [4-1:0] node27509;
	wire [4-1:0] node27511;
	wire [4-1:0] node27512;
	wire [4-1:0] node27515;
	wire [4-1:0] node27518;
	wire [4-1:0] node27520;
	wire [4-1:0] node27523;
	wire [4-1:0] node27524;
	wire [4-1:0] node27525;
	wire [4-1:0] node27528;
	wire [4-1:0] node27531;
	wire [4-1:0] node27533;
	wire [4-1:0] node27534;
	wire [4-1:0] node27535;
	wire [4-1:0] node27538;
	wire [4-1:0] node27542;
	wire [4-1:0] node27543;
	wire [4-1:0] node27544;
	wire [4-1:0] node27545;
	wire [4-1:0] node27547;
	wire [4-1:0] node27550;
	wire [4-1:0] node27551;
	wire [4-1:0] node27552;
	wire [4-1:0] node27556;
	wire [4-1:0] node27558;
	wire [4-1:0] node27561;
	wire [4-1:0] node27562;
	wire [4-1:0] node27566;
	wire [4-1:0] node27567;
	wire [4-1:0] node27568;
	wire [4-1:0] node27571;
	wire [4-1:0] node27572;
	wire [4-1:0] node27575;
	wire [4-1:0] node27576;
	wire [4-1:0] node27581;
	wire [4-1:0] node27582;
	wire [4-1:0] node27583;
	wire [4-1:0] node27584;
	wire [4-1:0] node27585;
	wire [4-1:0] node27586;
	wire [4-1:0] node27587;
	wire [4-1:0] node27588;
	wire [4-1:0] node27591;
	wire [4-1:0] node27594;
	wire [4-1:0] node27596;
	wire [4-1:0] node27599;
	wire [4-1:0] node27600;
	wire [4-1:0] node27601;
	wire [4-1:0] node27603;
	wire [4-1:0] node27606;
	wire [4-1:0] node27608;
	wire [4-1:0] node27611;
	wire [4-1:0] node27612;
	wire [4-1:0] node27615;
	wire [4-1:0] node27617;
	wire [4-1:0] node27620;
	wire [4-1:0] node27621;
	wire [4-1:0] node27622;
	wire [4-1:0] node27623;
	wire [4-1:0] node27624;
	wire [4-1:0] node27627;
	wire [4-1:0] node27631;
	wire [4-1:0] node27632;
	wire [4-1:0] node27633;
	wire [4-1:0] node27634;
	wire [4-1:0] node27638;
	wire [4-1:0] node27641;
	wire [4-1:0] node27643;
	wire [4-1:0] node27644;
	wire [4-1:0] node27647;
	wire [4-1:0] node27650;
	wire [4-1:0] node27651;
	wire [4-1:0] node27654;
	wire [4-1:0] node27655;
	wire [4-1:0] node27657;
	wire [4-1:0] node27660;
	wire [4-1:0] node27662;
	wire [4-1:0] node27665;
	wire [4-1:0] node27666;
	wire [4-1:0] node27667;
	wire [4-1:0] node27668;
	wire [4-1:0] node27669;
	wire [4-1:0] node27673;
	wire [4-1:0] node27674;
	wire [4-1:0] node27675;
	wire [4-1:0] node27680;
	wire [4-1:0] node27681;
	wire [4-1:0] node27682;
	wire [4-1:0] node27685;
	wire [4-1:0] node27688;
	wire [4-1:0] node27690;
	wire [4-1:0] node27692;
	wire [4-1:0] node27694;
	wire [4-1:0] node27697;
	wire [4-1:0] node27698;
	wire [4-1:0] node27700;
	wire [4-1:0] node27701;
	wire [4-1:0] node27702;
	wire [4-1:0] node27704;
	wire [4-1:0] node27708;
	wire [4-1:0] node27710;
	wire [4-1:0] node27711;
	wire [4-1:0] node27714;
	wire [4-1:0] node27717;
	wire [4-1:0] node27718;
	wire [4-1:0] node27719;
	wire [4-1:0] node27722;
	wire [4-1:0] node27724;
	wire [4-1:0] node27728;
	wire [4-1:0] node27729;
	wire [4-1:0] node27730;
	wire [4-1:0] node27731;
	wire [4-1:0] node27732;
	wire [4-1:0] node27733;
	wire [4-1:0] node27736;
	wire [4-1:0] node27739;
	wire [4-1:0] node27741;
	wire [4-1:0] node27744;
	wire [4-1:0] node27745;
	wire [4-1:0] node27746;
	wire [4-1:0] node27749;
	wire [4-1:0] node27752;
	wire [4-1:0] node27754;
	wire [4-1:0] node27755;
	wire [4-1:0] node27759;
	wire [4-1:0] node27760;
	wire [4-1:0] node27761;
	wire [4-1:0] node27762;
	wire [4-1:0] node27765;
	wire [4-1:0] node27768;
	wire [4-1:0] node27769;
	wire [4-1:0] node27772;
	wire [4-1:0] node27775;
	wire [4-1:0] node27776;
	wire [4-1:0] node27777;
	wire [4-1:0] node27779;
	wire [4-1:0] node27782;
	wire [4-1:0] node27783;
	wire [4-1:0] node27787;
	wire [4-1:0] node27790;
	wire [4-1:0] node27791;
	wire [4-1:0] node27792;
	wire [4-1:0] node27793;
	wire [4-1:0] node27794;
	wire [4-1:0] node27795;
	wire [4-1:0] node27799;
	wire [4-1:0] node27800;
	wire [4-1:0] node27802;
	wire [4-1:0] node27805;
	wire [4-1:0] node27807;
	wire [4-1:0] node27811;
	wire [4-1:0] node27812;
	wire [4-1:0] node27814;
	wire [4-1:0] node27815;
	wire [4-1:0] node27818;
	wire [4-1:0] node27819;
	wire [4-1:0] node27823;
	wire [4-1:0] node27824;
	wire [4-1:0] node27828;
	wire [4-1:0] node27829;
	wire [4-1:0] node27830;
	wire [4-1:0] node27831;
	wire [4-1:0] node27835;
	wire [4-1:0] node27836;
	wire [4-1:0] node27837;
	wire [4-1:0] node27841;
	wire [4-1:0] node27844;
	wire [4-1:0] node27845;
	wire [4-1:0] node27846;
	wire [4-1:0] node27847;
	wire [4-1:0] node27852;
	wire [4-1:0] node27853;
	wire [4-1:0] node27854;
	wire [4-1:0] node27858;
	wire [4-1:0] node27861;
	wire [4-1:0] node27862;
	wire [4-1:0] node27863;
	wire [4-1:0] node27864;
	wire [4-1:0] node27865;
	wire [4-1:0] node27866;
	wire [4-1:0] node27867;
	wire [4-1:0] node27868;
	wire [4-1:0] node27873;
	wire [4-1:0] node27874;
	wire [4-1:0] node27877;
	wire [4-1:0] node27878;
	wire [4-1:0] node27880;
	wire [4-1:0] node27883;
	wire [4-1:0] node27884;
	wire [4-1:0] node27888;
	wire [4-1:0] node27889;
	wire [4-1:0] node27890;
	wire [4-1:0] node27892;
	wire [4-1:0] node27895;
	wire [4-1:0] node27896;
	wire [4-1:0] node27897;
	wire [4-1:0] node27900;
	wire [4-1:0] node27904;
	wire [4-1:0] node27906;
	wire [4-1:0] node27908;
	wire [4-1:0] node27910;
	wire [4-1:0] node27913;
	wire [4-1:0] node27914;
	wire [4-1:0] node27915;
	wire [4-1:0] node27917;
	wire [4-1:0] node27920;
	wire [4-1:0] node27922;
	wire [4-1:0] node27925;
	wire [4-1:0] node27927;
	wire [4-1:0] node27928;
	wire [4-1:0] node27931;
	wire [4-1:0] node27934;
	wire [4-1:0] node27935;
	wire [4-1:0] node27936;
	wire [4-1:0] node27937;
	wire [4-1:0] node27938;
	wire [4-1:0] node27941;
	wire [4-1:0] node27944;
	wire [4-1:0] node27946;
	wire [4-1:0] node27949;
	wire [4-1:0] node27950;
	wire [4-1:0] node27951;
	wire [4-1:0] node27952;
	wire [4-1:0] node27955;
	wire [4-1:0] node27958;
	wire [4-1:0] node27959;
	wire [4-1:0] node27963;
	wire [4-1:0] node27964;
	wire [4-1:0] node27965;
	wire [4-1:0] node27968;
	wire [4-1:0] node27971;
	wire [4-1:0] node27972;
	wire [4-1:0] node27973;
	wire [4-1:0] node27977;
	wire [4-1:0] node27979;
	wire [4-1:0] node27982;
	wire [4-1:0] node27983;
	wire [4-1:0] node27985;
	wire [4-1:0] node27986;
	wire [4-1:0] node27987;
	wire [4-1:0] node27991;
	wire [4-1:0] node27992;
	wire [4-1:0] node27996;
	wire [4-1:0] node27997;
	wire [4-1:0] node27998;
	wire [4-1:0] node27999;
	wire [4-1:0] node28002;
	wire [4-1:0] node28006;
	wire [4-1:0] node28007;
	wire [4-1:0] node28008;
	wire [4-1:0] node28012;
	wire [4-1:0] node28015;
	wire [4-1:0] node28016;
	wire [4-1:0] node28017;
	wire [4-1:0] node28018;
	wire [4-1:0] node28019;
	wire [4-1:0] node28020;
	wire [4-1:0] node28023;
	wire [4-1:0] node28026;
	wire [4-1:0] node28027;
	wire [4-1:0] node28029;
	wire [4-1:0] node28030;
	wire [4-1:0] node28035;
	wire [4-1:0] node28036;
	wire [4-1:0] node28038;
	wire [4-1:0] node28039;
	wire [4-1:0] node28042;
	wire [4-1:0] node28045;
	wire [4-1:0] node28047;
	wire [4-1:0] node28048;
	wire [4-1:0] node28051;
	wire [4-1:0] node28054;
	wire [4-1:0] node28055;
	wire [4-1:0] node28056;
	wire [4-1:0] node28057;
	wire [4-1:0] node28061;
	wire [4-1:0] node28062;
	wire [4-1:0] node28066;
	wire [4-1:0] node28067;
	wire [4-1:0] node28068;
	wire [4-1:0] node28072;
	wire [4-1:0] node28073;
	wire [4-1:0] node28077;
	wire [4-1:0] node28078;
	wire [4-1:0] node28079;
	wire [4-1:0] node28080;
	wire [4-1:0] node28083;
	wire [4-1:0] node28084;
	wire [4-1:0] node28085;
	wire [4-1:0] node28089;
	wire [4-1:0] node28090;
	wire [4-1:0] node28094;
	wire [4-1:0] node28095;
	wire [4-1:0] node28096;
	wire [4-1:0] node28097;
	wire [4-1:0] node28101;
	wire [4-1:0] node28104;
	wire [4-1:0] node28105;
	wire [4-1:0] node28106;
	wire [4-1:0] node28107;
	wire [4-1:0] node28111;
	wire [4-1:0] node28115;
	wire [4-1:0] node28116;
	wire [4-1:0] node28117;
	wire [4-1:0] node28118;
	wire [4-1:0] node28122;
	wire [4-1:0] node28123;
	wire [4-1:0] node28127;
	wire [4-1:0] node28128;
	wire [4-1:0] node28129;
	wire [4-1:0] node28133;
	wire [4-1:0] node28134;
	wire [4-1:0] node28138;
	wire [4-1:0] node28139;
	wire [4-1:0] node28140;
	wire [4-1:0] node28141;
	wire [4-1:0] node28142;
	wire [4-1:0] node28143;
	wire [4-1:0] node28144;
	wire [4-1:0] node28145;
	wire [4-1:0] node28146;
	wire [4-1:0] node28147;
	wire [4-1:0] node28150;
	wire [4-1:0] node28153;
	wire [4-1:0] node28155;
	wire [4-1:0] node28156;
	wire [4-1:0] node28160;
	wire [4-1:0] node28161;
	wire [4-1:0] node28162;
	wire [4-1:0] node28166;
	wire [4-1:0] node28167;
	wire [4-1:0] node28168;
	wire [4-1:0] node28173;
	wire [4-1:0] node28174;
	wire [4-1:0] node28176;
	wire [4-1:0] node28179;
	wire [4-1:0] node28180;
	wire [4-1:0] node28182;
	wire [4-1:0] node28185;
	wire [4-1:0] node28186;
	wire [4-1:0] node28189;
	wire [4-1:0] node28192;
	wire [4-1:0] node28193;
	wire [4-1:0] node28194;
	wire [4-1:0] node28196;
	wire [4-1:0] node28199;
	wire [4-1:0] node28201;
	wire [4-1:0] node28202;
	wire [4-1:0] node28205;
	wire [4-1:0] node28208;
	wire [4-1:0] node28209;
	wire [4-1:0] node28210;
	wire [4-1:0] node28211;
	wire [4-1:0] node28214;
	wire [4-1:0] node28217;
	wire [4-1:0] node28219;
	wire [4-1:0] node28220;
	wire [4-1:0] node28223;
	wire [4-1:0] node28226;
	wire [4-1:0] node28228;
	wire [4-1:0] node28230;
	wire [4-1:0] node28231;
	wire [4-1:0] node28235;
	wire [4-1:0] node28236;
	wire [4-1:0] node28237;
	wire [4-1:0] node28238;
	wire [4-1:0] node28239;
	wire [4-1:0] node28240;
	wire [4-1:0] node28243;
	wire [4-1:0] node28247;
	wire [4-1:0] node28248;
	wire [4-1:0] node28249;
	wire [4-1:0] node28253;
	wire [4-1:0] node28255;
	wire [4-1:0] node28257;
	wire [4-1:0] node28260;
	wire [4-1:0] node28261;
	wire [4-1:0] node28262;
	wire [4-1:0] node28263;
	wire [4-1:0] node28266;
	wire [4-1:0] node28270;
	wire [4-1:0] node28272;
	wire [4-1:0] node28275;
	wire [4-1:0] node28276;
	wire [4-1:0] node28277;
	wire [4-1:0] node28279;
	wire [4-1:0] node28282;
	wire [4-1:0] node28284;
	wire [4-1:0] node28287;
	wire [4-1:0] node28288;
	wire [4-1:0] node28290;
	wire [4-1:0] node28293;
	wire [4-1:0] node28295;
	wire [4-1:0] node28298;
	wire [4-1:0] node28299;
	wire [4-1:0] node28300;
	wire [4-1:0] node28301;
	wire [4-1:0] node28302;
	wire [4-1:0] node28303;
	wire [4-1:0] node28307;
	wire [4-1:0] node28308;
	wire [4-1:0] node28311;
	wire [4-1:0] node28313;
	wire [4-1:0] node28316;
	wire [4-1:0] node28317;
	wire [4-1:0] node28318;
	wire [4-1:0] node28319;
	wire [4-1:0] node28322;
	wire [4-1:0] node28325;
	wire [4-1:0] node28326;
	wire [4-1:0] node28327;
	wire [4-1:0] node28330;
	wire [4-1:0] node28334;
	wire [4-1:0] node28335;
	wire [4-1:0] node28339;
	wire [4-1:0] node28340;
	wire [4-1:0] node28341;
	wire [4-1:0] node28342;
	wire [4-1:0] node28346;
	wire [4-1:0] node28347;
	wire [4-1:0] node28351;
	wire [4-1:0] node28352;
	wire [4-1:0] node28353;
	wire [4-1:0] node28357;
	wire [4-1:0] node28358;
	wire [4-1:0] node28362;
	wire [4-1:0] node28363;
	wire [4-1:0] node28364;
	wire [4-1:0] node28365;
	wire [4-1:0] node28366;
	wire [4-1:0] node28367;
	wire [4-1:0] node28370;
	wire [4-1:0] node28373;
	wire [4-1:0] node28374;
	wire [4-1:0] node28378;
	wire [4-1:0] node28379;
	wire [4-1:0] node28380;
	wire [4-1:0] node28384;
	wire [4-1:0] node28385;
	wire [4-1:0] node28386;
	wire [4-1:0] node28389;
	wire [4-1:0] node28392;
	wire [4-1:0] node28393;
	wire [4-1:0] node28396;
	wire [4-1:0] node28399;
	wire [4-1:0] node28400;
	wire [4-1:0] node28402;
	wire [4-1:0] node28403;
	wire [4-1:0] node28405;
	wire [4-1:0] node28408;
	wire [4-1:0] node28409;
	wire [4-1:0] node28413;
	wire [4-1:0] node28414;
	wire [4-1:0] node28416;
	wire [4-1:0] node28419;
	wire [4-1:0] node28420;
	wire [4-1:0] node28421;
	wire [4-1:0] node28426;
	wire [4-1:0] node28427;
	wire [4-1:0] node28428;
	wire [4-1:0] node28429;
	wire [4-1:0] node28430;
	wire [4-1:0] node28433;
	wire [4-1:0] node28436;
	wire [4-1:0] node28437;
	wire [4-1:0] node28440;
	wire [4-1:0] node28443;
	wire [4-1:0] node28444;
	wire [4-1:0] node28447;
	wire [4-1:0] node28450;
	wire [4-1:0] node28451;
	wire [4-1:0] node28452;
	wire [4-1:0] node28456;
	wire [4-1:0] node28457;
	wire [4-1:0] node28460;
	wire [4-1:0] node28463;
	wire [4-1:0] node28464;
	wire [4-1:0] node28465;
	wire [4-1:0] node28466;
	wire [4-1:0] node28467;
	wire [4-1:0] node28468;
	wire [4-1:0] node28470;
	wire [4-1:0] node28473;
	wire [4-1:0] node28475;
	wire [4-1:0] node28478;
	wire [4-1:0] node28479;
	wire [4-1:0] node28481;
	wire [4-1:0] node28484;
	wire [4-1:0] node28486;
	wire [4-1:0] node28489;
	wire [4-1:0] node28490;
	wire [4-1:0] node28492;
	wire [4-1:0] node28493;
	wire [4-1:0] node28495;
	wire [4-1:0] node28496;
	wire [4-1:0] node28499;
	wire [4-1:0] node28502;
	wire [4-1:0] node28503;
	wire [4-1:0] node28507;
	wire [4-1:0] node28508;
	wire [4-1:0] node28509;
	wire [4-1:0] node28510;
	wire [4-1:0] node28515;
	wire [4-1:0] node28516;
	wire [4-1:0] node28519;
	wire [4-1:0] node28522;
	wire [4-1:0] node28523;
	wire [4-1:0] node28524;
	wire [4-1:0] node28525;
	wire [4-1:0] node28526;
	wire [4-1:0] node28527;
	wire [4-1:0] node28530;
	wire [4-1:0] node28533;
	wire [4-1:0] node28536;
	wire [4-1:0] node28537;
	wire [4-1:0] node28539;
	wire [4-1:0] node28543;
	wire [4-1:0] node28544;
	wire [4-1:0] node28545;
	wire [4-1:0] node28546;
	wire [4-1:0] node28549;
	wire [4-1:0] node28550;
	wire [4-1:0] node28555;
	wire [4-1:0] node28556;
	wire [4-1:0] node28558;
	wire [4-1:0] node28561;
	wire [4-1:0] node28562;
	wire [4-1:0] node28566;
	wire [4-1:0] node28567;
	wire [4-1:0] node28568;
	wire [4-1:0] node28569;
	wire [4-1:0] node28572;
	wire [4-1:0] node28575;
	wire [4-1:0] node28576;
	wire [4-1:0] node28579;
	wire [4-1:0] node28582;
	wire [4-1:0] node28584;
	wire [4-1:0] node28585;
	wire [4-1:0] node28588;
	wire [4-1:0] node28591;
	wire [4-1:0] node28592;
	wire [4-1:0] node28593;
	wire [4-1:0] node28594;
	wire [4-1:0] node28595;
	wire [4-1:0] node28596;
	wire [4-1:0] node28597;
	wire [4-1:0] node28598;
	wire [4-1:0] node28601;
	wire [4-1:0] node28606;
	wire [4-1:0] node28607;
	wire [4-1:0] node28608;
	wire [4-1:0] node28612;
	wire [4-1:0] node28613;
	wire [4-1:0] node28617;
	wire [4-1:0] node28618;
	wire [4-1:0] node28619;
	wire [4-1:0] node28621;
	wire [4-1:0] node28624;
	wire [4-1:0] node28625;
	wire [4-1:0] node28626;
	wire [4-1:0] node28630;
	wire [4-1:0] node28633;
	wire [4-1:0] node28634;
	wire [4-1:0] node28635;
	wire [4-1:0] node28640;
	wire [4-1:0] node28641;
	wire [4-1:0] node28642;
	wire [4-1:0] node28643;
	wire [4-1:0] node28647;
	wire [4-1:0] node28648;
	wire [4-1:0] node28652;
	wire [4-1:0] node28653;
	wire [4-1:0] node28654;
	wire [4-1:0] node28658;
	wire [4-1:0] node28659;
	wire [4-1:0] node28663;
	wire [4-1:0] node28664;
	wire [4-1:0] node28665;
	wire [4-1:0] node28666;
	wire [4-1:0] node28667;
	wire [4-1:0] node28671;
	wire [4-1:0] node28672;
	wire [4-1:0] node28676;
	wire [4-1:0] node28677;
	wire [4-1:0] node28678;
	wire [4-1:0] node28682;
	wire [4-1:0] node28683;
	wire [4-1:0] node28687;
	wire [4-1:0] node28688;
	wire [4-1:0] node28689;
	wire [4-1:0] node28690;
	wire [4-1:0] node28694;
	wire [4-1:0] node28695;
	wire [4-1:0] node28699;
	wire [4-1:0] node28700;
	wire [4-1:0] node28703;
	wire [4-1:0] node28704;
	wire [4-1:0] node28708;
	wire [4-1:0] node28709;
	wire [4-1:0] node28710;
	wire [4-1:0] node28711;
	wire [4-1:0] node28712;
	wire [4-1:0] node28713;
	wire [4-1:0] node28714;
	wire [4-1:0] node28716;
	wire [4-1:0] node28717;
	wire [4-1:0] node28721;
	wire [4-1:0] node28722;
	wire [4-1:0] node28723;
	wire [4-1:0] node28726;
	wire [4-1:0] node28728;
	wire [4-1:0] node28731;
	wire [4-1:0] node28732;
	wire [4-1:0] node28735;
	wire [4-1:0] node28738;
	wire [4-1:0] node28739;
	wire [4-1:0] node28742;
	wire [4-1:0] node28744;
	wire [4-1:0] node28746;
	wire [4-1:0] node28747;
	wire [4-1:0] node28750;
	wire [4-1:0] node28753;
	wire [4-1:0] node28754;
	wire [4-1:0] node28755;
	wire [4-1:0] node28757;
	wire [4-1:0] node28758;
	wire [4-1:0] node28761;
	wire [4-1:0] node28764;
	wire [4-1:0] node28766;
	wire [4-1:0] node28767;
	wire [4-1:0] node28771;
	wire [4-1:0] node28772;
	wire [4-1:0] node28773;
	wire [4-1:0] node28774;
	wire [4-1:0] node28778;
	wire [4-1:0] node28779;
	wire [4-1:0] node28783;
	wire [4-1:0] node28784;
	wire [4-1:0] node28785;
	wire [4-1:0] node28788;
	wire [4-1:0] node28791;
	wire [4-1:0] node28793;
	wire [4-1:0] node28796;
	wire [4-1:0] node28797;
	wire [4-1:0] node28798;
	wire [4-1:0] node28799;
	wire [4-1:0] node28802;
	wire [4-1:0] node28803;
	wire [4-1:0] node28805;
	wire [4-1:0] node28807;
	wire [4-1:0] node28811;
	wire [4-1:0] node28812;
	wire [4-1:0] node28813;
	wire [4-1:0] node28814;
	wire [4-1:0] node28817;
	wire [4-1:0] node28820;
	wire [4-1:0] node28821;
	wire [4-1:0] node28822;
	wire [4-1:0] node28826;
	wire [4-1:0] node28827;
	wire [4-1:0] node28831;
	wire [4-1:0] node28834;
	wire [4-1:0] node28835;
	wire [4-1:0] node28836;
	wire [4-1:0] node28837;
	wire [4-1:0] node28838;
	wire [4-1:0] node28842;
	wire [4-1:0] node28843;
	wire [4-1:0] node28845;
	wire [4-1:0] node28849;
	wire [4-1:0] node28850;
	wire [4-1:0] node28853;
	wire [4-1:0] node28856;
	wire [4-1:0] node28857;
	wire [4-1:0] node28858;
	wire [4-1:0] node28859;
	wire [4-1:0] node28862;
	wire [4-1:0] node28865;
	wire [4-1:0] node28866;
	wire [4-1:0] node28870;
	wire [4-1:0] node28871;
	wire [4-1:0] node28874;
	wire [4-1:0] node28877;
	wire [4-1:0] node28878;
	wire [4-1:0] node28879;
	wire [4-1:0] node28880;
	wire [4-1:0] node28881;
	wire [4-1:0] node28882;
	wire [4-1:0] node28883;
	wire [4-1:0] node28887;
	wire [4-1:0] node28889;
	wire [4-1:0] node28892;
	wire [4-1:0] node28893;
	wire [4-1:0] node28895;
	wire [4-1:0] node28898;
	wire [4-1:0] node28901;
	wire [4-1:0] node28902;
	wire [4-1:0] node28903;
	wire [4-1:0] node28905;
	wire [4-1:0] node28908;
	wire [4-1:0] node28909;
	wire [4-1:0] node28910;
	wire [4-1:0] node28914;
	wire [4-1:0] node28917;
	wire [4-1:0] node28919;
	wire [4-1:0] node28920;
	wire [4-1:0] node28923;
	wire [4-1:0] node28926;
	wire [4-1:0] node28927;
	wire [4-1:0] node28928;
	wire [4-1:0] node28929;
	wire [4-1:0] node28930;
	wire [4-1:0] node28934;
	wire [4-1:0] node28936;
	wire [4-1:0] node28939;
	wire [4-1:0] node28940;
	wire [4-1:0] node28941;
	wire [4-1:0] node28945;
	wire [4-1:0] node28948;
	wire [4-1:0] node28949;
	wire [4-1:0] node28950;
	wire [4-1:0] node28951;
	wire [4-1:0] node28954;
	wire [4-1:0] node28957;
	wire [4-1:0] node28958;
	wire [4-1:0] node28961;
	wire [4-1:0] node28964;
	wire [4-1:0] node28965;
	wire [4-1:0] node28967;
	wire [4-1:0] node28970;
	wire [4-1:0] node28971;
	wire [4-1:0] node28975;
	wire [4-1:0] node28976;
	wire [4-1:0] node28977;
	wire [4-1:0] node28978;
	wire [4-1:0] node28979;
	wire [4-1:0] node28980;
	wire [4-1:0] node28983;
	wire [4-1:0] node28986;
	wire [4-1:0] node28987;
	wire [4-1:0] node28991;
	wire [4-1:0] node28992;
	wire [4-1:0] node28996;
	wire [4-1:0] node28997;
	wire [4-1:0] node28998;
	wire [4-1:0] node29001;
	wire [4-1:0] node29004;
	wire [4-1:0] node29005;
	wire [4-1:0] node29006;
	wire [4-1:0] node29010;
	wire [4-1:0] node29012;
	wire [4-1:0] node29015;
	wire [4-1:0] node29016;
	wire [4-1:0] node29017;
	wire [4-1:0] node29019;
	wire [4-1:0] node29020;
	wire [4-1:0] node29024;
	wire [4-1:0] node29025;
	wire [4-1:0] node29027;
	wire [4-1:0] node29029;
	wire [4-1:0] node29032;
	wire [4-1:0] node29034;
	wire [4-1:0] node29037;
	wire [4-1:0] node29038;
	wire [4-1:0] node29039;
	wire [4-1:0] node29041;
	wire [4-1:0] node29042;
	wire [4-1:0] node29045;
	wire [4-1:0] node29048;
	wire [4-1:0] node29049;
	wire [4-1:0] node29052;
	wire [4-1:0] node29054;
	wire [4-1:0] node29057;
	wire [4-1:0] node29058;
	wire [4-1:0] node29059;
	wire [4-1:0] node29061;
	wire [4-1:0] node29065;
	wire [4-1:0] node29067;
	wire [4-1:0] node29069;
	wire [4-1:0] node29072;
	wire [4-1:0] node29073;
	wire [4-1:0] node29074;
	wire [4-1:0] node29075;
	wire [4-1:0] node29076;
	wire [4-1:0] node29077;
	wire [4-1:0] node29078;
	wire [4-1:0] node29079;
	wire [4-1:0] node29083;
	wire [4-1:0] node29084;
	wire [4-1:0] node29085;
	wire [4-1:0] node29091;
	wire [4-1:0] node29092;
	wire [4-1:0] node29095;
	wire [4-1:0] node29096;
	wire [4-1:0] node29100;
	wire [4-1:0] node29101;
	wire [4-1:0] node29102;
	wire [4-1:0] node29103;
	wire [4-1:0] node29107;
	wire [4-1:0] node29108;
	wire [4-1:0] node29111;
	wire [4-1:0] node29114;
	wire [4-1:0] node29115;
	wire [4-1:0] node29116;
	wire [4-1:0] node29117;
	wire [4-1:0] node29120;
	wire [4-1:0] node29123;
	wire [4-1:0] node29125;
	wire [4-1:0] node29127;
	wire [4-1:0] node29130;
	wire [4-1:0] node29131;
	wire [4-1:0] node29132;
	wire [4-1:0] node29137;
	wire [4-1:0] node29138;
	wire [4-1:0] node29139;
	wire [4-1:0] node29140;
	wire [4-1:0] node29141;
	wire [4-1:0] node29143;
	wire [4-1:0] node29147;
	wire [4-1:0] node29148;
	wire [4-1:0] node29150;
	wire [4-1:0] node29153;
	wire [4-1:0] node29156;
	wire [4-1:0] node29157;
	wire [4-1:0] node29159;
	wire [4-1:0] node29162;
	wire [4-1:0] node29164;
	wire [4-1:0] node29167;
	wire [4-1:0] node29168;
	wire [4-1:0] node29169;
	wire [4-1:0] node29171;
	wire [4-1:0] node29174;
	wire [4-1:0] node29175;
	wire [4-1:0] node29176;
	wire [4-1:0] node29179;
	wire [4-1:0] node29182;
	wire [4-1:0] node29183;
	wire [4-1:0] node29185;
	wire [4-1:0] node29188;
	wire [4-1:0] node29189;
	wire [4-1:0] node29193;
	wire [4-1:0] node29194;
	wire [4-1:0] node29197;
	wire [4-1:0] node29200;
	wire [4-1:0] node29201;
	wire [4-1:0] node29202;
	wire [4-1:0] node29203;
	wire [4-1:0] node29204;
	wire [4-1:0] node29205;
	wire [4-1:0] node29209;
	wire [4-1:0] node29210;
	wire [4-1:0] node29212;
	wire [4-1:0] node29215;
	wire [4-1:0] node29218;
	wire [4-1:0] node29219;
	wire [4-1:0] node29221;
	wire [4-1:0] node29222;
	wire [4-1:0] node29226;
	wire [4-1:0] node29227;
	wire [4-1:0] node29231;
	wire [4-1:0] node29232;
	wire [4-1:0] node29233;
	wire [4-1:0] node29234;
	wire [4-1:0] node29235;
	wire [4-1:0] node29238;
	wire [4-1:0] node29241;
	wire [4-1:0] node29243;
	wire [4-1:0] node29246;
	wire [4-1:0] node29248;
	wire [4-1:0] node29249;
	wire [4-1:0] node29252;
	wire [4-1:0] node29255;
	wire [4-1:0] node29256;
	wire [4-1:0] node29257;
	wire [4-1:0] node29258;
	wire [4-1:0] node29261;
	wire [4-1:0] node29265;
	wire [4-1:0] node29266;
	wire [4-1:0] node29269;
	wire [4-1:0] node29272;
	wire [4-1:0] node29273;
	wire [4-1:0] node29274;
	wire [4-1:0] node29275;
	wire [4-1:0] node29277;
	wire [4-1:0] node29280;
	wire [4-1:0] node29281;
	wire [4-1:0] node29282;
	wire [4-1:0] node29286;
	wire [4-1:0] node29289;
	wire [4-1:0] node29290;
	wire [4-1:0] node29291;
	wire [4-1:0] node29293;
	wire [4-1:0] node29296;
	wire [4-1:0] node29299;
	wire [4-1:0] node29301;
	wire [4-1:0] node29302;
	wire [4-1:0] node29306;
	wire [4-1:0] node29307;
	wire [4-1:0] node29308;
	wire [4-1:0] node29309;
	wire [4-1:0] node29313;
	wire [4-1:0] node29314;
	wire [4-1:0] node29318;
	wire [4-1:0] node29319;
	wire [4-1:0] node29321;
	wire [4-1:0] node29324;
	wire [4-1:0] node29327;
	wire [4-1:0] node29328;
	wire [4-1:0] node29329;
	wire [4-1:0] node29330;
	wire [4-1:0] node29331;
	wire [4-1:0] node29332;
	wire [4-1:0] node29333;
	wire [4-1:0] node29334;
	wire [4-1:0] node29335;
	wire [4-1:0] node29336;
	wire [4-1:0] node29338;
	wire [4-1:0] node29341;
	wire [4-1:0] node29343;
	wire [4-1:0] node29346;
	wire [4-1:0] node29347;
	wire [4-1:0] node29349;
	wire [4-1:0] node29351;
	wire [4-1:0] node29354;
	wire [4-1:0] node29357;
	wire [4-1:0] node29358;
	wire [4-1:0] node29359;
	wire [4-1:0] node29360;
	wire [4-1:0] node29361;
	wire [4-1:0] node29365;
	wire [4-1:0] node29368;
	wire [4-1:0] node29370;
	wire [4-1:0] node29372;
	wire [4-1:0] node29375;
	wire [4-1:0] node29376;
	wire [4-1:0] node29377;
	wire [4-1:0] node29380;
	wire [4-1:0] node29383;
	wire [4-1:0] node29384;
	wire [4-1:0] node29386;
	wire [4-1:0] node29390;
	wire [4-1:0] node29391;
	wire [4-1:0] node29392;
	wire [4-1:0] node29393;
	wire [4-1:0] node29394;
	wire [4-1:0] node29397;
	wire [4-1:0] node29400;
	wire [4-1:0] node29401;
	wire [4-1:0] node29402;
	wire [4-1:0] node29403;
	wire [4-1:0] node29406;
	wire [4-1:0] node29409;
	wire [4-1:0] node29411;
	wire [4-1:0] node29415;
	wire [4-1:0] node29416;
	wire [4-1:0] node29417;
	wire [4-1:0] node29419;
	wire [4-1:0] node29423;
	wire [4-1:0] node29424;
	wire [4-1:0] node29427;
	wire [4-1:0] node29428;
	wire [4-1:0] node29430;
	wire [4-1:0] node29434;
	wire [4-1:0] node29435;
	wire [4-1:0] node29436;
	wire [4-1:0] node29437;
	wire [4-1:0] node29441;
	wire [4-1:0] node29442;
	wire [4-1:0] node29443;
	wire [4-1:0] node29447;
	wire [4-1:0] node29450;
	wire [4-1:0] node29451;
	wire [4-1:0] node29454;
	wire [4-1:0] node29455;
	wire [4-1:0] node29457;
	wire [4-1:0] node29460;
	wire [4-1:0] node29462;
	wire [4-1:0] node29465;
	wire [4-1:0] node29466;
	wire [4-1:0] node29467;
	wire [4-1:0] node29468;
	wire [4-1:0] node29469;
	wire [4-1:0] node29470;
	wire [4-1:0] node29473;
	wire [4-1:0] node29475;
	wire [4-1:0] node29478;
	wire [4-1:0] node29479;
	wire [4-1:0] node29482;
	wire [4-1:0] node29484;
	wire [4-1:0] node29487;
	wire [4-1:0] node29488;
	wire [4-1:0] node29489;
	wire [4-1:0] node29492;
	wire [4-1:0] node29494;
	wire [4-1:0] node29497;
	wire [4-1:0] node29499;
	wire [4-1:0] node29502;
	wire [4-1:0] node29503;
	wire [4-1:0] node29504;
	wire [4-1:0] node29505;
	wire [4-1:0] node29508;
	wire [4-1:0] node29510;
	wire [4-1:0] node29513;
	wire [4-1:0] node29514;
	wire [4-1:0] node29517;
	wire [4-1:0] node29519;
	wire [4-1:0] node29522;
	wire [4-1:0] node29524;
	wire [4-1:0] node29525;
	wire [4-1:0] node29526;
	wire [4-1:0] node29529;
	wire [4-1:0] node29532;
	wire [4-1:0] node29534;
	wire [4-1:0] node29537;
	wire [4-1:0] node29538;
	wire [4-1:0] node29539;
	wire [4-1:0] node29540;
	wire [4-1:0] node29541;
	wire [4-1:0] node29542;
	wire [4-1:0] node29545;
	wire [4-1:0] node29549;
	wire [4-1:0] node29551;
	wire [4-1:0] node29552;
	wire [4-1:0] node29553;
	wire [4-1:0] node29556;
	wire [4-1:0] node29559;
	wire [4-1:0] node29560;
	wire [4-1:0] node29564;
	wire [4-1:0] node29565;
	wire [4-1:0] node29566;
	wire [4-1:0] node29570;
	wire [4-1:0] node29571;
	wire [4-1:0] node29572;
	wire [4-1:0] node29577;
	wire [4-1:0] node29578;
	wire [4-1:0] node29579;
	wire [4-1:0] node29580;
	wire [4-1:0] node29583;
	wire [4-1:0] node29586;
	wire [4-1:0] node29587;
	wire [4-1:0] node29590;
	wire [4-1:0] node29593;
	wire [4-1:0] node29594;
	wire [4-1:0] node29596;
	wire [4-1:0] node29599;
	wire [4-1:0] node29601;
	wire [4-1:0] node29603;
	wire [4-1:0] node29604;
	wire [4-1:0] node29607;
	wire [4-1:0] node29610;
	wire [4-1:0] node29611;
	wire [4-1:0] node29612;
	wire [4-1:0] node29613;
	wire [4-1:0] node29614;
	wire [4-1:0] node29615;
	wire [4-1:0] node29616;
	wire [4-1:0] node29617;
	wire [4-1:0] node29620;
	wire [4-1:0] node29624;
	wire [4-1:0] node29625;
	wire [4-1:0] node29627;
	wire [4-1:0] node29628;
	wire [4-1:0] node29631;
	wire [4-1:0] node29635;
	wire [4-1:0] node29636;
	wire [4-1:0] node29637;
	wire [4-1:0] node29642;
	wire [4-1:0] node29643;
	wire [4-1:0] node29645;
	wire [4-1:0] node29646;
	wire [4-1:0] node29648;
	wire [4-1:0] node29649;
	wire [4-1:0] node29653;
	wire [4-1:0] node29654;
	wire [4-1:0] node29658;
	wire [4-1:0] node29659;
	wire [4-1:0] node29660;
	wire [4-1:0] node29662;
	wire [4-1:0] node29663;
	wire [4-1:0] node29667;
	wire [4-1:0] node29669;
	wire [4-1:0] node29672;
	wire [4-1:0] node29673;
	wire [4-1:0] node29674;
	wire [4-1:0] node29677;
	wire [4-1:0] node29679;
	wire [4-1:0] node29682;
	wire [4-1:0] node29683;
	wire [4-1:0] node29687;
	wire [4-1:0] node29688;
	wire [4-1:0] node29689;
	wire [4-1:0] node29690;
	wire [4-1:0] node29691;
	wire [4-1:0] node29692;
	wire [4-1:0] node29697;
	wire [4-1:0] node29699;
	wire [4-1:0] node29700;
	wire [4-1:0] node29702;
	wire [4-1:0] node29706;
	wire [4-1:0] node29707;
	wire [4-1:0] node29709;
	wire [4-1:0] node29712;
	wire [4-1:0] node29713;
	wire [4-1:0] node29714;
	wire [4-1:0] node29718;
	wire [4-1:0] node29721;
	wire [4-1:0] node29722;
	wire [4-1:0] node29723;
	wire [4-1:0] node29724;
	wire [4-1:0] node29725;
	wire [4-1:0] node29727;
	wire [4-1:0] node29730;
	wire [4-1:0] node29731;
	wire [4-1:0] node29734;
	wire [4-1:0] node29737;
	wire [4-1:0] node29738;
	wire [4-1:0] node29742;
	wire [4-1:0] node29743;
	wire [4-1:0] node29746;
	wire [4-1:0] node29749;
	wire [4-1:0] node29750;
	wire [4-1:0] node29751;
	wire [4-1:0] node29752;
	wire [4-1:0] node29757;
	wire [4-1:0] node29760;
	wire [4-1:0] node29761;
	wire [4-1:0] node29762;
	wire [4-1:0] node29763;
	wire [4-1:0] node29764;
	wire [4-1:0] node29765;
	wire [4-1:0] node29767;
	wire [4-1:0] node29768;
	wire [4-1:0] node29771;
	wire [4-1:0] node29774;
	wire [4-1:0] node29775;
	wire [4-1:0] node29777;
	wire [4-1:0] node29781;
	wire [4-1:0] node29784;
	wire [4-1:0] node29785;
	wire [4-1:0] node29786;
	wire [4-1:0] node29787;
	wire [4-1:0] node29791;
	wire [4-1:0] node29794;
	wire [4-1:0] node29795;
	wire [4-1:0] node29796;
	wire [4-1:0] node29799;
	wire [4-1:0] node29802;
	wire [4-1:0] node29804;
	wire [4-1:0] node29805;
	wire [4-1:0] node29808;
	wire [4-1:0] node29811;
	wire [4-1:0] node29812;
	wire [4-1:0] node29813;
	wire [4-1:0] node29814;
	wire [4-1:0] node29816;
	wire [4-1:0] node29819;
	wire [4-1:0] node29821;
	wire [4-1:0] node29824;
	wire [4-1:0] node29826;
	wire [4-1:0] node29828;
	wire [4-1:0] node29831;
	wire [4-1:0] node29832;
	wire [4-1:0] node29833;
	wire [4-1:0] node29837;
	wire [4-1:0] node29838;
	wire [4-1:0] node29839;
	wire [4-1:0] node29840;
	wire [4-1:0] node29846;
	wire [4-1:0] node29847;
	wire [4-1:0] node29848;
	wire [4-1:0] node29849;
	wire [4-1:0] node29850;
	wire [4-1:0] node29852;
	wire [4-1:0] node29855;
	wire [4-1:0] node29856;
	wire [4-1:0] node29860;
	wire [4-1:0] node29861;
	wire [4-1:0] node29865;
	wire [4-1:0] node29866;
	wire [4-1:0] node29867;
	wire [4-1:0] node29869;
	wire [4-1:0] node29872;
	wire [4-1:0] node29875;
	wire [4-1:0] node29876;
	wire [4-1:0] node29879;
	wire [4-1:0] node29880;
	wire [4-1:0] node29881;
	wire [4-1:0] node29885;
	wire [4-1:0] node29888;
	wire [4-1:0] node29889;
	wire [4-1:0] node29890;
	wire [4-1:0] node29891;
	wire [4-1:0] node29892;
	wire [4-1:0] node29893;
	wire [4-1:0] node29897;
	wire [4-1:0] node29898;
	wire [4-1:0] node29903;
	wire [4-1:0] node29904;
	wire [4-1:0] node29907;
	wire [4-1:0] node29910;
	wire [4-1:0] node29911;
	wire [4-1:0] node29912;
	wire [4-1:0] node29913;
	wire [4-1:0] node29914;
	wire [4-1:0] node29920;
	wire [4-1:0] node29921;
	wire [4-1:0] node29925;
	wire [4-1:0] node29926;
	wire [4-1:0] node29927;
	wire [4-1:0] node29928;
	wire [4-1:0] node29929;
	wire [4-1:0] node29930;
	wire [4-1:0] node29932;
	wire [4-1:0] node29935;
	wire [4-1:0] node29937;
	wire [4-1:0] node29939;
	wire [4-1:0] node29942;
	wire [4-1:0] node29943;
	wire [4-1:0] node29945;
	wire [4-1:0] node29947;
	wire [4-1:0] node29949;
	wire [4-1:0] node29952;
	wire [4-1:0] node29953;
	wire [4-1:0] node29955;
	wire [4-1:0] node29958;
	wire [4-1:0] node29960;
	wire [4-1:0] node29963;
	wire [4-1:0] node29964;
	wire [4-1:0] node29965;
	wire [4-1:0] node29966;
	wire [4-1:0] node29968;
	wire [4-1:0] node29971;
	wire [4-1:0] node29973;
	wire [4-1:0] node29976;
	wire [4-1:0] node29977;
	wire [4-1:0] node29979;
	wire [4-1:0] node29982;
	wire [4-1:0] node29984;
	wire [4-1:0] node29987;
	wire [4-1:0] node29988;
	wire [4-1:0] node29989;
	wire [4-1:0] node29991;
	wire [4-1:0] node29994;
	wire [4-1:0] node29995;
	wire [4-1:0] node29996;
	wire [4-1:0] node30000;
	wire [4-1:0] node30001;
	wire [4-1:0] node30004;
	wire [4-1:0] node30007;
	wire [4-1:0] node30008;
	wire [4-1:0] node30009;
	wire [4-1:0] node30013;
	wire [4-1:0] node30014;
	wire [4-1:0] node30018;
	wire [4-1:0] node30019;
	wire [4-1:0] node30020;
	wire [4-1:0] node30021;
	wire [4-1:0] node30022;
	wire [4-1:0] node30025;
	wire [4-1:0] node30026;
	wire [4-1:0] node30027;
	wire [4-1:0] node30028;
	wire [4-1:0] node30031;
	wire [4-1:0] node30035;
	wire [4-1:0] node30037;
	wire [4-1:0] node30040;
	wire [4-1:0] node30041;
	wire [4-1:0] node30043;
	wire [4-1:0] node30046;
	wire [4-1:0] node30048;
	wire [4-1:0] node30051;
	wire [4-1:0] node30052;
	wire [4-1:0] node30053;
	wire [4-1:0] node30055;
	wire [4-1:0] node30059;
	wire [4-1:0] node30060;
	wire [4-1:0] node30062;
	wire [4-1:0] node30065;
	wire [4-1:0] node30068;
	wire [4-1:0] node30069;
	wire [4-1:0] node30070;
	wire [4-1:0] node30071;
	wire [4-1:0] node30073;
	wire [4-1:0] node30076;
	wire [4-1:0] node30078;
	wire [4-1:0] node30081;
	wire [4-1:0] node30082;
	wire [4-1:0] node30084;
	wire [4-1:0] node30088;
	wire [4-1:0] node30089;
	wire [4-1:0] node30090;
	wire [4-1:0] node30091;
	wire [4-1:0] node30095;
	wire [4-1:0] node30096;
	wire [4-1:0] node30099;
	wire [4-1:0] node30101;
	wire [4-1:0] node30104;
	wire [4-1:0] node30105;
	wire [4-1:0] node30106;
	wire [4-1:0] node30108;
	wire [4-1:0] node30111;
	wire [4-1:0] node30113;
	wire [4-1:0] node30116;
	wire [4-1:0] node30117;
	wire [4-1:0] node30121;
	wire [4-1:0] node30122;
	wire [4-1:0] node30123;
	wire [4-1:0] node30124;
	wire [4-1:0] node30125;
	wire [4-1:0] node30126;
	wire [4-1:0] node30127;
	wire [4-1:0] node30128;
	wire [4-1:0] node30132;
	wire [4-1:0] node30135;
	wire [4-1:0] node30136;
	wire [4-1:0] node30137;
	wire [4-1:0] node30141;
	wire [4-1:0] node30142;
	wire [4-1:0] node30145;
	wire [4-1:0] node30148;
	wire [4-1:0] node30149;
	wire [4-1:0] node30150;
	wire [4-1:0] node30152;
	wire [4-1:0] node30155;
	wire [4-1:0] node30157;
	wire [4-1:0] node30160;
	wire [4-1:0] node30162;
	wire [4-1:0] node30165;
	wire [4-1:0] node30166;
	wire [4-1:0] node30168;
	wire [4-1:0] node30170;
	wire [4-1:0] node30173;
	wire [4-1:0] node30174;
	wire [4-1:0] node30177;
	wire [4-1:0] node30179;
	wire [4-1:0] node30182;
	wire [4-1:0] node30183;
	wire [4-1:0] node30184;
	wire [4-1:0] node30185;
	wire [4-1:0] node30188;
	wire [4-1:0] node30190;
	wire [4-1:0] node30193;
	wire [4-1:0] node30194;
	wire [4-1:0] node30196;
	wire [4-1:0] node30199;
	wire [4-1:0] node30201;
	wire [4-1:0] node30204;
	wire [4-1:0] node30205;
	wire [4-1:0] node30206;
	wire [4-1:0] node30207;
	wire [4-1:0] node30208;
	wire [4-1:0] node30209;
	wire [4-1:0] node30213;
	wire [4-1:0] node30216;
	wire [4-1:0] node30217;
	wire [4-1:0] node30221;
	wire [4-1:0] node30222;
	wire [4-1:0] node30225;
	wire [4-1:0] node30228;
	wire [4-1:0] node30229;
	wire [4-1:0] node30232;
	wire [4-1:0] node30234;
	wire [4-1:0] node30237;
	wire [4-1:0] node30238;
	wire [4-1:0] node30239;
	wire [4-1:0] node30240;
	wire [4-1:0] node30242;
	wire [4-1:0] node30243;
	wire [4-1:0] node30246;
	wire [4-1:0] node30249;
	wire [4-1:0] node30250;
	wire [4-1:0] node30252;
	wire [4-1:0] node30255;
	wire [4-1:0] node30257;
	wire [4-1:0] node30260;
	wire [4-1:0] node30261;
	wire [4-1:0] node30262;
	wire [4-1:0] node30264;
	wire [4-1:0] node30267;
	wire [4-1:0] node30269;
	wire [4-1:0] node30272;
	wire [4-1:0] node30273;
	wire [4-1:0] node30275;
	wire [4-1:0] node30278;
	wire [4-1:0] node30280;
	wire [4-1:0] node30283;
	wire [4-1:0] node30284;
	wire [4-1:0] node30285;
	wire [4-1:0] node30286;
	wire [4-1:0] node30290;
	wire [4-1:0] node30291;
	wire [4-1:0] node30293;
	wire [4-1:0] node30296;
	wire [4-1:0] node30298;
	wire [4-1:0] node30301;
	wire [4-1:0] node30302;
	wire [4-1:0] node30303;
	wire [4-1:0] node30304;
	wire [4-1:0] node30306;
	wire [4-1:0] node30309;
	wire [4-1:0] node30311;
	wire [4-1:0] node30314;
	wire [4-1:0] node30315;
	wire [4-1:0] node30317;
	wire [4-1:0] node30320;
	wire [4-1:0] node30322;
	wire [4-1:0] node30325;
	wire [4-1:0] node30326;
	wire [4-1:0] node30327;
	wire [4-1:0] node30328;
	wire [4-1:0] node30332;
	wire [4-1:0] node30334;
	wire [4-1:0] node30335;
	wire [4-1:0] node30338;
	wire [4-1:0] node30341;
	wire [4-1:0] node30342;
	wire [4-1:0] node30343;
	wire [4-1:0] node30347;
	wire [4-1:0] node30349;
	wire [4-1:0] node30350;
	wire [4-1:0] node30353;
	wire [4-1:0] node30356;
	wire [4-1:0] node30357;
	wire [4-1:0] node30358;
	wire [4-1:0] node30359;
	wire [4-1:0] node30360;
	wire [4-1:0] node30361;
	wire [4-1:0] node30362;
	wire [4-1:0] node30363;
	wire [4-1:0] node30365;
	wire [4-1:0] node30368;
	wire [4-1:0] node30370;
	wire [4-1:0] node30371;
	wire [4-1:0] node30372;
	wire [4-1:0] node30376;
	wire [4-1:0] node30378;
	wire [4-1:0] node30381;
	wire [4-1:0] node30382;
	wire [4-1:0] node30383;
	wire [4-1:0] node30385;
	wire [4-1:0] node30388;
	wire [4-1:0] node30389;
	wire [4-1:0] node30392;
	wire [4-1:0] node30395;
	wire [4-1:0] node30396;
	wire [4-1:0] node30398;
	wire [4-1:0] node30400;
	wire [4-1:0] node30403;
	wire [4-1:0] node30404;
	wire [4-1:0] node30408;
	wire [4-1:0] node30409;
	wire [4-1:0] node30410;
	wire [4-1:0] node30411;
	wire [4-1:0] node30413;
	wire [4-1:0] node30416;
	wire [4-1:0] node30417;
	wire [4-1:0] node30420;
	wire [4-1:0] node30423;
	wire [4-1:0] node30424;
	wire [4-1:0] node30426;
	wire [4-1:0] node30429;
	wire [4-1:0] node30430;
	wire [4-1:0] node30431;
	wire [4-1:0] node30434;
	wire [4-1:0] node30437;
	wire [4-1:0] node30438;
	wire [4-1:0] node30441;
	wire [4-1:0] node30444;
	wire [4-1:0] node30445;
	wire [4-1:0] node30446;
	wire [4-1:0] node30448;
	wire [4-1:0] node30451;
	wire [4-1:0] node30452;
	wire [4-1:0] node30455;
	wire [4-1:0] node30458;
	wire [4-1:0] node30460;
	wire [4-1:0] node30462;
	wire [4-1:0] node30465;
	wire [4-1:0] node30466;
	wire [4-1:0] node30467;
	wire [4-1:0] node30468;
	wire [4-1:0] node30469;
	wire [4-1:0] node30470;
	wire [4-1:0] node30475;
	wire [4-1:0] node30476;
	wire [4-1:0] node30478;
	wire [4-1:0] node30481;
	wire [4-1:0] node30483;
	wire [4-1:0] node30486;
	wire [4-1:0] node30487;
	wire [4-1:0] node30488;
	wire [4-1:0] node30492;
	wire [4-1:0] node30493;
	wire [4-1:0] node30496;
	wire [4-1:0] node30499;
	wire [4-1:0] node30500;
	wire [4-1:0] node30501;
	wire [4-1:0] node30502;
	wire [4-1:0] node30505;
	wire [4-1:0] node30508;
	wire [4-1:0] node30510;
	wire [4-1:0] node30513;
	wire [4-1:0] node30514;
	wire [4-1:0] node30515;
	wire [4-1:0] node30519;
	wire [4-1:0] node30520;
	wire [4-1:0] node30523;
	wire [4-1:0] node30526;
	wire [4-1:0] node30527;
	wire [4-1:0] node30528;
	wire [4-1:0] node30529;
	wire [4-1:0] node30530;
	wire [4-1:0] node30532;
	wire [4-1:0] node30533;
	wire [4-1:0] node30537;
	wire [4-1:0] node30538;
	wire [4-1:0] node30541;
	wire [4-1:0] node30544;
	wire [4-1:0] node30545;
	wire [4-1:0] node30546;
	wire [4-1:0] node30548;
	wire [4-1:0] node30552;
	wire [4-1:0] node30553;
	wire [4-1:0] node30554;
	wire [4-1:0] node30557;
	wire [4-1:0] node30560;
	wire [4-1:0] node30561;
	wire [4-1:0] node30564;
	wire [4-1:0] node30567;
	wire [4-1:0] node30568;
	wire [4-1:0] node30569;
	wire [4-1:0] node30570;
	wire [4-1:0] node30573;
	wire [4-1:0] node30576;
	wire [4-1:0] node30577;
	wire [4-1:0] node30578;
	wire [4-1:0] node30582;
	wire [4-1:0] node30583;
	wire [4-1:0] node30586;
	wire [4-1:0] node30589;
	wire [4-1:0] node30590;
	wire [4-1:0] node30591;
	wire [4-1:0] node30592;
	wire [4-1:0] node30595;
	wire [4-1:0] node30598;
	wire [4-1:0] node30601;
	wire [4-1:0] node30603;
	wire [4-1:0] node30604;
	wire [4-1:0] node30608;
	wire [4-1:0] node30609;
	wire [4-1:0] node30610;
	wire [4-1:0] node30611;
	wire [4-1:0] node30612;
	wire [4-1:0] node30614;
	wire [4-1:0] node30615;
	wire [4-1:0] node30618;
	wire [4-1:0] node30621;
	wire [4-1:0] node30622;
	wire [4-1:0] node30624;
	wire [4-1:0] node30627;
	wire [4-1:0] node30630;
	wire [4-1:0] node30631;
	wire [4-1:0] node30632;
	wire [4-1:0] node30635;
	wire [4-1:0] node30637;
	wire [4-1:0] node30640;
	wire [4-1:0] node30642;
	wire [4-1:0] node30644;
	wire [4-1:0] node30647;
	wire [4-1:0] node30648;
	wire [4-1:0] node30650;
	wire [4-1:0] node30653;
	wire [4-1:0] node30654;
	wire [4-1:0] node30656;
	wire [4-1:0] node30660;
	wire [4-1:0] node30661;
	wire [4-1:0] node30662;
	wire [4-1:0] node30663;
	wire [4-1:0] node30664;
	wire [4-1:0] node30667;
	wire [4-1:0] node30669;
	wire [4-1:0] node30672;
	wire [4-1:0] node30673;
	wire [4-1:0] node30674;
	wire [4-1:0] node30677;
	wire [4-1:0] node30680;
	wire [4-1:0] node30681;
	wire [4-1:0] node30685;
	wire [4-1:0] node30686;
	wire [4-1:0] node30687;
	wire [4-1:0] node30690;
	wire [4-1:0] node30693;
	wire [4-1:0] node30694;
	wire [4-1:0] node30698;
	wire [4-1:0] node30699;
	wire [4-1:0] node30700;
	wire [4-1:0] node30701;
	wire [4-1:0] node30705;
	wire [4-1:0] node30707;
	wire [4-1:0] node30709;
	wire [4-1:0] node30712;
	wire [4-1:0] node30713;
	wire [4-1:0] node30714;
	wire [4-1:0] node30716;
	wire [4-1:0] node30719;
	wire [4-1:0] node30722;
	wire [4-1:0] node30724;
	wire [4-1:0] node30725;
	wire [4-1:0] node30729;
	wire [4-1:0] node30730;
	wire [4-1:0] node30731;
	wire [4-1:0] node30732;
	wire [4-1:0] node30733;
	wire [4-1:0] node30734;
	wire [4-1:0] node30735;
	wire [4-1:0] node30739;
	wire [4-1:0] node30741;
	wire [4-1:0] node30742;
	wire [4-1:0] node30746;
	wire [4-1:0] node30747;
	wire [4-1:0] node30748;
	wire [4-1:0] node30749;
	wire [4-1:0] node30754;
	wire [4-1:0] node30755;
	wire [4-1:0] node30759;
	wire [4-1:0] node30760;
	wire [4-1:0] node30761;
	wire [4-1:0] node30762;
	wire [4-1:0] node30767;
	wire [4-1:0] node30769;
	wire [4-1:0] node30770;
	wire [4-1:0] node30773;
	wire [4-1:0] node30774;
	wire [4-1:0] node30778;
	wire [4-1:0] node30779;
	wire [4-1:0] node30780;
	wire [4-1:0] node30781;
	wire [4-1:0] node30782;
	wire [4-1:0] node30783;
	wire [4-1:0] node30784;
	wire [4-1:0] node30787;
	wire [4-1:0] node30791;
	wire [4-1:0] node30792;
	wire [4-1:0] node30796;
	wire [4-1:0] node30797;
	wire [4-1:0] node30800;
	wire [4-1:0] node30803;
	wire [4-1:0] node30804;
	wire [4-1:0] node30805;
	wire [4-1:0] node30806;
	wire [4-1:0] node30807;
	wire [4-1:0] node30812;
	wire [4-1:0] node30815;
	wire [4-1:0] node30816;
	wire [4-1:0] node30817;
	wire [4-1:0] node30822;
	wire [4-1:0] node30823;
	wire [4-1:0] node30824;
	wire [4-1:0] node30825;
	wire [4-1:0] node30827;
	wire [4-1:0] node30830;
	wire [4-1:0] node30831;
	wire [4-1:0] node30833;
	wire [4-1:0] node30837;
	wire [4-1:0] node30839;
	wire [4-1:0] node30842;
	wire [4-1:0] node30843;
	wire [4-1:0] node30845;
	wire [4-1:0] node30848;
	wire [4-1:0] node30850;
	wire [4-1:0] node30853;
	wire [4-1:0] node30854;
	wire [4-1:0] node30855;
	wire [4-1:0] node30856;
	wire [4-1:0] node30857;
	wire [4-1:0] node30859;
	wire [4-1:0] node30860;
	wire [4-1:0] node30863;
	wire [4-1:0] node30866;
	wire [4-1:0] node30868;
	wire [4-1:0] node30870;
	wire [4-1:0] node30872;
	wire [4-1:0] node30875;
	wire [4-1:0] node30876;
	wire [4-1:0] node30878;
	wire [4-1:0] node30879;
	wire [4-1:0] node30880;
	wire [4-1:0] node30883;
	wire [4-1:0] node30886;
	wire [4-1:0] node30887;
	wire [4-1:0] node30890;
	wire [4-1:0] node30893;
	wire [4-1:0] node30895;
	wire [4-1:0] node30897;
	wire [4-1:0] node30900;
	wire [4-1:0] node30901;
	wire [4-1:0] node30902;
	wire [4-1:0] node30904;
	wire [4-1:0] node30905;
	wire [4-1:0] node30908;
	wire [4-1:0] node30909;
	wire [4-1:0] node30913;
	wire [4-1:0] node30914;
	wire [4-1:0] node30915;
	wire [4-1:0] node30919;
	wire [4-1:0] node30920;
	wire [4-1:0] node30923;
	wire [4-1:0] node30926;
	wire [4-1:0] node30927;
	wire [4-1:0] node30930;
	wire [4-1:0] node30933;
	wire [4-1:0] node30934;
	wire [4-1:0] node30935;
	wire [4-1:0] node30936;
	wire [4-1:0] node30937;
	wire [4-1:0] node30938;
	wire [4-1:0] node30942;
	wire [4-1:0] node30943;
	wire [4-1:0] node30947;
	wire [4-1:0] node30949;
	wire [4-1:0] node30950;
	wire [4-1:0] node30954;
	wire [4-1:0] node30955;
	wire [4-1:0] node30957;
	wire [4-1:0] node30960;
	wire [4-1:0] node30961;
	wire [4-1:0] node30963;
	wire [4-1:0] node30966;
	wire [4-1:0] node30967;
	wire [4-1:0] node30970;
	wire [4-1:0] node30973;
	wire [4-1:0] node30974;
	wire [4-1:0] node30975;
	wire [4-1:0] node30977;
	wire [4-1:0] node30978;
	wire [4-1:0] node30982;
	wire [4-1:0] node30983;
	wire [4-1:0] node30985;
	wire [4-1:0] node30986;
	wire [4-1:0] node30990;
	wire [4-1:0] node30991;
	wire [4-1:0] node30995;
	wire [4-1:0] node30996;
	wire [4-1:0] node30997;
	wire [4-1:0] node31000;
	wire [4-1:0] node31003;
	wire [4-1:0] node31004;
	wire [4-1:0] node31005;
	wire [4-1:0] node31008;
	wire [4-1:0] node31011;
	wire [4-1:0] node31012;
	wire [4-1:0] node31015;
	wire [4-1:0] node31018;
	wire [4-1:0] node31019;
	wire [4-1:0] node31020;
	wire [4-1:0] node31021;
	wire [4-1:0] node31022;
	wire [4-1:0] node31023;
	wire [4-1:0] node31024;
	wire [4-1:0] node31025;
	wire [4-1:0] node31026;
	wire [4-1:0] node31030;
	wire [4-1:0] node31034;
	wire [4-1:0] node31035;
	wire [4-1:0] node31036;
	wire [4-1:0] node31040;
	wire [4-1:0] node31041;
	wire [4-1:0] node31045;
	wire [4-1:0] node31046;
	wire [4-1:0] node31047;
	wire [4-1:0] node31048;
	wire [4-1:0] node31052;
	wire [4-1:0] node31053;
	wire [4-1:0] node31057;
	wire [4-1:0] node31059;
	wire [4-1:0] node31060;
	wire [4-1:0] node31064;
	wire [4-1:0] node31065;
	wire [4-1:0] node31066;
	wire [4-1:0] node31067;
	wire [4-1:0] node31068;
	wire [4-1:0] node31072;
	wire [4-1:0] node31073;
	wire [4-1:0] node31077;
	wire [4-1:0] node31078;
	wire [4-1:0] node31079;
	wire [4-1:0] node31083;
	wire [4-1:0] node31086;
	wire [4-1:0] node31087;
	wire [4-1:0] node31088;
	wire [4-1:0] node31089;
	wire [4-1:0] node31093;
	wire [4-1:0] node31094;
	wire [4-1:0] node31098;
	wire [4-1:0] node31099;
	wire [4-1:0] node31100;
	wire [4-1:0] node31104;
	wire [4-1:0] node31106;
	wire [4-1:0] node31109;
	wire [4-1:0] node31110;
	wire [4-1:0] node31111;
	wire [4-1:0] node31112;
	wire [4-1:0] node31113;
	wire [4-1:0] node31114;
	wire [4-1:0] node31118;
	wire [4-1:0] node31119;
	wire [4-1:0] node31123;
	wire [4-1:0] node31124;
	wire [4-1:0] node31125;
	wire [4-1:0] node31129;
	wire [4-1:0] node31132;
	wire [4-1:0] node31133;
	wire [4-1:0] node31134;
	wire [4-1:0] node31135;
	wire [4-1:0] node31139;
	wire [4-1:0] node31140;
	wire [4-1:0] node31144;
	wire [4-1:0] node31145;
	wire [4-1:0] node31146;
	wire [4-1:0] node31150;
	wire [4-1:0] node31151;
	wire [4-1:0] node31155;
	wire [4-1:0] node31156;
	wire [4-1:0] node31157;
	wire [4-1:0] node31158;
	wire [4-1:0] node31159;
	wire [4-1:0] node31163;
	wire [4-1:0] node31164;
	wire [4-1:0] node31168;
	wire [4-1:0] node31169;
	wire [4-1:0] node31170;
	wire [4-1:0] node31175;
	wire [4-1:0] node31176;
	wire [4-1:0] node31177;
	wire [4-1:0] node31179;
	wire [4-1:0] node31180;
	wire [4-1:0] node31184;
	wire [4-1:0] node31186;
	wire [4-1:0] node31189;
	wire [4-1:0] node31190;
	wire [4-1:0] node31192;
	wire [4-1:0] node31195;
	wire [4-1:0] node31196;
	wire [4-1:0] node31197;
	wire [4-1:0] node31202;
	wire [4-1:0] node31203;
	wire [4-1:0] node31204;
	wire [4-1:0] node31205;
	wire [4-1:0] node31206;
	wire [4-1:0] node31207;
	wire [4-1:0] node31209;
	wire [4-1:0] node31213;
	wire [4-1:0] node31214;
	wire [4-1:0] node31216;
	wire [4-1:0] node31219;
	wire [4-1:0] node31220;
	wire [4-1:0] node31224;
	wire [4-1:0] node31225;
	wire [4-1:0] node31226;
	wire [4-1:0] node31228;
	wire [4-1:0] node31232;
	wire [4-1:0] node31234;
	wire [4-1:0] node31237;
	wire [4-1:0] node31238;
	wire [4-1:0] node31239;
	wire [4-1:0] node31240;
	wire [4-1:0] node31242;
	wire [4-1:0] node31245;
	wire [4-1:0] node31247;
	wire [4-1:0] node31250;
	wire [4-1:0] node31251;
	wire [4-1:0] node31252;
	wire [4-1:0] node31256;
	wire [4-1:0] node31257;
	wire [4-1:0] node31261;
	wire [4-1:0] node31262;
	wire [4-1:0] node31263;
	wire [4-1:0] node31267;
	wire [4-1:0] node31268;
	wire [4-1:0] node31272;
	wire [4-1:0] node31273;
	wire [4-1:0] node31274;
	wire [4-1:0] node31275;
	wire [4-1:0] node31276;
	wire [4-1:0] node31277;
	wire [4-1:0] node31281;
	wire [4-1:0] node31283;
	wire [4-1:0] node31286;
	wire [4-1:0] node31287;
	wire [4-1:0] node31288;
	wire [4-1:0] node31290;
	wire [4-1:0] node31293;
	wire [4-1:0] node31294;
	wire [4-1:0] node31295;
	wire [4-1:0] node31298;
	wire [4-1:0] node31301;
	wire [4-1:0] node31302;
	wire [4-1:0] node31305;
	wire [4-1:0] node31309;
	wire [4-1:0] node31310;
	wire [4-1:0] node31311;
	wire [4-1:0] node31315;
	wire [4-1:0] node31317;
	wire [4-1:0] node31320;
	wire [4-1:0] node31321;
	wire [4-1:0] node31322;
	wire [4-1:0] node31323;
	wire [4-1:0] node31324;
	wire [4-1:0] node31328;
	wire [4-1:0] node31329;
	wire [4-1:0] node31333;
	wire [4-1:0] node31334;
	wire [4-1:0] node31338;
	wire [4-1:0] node31339;
	wire [4-1:0] node31341;
	wire [4-1:0] node31342;
	wire [4-1:0] node31346;
	wire [4-1:0] node31347;
	wire [4-1:0] node31351;
	wire [4-1:0] node31352;
	wire [4-1:0] node31353;
	wire [4-1:0] node31354;
	wire [4-1:0] node31355;
	wire [4-1:0] node31356;
	wire [4-1:0] node31357;
	wire [4-1:0] node31358;
	wire [4-1:0] node31359;
	wire [4-1:0] node31360;
	wire [4-1:0] node31363;
	wire [4-1:0] node31366;
	wire [4-1:0] node31367;
	wire [4-1:0] node31369;
	wire [4-1:0] node31372;
	wire [4-1:0] node31373;
	wire [4-1:0] node31377;
	wire [4-1:0] node31378;
	wire [4-1:0] node31379;
	wire [4-1:0] node31381;
	wire [4-1:0] node31384;
	wire [4-1:0] node31387;
	wire [4-1:0] node31388;
	wire [4-1:0] node31390;
	wire [4-1:0] node31393;
	wire [4-1:0] node31395;
	wire [4-1:0] node31398;
	wire [4-1:0] node31399;
	wire [4-1:0] node31400;
	wire [4-1:0] node31402;
	wire [4-1:0] node31403;
	wire [4-1:0] node31406;
	wire [4-1:0] node31409;
	wire [4-1:0] node31410;
	wire [4-1:0] node31412;
	wire [4-1:0] node31416;
	wire [4-1:0] node31417;
	wire [4-1:0] node31418;
	wire [4-1:0] node31421;
	wire [4-1:0] node31424;
	wire [4-1:0] node31425;
	wire [4-1:0] node31427;
	wire [4-1:0] node31431;
	wire [4-1:0] node31432;
	wire [4-1:0] node31433;
	wire [4-1:0] node31434;
	wire [4-1:0] node31435;
	wire [4-1:0] node31438;
	wire [4-1:0] node31440;
	wire [4-1:0] node31443;
	wire [4-1:0] node31444;
	wire [4-1:0] node31446;
	wire [4-1:0] node31450;
	wire [4-1:0] node31451;
	wire [4-1:0] node31452;
	wire [4-1:0] node31453;
	wire [4-1:0] node31456;
	wire [4-1:0] node31459;
	wire [4-1:0] node31460;
	wire [4-1:0] node31465;
	wire [4-1:0] node31466;
	wire [4-1:0] node31467;
	wire [4-1:0] node31468;
	wire [4-1:0] node31471;
	wire [4-1:0] node31473;
	wire [4-1:0] node31476;
	wire [4-1:0] node31477;
	wire [4-1:0] node31481;
	wire [4-1:0] node31482;
	wire [4-1:0] node31484;
	wire [4-1:0] node31485;
	wire [4-1:0] node31488;
	wire [4-1:0] node31491;
	wire [4-1:0] node31492;
	wire [4-1:0] node31495;
	wire [4-1:0] node31497;
	wire [4-1:0] node31500;
	wire [4-1:0] node31501;
	wire [4-1:0] node31502;
	wire [4-1:0] node31503;
	wire [4-1:0] node31504;
	wire [4-1:0] node31505;
	wire [4-1:0] node31507;
	wire [4-1:0] node31511;
	wire [4-1:0] node31512;
	wire [4-1:0] node31514;
	wire [4-1:0] node31517;
	wire [4-1:0] node31520;
	wire [4-1:0] node31521;
	wire [4-1:0] node31522;
	wire [4-1:0] node31524;
	wire [4-1:0] node31527;
	wire [4-1:0] node31529;
	wire [4-1:0] node31532;
	wire [4-1:0] node31534;
	wire [4-1:0] node31537;
	wire [4-1:0] node31538;
	wire [4-1:0] node31539;
	wire [4-1:0] node31540;
	wire [4-1:0] node31543;
	wire [4-1:0] node31545;
	wire [4-1:0] node31548;
	wire [4-1:0] node31549;
	wire [4-1:0] node31552;
	wire [4-1:0] node31554;
	wire [4-1:0] node31557;
	wire [4-1:0] node31558;
	wire [4-1:0] node31559;
	wire [4-1:0] node31560;
	wire [4-1:0] node31563;
	wire [4-1:0] node31567;
	wire [4-1:0] node31568;
	wire [4-1:0] node31570;
	wire [4-1:0] node31572;
	wire [4-1:0] node31575;
	wire [4-1:0] node31578;
	wire [4-1:0] node31579;
	wire [4-1:0] node31580;
	wire [4-1:0] node31581;
	wire [4-1:0] node31582;
	wire [4-1:0] node31584;
	wire [4-1:0] node31588;
	wire [4-1:0] node31590;
	wire [4-1:0] node31591;
	wire [4-1:0] node31594;
	wire [4-1:0] node31597;
	wire [4-1:0] node31598;
	wire [4-1:0] node31599;
	wire [4-1:0] node31601;
	wire [4-1:0] node31604;
	wire [4-1:0] node31605;
	wire [4-1:0] node31609;
	wire [4-1:0] node31610;
	wire [4-1:0] node31611;
	wire [4-1:0] node31615;
	wire [4-1:0] node31617;
	wire [4-1:0] node31618;
	wire [4-1:0] node31622;
	wire [4-1:0] node31623;
	wire [4-1:0] node31624;
	wire [4-1:0] node31625;
	wire [4-1:0] node31628;
	wire [4-1:0] node31630;
	wire [4-1:0] node31633;
	wire [4-1:0] node31634;
	wire [4-1:0] node31637;
	wire [4-1:0] node31639;
	wire [4-1:0] node31642;
	wire [4-1:0] node31643;
	wire [4-1:0] node31646;
	wire [4-1:0] node31647;
	wire [4-1:0] node31648;
	wire [4-1:0] node31653;
	wire [4-1:0] node31654;
	wire [4-1:0] node31655;
	wire [4-1:0] node31656;
	wire [4-1:0] node31657;
	wire [4-1:0] node31658;
	wire [4-1:0] node31659;
	wire [4-1:0] node31662;
	wire [4-1:0] node31665;
	wire [4-1:0] node31666;
	wire [4-1:0] node31667;
	wire [4-1:0] node31668;
	wire [4-1:0] node31672;
	wire [4-1:0] node31673;
	wire [4-1:0] node31676;
	wire [4-1:0] node31680;
	wire [4-1:0] node31681;
	wire [4-1:0] node31683;
	wire [4-1:0] node31685;
	wire [4-1:0] node31688;
	wire [4-1:0] node31691;
	wire [4-1:0] node31692;
	wire [4-1:0] node31693;
	wire [4-1:0] node31696;
	wire [4-1:0] node31699;
	wire [4-1:0] node31700;
	wire [4-1:0] node31701;
	wire [4-1:0] node31703;
	wire [4-1:0] node31706;
	wire [4-1:0] node31708;
	wire [4-1:0] node31709;
	wire [4-1:0] node31712;
	wire [4-1:0] node31715;
	wire [4-1:0] node31716;
	wire [4-1:0] node31718;
	wire [4-1:0] node31722;
	wire [4-1:0] node31723;
	wire [4-1:0] node31724;
	wire [4-1:0] node31725;
	wire [4-1:0] node31728;
	wire [4-1:0] node31730;
	wire [4-1:0] node31732;
	wire [4-1:0] node31735;
	wire [4-1:0] node31736;
	wire [4-1:0] node31737;
	wire [4-1:0] node31738;
	wire [4-1:0] node31740;
	wire [4-1:0] node31745;
	wire [4-1:0] node31747;
	wire [4-1:0] node31748;
	wire [4-1:0] node31752;
	wire [4-1:0] node31753;
	wire [4-1:0] node31754;
	wire [4-1:0] node31755;
	wire [4-1:0] node31756;
	wire [4-1:0] node31759;
	wire [4-1:0] node31762;
	wire [4-1:0] node31763;
	wire [4-1:0] node31766;
	wire [4-1:0] node31769;
	wire [4-1:0] node31771;
	wire [4-1:0] node31772;
	wire [4-1:0] node31775;
	wire [4-1:0] node31778;
	wire [4-1:0] node31780;
	wire [4-1:0] node31781;
	wire [4-1:0] node31782;
	wire [4-1:0] node31783;
	wire [4-1:0] node31787;
	wire [4-1:0] node31790;
	wire [4-1:0] node31792;
	wire [4-1:0] node31795;
	wire [4-1:0] node31796;
	wire [4-1:0] node31797;
	wire [4-1:0] node31798;
	wire [4-1:0] node31799;
	wire [4-1:0] node31800;
	wire [4-1:0] node31804;
	wire [4-1:0] node31805;
	wire [4-1:0] node31809;
	wire [4-1:0] node31810;
	wire [4-1:0] node31811;
	wire [4-1:0] node31813;
	wire [4-1:0] node31816;
	wire [4-1:0] node31818;
	wire [4-1:0] node31821;
	wire [4-1:0] node31822;
	wire [4-1:0] node31826;
	wire [4-1:0] node31827;
	wire [4-1:0] node31828;
	wire [4-1:0] node31829;
	wire [4-1:0] node31830;
	wire [4-1:0] node31834;
	wire [4-1:0] node31835;
	wire [4-1:0] node31839;
	wire [4-1:0] node31841;
	wire [4-1:0] node31844;
	wire [4-1:0] node31845;
	wire [4-1:0] node31846;
	wire [4-1:0] node31849;
	wire [4-1:0] node31850;
	wire [4-1:0] node31854;
	wire [4-1:0] node31855;
	wire [4-1:0] node31856;
	wire [4-1:0] node31859;
	wire [4-1:0] node31863;
	wire [4-1:0] node31864;
	wire [4-1:0] node31865;
	wire [4-1:0] node31866;
	wire [4-1:0] node31868;
	wire [4-1:0] node31871;
	wire [4-1:0] node31873;
	wire [4-1:0] node31876;
	wire [4-1:0] node31877;
	wire [4-1:0] node31878;
	wire [4-1:0] node31879;
	wire [4-1:0] node31882;
	wire [4-1:0] node31885;
	wire [4-1:0] node31887;
	wire [4-1:0] node31890;
	wire [4-1:0] node31891;
	wire [4-1:0] node31894;
	wire [4-1:0] node31897;
	wire [4-1:0] node31898;
	wire [4-1:0] node31899;
	wire [4-1:0] node31900;
	wire [4-1:0] node31903;
	wire [4-1:0] node31904;
	wire [4-1:0] node31908;
	wire [4-1:0] node31909;
	wire [4-1:0] node31912;
	wire [4-1:0] node31913;
	wire [4-1:0] node31917;
	wire [4-1:0] node31918;
	wire [4-1:0] node31919;
	wire [4-1:0] node31921;
	wire [4-1:0] node31925;
	wire [4-1:0] node31926;
	wire [4-1:0] node31930;
	wire [4-1:0] node31931;
	wire [4-1:0] node31932;
	wire [4-1:0] node31933;
	wire [4-1:0] node31934;
	wire [4-1:0] node31935;
	wire [4-1:0] node31936;
	wire [4-1:0] node31937;
	wire [4-1:0] node31940;
	wire [4-1:0] node31942;
	wire [4-1:0] node31945;
	wire [4-1:0] node31947;
	wire [4-1:0] node31949;
	wire [4-1:0] node31952;
	wire [4-1:0] node31953;
	wire [4-1:0] node31954;
	wire [4-1:0] node31956;
	wire [4-1:0] node31959;
	wire [4-1:0] node31961;
	wire [4-1:0] node31964;
	wire [4-1:0] node31966;
	wire [4-1:0] node31969;
	wire [4-1:0] node31970;
	wire [4-1:0] node31971;
	wire [4-1:0] node31973;
	wire [4-1:0] node31976;
	wire [4-1:0] node31977;
	wire [4-1:0] node31978;
	wire [4-1:0] node31982;
	wire [4-1:0] node31984;
	wire [4-1:0] node31987;
	wire [4-1:0] node31988;
	wire [4-1:0] node31989;
	wire [4-1:0] node31991;
	wire [4-1:0] node31995;
	wire [4-1:0] node31997;
	wire [4-1:0] node31998;
	wire [4-1:0] node32002;
	wire [4-1:0] node32003;
	wire [4-1:0] node32004;
	wire [4-1:0] node32005;
	wire [4-1:0] node32007;
	wire [4-1:0] node32009;
	wire [4-1:0] node32012;
	wire [4-1:0] node32014;
	wire [4-1:0] node32015;
	wire [4-1:0] node32018;
	wire [4-1:0] node32019;
	wire [4-1:0] node32023;
	wire [4-1:0] node32024;
	wire [4-1:0] node32025;
	wire [4-1:0] node32027;
	wire [4-1:0] node32030;
	wire [4-1:0] node32032;
	wire [4-1:0] node32035;
	wire [4-1:0] node32038;
	wire [4-1:0] node32039;
	wire [4-1:0] node32040;
	wire [4-1:0] node32041;
	wire [4-1:0] node32042;
	wire [4-1:0] node32047;
	wire [4-1:0] node32048;
	wire [4-1:0] node32050;
	wire [4-1:0] node32053;
	wire [4-1:0] node32055;
	wire [4-1:0] node32056;
	wire [4-1:0] node32060;
	wire [4-1:0] node32061;
	wire [4-1:0] node32062;
	wire [4-1:0] node32063;
	wire [4-1:0] node32066;
	wire [4-1:0] node32070;
	wire [4-1:0] node32071;
	wire [4-1:0] node32074;
	wire [4-1:0] node32077;
	wire [4-1:0] node32078;
	wire [4-1:0] node32079;
	wire [4-1:0] node32080;
	wire [4-1:0] node32081;
	wire [4-1:0] node32082;
	wire [4-1:0] node32084;
	wire [4-1:0] node32085;
	wire [4-1:0] node32090;
	wire [4-1:0] node32091;
	wire [4-1:0] node32092;
	wire [4-1:0] node32096;
	wire [4-1:0] node32097;
	wire [4-1:0] node32099;
	wire [4-1:0] node32102;
	wire [4-1:0] node32104;
	wire [4-1:0] node32107;
	wire [4-1:0] node32108;
	wire [4-1:0] node32109;
	wire [4-1:0] node32111;
	wire [4-1:0] node32114;
	wire [4-1:0] node32116;
	wire [4-1:0] node32119;
	wire [4-1:0] node32120;
	wire [4-1:0] node32124;
	wire [4-1:0] node32125;
	wire [4-1:0] node32126;
	wire [4-1:0] node32129;
	wire [4-1:0] node32130;
	wire [4-1:0] node32134;
	wire [4-1:0] node32135;
	wire [4-1:0] node32136;
	wire [4-1:0] node32140;
	wire [4-1:0] node32143;
	wire [4-1:0] node32144;
	wire [4-1:0] node32145;
	wire [4-1:0] node32146;
	wire [4-1:0] node32148;
	wire [4-1:0] node32149;
	wire [4-1:0] node32152;
	wire [4-1:0] node32155;
	wire [4-1:0] node32156;
	wire [4-1:0] node32157;
	wire [4-1:0] node32160;
	wire [4-1:0] node32163;
	wire [4-1:0] node32164;
	wire [4-1:0] node32168;
	wire [4-1:0] node32169;
	wire [4-1:0] node32171;
	wire [4-1:0] node32172;
	wire [4-1:0] node32175;
	wire [4-1:0] node32178;
	wire [4-1:0] node32179;
	wire [4-1:0] node32182;
	wire [4-1:0] node32185;
	wire [4-1:0] node32186;
	wire [4-1:0] node32187;
	wire [4-1:0] node32188;
	wire [4-1:0] node32190;
	wire [4-1:0] node32191;
	wire [4-1:0] node32194;
	wire [4-1:0] node32197;
	wire [4-1:0] node32198;
	wire [4-1:0] node32199;
	wire [4-1:0] node32202;
	wire [4-1:0] node32206;
	wire [4-1:0] node32207;
	wire [4-1:0] node32210;
	wire [4-1:0] node32213;
	wire [4-1:0] node32214;
	wire [4-1:0] node32216;
	wire [4-1:0] node32219;
	wire [4-1:0] node32220;
	wire [4-1:0] node32224;
	wire [4-1:0] node32225;
	wire [4-1:0] node32226;
	wire [4-1:0] node32227;
	wire [4-1:0] node32228;
	wire [4-1:0] node32229;
	wire [4-1:0] node32231;
	wire [4-1:0] node32235;
	wire [4-1:0] node32236;
	wire [4-1:0] node32237;
	wire [4-1:0] node32238;
	wire [4-1:0] node32240;
	wire [4-1:0] node32243;
	wire [4-1:0] node32245;
	wire [4-1:0] node32249;
	wire [4-1:0] node32251;
	wire [4-1:0] node32254;
	wire [4-1:0] node32255;
	wire [4-1:0] node32256;
	wire [4-1:0] node32257;
	wire [4-1:0] node32258;
	wire [4-1:0] node32262;
	wire [4-1:0] node32263;
	wire [4-1:0] node32266;
	wire [4-1:0] node32269;
	wire [4-1:0] node32270;
	wire [4-1:0] node32273;
	wire [4-1:0] node32274;
	wire [4-1:0] node32278;
	wire [4-1:0] node32279;
	wire [4-1:0] node32280;
	wire [4-1:0] node32281;
	wire [4-1:0] node32284;
	wire [4-1:0] node32287;
	wire [4-1:0] node32288;
	wire [4-1:0] node32292;
	wire [4-1:0] node32294;
	wire [4-1:0] node32297;
	wire [4-1:0] node32298;
	wire [4-1:0] node32299;
	wire [4-1:0] node32300;
	wire [4-1:0] node32301;
	wire [4-1:0] node32305;
	wire [4-1:0] node32306;
	wire [4-1:0] node32307;
	wire [4-1:0] node32310;
	wire [4-1:0] node32313;
	wire [4-1:0] node32314;
	wire [4-1:0] node32316;
	wire [4-1:0] node32319;
	wire [4-1:0] node32320;
	wire [4-1:0] node32323;
	wire [4-1:0] node32326;
	wire [4-1:0] node32327;
	wire [4-1:0] node32328;
	wire [4-1:0] node32331;
	wire [4-1:0] node32334;
	wire [4-1:0] node32335;
	wire [4-1:0] node32336;
	wire [4-1:0] node32340;
	wire [4-1:0] node32341;
	wire [4-1:0] node32345;
	wire [4-1:0] node32346;
	wire [4-1:0] node32349;
	wire [4-1:0] node32352;
	wire [4-1:0] node32353;
	wire [4-1:0] node32354;
	wire [4-1:0] node32355;
	wire [4-1:0] node32356;
	wire [4-1:0] node32357;
	wire [4-1:0] node32359;
	wire [4-1:0] node32363;
	wire [4-1:0] node32364;
	wire [4-1:0] node32365;
	wire [4-1:0] node32368;
	wire [4-1:0] node32372;
	wire [4-1:0] node32373;
	wire [4-1:0] node32374;
	wire [4-1:0] node32375;
	wire [4-1:0] node32378;
	wire [4-1:0] node32381;
	wire [4-1:0] node32382;
	wire [4-1:0] node32385;
	wire [4-1:0] node32388;
	wire [4-1:0] node32389;
	wire [4-1:0] node32390;
	wire [4-1:0] node32391;
	wire [4-1:0] node32395;
	wire [4-1:0] node32397;
	wire [4-1:0] node32400;
	wire [4-1:0] node32401;
	wire [4-1:0] node32405;
	wire [4-1:0] node32406;
	wire [4-1:0] node32409;
	wire [4-1:0] node32412;
	wire [4-1:0] node32413;
	wire [4-1:0] node32414;
	wire [4-1:0] node32415;
	wire [4-1:0] node32416;
	wire [4-1:0] node32419;
	wire [4-1:0] node32422;
	wire [4-1:0] node32423;
	wire [4-1:0] node32427;
	wire [4-1:0] node32428;
	wire [4-1:0] node32429;
	wire [4-1:0] node32432;
	wire [4-1:0] node32435;
	wire [4-1:0] node32437;
	wire [4-1:0] node32440;
	wire [4-1:0] node32441;
	wire [4-1:0] node32442;
	wire [4-1:0] node32445;
	wire [4-1:0] node32448;
	wire [4-1:0] node32449;
	wire [4-1:0] node32450;
	wire [4-1:0] node32452;
	wire [4-1:0] node32454;
	wire [4-1:0] node32457;
	wire [4-1:0] node32460;
	wire [4-1:0] node32461;
	wire [4-1:0] node32463;
	wire [4-1:0] node32467;
	wire [4-1:0] node32468;
	wire [4-1:0] node32469;
	wire [4-1:0] node32470;
	wire [4-1:0] node32471;
	wire [4-1:0] node32472;
	wire [4-1:0] node32473;
	wire [4-1:0] node32474;
	wire [4-1:0] node32475;
	wire [4-1:0] node32478;
	wire [4-1:0] node32479;
	wire [4-1:0] node32480;
	wire [4-1:0] node32484;
	wire [4-1:0] node32487;
	wire [4-1:0] node32489;
	wire [4-1:0] node32490;
	wire [4-1:0] node32493;
	wire [4-1:0] node32496;
	wire [4-1:0] node32497;
	wire [4-1:0] node32498;
	wire [4-1:0] node32501;
	wire [4-1:0] node32505;
	wire [4-1:0] node32506;
	wire [4-1:0] node32507;
	wire [4-1:0] node32508;
	wire [4-1:0] node32509;
	wire [4-1:0] node32513;
	wire [4-1:0] node32516;
	wire [4-1:0] node32517;
	wire [4-1:0] node32518;
	wire [4-1:0] node32522;
	wire [4-1:0] node32523;
	wire [4-1:0] node32526;
	wire [4-1:0] node32529;
	wire [4-1:0] node32530;
	wire [4-1:0] node32531;
	wire [4-1:0] node32534;
	wire [4-1:0] node32535;
	wire [4-1:0] node32537;
	wire [4-1:0] node32542;
	wire [4-1:0] node32543;
	wire [4-1:0] node32544;
	wire [4-1:0] node32545;
	wire [4-1:0] node32547;
	wire [4-1:0] node32550;
	wire [4-1:0] node32551;
	wire [4-1:0] node32553;
	wire [4-1:0] node32556;
	wire [4-1:0] node32558;
	wire [4-1:0] node32561;
	wire [4-1:0] node32562;
	wire [4-1:0] node32564;
	wire [4-1:0] node32567;
	wire [4-1:0] node32569;
	wire [4-1:0] node32570;
	wire [4-1:0] node32573;
	wire [4-1:0] node32576;
	wire [4-1:0] node32577;
	wire [4-1:0] node32578;
	wire [4-1:0] node32579;
	wire [4-1:0] node32580;
	wire [4-1:0] node32583;
	wire [4-1:0] node32586;
	wire [4-1:0] node32587;
	wire [4-1:0] node32591;
	wire [4-1:0] node32593;
	wire [4-1:0] node32595;
	wire [4-1:0] node32597;
	wire [4-1:0] node32600;
	wire [4-1:0] node32601;
	wire [4-1:0] node32602;
	wire [4-1:0] node32605;
	wire [4-1:0] node32608;
	wire [4-1:0] node32609;
	wire [4-1:0] node32613;
	wire [4-1:0] node32614;
	wire [4-1:0] node32615;
	wire [4-1:0] node32616;
	wire [4-1:0] node32617;
	wire [4-1:0] node32618;
	wire [4-1:0] node32619;
	wire [4-1:0] node32623;
	wire [4-1:0] node32624;
	wire [4-1:0] node32627;
	wire [4-1:0] node32630;
	wire [4-1:0] node32631;
	wire [4-1:0] node32632;
	wire [4-1:0] node32636;
	wire [4-1:0] node32637;
	wire [4-1:0] node32640;
	wire [4-1:0] node32643;
	wire [4-1:0] node32644;
	wire [4-1:0] node32645;
	wire [4-1:0] node32649;
	wire [4-1:0] node32651;
	wire [4-1:0] node32654;
	wire [4-1:0] node32655;
	wire [4-1:0] node32657;
	wire [4-1:0] node32658;
	wire [4-1:0] node32662;
	wire [4-1:0] node32664;
	wire [4-1:0] node32665;
	wire [4-1:0] node32669;
	wire [4-1:0] node32670;
	wire [4-1:0] node32671;
	wire [4-1:0] node32672;
	wire [4-1:0] node32673;
	wire [4-1:0] node32675;
	wire [4-1:0] node32678;
	wire [4-1:0] node32679;
	wire [4-1:0] node32680;
	wire [4-1:0] node32685;
	wire [4-1:0] node32687;
	wire [4-1:0] node32690;
	wire [4-1:0] node32691;
	wire [4-1:0] node32693;
	wire [4-1:0] node32696;
	wire [4-1:0] node32697;
	wire [4-1:0] node32699;
	wire [4-1:0] node32700;
	wire [4-1:0] node32704;
	wire [4-1:0] node32705;
	wire [4-1:0] node32708;
	wire [4-1:0] node32711;
	wire [4-1:0] node32712;
	wire [4-1:0] node32713;
	wire [4-1:0] node32715;
	wire [4-1:0] node32717;
	wire [4-1:0] node32720;
	wire [4-1:0] node32722;
	wire [4-1:0] node32723;
	wire [4-1:0] node32725;
	wire [4-1:0] node32728;
	wire [4-1:0] node32731;
	wire [4-1:0] node32732;
	wire [4-1:0] node32735;
	wire [4-1:0] node32738;
	wire [4-1:0] node32739;
	wire [4-1:0] node32740;
	wire [4-1:0] node32741;
	wire [4-1:0] node32742;
	wire [4-1:0] node32743;
	wire [4-1:0] node32744;
	wire [4-1:0] node32746;
	wire [4-1:0] node32747;
	wire [4-1:0] node32751;
	wire [4-1:0] node32752;
	wire [4-1:0] node32755;
	wire [4-1:0] node32758;
	wire [4-1:0] node32759;
	wire [4-1:0] node32760;
	wire [4-1:0] node32763;
	wire [4-1:0] node32766;
	wire [4-1:0] node32768;
	wire [4-1:0] node32771;
	wire [4-1:0] node32772;
	wire [4-1:0] node32773;
	wire [4-1:0] node32776;
	wire [4-1:0] node32778;
	wire [4-1:0] node32781;
	wire [4-1:0] node32782;
	wire [4-1:0] node32784;
	wire [4-1:0] node32786;
	wire [4-1:0] node32790;
	wire [4-1:0] node32791;
	wire [4-1:0] node32792;
	wire [4-1:0] node32795;
	wire [4-1:0] node32798;
	wire [4-1:0] node32799;
	wire [4-1:0] node32800;
	wire [4-1:0] node32802;
	wire [4-1:0] node32805;
	wire [4-1:0] node32806;
	wire [4-1:0] node32809;
	wire [4-1:0] node32810;
	wire [4-1:0] node32814;
	wire [4-1:0] node32815;
	wire [4-1:0] node32816;
	wire [4-1:0] node32819;
	wire [4-1:0] node32823;
	wire [4-1:0] node32824;
	wire [4-1:0] node32825;
	wire [4-1:0] node32826;
	wire [4-1:0] node32828;
	wire [4-1:0] node32831;
	wire [4-1:0] node32832;
	wire [4-1:0] node32833;
	wire [4-1:0] node32836;
	wire [4-1:0] node32839;
	wire [4-1:0] node32840;
	wire [4-1:0] node32844;
	wire [4-1:0] node32845;
	wire [4-1:0] node32846;
	wire [4-1:0] node32849;
	wire [4-1:0] node32850;
	wire [4-1:0] node32854;
	wire [4-1:0] node32857;
	wire [4-1:0] node32858;
	wire [4-1:0] node32859;
	wire [4-1:0] node32860;
	wire [4-1:0] node32864;
	wire [4-1:0] node32865;
	wire [4-1:0] node32868;
	wire [4-1:0] node32871;
	wire [4-1:0] node32872;
	wire [4-1:0] node32875;
	wire [4-1:0] node32876;
	wire [4-1:0] node32877;
	wire [4-1:0] node32881;
	wire [4-1:0] node32882;
	wire [4-1:0] node32886;
	wire [4-1:0] node32887;
	wire [4-1:0] node32888;
	wire [4-1:0] node32889;
	wire [4-1:0] node32890;
	wire [4-1:0] node32892;
	wire [4-1:0] node32895;
	wire [4-1:0] node32896;
	wire [4-1:0] node32897;
	wire [4-1:0] node32899;
	wire [4-1:0] node32902;
	wire [4-1:0] node32904;
	wire [4-1:0] node32908;
	wire [4-1:0] node32909;
	wire [4-1:0] node32910;
	wire [4-1:0] node32911;
	wire [4-1:0] node32915;
	wire [4-1:0] node32916;
	wire [4-1:0] node32920;
	wire [4-1:0] node32922;
	wire [4-1:0] node32923;
	wire [4-1:0] node32927;
	wire [4-1:0] node32928;
	wire [4-1:0] node32929;
	wire [4-1:0] node32932;
	wire [4-1:0] node32933;
	wire [4-1:0] node32936;
	wire [4-1:0] node32937;
	wire [4-1:0] node32941;
	wire [4-1:0] node32942;
	wire [4-1:0] node32943;
	wire [4-1:0] node32944;
	wire [4-1:0] node32948;
	wire [4-1:0] node32951;
	wire [4-1:0] node32952;
	wire [4-1:0] node32955;
	wire [4-1:0] node32956;
	wire [4-1:0] node32960;
	wire [4-1:0] node32961;
	wire [4-1:0] node32962;
	wire [4-1:0] node32963;
	wire [4-1:0] node32965;
	wire [4-1:0] node32968;
	wire [4-1:0] node32970;
	wire [4-1:0] node32973;
	wire [4-1:0] node32974;
	wire [4-1:0] node32975;
	wire [4-1:0] node32977;
	wire [4-1:0] node32980;
	wire [4-1:0] node32982;
	wire [4-1:0] node32985;
	wire [4-1:0] node32987;
	wire [4-1:0] node32990;
	wire [4-1:0] node32991;
	wire [4-1:0] node32993;
	wire [4-1:0] node32996;
	wire [4-1:0] node32997;
	wire [4-1:0] node32998;
	wire [4-1:0] node33002;
	wire [4-1:0] node33003;
	wire [4-1:0] node33007;
	wire [4-1:0] node33008;
	wire [4-1:0] node33009;
	wire [4-1:0] node33010;
	wire [4-1:0] node33011;
	wire [4-1:0] node33012;
	wire [4-1:0] node33013;
	wire [4-1:0] node33014;
	wire [4-1:0] node33015;
	wire [4-1:0] node33017;
	wire [4-1:0] node33020;
	wire [4-1:0] node33021;
	wire [4-1:0] node33025;
	wire [4-1:0] node33026;
	wire [4-1:0] node33029;
	wire [4-1:0] node33032;
	wire [4-1:0] node33033;
	wire [4-1:0] node33035;
	wire [4-1:0] node33039;
	wire [4-1:0] node33040;
	wire [4-1:0] node33041;
	wire [4-1:0] node33042;
	wire [4-1:0] node33046;
	wire [4-1:0] node33047;
	wire [4-1:0] node33051;
	wire [4-1:0] node33052;
	wire [4-1:0] node33054;
	wire [4-1:0] node33057;
	wire [4-1:0] node33058;
	wire [4-1:0] node33062;
	wire [4-1:0] node33063;
	wire [4-1:0] node33064;
	wire [4-1:0] node33066;
	wire [4-1:0] node33068;
	wire [4-1:0] node33071;
	wire [4-1:0] node33072;
	wire [4-1:0] node33074;
	wire [4-1:0] node33075;
	wire [4-1:0] node33079;
	wire [4-1:0] node33080;
	wire [4-1:0] node33083;
	wire [4-1:0] node33086;
	wire [4-1:0] node33087;
	wire [4-1:0] node33089;
	wire [4-1:0] node33090;
	wire [4-1:0] node33093;
	wire [4-1:0] node33096;
	wire [4-1:0] node33097;
	wire [4-1:0] node33098;
	wire [4-1:0] node33101;
	wire [4-1:0] node33104;
	wire [4-1:0] node33107;
	wire [4-1:0] node33108;
	wire [4-1:0] node33109;
	wire [4-1:0] node33110;
	wire [4-1:0] node33111;
	wire [4-1:0] node33113;
	wire [4-1:0] node33116;
	wire [4-1:0] node33117;
	wire [4-1:0] node33118;
	wire [4-1:0] node33123;
	wire [4-1:0] node33124;
	wire [4-1:0] node33125;
	wire [4-1:0] node33129;
	wire [4-1:0] node33131;
	wire [4-1:0] node33132;
	wire [4-1:0] node33135;
	wire [4-1:0] node33138;
	wire [4-1:0] node33139;
	wire [4-1:0] node33140;
	wire [4-1:0] node33143;
	wire [4-1:0] node33144;
	wire [4-1:0] node33147;
	wire [4-1:0] node33148;
	wire [4-1:0] node33152;
	wire [4-1:0] node33153;
	wire [4-1:0] node33155;
	wire [4-1:0] node33158;
	wire [4-1:0] node33160;
	wire [4-1:0] node33162;
	wire [4-1:0] node33165;
	wire [4-1:0] node33166;
	wire [4-1:0] node33167;
	wire [4-1:0] node33168;
	wire [4-1:0] node33169;
	wire [4-1:0] node33170;
	wire [4-1:0] node33173;
	wire [4-1:0] node33177;
	wire [4-1:0] node33180;
	wire [4-1:0] node33181;
	wire [4-1:0] node33182;
	wire [4-1:0] node33183;
	wire [4-1:0] node33186;
	wire [4-1:0] node33189;
	wire [4-1:0] node33190;
	wire [4-1:0] node33194;
	wire [4-1:0] node33195;
	wire [4-1:0] node33198;
	wire [4-1:0] node33201;
	wire [4-1:0] node33202;
	wire [4-1:0] node33203;
	wire [4-1:0] node33204;
	wire [4-1:0] node33206;
	wire [4-1:0] node33210;
	wire [4-1:0] node33211;
	wire [4-1:0] node33215;
	wire [4-1:0] node33216;
	wire [4-1:0] node33220;
	wire [4-1:0] node33221;
	wire [4-1:0] node33222;
	wire [4-1:0] node33223;
	wire [4-1:0] node33224;
	wire [4-1:0] node33225;
	wire [4-1:0] node33228;
	wire [4-1:0] node33231;
	wire [4-1:0] node33232;
	wire [4-1:0] node33233;
	wire [4-1:0] node33236;
	wire [4-1:0] node33238;
	wire [4-1:0] node33242;
	wire [4-1:0] node33243;
	wire [4-1:0] node33246;
	wire [4-1:0] node33249;
	wire [4-1:0] node33250;
	wire [4-1:0] node33251;
	wire [4-1:0] node33254;
	wire [4-1:0] node33257;
	wire [4-1:0] node33258;
	wire [4-1:0] node33261;
	wire [4-1:0] node33264;
	wire [4-1:0] node33265;
	wire [4-1:0] node33266;
	wire [4-1:0] node33267;
	wire [4-1:0] node33270;
	wire [4-1:0] node33273;
	wire [4-1:0] node33274;
	wire [4-1:0] node33275;
	wire [4-1:0] node33278;
	wire [4-1:0] node33282;
	wire [4-1:0] node33283;
	wire [4-1:0] node33284;
	wire [4-1:0] node33286;
	wire [4-1:0] node33288;
	wire [4-1:0] node33291;
	wire [4-1:0] node33292;
	wire [4-1:0] node33295;
	wire [4-1:0] node33298;
	wire [4-1:0] node33299;
	wire [4-1:0] node33302;
	wire [4-1:0] node33305;
	wire [4-1:0] node33306;
	wire [4-1:0] node33307;
	wire [4-1:0] node33308;
	wire [4-1:0] node33309;
	wire [4-1:0] node33310;
	wire [4-1:0] node33311;
	wire [4-1:0] node33312;
	wire [4-1:0] node33316;
	wire [4-1:0] node33318;
	wire [4-1:0] node33321;
	wire [4-1:0] node33322;
	wire [4-1:0] node33323;
	wire [4-1:0] node33325;
	wire [4-1:0] node33330;
	wire [4-1:0] node33331;
	wire [4-1:0] node33332;
	wire [4-1:0] node33333;
	wire [4-1:0] node33334;
	wire [4-1:0] node33337;
	wire [4-1:0] node33341;
	wire [4-1:0] node33343;
	wire [4-1:0] node33346;
	wire [4-1:0] node33348;
	wire [4-1:0] node33350;
	wire [4-1:0] node33351;
	wire [4-1:0] node33354;
	wire [4-1:0] node33357;
	wire [4-1:0] node33358;
	wire [4-1:0] node33359;
	wire [4-1:0] node33360;
	wire [4-1:0] node33361;
	wire [4-1:0] node33365;
	wire [4-1:0] node33367;
	wire [4-1:0] node33370;
	wire [4-1:0] node33371;
	wire [4-1:0] node33372;
	wire [4-1:0] node33373;
	wire [4-1:0] node33378;
	wire [4-1:0] node33379;
	wire [4-1:0] node33381;
	wire [4-1:0] node33384;
	wire [4-1:0] node33387;
	wire [4-1:0] node33388;
	wire [4-1:0] node33390;
	wire [4-1:0] node33391;
	wire [4-1:0] node33395;
	wire [4-1:0] node33396;
	wire [4-1:0] node33398;
	wire [4-1:0] node33401;
	wire [4-1:0] node33402;
	wire [4-1:0] node33405;
	wire [4-1:0] node33408;
	wire [4-1:0] node33409;
	wire [4-1:0] node33410;
	wire [4-1:0] node33411;
	wire [4-1:0] node33412;
	wire [4-1:0] node33414;
	wire [4-1:0] node33417;
	wire [4-1:0] node33418;
	wire [4-1:0] node33421;
	wire [4-1:0] node33424;
	wire [4-1:0] node33425;
	wire [4-1:0] node33426;
	wire [4-1:0] node33430;
	wire [4-1:0] node33433;
	wire [4-1:0] node33434;
	wire [4-1:0] node33435;
	wire [4-1:0] node33436;
	wire [4-1:0] node33439;
	wire [4-1:0] node33443;
	wire [4-1:0] node33444;
	wire [4-1:0] node33445;
	wire [4-1:0] node33449;
	wire [4-1:0] node33452;
	wire [4-1:0] node33453;
	wire [4-1:0] node33455;
	wire [4-1:0] node33456;
	wire [4-1:0] node33459;
	wire [4-1:0] node33460;
	wire [4-1:0] node33463;
	wire [4-1:0] node33466;
	wire [4-1:0] node33467;
	wire [4-1:0] node33468;
	wire [4-1:0] node33470;
	wire [4-1:0] node33473;
	wire [4-1:0] node33476;
	wire [4-1:0] node33477;
	wire [4-1:0] node33479;
	wire [4-1:0] node33481;
	wire [4-1:0] node33484;
	wire [4-1:0] node33485;
	wire [4-1:0] node33489;
	wire [4-1:0] node33490;
	wire [4-1:0] node33491;
	wire [4-1:0] node33492;
	wire [4-1:0] node33493;
	wire [4-1:0] node33495;
	wire [4-1:0] node33496;
	wire [4-1:0] node33500;
	wire [4-1:0] node33501;
	wire [4-1:0] node33505;
	wire [4-1:0] node33506;
	wire [4-1:0] node33507;
	wire [4-1:0] node33508;
	wire [4-1:0] node33511;
	wire [4-1:0] node33514;
	wire [4-1:0] node33516;
	wire [4-1:0] node33519;
	wire [4-1:0] node33521;
	wire [4-1:0] node33524;
	wire [4-1:0] node33525;
	wire [4-1:0] node33526;
	wire [4-1:0] node33527;
	wire [4-1:0] node33528;
	wire [4-1:0] node33529;
	wire [4-1:0] node33533;
	wire [4-1:0] node33535;
	wire [4-1:0] node33538;
	wire [4-1:0] node33541;
	wire [4-1:0] node33542;
	wire [4-1:0] node33546;
	wire [4-1:0] node33547;
	wire [4-1:0] node33548;
	wire [4-1:0] node33551;
	wire [4-1:0] node33554;
	wire [4-1:0] node33555;
	wire [4-1:0] node33558;
	wire [4-1:0] node33561;
	wire [4-1:0] node33562;
	wire [4-1:0] node33563;
	wire [4-1:0] node33565;
	wire [4-1:0] node33566;
	wire [4-1:0] node33569;
	wire [4-1:0] node33572;
	wire [4-1:0] node33573;
	wire [4-1:0] node33576;
	wire [4-1:0] node33579;
	wire [4-1:0] node33580;
	wire [4-1:0] node33581;
	wire [4-1:0] node33582;
	wire [4-1:0] node33585;
	wire [4-1:0] node33588;
	wire [4-1:0] node33589;
	wire [4-1:0] node33590;
	wire [4-1:0] node33593;
	wire [4-1:0] node33596;
	wire [4-1:0] node33598;
	wire [4-1:0] node33601;
	wire [4-1:0] node33602;
	wire [4-1:0] node33604;
	wire [4-1:0] node33607;
	wire [4-1:0] node33608;
	wire [4-1:0] node33612;
	wire [4-1:0] node33613;
	wire [4-1:0] node33614;
	wire [4-1:0] node33615;
	wire [4-1:0] node33616;
	wire [4-1:0] node33617;
	wire [4-1:0] node33618;
	wire [4-1:0] node33619;
	wire [4-1:0] node33620;
	wire [4-1:0] node33621;
	wire [4-1:0] node33622;
	wire [4-1:0] node33623;
	wire [4-1:0] node33627;
	wire [4-1:0] node33628;
	wire [4-1:0] node33630;
	wire [4-1:0] node33633;
	wire [4-1:0] node33635;
	wire [4-1:0] node33636;
	wire [4-1:0] node33640;
	wire [4-1:0] node33641;
	wire [4-1:0] node33642;
	wire [4-1:0] node33645;
	wire [4-1:0] node33648;
	wire [4-1:0] node33651;
	wire [4-1:0] node33652;
	wire [4-1:0] node33653;
	wire [4-1:0] node33654;
	wire [4-1:0] node33657;
	wire [4-1:0] node33660;
	wire [4-1:0] node33661;
	wire [4-1:0] node33662;
	wire [4-1:0] node33664;
	wire [4-1:0] node33669;
	wire [4-1:0] node33670;
	wire [4-1:0] node33671;
	wire [4-1:0] node33672;
	wire [4-1:0] node33673;
	wire [4-1:0] node33676;
	wire [4-1:0] node33679;
	wire [4-1:0] node33681;
	wire [4-1:0] node33685;
	wire [4-1:0] node33686;
	wire [4-1:0] node33688;
	wire [4-1:0] node33689;
	wire [4-1:0] node33692;
	wire [4-1:0] node33695;
	wire [4-1:0] node33696;
	wire [4-1:0] node33699;
	wire [4-1:0] node33702;
	wire [4-1:0] node33703;
	wire [4-1:0] node33704;
	wire [4-1:0] node33705;
	wire [4-1:0] node33706;
	wire [4-1:0] node33708;
	wire [4-1:0] node33711;
	wire [4-1:0] node33713;
	wire [4-1:0] node33716;
	wire [4-1:0] node33717;
	wire [4-1:0] node33718;
	wire [4-1:0] node33722;
	wire [4-1:0] node33723;
	wire [4-1:0] node33726;
	wire [4-1:0] node33729;
	wire [4-1:0] node33730;
	wire [4-1:0] node33731;
	wire [4-1:0] node33734;
	wire [4-1:0] node33736;
	wire [4-1:0] node33739;
	wire [4-1:0] node33740;
	wire [4-1:0] node33743;
	wire [4-1:0] node33746;
	wire [4-1:0] node33747;
	wire [4-1:0] node33748;
	wire [4-1:0] node33749;
	wire [4-1:0] node33750;
	wire [4-1:0] node33754;
	wire [4-1:0] node33756;
	wire [4-1:0] node33758;
	wire [4-1:0] node33761;
	wire [4-1:0] node33762;
	wire [4-1:0] node33763;
	wire [4-1:0] node33766;
	wire [4-1:0] node33770;
	wire [4-1:0] node33771;
	wire [4-1:0] node33772;
	wire [4-1:0] node33775;
	wire [4-1:0] node33777;
	wire [4-1:0] node33780;
	wire [4-1:0] node33781;
	wire [4-1:0] node33784;
	wire [4-1:0] node33786;
	wire [4-1:0] node33787;
	wire [4-1:0] node33791;
	wire [4-1:0] node33792;
	wire [4-1:0] node33793;
	wire [4-1:0] node33794;
	wire [4-1:0] node33795;
	wire [4-1:0] node33796;
	wire [4-1:0] node33800;
	wire [4-1:0] node33801;
	wire [4-1:0] node33802;
	wire [4-1:0] node33805;
	wire [4-1:0] node33808;
	wire [4-1:0] node33810;
	wire [4-1:0] node33811;
	wire [4-1:0] node33814;
	wire [4-1:0] node33817;
	wire [4-1:0] node33818;
	wire [4-1:0] node33821;
	wire [4-1:0] node33822;
	wire [4-1:0] node33824;
	wire [4-1:0] node33827;
	wire [4-1:0] node33828;
	wire [4-1:0] node33832;
	wire [4-1:0] node33833;
	wire [4-1:0] node33834;
	wire [4-1:0] node33835;
	wire [4-1:0] node33837;
	wire [4-1:0] node33840;
	wire [4-1:0] node33841;
	wire [4-1:0] node33845;
	wire [4-1:0] node33846;
	wire [4-1:0] node33847;
	wire [4-1:0] node33852;
	wire [4-1:0] node33853;
	wire [4-1:0] node33855;
	wire [4-1:0] node33856;
	wire [4-1:0] node33860;
	wire [4-1:0] node33862;
	wire [4-1:0] node33864;
	wire [4-1:0] node33865;
	wire [4-1:0] node33869;
	wire [4-1:0] node33870;
	wire [4-1:0] node33871;
	wire [4-1:0] node33872;
	wire [4-1:0] node33873;
	wire [4-1:0] node33874;
	wire [4-1:0] node33878;
	wire [4-1:0] node33879;
	wire [4-1:0] node33882;
	wire [4-1:0] node33885;
	wire [4-1:0] node33886;
	wire [4-1:0] node33889;
	wire [4-1:0] node33892;
	wire [4-1:0] node33893;
	wire [4-1:0] node33894;
	wire [4-1:0] node33896;
	wire [4-1:0] node33897;
	wire [4-1:0] node33901;
	wire [4-1:0] node33903;
	wire [4-1:0] node33904;
	wire [4-1:0] node33907;
	wire [4-1:0] node33910;
	wire [4-1:0] node33911;
	wire [4-1:0] node33912;
	wire [4-1:0] node33916;
	wire [4-1:0] node33917;
	wire [4-1:0] node33918;
	wire [4-1:0] node33921;
	wire [4-1:0] node33925;
	wire [4-1:0] node33926;
	wire [4-1:0] node33927;
	wire [4-1:0] node33928;
	wire [4-1:0] node33931;
	wire [4-1:0] node33934;
	wire [4-1:0] node33935;
	wire [4-1:0] node33936;
	wire [4-1:0] node33940;
	wire [4-1:0] node33943;
	wire [4-1:0] node33944;
	wire [4-1:0] node33945;
	wire [4-1:0] node33946;
	wire [4-1:0] node33950;
	wire [4-1:0] node33952;
	wire [4-1:0] node33955;
	wire [4-1:0] node33956;
	wire [4-1:0] node33958;
	wire [4-1:0] node33959;
	wire [4-1:0] node33962;
	wire [4-1:0] node33966;
	wire [4-1:0] node33967;
	wire [4-1:0] node33968;
	wire [4-1:0] node33969;
	wire [4-1:0] node33970;
	wire [4-1:0] node33971;
	wire [4-1:0] node33973;
	wire [4-1:0] node33974;
	wire [4-1:0] node33977;
	wire [4-1:0] node33980;
	wire [4-1:0] node33982;
	wire [4-1:0] node33984;
	wire [4-1:0] node33987;
	wire [4-1:0] node33988;
	wire [4-1:0] node33989;
	wire [4-1:0] node33992;
	wire [4-1:0] node33993;
	wire [4-1:0] node33997;
	wire [4-1:0] node33998;
	wire [4-1:0] node33999;
	wire [4-1:0] node34002;
	wire [4-1:0] node34005;
	wire [4-1:0] node34006;
	wire [4-1:0] node34009;
	wire [4-1:0] node34012;
	wire [4-1:0] node34013;
	wire [4-1:0] node34014;
	wire [4-1:0] node34016;
	wire [4-1:0] node34017;
	wire [4-1:0] node34020;
	wire [4-1:0] node34023;
	wire [4-1:0] node34024;
	wire [4-1:0] node34025;
	wire [4-1:0] node34029;
	wire [4-1:0] node34032;
	wire [4-1:0] node34033;
	wire [4-1:0] node34036;
	wire [4-1:0] node34038;
	wire [4-1:0] node34039;
	wire [4-1:0] node34043;
	wire [4-1:0] node34044;
	wire [4-1:0] node34045;
	wire [4-1:0] node34046;
	wire [4-1:0] node34047;
	wire [4-1:0] node34050;
	wire [4-1:0] node34053;
	wire [4-1:0] node34054;
	wire [4-1:0] node34057;
	wire [4-1:0] node34059;
	wire [4-1:0] node34062;
	wire [4-1:0] node34063;
	wire [4-1:0] node34065;
	wire [4-1:0] node34066;
	wire [4-1:0] node34069;
	wire [4-1:0] node34072;
	wire [4-1:0] node34073;
	wire [4-1:0] node34074;
	wire [4-1:0] node34077;
	wire [4-1:0] node34081;
	wire [4-1:0] node34082;
	wire [4-1:0] node34083;
	wire [4-1:0] node34084;
	wire [4-1:0] node34088;
	wire [4-1:0] node34089;
	wire [4-1:0] node34090;
	wire [4-1:0] node34094;
	wire [4-1:0] node34095;
	wire [4-1:0] node34099;
	wire [4-1:0] node34100;
	wire [4-1:0] node34101;
	wire [4-1:0] node34104;
	wire [4-1:0] node34107;
	wire [4-1:0] node34108;
	wire [4-1:0] node34109;
	wire [4-1:0] node34110;
	wire [4-1:0] node34114;
	wire [4-1:0] node34115;
	wire [4-1:0] node34119;
	wire [4-1:0] node34122;
	wire [4-1:0] node34123;
	wire [4-1:0] node34124;
	wire [4-1:0] node34125;
	wire [4-1:0] node34127;
	wire [4-1:0] node34128;
	wire [4-1:0] node34131;
	wire [4-1:0] node34134;
	wire [4-1:0] node34135;
	wire [4-1:0] node34136;
	wire [4-1:0] node34137;
	wire [4-1:0] node34140;
	wire [4-1:0] node34141;
	wire [4-1:0] node34145;
	wire [4-1:0] node34147;
	wire [4-1:0] node34150;
	wire [4-1:0] node34151;
	wire [4-1:0] node34154;
	wire [4-1:0] node34155;
	wire [4-1:0] node34156;
	wire [4-1:0] node34160;
	wire [4-1:0] node34163;
	wire [4-1:0] node34164;
	wire [4-1:0] node34165;
	wire [4-1:0] node34166;
	wire [4-1:0] node34167;
	wire [4-1:0] node34170;
	wire [4-1:0] node34173;
	wire [4-1:0] node34174;
	wire [4-1:0] node34177;
	wire [4-1:0] node34180;
	wire [4-1:0] node34181;
	wire [4-1:0] node34184;
	wire [4-1:0] node34186;
	wire [4-1:0] node34189;
	wire [4-1:0] node34190;
	wire [4-1:0] node34191;
	wire [4-1:0] node34194;
	wire [4-1:0] node34197;
	wire [4-1:0] node34198;
	wire [4-1:0] node34201;
	wire [4-1:0] node34204;
	wire [4-1:0] node34205;
	wire [4-1:0] node34206;
	wire [4-1:0] node34207;
	wire [4-1:0] node34208;
	wire [4-1:0] node34209;
	wire [4-1:0] node34213;
	wire [4-1:0] node34214;
	wire [4-1:0] node34217;
	wire [4-1:0] node34218;
	wire [4-1:0] node34222;
	wire [4-1:0] node34223;
	wire [4-1:0] node34227;
	wire [4-1:0] node34228;
	wire [4-1:0] node34230;
	wire [4-1:0] node34232;
	wire [4-1:0] node34235;
	wire [4-1:0] node34236;
	wire [4-1:0] node34237;
	wire [4-1:0] node34239;
	wire [4-1:0] node34243;
	wire [4-1:0] node34244;
	wire [4-1:0] node34246;
	wire [4-1:0] node34249;
	wire [4-1:0] node34250;
	wire [4-1:0] node34253;
	wire [4-1:0] node34256;
	wire [4-1:0] node34257;
	wire [4-1:0] node34258;
	wire [4-1:0] node34262;
	wire [4-1:0] node34263;
	wire [4-1:0] node34265;
	wire [4-1:0] node34268;
	wire [4-1:0] node34271;
	wire [4-1:0] node34272;
	wire [4-1:0] node34273;
	wire [4-1:0] node34274;
	wire [4-1:0] node34275;
	wire [4-1:0] node34276;
	wire [4-1:0] node34277;
	wire [4-1:0] node34278;
	wire [4-1:0] node34280;
	wire [4-1:0] node34283;
	wire [4-1:0] node34285;
	wire [4-1:0] node34288;
	wire [4-1:0] node34289;
	wire [4-1:0] node34292;
	wire [4-1:0] node34293;
	wire [4-1:0] node34294;
	wire [4-1:0] node34299;
	wire [4-1:0] node34300;
	wire [4-1:0] node34301;
	wire [4-1:0] node34302;
	wire [4-1:0] node34306;
	wire [4-1:0] node34308;
	wire [4-1:0] node34311;
	wire [4-1:0] node34312;
	wire [4-1:0] node34314;
	wire [4-1:0] node34315;
	wire [4-1:0] node34319;
	wire [4-1:0] node34320;
	wire [4-1:0] node34321;
	wire [4-1:0] node34324;
	wire [4-1:0] node34327;
	wire [4-1:0] node34329;
	wire [4-1:0] node34332;
	wire [4-1:0] node34333;
	wire [4-1:0] node34334;
	wire [4-1:0] node34335;
	wire [4-1:0] node34337;
	wire [4-1:0] node34338;
	wire [4-1:0] node34341;
	wire [4-1:0] node34344;
	wire [4-1:0] node34345;
	wire [4-1:0] node34346;
	wire [4-1:0] node34350;
	wire [4-1:0] node34351;
	wire [4-1:0] node34354;
	wire [4-1:0] node34357;
	wire [4-1:0] node34358;
	wire [4-1:0] node34359;
	wire [4-1:0] node34364;
	wire [4-1:0] node34365;
	wire [4-1:0] node34366;
	wire [4-1:0] node34367;
	wire [4-1:0] node34371;
	wire [4-1:0] node34372;
	wire [4-1:0] node34376;
	wire [4-1:0] node34377;
	wire [4-1:0] node34378;
	wire [4-1:0] node34379;
	wire [4-1:0] node34385;
	wire [4-1:0] node34386;
	wire [4-1:0] node34387;
	wire [4-1:0] node34388;
	wire [4-1:0] node34390;
	wire [4-1:0] node34393;
	wire [4-1:0] node34394;
	wire [4-1:0] node34395;
	wire [4-1:0] node34398;
	wire [4-1:0] node34402;
	wire [4-1:0] node34403;
	wire [4-1:0] node34405;
	wire [4-1:0] node34407;
	wire [4-1:0] node34408;
	wire [4-1:0] node34413;
	wire [4-1:0] node34414;
	wire [4-1:0] node34415;
	wire [4-1:0] node34416;
	wire [4-1:0] node34417;
	wire [4-1:0] node34420;
	wire [4-1:0] node34423;
	wire [4-1:0] node34424;
	wire [4-1:0] node34427;
	wire [4-1:0] node34430;
	wire [4-1:0] node34432;
	wire [4-1:0] node34433;
	wire [4-1:0] node34437;
	wire [4-1:0] node34438;
	wire [4-1:0] node34439;
	wire [4-1:0] node34440;
	wire [4-1:0] node34445;
	wire [4-1:0] node34446;
	wire [4-1:0] node34448;
	wire [4-1:0] node34452;
	wire [4-1:0] node34453;
	wire [4-1:0] node34454;
	wire [4-1:0] node34455;
	wire [4-1:0] node34456;
	wire [4-1:0] node34457;
	wire [4-1:0] node34459;
	wire [4-1:0] node34462;
	wire [4-1:0] node34463;
	wire [4-1:0] node34466;
	wire [4-1:0] node34469;
	wire [4-1:0] node34470;
	wire [4-1:0] node34471;
	wire [4-1:0] node34474;
	wire [4-1:0] node34478;
	wire [4-1:0] node34479;
	wire [4-1:0] node34481;
	wire [4-1:0] node34482;
	wire [4-1:0] node34486;
	wire [4-1:0] node34488;
	wire [4-1:0] node34489;
	wire [4-1:0] node34493;
	wire [4-1:0] node34494;
	wire [4-1:0] node34495;
	wire [4-1:0] node34496;
	wire [4-1:0] node34497;
	wire [4-1:0] node34502;
	wire [4-1:0] node34503;
	wire [4-1:0] node34504;
	wire [4-1:0] node34507;
	wire [4-1:0] node34510;
	wire [4-1:0] node34512;
	wire [4-1:0] node34515;
	wire [4-1:0] node34516;
	wire [4-1:0] node34517;
	wire [4-1:0] node34518;
	wire [4-1:0] node34522;
	wire [4-1:0] node34523;
	wire [4-1:0] node34526;
	wire [4-1:0] node34529;
	wire [4-1:0] node34530;
	wire [4-1:0] node34531;
	wire [4-1:0] node34535;
	wire [4-1:0] node34536;
	wire [4-1:0] node34539;
	wire [4-1:0] node34542;
	wire [4-1:0] node34543;
	wire [4-1:0] node34544;
	wire [4-1:0] node34545;
	wire [4-1:0] node34546;
	wire [4-1:0] node34548;
	wire [4-1:0] node34549;
	wire [4-1:0] node34552;
	wire [4-1:0] node34555;
	wire [4-1:0] node34556;
	wire [4-1:0] node34559;
	wire [4-1:0] node34562;
	wire [4-1:0] node34563;
	wire [4-1:0] node34565;
	wire [4-1:0] node34568;
	wire [4-1:0] node34569;
	wire [4-1:0] node34572;
	wire [4-1:0] node34575;
	wire [4-1:0] node34576;
	wire [4-1:0] node34577;
	wire [4-1:0] node34581;
	wire [4-1:0] node34582;
	wire [4-1:0] node34583;
	wire [4-1:0] node34584;
	wire [4-1:0] node34589;
	wire [4-1:0] node34590;
	wire [4-1:0] node34592;
	wire [4-1:0] node34595;
	wire [4-1:0] node34596;
	wire [4-1:0] node34600;
	wire [4-1:0] node34601;
	wire [4-1:0] node34602;
	wire [4-1:0] node34604;
	wire [4-1:0] node34605;
	wire [4-1:0] node34607;
	wire [4-1:0] node34611;
	wire [4-1:0] node34612;
	wire [4-1:0] node34613;
	wire [4-1:0] node34617;
	wire [4-1:0] node34618;
	wire [4-1:0] node34620;
	wire [4-1:0] node34624;
	wire [4-1:0] node34625;
	wire [4-1:0] node34626;
	wire [4-1:0] node34627;
	wire [4-1:0] node34631;
	wire [4-1:0] node34633;
	wire [4-1:0] node34636;
	wire [4-1:0] node34637;
	wire [4-1:0] node34638;
	wire [4-1:0] node34639;
	wire [4-1:0] node34643;
	wire [4-1:0] node34646;
	wire [4-1:0] node34647;
	wire [4-1:0] node34648;
	wire [4-1:0] node34653;
	wire [4-1:0] node34654;
	wire [4-1:0] node34655;
	wire [4-1:0] node34656;
	wire [4-1:0] node34657;
	wire [4-1:0] node34658;
	wire [4-1:0] node34659;
	wire [4-1:0] node34661;
	wire [4-1:0] node34664;
	wire [4-1:0] node34666;
	wire [4-1:0] node34668;
	wire [4-1:0] node34671;
	wire [4-1:0] node34672;
	wire [4-1:0] node34673;
	wire [4-1:0] node34674;
	wire [4-1:0] node34677;
	wire [4-1:0] node34680;
	wire [4-1:0] node34682;
	wire [4-1:0] node34685;
	wire [4-1:0] node34686;
	wire [4-1:0] node34687;
	wire [4-1:0] node34690;
	wire [4-1:0] node34694;
	wire [4-1:0] node34695;
	wire [4-1:0] node34697;
	wire [4-1:0] node34698;
	wire [4-1:0] node34701;
	wire [4-1:0] node34704;
	wire [4-1:0] node34705;
	wire [4-1:0] node34707;
	wire [4-1:0] node34710;
	wire [4-1:0] node34711;
	wire [4-1:0] node34715;
	wire [4-1:0] node34716;
	wire [4-1:0] node34717;
	wire [4-1:0] node34718;
	wire [4-1:0] node34719;
	wire [4-1:0] node34724;
	wire [4-1:0] node34725;
	wire [4-1:0] node34726;
	wire [4-1:0] node34728;
	wire [4-1:0] node34733;
	wire [4-1:0] node34734;
	wire [4-1:0] node34736;
	wire [4-1:0] node34737;
	wire [4-1:0] node34740;
	wire [4-1:0] node34743;
	wire [4-1:0] node34744;
	wire [4-1:0] node34745;
	wire [4-1:0] node34748;
	wire [4-1:0] node34751;
	wire [4-1:0] node34754;
	wire [4-1:0] node34755;
	wire [4-1:0] node34756;
	wire [4-1:0] node34757;
	wire [4-1:0] node34760;
	wire [4-1:0] node34761;
	wire [4-1:0] node34762;
	wire [4-1:0] node34764;
	wire [4-1:0] node34767;
	wire [4-1:0] node34768;
	wire [4-1:0] node34771;
	wire [4-1:0] node34774;
	wire [4-1:0] node34775;
	wire [4-1:0] node34779;
	wire [4-1:0] node34780;
	wire [4-1:0] node34781;
	wire [4-1:0] node34782;
	wire [4-1:0] node34785;
	wire [4-1:0] node34788;
	wire [4-1:0] node34789;
	wire [4-1:0] node34793;
	wire [4-1:0] node34794;
	wire [4-1:0] node34796;
	wire [4-1:0] node34799;
	wire [4-1:0] node34800;
	wire [4-1:0] node34804;
	wire [4-1:0] node34805;
	wire [4-1:0] node34806;
	wire [4-1:0] node34807;
	wire [4-1:0] node34808;
	wire [4-1:0] node34810;
	wire [4-1:0] node34814;
	wire [4-1:0] node34815;
	wire [4-1:0] node34818;
	wire [4-1:0] node34819;
	wire [4-1:0] node34823;
	wire [4-1:0] node34824;
	wire [4-1:0] node34825;
	wire [4-1:0] node34826;
	wire [4-1:0] node34831;
	wire [4-1:0] node34832;
	wire [4-1:0] node34836;
	wire [4-1:0] node34837;
	wire [4-1:0] node34838;
	wire [4-1:0] node34841;
	wire [4-1:0] node34844;
	wire [4-1:0] node34845;
	wire [4-1:0] node34848;
	wire [4-1:0] node34851;
	wire [4-1:0] node34852;
	wire [4-1:0] node34853;
	wire [4-1:0] node34854;
	wire [4-1:0] node34855;
	wire [4-1:0] node34856;
	wire [4-1:0] node34858;
	wire [4-1:0] node34862;
	wire [4-1:0] node34863;
	wire [4-1:0] node34864;
	wire [4-1:0] node34867;
	wire [4-1:0] node34870;
	wire [4-1:0] node34872;
	wire [4-1:0] node34875;
	wire [4-1:0] node34876;
	wire [4-1:0] node34877;
	wire [4-1:0] node34878;
	wire [4-1:0] node34882;
	wire [4-1:0] node34884;
	wire [4-1:0] node34887;
	wire [4-1:0] node34888;
	wire [4-1:0] node34889;
	wire [4-1:0] node34893;
	wire [4-1:0] node34896;
	wire [4-1:0] node34897;
	wire [4-1:0] node34898;
	wire [4-1:0] node34900;
	wire [4-1:0] node34903;
	wire [4-1:0] node34904;
	wire [4-1:0] node34908;
	wire [4-1:0] node34909;
	wire [4-1:0] node34910;
	wire [4-1:0] node34912;
	wire [4-1:0] node34915;
	wire [4-1:0] node34916;
	wire [4-1:0] node34919;
	wire [4-1:0] node34921;
	wire [4-1:0] node34924;
	wire [4-1:0] node34926;
	wire [4-1:0] node34929;
	wire [4-1:0] node34930;
	wire [4-1:0] node34931;
	wire [4-1:0] node34932;
	wire [4-1:0] node34933;
	wire [4-1:0] node34936;
	wire [4-1:0] node34939;
	wire [4-1:0] node34940;
	wire [4-1:0] node34941;
	wire [4-1:0] node34945;
	wire [4-1:0] node34948;
	wire [4-1:0] node34949;
	wire [4-1:0] node34950;
	wire [4-1:0] node34953;
	wire [4-1:0] node34956;
	wire [4-1:0] node34958;
	wire [4-1:0] node34960;
	wire [4-1:0] node34963;
	wire [4-1:0] node34964;
	wire [4-1:0] node34965;
	wire [4-1:0] node34966;
	wire [4-1:0] node34967;
	wire [4-1:0] node34971;
	wire [4-1:0] node34973;
	wire [4-1:0] node34976;
	wire [4-1:0] node34977;
	wire [4-1:0] node34978;
	wire [4-1:0] node34980;
	wire [4-1:0] node34983;
	wire [4-1:0] node34984;
	wire [4-1:0] node34987;
	wire [4-1:0] node34990;
	wire [4-1:0] node34991;
	wire [4-1:0] node34992;
	wire [4-1:0] node34995;
	wire [4-1:0] node34998;
	wire [4-1:0] node34999;
	wire [4-1:0] node35002;
	wire [4-1:0] node35005;
	wire [4-1:0] node35006;
	wire [4-1:0] node35007;
	wire [4-1:0] node35008;
	wire [4-1:0] node35011;
	wire [4-1:0] node35014;
	wire [4-1:0] node35015;
	wire [4-1:0] node35016;
	wire [4-1:0] node35019;
	wire [4-1:0] node35023;
	wire [4-1:0] node35025;
	wire [4-1:0] node35028;
	wire [4-1:0] node35029;
	wire [4-1:0] node35030;
	wire [4-1:0] node35031;
	wire [4-1:0] node35032;
	wire [4-1:0] node35033;
	wire [4-1:0] node35034;
	wire [4-1:0] node35035;
	wire [4-1:0] node35036;
	wire [4-1:0] node35037;
	wire [4-1:0] node35041;
	wire [4-1:0] node35043;
	wire [4-1:0] node35046;
	wire [4-1:0] node35048;
	wire [4-1:0] node35049;
	wire [4-1:0] node35051;
	wire [4-1:0] node35055;
	wire [4-1:0] node35056;
	wire [4-1:0] node35057;
	wire [4-1:0] node35058;
	wire [4-1:0] node35061;
	wire [4-1:0] node35063;
	wire [4-1:0] node35066;
	wire [4-1:0] node35068;
	wire [4-1:0] node35071;
	wire [4-1:0] node35072;
	wire [4-1:0] node35073;
	wire [4-1:0] node35077;
	wire [4-1:0] node35079;
	wire [4-1:0] node35082;
	wire [4-1:0] node35083;
	wire [4-1:0] node35084;
	wire [4-1:0] node35086;
	wire [4-1:0] node35089;
	wire [4-1:0] node35090;
	wire [4-1:0] node35091;
	wire [4-1:0] node35095;
	wire [4-1:0] node35096;
	wire [4-1:0] node35099;
	wire [4-1:0] node35102;
	wire [4-1:0] node35103;
	wire [4-1:0] node35104;
	wire [4-1:0] node35105;
	wire [4-1:0] node35109;
	wire [4-1:0] node35110;
	wire [4-1:0] node35114;
	wire [4-1:0] node35115;
	wire [4-1:0] node35116;
	wire [4-1:0] node35120;
	wire [4-1:0] node35122;
	wire [4-1:0] node35125;
	wire [4-1:0] node35126;
	wire [4-1:0] node35127;
	wire [4-1:0] node35128;
	wire [4-1:0] node35129;
	wire [4-1:0] node35130;
	wire [4-1:0] node35133;
	wire [4-1:0] node35136;
	wire [4-1:0] node35137;
	wire [4-1:0] node35141;
	wire [4-1:0] node35142;
	wire [4-1:0] node35143;
	wire [4-1:0] node35146;
	wire [4-1:0] node35149;
	wire [4-1:0] node35151;
	wire [4-1:0] node35154;
	wire [4-1:0] node35155;
	wire [4-1:0] node35156;
	wire [4-1:0] node35157;
	wire [4-1:0] node35160;
	wire [4-1:0] node35163;
	wire [4-1:0] node35165;
	wire [4-1:0] node35168;
	wire [4-1:0] node35170;
	wire [4-1:0] node35173;
	wire [4-1:0] node35174;
	wire [4-1:0] node35175;
	wire [4-1:0] node35176;
	wire [4-1:0] node35177;
	wire [4-1:0] node35180;
	wire [4-1:0] node35183;
	wire [4-1:0] node35184;
	wire [4-1:0] node35188;
	wire [4-1:0] node35189;
	wire [4-1:0] node35190;
	wire [4-1:0] node35193;
	wire [4-1:0] node35196;
	wire [4-1:0] node35199;
	wire [4-1:0] node35200;
	wire [4-1:0] node35202;
	wire [4-1:0] node35204;
	wire [4-1:0] node35207;
	wire [4-1:0] node35208;
	wire [4-1:0] node35209;
	wire [4-1:0] node35211;
	wire [4-1:0] node35214;
	wire [4-1:0] node35215;
	wire [4-1:0] node35219;
	wire [4-1:0] node35220;
	wire [4-1:0] node35224;
	wire [4-1:0] node35225;
	wire [4-1:0] node35226;
	wire [4-1:0] node35227;
	wire [4-1:0] node35228;
	wire [4-1:0] node35229;
	wire [4-1:0] node35230;
	wire [4-1:0] node35233;
	wire [4-1:0] node35235;
	wire [4-1:0] node35238;
	wire [4-1:0] node35239;
	wire [4-1:0] node35243;
	wire [4-1:0] node35244;
	wire [4-1:0] node35245;
	wire [4-1:0] node35249;
	wire [4-1:0] node35252;
	wire [4-1:0] node35253;
	wire [4-1:0] node35254;
	wire [4-1:0] node35255;
	wire [4-1:0] node35259;
	wire [4-1:0] node35261;
	wire [4-1:0] node35264;
	wire [4-1:0] node35265;
	wire [4-1:0] node35266;
	wire [4-1:0] node35269;
	wire [4-1:0] node35272;
	wire [4-1:0] node35274;
	wire [4-1:0] node35275;
	wire [4-1:0] node35278;
	wire [4-1:0] node35281;
	wire [4-1:0] node35282;
	wire [4-1:0] node35283;
	wire [4-1:0] node35284;
	wire [4-1:0] node35288;
	wire [4-1:0] node35289;
	wire [4-1:0] node35291;
	wire [4-1:0] node35294;
	wire [4-1:0] node35295;
	wire [4-1:0] node35299;
	wire [4-1:0] node35300;
	wire [4-1:0] node35301;
	wire [4-1:0] node35303;
	wire [4-1:0] node35306;
	wire [4-1:0] node35308;
	wire [4-1:0] node35311;
	wire [4-1:0] node35312;
	wire [4-1:0] node35313;
	wire [4-1:0] node35316;
	wire [4-1:0] node35320;
	wire [4-1:0] node35321;
	wire [4-1:0] node35322;
	wire [4-1:0] node35323;
	wire [4-1:0] node35324;
	wire [4-1:0] node35325;
	wire [4-1:0] node35329;
	wire [4-1:0] node35330;
	wire [4-1:0] node35333;
	wire [4-1:0] node35336;
	wire [4-1:0] node35337;
	wire [4-1:0] node35338;
	wire [4-1:0] node35341;
	wire [4-1:0] node35344;
	wire [4-1:0] node35347;
	wire [4-1:0] node35348;
	wire [4-1:0] node35349;
	wire [4-1:0] node35350;
	wire [4-1:0] node35351;
	wire [4-1:0] node35354;
	wire [4-1:0] node35357;
	wire [4-1:0] node35358;
	wire [4-1:0] node35362;
	wire [4-1:0] node35364;
	wire [4-1:0] node35365;
	wire [4-1:0] node35369;
	wire [4-1:0] node35370;
	wire [4-1:0] node35371;
	wire [4-1:0] node35375;
	wire [4-1:0] node35377;
	wire [4-1:0] node35380;
	wire [4-1:0] node35381;
	wire [4-1:0] node35382;
	wire [4-1:0] node35383;
	wire [4-1:0] node35386;
	wire [4-1:0] node35388;
	wire [4-1:0] node35390;
	wire [4-1:0] node35393;
	wire [4-1:0] node35394;
	wire [4-1:0] node35395;
	wire [4-1:0] node35398;
	wire [4-1:0] node35401;
	wire [4-1:0] node35402;
	wire [4-1:0] node35403;
	wire [4-1:0] node35406;
	wire [4-1:0] node35409;
	wire [4-1:0] node35412;
	wire [4-1:0] node35413;
	wire [4-1:0] node35414;
	wire [4-1:0] node35417;
	wire [4-1:0] node35420;
	wire [4-1:0] node35421;
	wire [4-1:0] node35424;
	wire [4-1:0] node35425;
	wire [4-1:0] node35427;
	wire [4-1:0] node35431;
	wire [4-1:0] node35432;
	wire [4-1:0] node35433;
	wire [4-1:0] node35434;
	wire [4-1:0] node35435;
	wire [4-1:0] node35436;
	wire [4-1:0] node35437;
	wire [4-1:0] node35441;
	wire [4-1:0] node35442;
	wire [4-1:0] node35444;
	wire [4-1:0] node35448;
	wire [4-1:0] node35449;
	wire [4-1:0] node35452;
	wire [4-1:0] node35453;
	wire [4-1:0] node35456;
	wire [4-1:0] node35457;
	wire [4-1:0] node35461;
	wire [4-1:0] node35462;
	wire [4-1:0] node35463;
	wire [4-1:0] node35464;
	wire [4-1:0] node35466;
	wire [4-1:0] node35469;
	wire [4-1:0] node35470;
	wire [4-1:0] node35474;
	wire [4-1:0] node35476;
	wire [4-1:0] node35477;
	wire [4-1:0] node35481;
	wire [4-1:0] node35482;
	wire [4-1:0] node35484;
	wire [4-1:0] node35487;
	wire [4-1:0] node35489;
	wire [4-1:0] node35490;
	wire [4-1:0] node35494;
	wire [4-1:0] node35495;
	wire [4-1:0] node35496;
	wire [4-1:0] node35497;
	wire [4-1:0] node35498;
	wire [4-1:0] node35499;
	wire [4-1:0] node35500;
	wire [4-1:0] node35506;
	wire [4-1:0] node35507;
	wire [4-1:0] node35509;
	wire [4-1:0] node35512;
	wire [4-1:0] node35513;
	wire [4-1:0] node35517;
	wire [4-1:0] node35518;
	wire [4-1:0] node35519;
	wire [4-1:0] node35520;
	wire [4-1:0] node35524;
	wire [4-1:0] node35526;
	wire [4-1:0] node35529;
	wire [4-1:0] node35530;
	wire [4-1:0] node35531;
	wire [4-1:0] node35534;
	wire [4-1:0] node35537;
	wire [4-1:0] node35538;
	wire [4-1:0] node35541;
	wire [4-1:0] node35544;
	wire [4-1:0] node35545;
	wire [4-1:0] node35546;
	wire [4-1:0] node35547;
	wire [4-1:0] node35548;
	wire [4-1:0] node35551;
	wire [4-1:0] node35554;
	wire [4-1:0] node35555;
	wire [4-1:0] node35556;
	wire [4-1:0] node35559;
	wire [4-1:0] node35564;
	wire [4-1:0] node35565;
	wire [4-1:0] node35566;
	wire [4-1:0] node35567;
	wire [4-1:0] node35570;
	wire [4-1:0] node35574;
	wire [4-1:0] node35575;
	wire [4-1:0] node35577;
	wire [4-1:0] node35581;
	wire [4-1:0] node35582;
	wire [4-1:0] node35583;
	wire [4-1:0] node35584;
	wire [4-1:0] node35585;
	wire [4-1:0] node35586;
	wire [4-1:0] node35588;
	wire [4-1:0] node35591;
	wire [4-1:0] node35594;
	wire [4-1:0] node35596;
	wire [4-1:0] node35599;
	wire [4-1:0] node35600;
	wire [4-1:0] node35601;
	wire [4-1:0] node35602;
	wire [4-1:0] node35603;
	wire [4-1:0] node35608;
	wire [4-1:0] node35609;
	wire [4-1:0] node35613;
	wire [4-1:0] node35614;
	wire [4-1:0] node35617;
	wire [4-1:0] node35620;
	wire [4-1:0] node35621;
	wire [4-1:0] node35622;
	wire [4-1:0] node35624;
	wire [4-1:0] node35626;
	wire [4-1:0] node35629;
	wire [4-1:0] node35630;
	wire [4-1:0] node35632;
	wire [4-1:0] node35633;
	wire [4-1:0] node35636;
	wire [4-1:0] node35639;
	wire [4-1:0] node35640;
	wire [4-1:0] node35644;
	wire [4-1:0] node35645;
	wire [4-1:0] node35647;
	wire [4-1:0] node35649;
	wire [4-1:0] node35652;
	wire [4-1:0] node35653;
	wire [4-1:0] node35657;
	wire [4-1:0] node35658;
	wire [4-1:0] node35659;
	wire [4-1:0] node35660;
	wire [4-1:0] node35661;
	wire [4-1:0] node35662;
	wire [4-1:0] node35666;
	wire [4-1:0] node35668;
	wire [4-1:0] node35671;
	wire [4-1:0] node35672;
	wire [4-1:0] node35673;
	wire [4-1:0] node35675;
	wire [4-1:0] node35679;
	wire [4-1:0] node35680;
	wire [4-1:0] node35683;
	wire [4-1:0] node35686;
	wire [4-1:0] node35687;
	wire [4-1:0] node35688;
	wire [4-1:0] node35689;
	wire [4-1:0] node35691;
	wire [4-1:0] node35694;
	wire [4-1:0] node35698;
	wire [4-1:0] node35699;
	wire [4-1:0] node35702;
	wire [4-1:0] node35704;
	wire [4-1:0] node35707;
	wire [4-1:0] node35708;
	wire [4-1:0] node35709;
	wire [4-1:0] node35711;
	wire [4-1:0] node35712;
	wire [4-1:0] node35715;
	wire [4-1:0] node35718;
	wire [4-1:0] node35719;
	wire [4-1:0] node35721;
	wire [4-1:0] node35724;
	wire [4-1:0] node35725;
	wire [4-1:0] node35728;
	wire [4-1:0] node35731;
	wire [4-1:0] node35732;
	wire [4-1:0] node35733;
	wire [4-1:0] node35734;
	wire [4-1:0] node35738;
	wire [4-1:0] node35739;
	wire [4-1:0] node35743;
	wire [4-1:0] node35745;
	wire [4-1:0] node35746;
	wire [4-1:0] node35747;
	wire [4-1:0] node35752;
	wire [4-1:0] node35753;
	wire [4-1:0] node35754;
	wire [4-1:0] node35755;
	wire [4-1:0] node35756;
	wire [4-1:0] node35757;
	wire [4-1:0] node35758;
	wire [4-1:0] node35759;
	wire [4-1:0] node35762;
	wire [4-1:0] node35764;
	wire [4-1:0] node35767;
	wire [4-1:0] node35768;
	wire [4-1:0] node35769;
	wire [4-1:0] node35772;
	wire [4-1:0] node35775;
	wire [4-1:0] node35776;
	wire [4-1:0] node35778;
	wire [4-1:0] node35781;
	wire [4-1:0] node35783;
	wire [4-1:0] node35786;
	wire [4-1:0] node35787;
	wire [4-1:0] node35789;
	wire [4-1:0] node35792;
	wire [4-1:0] node35793;
	wire [4-1:0] node35796;
	wire [4-1:0] node35798;
	wire [4-1:0] node35801;
	wire [4-1:0] node35802;
	wire [4-1:0] node35803;
	wire [4-1:0] node35804;
	wire [4-1:0] node35806;
	wire [4-1:0] node35809;
	wire [4-1:0] node35811;
	wire [4-1:0] node35814;
	wire [4-1:0] node35815;
	wire [4-1:0] node35817;
	wire [4-1:0] node35820;
	wire [4-1:0] node35823;
	wire [4-1:0] node35824;
	wire [4-1:0] node35825;
	wire [4-1:0] node35826;
	wire [4-1:0] node35830;
	wire [4-1:0] node35831;
	wire [4-1:0] node35835;
	wire [4-1:0] node35836;
	wire [4-1:0] node35837;
	wire [4-1:0] node35841;
	wire [4-1:0] node35842;
	wire [4-1:0] node35846;
	wire [4-1:0] node35847;
	wire [4-1:0] node35848;
	wire [4-1:0] node35849;
	wire [4-1:0] node35850;
	wire [4-1:0] node35851;
	wire [4-1:0] node35853;
	wire [4-1:0] node35856;
	wire [4-1:0] node35857;
	wire [4-1:0] node35861;
	wire [4-1:0] node35862;
	wire [4-1:0] node35866;
	wire [4-1:0] node35867;
	wire [4-1:0] node35869;
	wire [4-1:0] node35870;
	wire [4-1:0] node35873;
	wire [4-1:0] node35876;
	wire [4-1:0] node35877;
	wire [4-1:0] node35878;
	wire [4-1:0] node35881;
	wire [4-1:0] node35885;
	wire [4-1:0] node35886;
	wire [4-1:0] node35888;
	wire [4-1:0] node35889;
	wire [4-1:0] node35892;
	wire [4-1:0] node35895;
	wire [4-1:0] node35896;
	wire [4-1:0] node35899;
	wire [4-1:0] node35901;
	wire [4-1:0] node35903;
	wire [4-1:0] node35906;
	wire [4-1:0] node35907;
	wire [4-1:0] node35908;
	wire [4-1:0] node35910;
	wire [4-1:0] node35911;
	wire [4-1:0] node35913;
	wire [4-1:0] node35916;
	wire [4-1:0] node35918;
	wire [4-1:0] node35921;
	wire [4-1:0] node35922;
	wire [4-1:0] node35923;
	wire [4-1:0] node35924;
	wire [4-1:0] node35930;
	wire [4-1:0] node35931;
	wire [4-1:0] node35932;
	wire [4-1:0] node35935;
	wire [4-1:0] node35937;
	wire [4-1:0] node35938;
	wire [4-1:0] node35942;
	wire [4-1:0] node35943;
	wire [4-1:0] node35944;
	wire [4-1:0] node35948;
	wire [4-1:0] node35951;
	wire [4-1:0] node35952;
	wire [4-1:0] node35953;
	wire [4-1:0] node35954;
	wire [4-1:0] node35955;
	wire [4-1:0] node35956;
	wire [4-1:0] node35957;
	wire [4-1:0] node35958;
	wire [4-1:0] node35962;
	wire [4-1:0] node35963;
	wire [4-1:0] node35967;
	wire [4-1:0] node35969;
	wire [4-1:0] node35972;
	wire [4-1:0] node35973;
	wire [4-1:0] node35976;
	wire [4-1:0] node35979;
	wire [4-1:0] node35980;
	wire [4-1:0] node35982;
	wire [4-1:0] node35985;
	wire [4-1:0] node35987;
	wire [4-1:0] node35988;
	wire [4-1:0] node35991;
	wire [4-1:0] node35994;
	wire [4-1:0] node35995;
	wire [4-1:0] node35996;
	wire [4-1:0] node35997;
	wire [4-1:0] node35998;
	wire [4-1:0] node36001;
	wire [4-1:0] node36004;
	wire [4-1:0] node36005;
	wire [4-1:0] node36009;
	wire [4-1:0] node36010;
	wire [4-1:0] node36013;
	wire [4-1:0] node36016;
	wire [4-1:0] node36017;
	wire [4-1:0] node36018;
	wire [4-1:0] node36021;
	wire [4-1:0] node36024;
	wire [4-1:0] node36025;
	wire [4-1:0] node36029;
	wire [4-1:0] node36030;
	wire [4-1:0] node36031;
	wire [4-1:0] node36032;
	wire [4-1:0] node36033;
	wire [4-1:0] node36036;
	wire [4-1:0] node36038;
	wire [4-1:0] node36041;
	wire [4-1:0] node36042;
	wire [4-1:0] node36046;
	wire [4-1:0] node36047;
	wire [4-1:0] node36049;
	wire [4-1:0] node36050;
	wire [4-1:0] node36053;
	wire [4-1:0] node36056;
	wire [4-1:0] node36057;
	wire [4-1:0] node36060;
	wire [4-1:0] node36063;
	wire [4-1:0] node36064;
	wire [4-1:0] node36065;
	wire [4-1:0] node36066;
	wire [4-1:0] node36070;
	wire [4-1:0] node36071;
	wire [4-1:0] node36074;
	wire [4-1:0] node36077;
	wire [4-1:0] node36078;
	wire [4-1:0] node36079;
	wire [4-1:0] node36082;
	wire [4-1:0] node36085;
	wire [4-1:0] node36087;
	wire [4-1:0] node36090;
	wire [4-1:0] node36091;
	wire [4-1:0] node36092;
	wire [4-1:0] node36093;
	wire [4-1:0] node36094;
	wire [4-1:0] node36095;
	wire [4-1:0] node36096;
	wire [4-1:0] node36099;
	wire [4-1:0] node36101;
	wire [4-1:0] node36104;
	wire [4-1:0] node36106;
	wire [4-1:0] node36108;
	wire [4-1:0] node36111;
	wire [4-1:0] node36112;
	wire [4-1:0] node36113;
	wire [4-1:0] node36116;
	wire [4-1:0] node36117;
	wire [4-1:0] node36120;
	wire [4-1:0] node36123;
	wire [4-1:0] node36124;
	wire [4-1:0] node36125;
	wire [4-1:0] node36126;
	wire [4-1:0] node36131;
	wire [4-1:0] node36132;
	wire [4-1:0] node36136;
	wire [4-1:0] node36137;
	wire [4-1:0] node36138;
	wire [4-1:0] node36139;
	wire [4-1:0] node36142;
	wire [4-1:0] node36145;
	wire [4-1:0] node36146;
	wire [4-1:0] node36147;
	wire [4-1:0] node36150;
	wire [4-1:0] node36153;
	wire [4-1:0] node36154;
	wire [4-1:0] node36158;
	wire [4-1:0] node36159;
	wire [4-1:0] node36160;
	wire [4-1:0] node36161;
	wire [4-1:0] node36163;
	wire [4-1:0] node36167;
	wire [4-1:0] node36170;
	wire [4-1:0] node36171;
	wire [4-1:0] node36173;
	wire [4-1:0] node36174;
	wire [4-1:0] node36177;
	wire [4-1:0] node36180;
	wire [4-1:0] node36181;
	wire [4-1:0] node36183;
	wire [4-1:0] node36186;
	wire [4-1:0] node36187;
	wire [4-1:0] node36190;
	wire [4-1:0] node36193;
	wire [4-1:0] node36194;
	wire [4-1:0] node36195;
	wire [4-1:0] node36196;
	wire [4-1:0] node36197;
	wire [4-1:0] node36199;
	wire [4-1:0] node36202;
	wire [4-1:0] node36204;
	wire [4-1:0] node36206;
	wire [4-1:0] node36209;
	wire [4-1:0] node36210;
	wire [4-1:0] node36211;
	wire [4-1:0] node36215;
	wire [4-1:0] node36217;
	wire [4-1:0] node36220;
	wire [4-1:0] node36221;
	wire [4-1:0] node36222;
	wire [4-1:0] node36225;
	wire [4-1:0] node36226;
	wire [4-1:0] node36229;
	wire [4-1:0] node36232;
	wire [4-1:0] node36233;
	wire [4-1:0] node36234;
	wire [4-1:0] node36235;
	wire [4-1:0] node36238;
	wire [4-1:0] node36243;
	wire [4-1:0] node36244;
	wire [4-1:0] node36245;
	wire [4-1:0] node36246;
	wire [4-1:0] node36249;
	wire [4-1:0] node36252;
	wire [4-1:0] node36253;
	wire [4-1:0] node36254;
	wire [4-1:0] node36258;
	wire [4-1:0] node36259;
	wire [4-1:0] node36262;
	wire [4-1:0] node36265;
	wire [4-1:0] node36266;
	wire [4-1:0] node36267;
	wire [4-1:0] node36268;
	wire [4-1:0] node36271;
	wire [4-1:0] node36275;
	wire [4-1:0] node36276;
	wire [4-1:0] node36278;
	wire [4-1:0] node36281;
	wire [4-1:0] node36282;
	wire [4-1:0] node36285;
	wire [4-1:0] node36288;
	wire [4-1:0] node36289;
	wire [4-1:0] node36290;
	wire [4-1:0] node36291;
	wire [4-1:0] node36292;
	wire [4-1:0] node36293;
	wire [4-1:0] node36294;
	wire [4-1:0] node36295;
	wire [4-1:0] node36300;
	wire [4-1:0] node36301;
	wire [4-1:0] node36305;
	wire [4-1:0] node36307;
	wire [4-1:0] node36309;
	wire [4-1:0] node36312;
	wire [4-1:0] node36313;
	wire [4-1:0] node36314;
	wire [4-1:0] node36316;
	wire [4-1:0] node36318;
	wire [4-1:0] node36322;
	wire [4-1:0] node36323;
	wire [4-1:0] node36324;
	wire [4-1:0] node36326;
	wire [4-1:0] node36330;
	wire [4-1:0] node36332;
	wire [4-1:0] node36335;
	wire [4-1:0] node36336;
	wire [4-1:0] node36337;
	wire [4-1:0] node36338;
	wire [4-1:0] node36340;
	wire [4-1:0] node36343;
	wire [4-1:0] node36346;
	wire [4-1:0] node36348;
	wire [4-1:0] node36351;
	wire [4-1:0] node36352;
	wire [4-1:0] node36353;
	wire [4-1:0] node36355;
	wire [4-1:0] node36358;
	wire [4-1:0] node36360;
	wire [4-1:0] node36363;
	wire [4-1:0] node36364;
	wire [4-1:0] node36366;
	wire [4-1:0] node36368;
	wire [4-1:0] node36371;
	wire [4-1:0] node36372;
	wire [4-1:0] node36373;
	wire [4-1:0] node36376;
	wire [4-1:0] node36380;
	wire [4-1:0] node36381;
	wire [4-1:0] node36382;
	wire [4-1:0] node36383;
	wire [4-1:0] node36385;
	wire [4-1:0] node36386;
	wire [4-1:0] node36388;
	wire [4-1:0] node36391;
	wire [4-1:0] node36393;
	wire [4-1:0] node36396;
	wire [4-1:0] node36397;
	wire [4-1:0] node36398;
	wire [4-1:0] node36401;
	wire [4-1:0] node36404;
	wire [4-1:0] node36405;
	wire [4-1:0] node36408;
	wire [4-1:0] node36411;
	wire [4-1:0] node36412;
	wire [4-1:0] node36413;
	wire [4-1:0] node36414;
	wire [4-1:0] node36418;
	wire [4-1:0] node36419;
	wire [4-1:0] node36423;
	wire [4-1:0] node36424;
	wire [4-1:0] node36427;
	wire [4-1:0] node36430;
	wire [4-1:0] node36431;
	wire [4-1:0] node36432;
	wire [4-1:0] node36434;
	wire [4-1:0] node36435;
	wire [4-1:0] node36439;
	wire [4-1:0] node36440;
	wire [4-1:0] node36443;
	wire [4-1:0] node36446;
	wire [4-1:0] node36447;
	wire [4-1:0] node36448;
	wire [4-1:0] node36450;
	wire [4-1:0] node36453;
	wire [4-1:0] node36455;
	wire [4-1:0] node36458;
	wire [4-1:0] node36460;
	wire [4-1:0] node36461;
	wire [4-1:0] node36464;
	wire [4-1:0] node36467;
	wire [4-1:0] node36468;
	wire [4-1:0] node36469;
	wire [4-1:0] node36470;
	wire [4-1:0] node36471;
	wire [4-1:0] node36472;
	wire [4-1:0] node36473;
	wire [4-1:0] node36474;
	wire [4-1:0] node36475;
	wire [4-1:0] node36476;
	wire [4-1:0] node36477;
	wire [4-1:0] node36480;
	wire [4-1:0] node36483;
	wire [4-1:0] node36486;
	wire [4-1:0] node36487;
	wire [4-1:0] node36490;
	wire [4-1:0] node36492;
	wire [4-1:0] node36495;
	wire [4-1:0] node36496;
	wire [4-1:0] node36497;
	wire [4-1:0] node36500;
	wire [4-1:0] node36502;
	wire [4-1:0] node36505;
	wire [4-1:0] node36506;
	wire [4-1:0] node36507;
	wire [4-1:0] node36511;
	wire [4-1:0] node36512;
	wire [4-1:0] node36515;
	wire [4-1:0] node36518;
	wire [4-1:0] node36519;
	wire [4-1:0] node36520;
	wire [4-1:0] node36521;
	wire [4-1:0] node36522;
	wire [4-1:0] node36525;
	wire [4-1:0] node36528;
	wire [4-1:0] node36530;
	wire [4-1:0] node36533;
	wire [4-1:0] node36534;
	wire [4-1:0] node36538;
	wire [4-1:0] node36539;
	wire [4-1:0] node36540;
	wire [4-1:0] node36543;
	wire [4-1:0] node36546;
	wire [4-1:0] node36547;
	wire [4-1:0] node36550;
	wire [4-1:0] node36553;
	wire [4-1:0] node36554;
	wire [4-1:0] node36555;
	wire [4-1:0] node36556;
	wire [4-1:0] node36557;
	wire [4-1:0] node36559;
	wire [4-1:0] node36563;
	wire [4-1:0] node36564;
	wire [4-1:0] node36567;
	wire [4-1:0] node36570;
	wire [4-1:0] node36571;
	wire [4-1:0] node36572;
	wire [4-1:0] node36575;
	wire [4-1:0] node36579;
	wire [4-1:0] node36580;
	wire [4-1:0] node36581;
	wire [4-1:0] node36582;
	wire [4-1:0] node36583;
	wire [4-1:0] node36584;
	wire [4-1:0] node36589;
	wire [4-1:0] node36592;
	wire [4-1:0] node36594;
	wire [4-1:0] node36597;
	wire [4-1:0] node36598;
	wire [4-1:0] node36600;
	wire [4-1:0] node36603;
	wire [4-1:0] node36604;
	wire [4-1:0] node36606;
	wire [4-1:0] node36609;
	wire [4-1:0] node36611;
	wire [4-1:0] node36614;
	wire [4-1:0] node36615;
	wire [4-1:0] node36616;
	wire [4-1:0] node36617;
	wire [4-1:0] node36618;
	wire [4-1:0] node36619;
	wire [4-1:0] node36621;
	wire [4-1:0] node36624;
	wire [4-1:0] node36626;
	wire [4-1:0] node36627;
	wire [4-1:0] node36630;
	wire [4-1:0] node36633;
	wire [4-1:0] node36634;
	wire [4-1:0] node36637;
	wire [4-1:0] node36638;
	wire [4-1:0] node36642;
	wire [4-1:0] node36643;
	wire [4-1:0] node36644;
	wire [4-1:0] node36645;
	wire [4-1:0] node36649;
	wire [4-1:0] node36651;
	wire [4-1:0] node36653;
	wire [4-1:0] node36656;
	wire [4-1:0] node36657;
	wire [4-1:0] node36659;
	wire [4-1:0] node36662;
	wire [4-1:0] node36664;
	wire [4-1:0] node36666;
	wire [4-1:0] node36669;
	wire [4-1:0] node36670;
	wire [4-1:0] node36671;
	wire [4-1:0] node36674;
	wire [4-1:0] node36675;
	wire [4-1:0] node36676;
	wire [4-1:0] node36679;
	wire [4-1:0] node36680;
	wire [4-1:0] node36684;
	wire [4-1:0] node36685;
	wire [4-1:0] node36686;
	wire [4-1:0] node36691;
	wire [4-1:0] node36692;
	wire [4-1:0] node36694;
	wire [4-1:0] node36695;
	wire [4-1:0] node36696;
	wire [4-1:0] node36700;
	wire [4-1:0] node36702;
	wire [4-1:0] node36705;
	wire [4-1:0] node36706;
	wire [4-1:0] node36709;
	wire [4-1:0] node36710;
	wire [4-1:0] node36714;
	wire [4-1:0] node36715;
	wire [4-1:0] node36716;
	wire [4-1:0] node36717;
	wire [4-1:0] node36719;
	wire [4-1:0] node36721;
	wire [4-1:0] node36724;
	wire [4-1:0] node36726;
	wire [4-1:0] node36727;
	wire [4-1:0] node36730;
	wire [4-1:0] node36733;
	wire [4-1:0] node36734;
	wire [4-1:0] node36737;
	wire [4-1:0] node36740;
	wire [4-1:0] node36741;
	wire [4-1:0] node36742;
	wire [4-1:0] node36745;
	wire [4-1:0] node36748;
	wire [4-1:0] node36749;
	wire [4-1:0] node36750;
	wire [4-1:0] node36753;
	wire [4-1:0] node36756;
	wire [4-1:0] node36757;
	wire [4-1:0] node36761;
	wire [4-1:0] node36762;
	wire [4-1:0] node36763;
	wire [4-1:0] node36764;
	wire [4-1:0] node36765;
	wire [4-1:0] node36766;
	wire [4-1:0] node36767;
	wire [4-1:0] node36770;
	wire [4-1:0] node36773;
	wire [4-1:0] node36774;
	wire [4-1:0] node36775;
	wire [4-1:0] node36777;
	wire [4-1:0] node36780;
	wire [4-1:0] node36781;
	wire [4-1:0] node36784;
	wire [4-1:0] node36787;
	wire [4-1:0] node36789;
	wire [4-1:0] node36792;
	wire [4-1:0] node36793;
	wire [4-1:0] node36794;
	wire [4-1:0] node36796;
	wire [4-1:0] node36799;
	wire [4-1:0] node36800;
	wire [4-1:0] node36804;
	wire [4-1:0] node36805;
	wire [4-1:0] node36808;
	wire [4-1:0] node36811;
	wire [4-1:0] node36812;
	wire [4-1:0] node36813;
	wire [4-1:0] node36814;
	wire [4-1:0] node36817;
	wire [4-1:0] node36820;
	wire [4-1:0] node36821;
	wire [4-1:0] node36822;
	wire [4-1:0] node36826;
	wire [4-1:0] node36827;
	wire [4-1:0] node36829;
	wire [4-1:0] node36832;
	wire [4-1:0] node36833;
	wire [4-1:0] node36836;
	wire [4-1:0] node36839;
	wire [4-1:0] node36840;
	wire [4-1:0] node36841;
	wire [4-1:0] node36843;
	wire [4-1:0] node36847;
	wire [4-1:0] node36848;
	wire [4-1:0] node36852;
	wire [4-1:0] node36853;
	wire [4-1:0] node36854;
	wire [4-1:0] node36855;
	wire [4-1:0] node36856;
	wire [4-1:0] node36857;
	wire [4-1:0] node36860;
	wire [4-1:0] node36863;
	wire [4-1:0] node36864;
	wire [4-1:0] node36868;
	wire [4-1:0] node36869;
	wire [4-1:0] node36873;
	wire [4-1:0] node36874;
	wire [4-1:0] node36876;
	wire [4-1:0] node36879;
	wire [4-1:0] node36881;
	wire [4-1:0] node36884;
	wire [4-1:0] node36885;
	wire [4-1:0] node36886;
	wire [4-1:0] node36887;
	wire [4-1:0] node36889;
	wire [4-1:0] node36890;
	wire [4-1:0] node36893;
	wire [4-1:0] node36897;
	wire [4-1:0] node36898;
	wire [4-1:0] node36900;
	wire [4-1:0] node36903;
	wire [4-1:0] node36905;
	wire [4-1:0] node36906;
	wire [4-1:0] node36910;
	wire [4-1:0] node36911;
	wire [4-1:0] node36914;
	wire [4-1:0] node36917;
	wire [4-1:0] node36918;
	wire [4-1:0] node36919;
	wire [4-1:0] node36920;
	wire [4-1:0] node36921;
	wire [4-1:0] node36923;
	wire [4-1:0] node36924;
	wire [4-1:0] node36925;
	wire [4-1:0] node36929;
	wire [4-1:0] node36932;
	wire [4-1:0] node36933;
	wire [4-1:0] node36934;
	wire [4-1:0] node36937;
	wire [4-1:0] node36940;
	wire [4-1:0] node36942;
	wire [4-1:0] node36945;
	wire [4-1:0] node36946;
	wire [4-1:0] node36947;
	wire [4-1:0] node36948;
	wire [4-1:0] node36953;
	wire [4-1:0] node36954;
	wire [4-1:0] node36957;
	wire [4-1:0] node36960;
	wire [4-1:0] node36961;
	wire [4-1:0] node36962;
	wire [4-1:0] node36963;
	wire [4-1:0] node36964;
	wire [4-1:0] node36965;
	wire [4-1:0] node36968;
	wire [4-1:0] node36972;
	wire [4-1:0] node36973;
	wire [4-1:0] node36975;
	wire [4-1:0] node36978;
	wire [4-1:0] node36979;
	wire [4-1:0] node36982;
	wire [4-1:0] node36985;
	wire [4-1:0] node36987;
	wire [4-1:0] node36988;
	wire [4-1:0] node36991;
	wire [4-1:0] node36994;
	wire [4-1:0] node36995;
	wire [4-1:0] node36996;
	wire [4-1:0] node36999;
	wire [4-1:0] node37002;
	wire [4-1:0] node37003;
	wire [4-1:0] node37007;
	wire [4-1:0] node37008;
	wire [4-1:0] node37009;
	wire [4-1:0] node37010;
	wire [4-1:0] node37011;
	wire [4-1:0] node37015;
	wire [4-1:0] node37016;
	wire [4-1:0] node37018;
	wire [4-1:0] node37021;
	wire [4-1:0] node37022;
	wire [4-1:0] node37025;
	wire [4-1:0] node37028;
	wire [4-1:0] node37029;
	wire [4-1:0] node37030;
	wire [4-1:0] node37033;
	wire [4-1:0] node37036;
	wire [4-1:0] node37037;
	wire [4-1:0] node37040;
	wire [4-1:0] node37043;
	wire [4-1:0] node37044;
	wire [4-1:0] node37045;
	wire [4-1:0] node37047;
	wire [4-1:0] node37050;
	wire [4-1:0] node37051;
	wire [4-1:0] node37054;
	wire [4-1:0] node37055;
	wire [4-1:0] node37058;
	wire [4-1:0] node37061;
	wire [4-1:0] node37062;
	wire [4-1:0] node37064;
	wire [4-1:0] node37067;
	wire [4-1:0] node37068;
	wire [4-1:0] node37071;
	wire [4-1:0] node37074;
	wire [4-1:0] node37075;
	wire [4-1:0] node37076;
	wire [4-1:0] node37077;
	wire [4-1:0] node37078;
	wire [4-1:0] node37079;
	wire [4-1:0] node37080;
	wire [4-1:0] node37081;
	wire [4-1:0] node37082;
	wire [4-1:0] node37083;
	wire [4-1:0] node37087;
	wire [4-1:0] node37090;
	wire [4-1:0] node37091;
	wire [4-1:0] node37094;
	wire [4-1:0] node37097;
	wire [4-1:0] node37098;
	wire [4-1:0] node37100;
	wire [4-1:0] node37101;
	wire [4-1:0] node37106;
	wire [4-1:0] node37107;
	wire [4-1:0] node37108;
	wire [4-1:0] node37109;
	wire [4-1:0] node37112;
	wire [4-1:0] node37115;
	wire [4-1:0] node37117;
	wire [4-1:0] node37120;
	wire [4-1:0] node37121;
	wire [4-1:0] node37123;
	wire [4-1:0] node37126;
	wire [4-1:0] node37129;
	wire [4-1:0] node37130;
	wire [4-1:0] node37131;
	wire [4-1:0] node37132;
	wire [4-1:0] node37133;
	wire [4-1:0] node37135;
	wire [4-1:0] node37138;
	wire [4-1:0] node37141;
	wire [4-1:0] node37142;
	wire [4-1:0] node37146;
	wire [4-1:0] node37147;
	wire [4-1:0] node37148;
	wire [4-1:0] node37151;
	wire [4-1:0] node37154;
	wire [4-1:0] node37156;
	wire [4-1:0] node37159;
	wire [4-1:0] node37160;
	wire [4-1:0] node37162;
	wire [4-1:0] node37165;
	wire [4-1:0] node37166;
	wire [4-1:0] node37169;
	wire [4-1:0] node37172;
	wire [4-1:0] node37173;
	wire [4-1:0] node37174;
	wire [4-1:0] node37175;
	wire [4-1:0] node37176;
	wire [4-1:0] node37178;
	wire [4-1:0] node37181;
	wire [4-1:0] node37184;
	wire [4-1:0] node37185;
	wire [4-1:0] node37186;
	wire [4-1:0] node37190;
	wire [4-1:0] node37191;
	wire [4-1:0] node37194;
	wire [4-1:0] node37197;
	wire [4-1:0] node37198;
	wire [4-1:0] node37199;
	wire [4-1:0] node37202;
	wire [4-1:0] node37204;
	wire [4-1:0] node37207;
	wire [4-1:0] node37208;
	wire [4-1:0] node37210;
	wire [4-1:0] node37213;
	wire [4-1:0] node37214;
	wire [4-1:0] node37218;
	wire [4-1:0] node37219;
	wire [4-1:0] node37220;
	wire [4-1:0] node37221;
	wire [4-1:0] node37224;
	wire [4-1:0] node37225;
	wire [4-1:0] node37228;
	wire [4-1:0] node37231;
	wire [4-1:0] node37232;
	wire [4-1:0] node37233;
	wire [4-1:0] node37235;
	wire [4-1:0] node37239;
	wire [4-1:0] node37240;
	wire [4-1:0] node37243;
	wire [4-1:0] node37246;
	wire [4-1:0] node37247;
	wire [4-1:0] node37248;
	wire [4-1:0] node37249;
	wire [4-1:0] node37253;
	wire [4-1:0] node37255;
	wire [4-1:0] node37256;
	wire [4-1:0] node37259;
	wire [4-1:0] node37262;
	wire [4-1:0] node37263;
	wire [4-1:0] node37265;
	wire [4-1:0] node37268;
	wire [4-1:0] node37269;
	wire [4-1:0] node37272;
	wire [4-1:0] node37275;
	wire [4-1:0] node37276;
	wire [4-1:0] node37277;
	wire [4-1:0] node37278;
	wire [4-1:0] node37279;
	wire [4-1:0] node37281;
	wire [4-1:0] node37283;
	wire [4-1:0] node37284;
	wire [4-1:0] node37288;
	wire [4-1:0] node37290;
	wire [4-1:0] node37293;
	wire [4-1:0] node37294;
	wire [4-1:0] node37295;
	wire [4-1:0] node37298;
	wire [4-1:0] node37299;
	wire [4-1:0] node37302;
	wire [4-1:0] node37305;
	wire [4-1:0] node37306;
	wire [4-1:0] node37309;
	wire [4-1:0] node37312;
	wire [4-1:0] node37313;
	wire [4-1:0] node37314;
	wire [4-1:0] node37316;
	wire [4-1:0] node37319;
	wire [4-1:0] node37321;
	wire [4-1:0] node37322;
	wire [4-1:0] node37325;
	wire [4-1:0] node37328;
	wire [4-1:0] node37329;
	wire [4-1:0] node37330;
	wire [4-1:0] node37331;
	wire [4-1:0] node37332;
	wire [4-1:0] node37337;
	wire [4-1:0] node37338;
	wire [4-1:0] node37339;
	wire [4-1:0] node37343;
	wire [4-1:0] node37344;
	wire [4-1:0] node37347;
	wire [4-1:0] node37350;
	wire [4-1:0] node37351;
	wire [4-1:0] node37354;
	wire [4-1:0] node37356;
	wire [4-1:0] node37357;
	wire [4-1:0] node37360;
	wire [4-1:0] node37363;
	wire [4-1:0] node37364;
	wire [4-1:0] node37365;
	wire [4-1:0] node37366;
	wire [4-1:0] node37368;
	wire [4-1:0] node37369;
	wire [4-1:0] node37370;
	wire [4-1:0] node37373;
	wire [4-1:0] node37377;
	wire [4-1:0] node37378;
	wire [4-1:0] node37381;
	wire [4-1:0] node37383;
	wire [4-1:0] node37386;
	wire [4-1:0] node37387;
	wire [4-1:0] node37388;
	wire [4-1:0] node37389;
	wire [4-1:0] node37392;
	wire [4-1:0] node37396;
	wire [4-1:0] node37397;
	wire [4-1:0] node37399;
	wire [4-1:0] node37402;
	wire [4-1:0] node37404;
	wire [4-1:0] node37407;
	wire [4-1:0] node37408;
	wire [4-1:0] node37409;
	wire [4-1:0] node37410;
	wire [4-1:0] node37411;
	wire [4-1:0] node37415;
	wire [4-1:0] node37418;
	wire [4-1:0] node37419;
	wire [4-1:0] node37420;
	wire [4-1:0] node37425;
	wire [4-1:0] node37426;
	wire [4-1:0] node37427;
	wire [4-1:0] node37428;
	wire [4-1:0] node37432;
	wire [4-1:0] node37435;
	wire [4-1:0] node37436;
	wire [4-1:0] node37439;
	wire [4-1:0] node37442;
	wire [4-1:0] node37443;
	wire [4-1:0] node37444;
	wire [4-1:0] node37445;
	wire [4-1:0] node37446;
	wire [4-1:0] node37447;
	wire [4-1:0] node37448;
	wire [4-1:0] node37450;
	wire [4-1:0] node37453;
	wire [4-1:0] node37455;
	wire [4-1:0] node37458;
	wire [4-1:0] node37459;
	wire [4-1:0] node37461;
	wire [4-1:0] node37464;
	wire [4-1:0] node37466;
	wire [4-1:0] node37469;
	wire [4-1:0] node37470;
	wire [4-1:0] node37472;
	wire [4-1:0] node37475;
	wire [4-1:0] node37477;
	wire [4-1:0] node37480;
	wire [4-1:0] node37481;
	wire [4-1:0] node37482;
	wire [4-1:0] node37483;
	wire [4-1:0] node37485;
	wire [4-1:0] node37488;
	wire [4-1:0] node37490;
	wire [4-1:0] node37494;
	wire [4-1:0] node37495;
	wire [4-1:0] node37496;
	wire [4-1:0] node37498;
	wire [4-1:0] node37500;
	wire [4-1:0] node37503;
	wire [4-1:0] node37505;
	wire [4-1:0] node37508;
	wire [4-1:0] node37509;
	wire [4-1:0] node37513;
	wire [4-1:0] node37514;
	wire [4-1:0] node37515;
	wire [4-1:0] node37516;
	wire [4-1:0] node37517;
	wire [4-1:0] node37521;
	wire [4-1:0] node37522;
	wire [4-1:0] node37525;
	wire [4-1:0] node37527;
	wire [4-1:0] node37530;
	wire [4-1:0] node37531;
	wire [4-1:0] node37534;
	wire [4-1:0] node37535;
	wire [4-1:0] node37536;
	wire [4-1:0] node37540;
	wire [4-1:0] node37543;
	wire [4-1:0] node37544;
	wire [4-1:0] node37545;
	wire [4-1:0] node37546;
	wire [4-1:0] node37548;
	wire [4-1:0] node37549;
	wire [4-1:0] node37552;
	wire [4-1:0] node37556;
	wire [4-1:0] node37557;
	wire [4-1:0] node37560;
	wire [4-1:0] node37563;
	wire [4-1:0] node37564;
	wire [4-1:0] node37565;
	wire [4-1:0] node37567;
	wire [4-1:0] node37571;
	wire [4-1:0] node37572;
	wire [4-1:0] node37575;
	wire [4-1:0] node37578;
	wire [4-1:0] node37579;
	wire [4-1:0] node37580;
	wire [4-1:0] node37581;
	wire [4-1:0] node37582;
	wire [4-1:0] node37583;
	wire [4-1:0] node37585;
	wire [4-1:0] node37589;
	wire [4-1:0] node37590;
	wire [4-1:0] node37594;
	wire [4-1:0] node37595;
	wire [4-1:0] node37596;
	wire [4-1:0] node37597;
	wire [4-1:0] node37599;
	wire [4-1:0] node37604;
	wire [4-1:0] node37605;
	wire [4-1:0] node37606;
	wire [4-1:0] node37610;
	wire [4-1:0] node37611;
	wire [4-1:0] node37615;
	wire [4-1:0] node37616;
	wire [4-1:0] node37617;
	wire [4-1:0] node37618;
	wire [4-1:0] node37619;
	wire [4-1:0] node37623;
	wire [4-1:0] node37624;
	wire [4-1:0] node37628;
	wire [4-1:0] node37629;
	wire [4-1:0] node37630;
	wire [4-1:0] node37635;
	wire [4-1:0] node37636;
	wire [4-1:0] node37637;
	wire [4-1:0] node37639;
	wire [4-1:0] node37640;
	wire [4-1:0] node37645;
	wire [4-1:0] node37646;
	wire [4-1:0] node37648;
	wire [4-1:0] node37651;
	wire [4-1:0] node37652;
	wire [4-1:0] node37653;
	wire [4-1:0] node37657;
	wire [4-1:0] node37660;
	wire [4-1:0] node37661;
	wire [4-1:0] node37662;
	wire [4-1:0] node37663;
	wire [4-1:0] node37666;
	wire [4-1:0] node37667;
	wire [4-1:0] node37669;
	wire [4-1:0] node37670;
	wire [4-1:0] node37675;
	wire [4-1:0] node37676;
	wire [4-1:0] node37679;
	wire [4-1:0] node37680;
	wire [4-1:0] node37683;
	wire [4-1:0] node37686;
	wire [4-1:0] node37687;
	wire [4-1:0] node37688;
	wire [4-1:0] node37689;
	wire [4-1:0] node37690;
	wire [4-1:0] node37694;
	wire [4-1:0] node37697;
	wire [4-1:0] node37698;
	wire [4-1:0] node37699;
	wire [4-1:0] node37704;
	wire [4-1:0] node37705;
	wire [4-1:0] node37707;
	wire [4-1:0] node37708;
	wire [4-1:0] node37711;
	wire [4-1:0] node37714;
	wire [4-1:0] node37716;
	wire [4-1:0] node37719;
	wire [4-1:0] node37720;
	wire [4-1:0] node37721;
	wire [4-1:0] node37722;
	wire [4-1:0] node37723;
	wire [4-1:0] node37724;
	wire [4-1:0] node37725;
	wire [4-1:0] node37726;
	wire [4-1:0] node37727;
	wire [4-1:0] node37728;
	wire [4-1:0] node37731;
	wire [4-1:0] node37735;
	wire [4-1:0] node37736;
	wire [4-1:0] node37739;
	wire [4-1:0] node37742;
	wire [4-1:0] node37743;
	wire [4-1:0] node37744;
	wire [4-1:0] node37746;
	wire [4-1:0] node37750;
	wire [4-1:0] node37752;
	wire [4-1:0] node37755;
	wire [4-1:0] node37756;
	wire [4-1:0] node37757;
	wire [4-1:0] node37758;
	wire [4-1:0] node37759;
	wire [4-1:0] node37761;
	wire [4-1:0] node37765;
	wire [4-1:0] node37766;
	wire [4-1:0] node37769;
	wire [4-1:0] node37772;
	wire [4-1:0] node37774;
	wire [4-1:0] node37776;
	wire [4-1:0] node37779;
	wire [4-1:0] node37780;
	wire [4-1:0] node37781;
	wire [4-1:0] node37784;
	wire [4-1:0] node37785;
	wire [4-1:0] node37789;
	wire [4-1:0] node37790;
	wire [4-1:0] node37793;
	wire [4-1:0] node37796;
	wire [4-1:0] node37797;
	wire [4-1:0] node37798;
	wire [4-1:0] node37799;
	wire [4-1:0] node37801;
	wire [4-1:0] node37802;
	wire [4-1:0] node37803;
	wire [4-1:0] node37806;
	wire [4-1:0] node37811;
	wire [4-1:0] node37812;
	wire [4-1:0] node37815;
	wire [4-1:0] node37817;
	wire [4-1:0] node37819;
	wire [4-1:0] node37822;
	wire [4-1:0] node37823;
	wire [4-1:0] node37824;
	wire [4-1:0] node37825;
	wire [4-1:0] node37826;
	wire [4-1:0] node37828;
	wire [4-1:0] node37832;
	wire [4-1:0] node37833;
	wire [4-1:0] node37834;
	wire [4-1:0] node37839;
	wire [4-1:0] node37840;
	wire [4-1:0] node37841;
	wire [4-1:0] node37844;
	wire [4-1:0] node37847;
	wire [4-1:0] node37849;
	wire [4-1:0] node37850;
	wire [4-1:0] node37854;
	wire [4-1:0] node37856;
	wire [4-1:0] node37857;
	wire [4-1:0] node37860;
	wire [4-1:0] node37863;
	wire [4-1:0] node37864;
	wire [4-1:0] node37865;
	wire [4-1:0] node37866;
	wire [4-1:0] node37869;
	wire [4-1:0] node37872;
	wire [4-1:0] node37873;
	wire [4-1:0] node37874;
	wire [4-1:0] node37875;
	wire [4-1:0] node37877;
	wire [4-1:0] node37880;
	wire [4-1:0] node37881;
	wire [4-1:0] node37884;
	wire [4-1:0] node37887;
	wire [4-1:0] node37888;
	wire [4-1:0] node37891;
	wire [4-1:0] node37894;
	wire [4-1:0] node37895;
	wire [4-1:0] node37896;
	wire [4-1:0] node37900;
	wire [4-1:0] node37901;
	wire [4-1:0] node37904;
	wire [4-1:0] node37907;
	wire [4-1:0] node37908;
	wire [4-1:0] node37909;
	wire [4-1:0] node37910;
	wire [4-1:0] node37911;
	wire [4-1:0] node37913;
	wire [4-1:0] node37914;
	wire [4-1:0] node37917;
	wire [4-1:0] node37920;
	wire [4-1:0] node37921;
	wire [4-1:0] node37924;
	wire [4-1:0] node37927;
	wire [4-1:0] node37928;
	wire [4-1:0] node37931;
	wire [4-1:0] node37934;
	wire [4-1:0] node37935;
	wire [4-1:0] node37936;
	wire [4-1:0] node37938;
	wire [4-1:0] node37941;
	wire [4-1:0] node37943;
	wire [4-1:0] node37946;
	wire [4-1:0] node37947;
	wire [4-1:0] node37950;
	wire [4-1:0] node37953;
	wire [4-1:0] node37954;
	wire [4-1:0] node37955;
	wire [4-1:0] node37956;
	wire [4-1:0] node37958;
	wire [4-1:0] node37959;
	wire [4-1:0] node37962;
	wire [4-1:0] node37965;
	wire [4-1:0] node37966;
	wire [4-1:0] node37969;
	wire [4-1:0] node37972;
	wire [4-1:0] node37973;
	wire [4-1:0] node37974;
	wire [4-1:0] node37978;
	wire [4-1:0] node37979;
	wire [4-1:0] node37983;
	wire [4-1:0] node37984;
	wire [4-1:0] node37987;
	wire [4-1:0] node37990;
	wire [4-1:0] node37991;
	wire [4-1:0] node37992;
	wire [4-1:0] node37993;
	wire [4-1:0] node37994;
	wire [4-1:0] node37995;
	wire [4-1:0] node37996;
	wire [4-1:0] node37999;
	wire [4-1:0] node38002;
	wire [4-1:0] node38003;
	wire [4-1:0] node38004;
	wire [4-1:0] node38008;
	wire [4-1:0] node38009;
	wire [4-1:0] node38012;
	wire [4-1:0] node38015;
	wire [4-1:0] node38016;
	wire [4-1:0] node38017;
	wire [4-1:0] node38019;
	wire [4-1:0] node38022;
	wire [4-1:0] node38023;
	wire [4-1:0] node38025;
	wire [4-1:0] node38028;
	wire [4-1:0] node38031;
	wire [4-1:0] node38032;
	wire [4-1:0] node38036;
	wire [4-1:0] node38037;
	wire [4-1:0] node38038;
	wire [4-1:0] node38039;
	wire [4-1:0] node38040;
	wire [4-1:0] node38042;
	wire [4-1:0] node38045;
	wire [4-1:0] node38047;
	wire [4-1:0] node38050;
	wire [4-1:0] node38052;
	wire [4-1:0] node38055;
	wire [4-1:0] node38056;
	wire [4-1:0] node38057;
	wire [4-1:0] node38061;
	wire [4-1:0] node38062;
	wire [4-1:0] node38064;
	wire [4-1:0] node38068;
	wire [4-1:0] node38069;
	wire [4-1:0] node38070;
	wire [4-1:0] node38071;
	wire [4-1:0] node38074;
	wire [4-1:0] node38077;
	wire [4-1:0] node38080;
	wire [4-1:0] node38081;
	wire [4-1:0] node38082;
	wire [4-1:0] node38086;
	wire [4-1:0] node38088;
	wire [4-1:0] node38091;
	wire [4-1:0] node38092;
	wire [4-1:0] node38093;
	wire [4-1:0] node38094;
	wire [4-1:0] node38095;
	wire [4-1:0] node38098;
	wire [4-1:0] node38102;
	wire [4-1:0] node38103;
	wire [4-1:0] node38104;
	wire [4-1:0] node38106;
	wire [4-1:0] node38110;
	wire [4-1:0] node38111;
	wire [4-1:0] node38112;
	wire [4-1:0] node38116;
	wire [4-1:0] node38117;
	wire [4-1:0] node38118;
	wire [4-1:0] node38122;
	wire [4-1:0] node38124;
	wire [4-1:0] node38127;
	wire [4-1:0] node38128;
	wire [4-1:0] node38129;
	wire [4-1:0] node38130;
	wire [4-1:0] node38133;
	wire [4-1:0] node38135;
	wire [4-1:0] node38138;
	wire [4-1:0] node38140;
	wire [4-1:0] node38141;
	wire [4-1:0] node38144;
	wire [4-1:0] node38147;
	wire [4-1:0] node38148;
	wire [4-1:0] node38149;
	wire [4-1:0] node38152;
	wire [4-1:0] node38153;
	wire [4-1:0] node38155;
	wire [4-1:0] node38158;
	wire [4-1:0] node38159;
	wire [4-1:0] node38163;
	wire [4-1:0] node38164;
	wire [4-1:0] node38168;
	wire [4-1:0] node38169;
	wire [4-1:0] node38170;
	wire [4-1:0] node38171;
	wire [4-1:0] node38172;
	wire [4-1:0] node38173;
	wire [4-1:0] node38174;
	wire [4-1:0] node38177;
	wire [4-1:0] node38180;
	wire [4-1:0] node38181;
	wire [4-1:0] node38184;
	wire [4-1:0] node38187;
	wire [4-1:0] node38190;
	wire [4-1:0] node38191;
	wire [4-1:0] node38192;
	wire [4-1:0] node38195;
	wire [4-1:0] node38198;
	wire [4-1:0] node38199;
	wire [4-1:0] node38202;
	wire [4-1:0] node38205;
	wire [4-1:0] node38206;
	wire [4-1:0] node38207;
	wire [4-1:0] node38210;
	wire [4-1:0] node38211;
	wire [4-1:0] node38212;
	wire [4-1:0] node38215;
	wire [4-1:0] node38218;
	wire [4-1:0] node38219;
	wire [4-1:0] node38222;
	wire [4-1:0] node38225;
	wire [4-1:0] node38226;
	wire [4-1:0] node38227;
	wire [4-1:0] node38230;
	wire [4-1:0] node38234;
	wire [4-1:0] node38235;
	wire [4-1:0] node38236;
	wire [4-1:0] node38237;
	wire [4-1:0] node38239;
	wire [4-1:0] node38240;
	wire [4-1:0] node38243;
	wire [4-1:0] node38246;
	wire [4-1:0] node38247;
	wire [4-1:0] node38250;
	wire [4-1:0] node38253;
	wire [4-1:0] node38254;
	wire [4-1:0] node38257;
	wire [4-1:0] node38258;
	wire [4-1:0] node38262;
	wire [4-1:0] node38263;
	wire [4-1:0] node38264;
	wire [4-1:0] node38265;
	wire [4-1:0] node38268;
	wire [4-1:0] node38271;
	wire [4-1:0] node38272;
	wire [4-1:0] node38275;
	wire [4-1:0] node38278;
	wire [4-1:0] node38279;
	wire [4-1:0] node38280;
	wire [4-1:0] node38283;
	wire [4-1:0] node38286;
	wire [4-1:0] node38288;
	wire [4-1:0] node38289;
	wire [4-1:0] node38292;
	wire [4-1:0] node38295;
	wire [4-1:0] node38296;
	wire [4-1:0] node38297;
	wire [4-1:0] node38298;
	wire [4-1:0] node38299;
	wire [4-1:0] node38300;
	wire [4-1:0] node38301;
	wire [4-1:0] node38302;
	wire [4-1:0] node38303;
	wire [4-1:0] node38306;
	wire [4-1:0] node38309;
	wire [4-1:0] node38310;
	wire [4-1:0] node38313;
	wire [4-1:0] node38316;
	wire [4-1:0] node38317;
	wire [4-1:0] node38318;
	wire [4-1:0] node38322;
	wire [4-1:0] node38325;
	wire [4-1:0] node38326;
	wire [4-1:0] node38327;
	wire [4-1:0] node38328;
	wire [4-1:0] node38332;
	wire [4-1:0] node38335;
	wire [4-1:0] node38336;
	wire [4-1:0] node38338;
	wire [4-1:0] node38340;
	wire [4-1:0] node38343;
	wire [4-1:0] node38344;
	wire [4-1:0] node38348;
	wire [4-1:0] node38349;
	wire [4-1:0] node38350;
	wire [4-1:0] node38351;
	wire [4-1:0] node38353;
	wire [4-1:0] node38356;
	wire [4-1:0] node38357;
	wire [4-1:0] node38361;
	wire [4-1:0] node38362;
	wire [4-1:0] node38364;
	wire [4-1:0] node38367;
	wire [4-1:0] node38368;
	wire [4-1:0] node38371;
	wire [4-1:0] node38374;
	wire [4-1:0] node38375;
	wire [4-1:0] node38376;
	wire [4-1:0] node38377;
	wire [4-1:0] node38380;
	wire [4-1:0] node38383;
	wire [4-1:0] node38384;
	wire [4-1:0] node38388;
	wire [4-1:0] node38389;
	wire [4-1:0] node38390;
	wire [4-1:0] node38392;
	wire [4-1:0] node38396;
	wire [4-1:0] node38397;
	wire [4-1:0] node38400;
	wire [4-1:0] node38403;
	wire [4-1:0] node38404;
	wire [4-1:0] node38405;
	wire [4-1:0] node38406;
	wire [4-1:0] node38407;
	wire [4-1:0] node38408;
	wire [4-1:0] node38411;
	wire [4-1:0] node38415;
	wire [4-1:0] node38417;
	wire [4-1:0] node38418;
	wire [4-1:0] node38422;
	wire [4-1:0] node38423;
	wire [4-1:0] node38424;
	wire [4-1:0] node38425;
	wire [4-1:0] node38426;
	wire [4-1:0] node38431;
	wire [4-1:0] node38432;
	wire [4-1:0] node38435;
	wire [4-1:0] node38438;
	wire [4-1:0] node38440;
	wire [4-1:0] node38441;
	wire [4-1:0] node38442;
	wire [4-1:0] node38446;
	wire [4-1:0] node38449;
	wire [4-1:0] node38450;
	wire [4-1:0] node38451;
	wire [4-1:0] node38452;
	wire [4-1:0] node38453;
	wire [4-1:0] node38454;
	wire [4-1:0] node38458;
	wire [4-1:0] node38459;
	wire [4-1:0] node38463;
	wire [4-1:0] node38464;
	wire [4-1:0] node38465;
	wire [4-1:0] node38468;
	wire [4-1:0] node38471;
	wire [4-1:0] node38473;
	wire [4-1:0] node38476;
	wire [4-1:0] node38477;
	wire [4-1:0] node38479;
	wire [4-1:0] node38482;
	wire [4-1:0] node38485;
	wire [4-1:0] node38486;
	wire [4-1:0] node38487;
	wire [4-1:0] node38490;
	wire [4-1:0] node38492;
	wire [4-1:0] node38495;
	wire [4-1:0] node38497;
	wire [4-1:0] node38499;
	wire [4-1:0] node38502;
	wire [4-1:0] node38503;
	wire [4-1:0] node38504;
	wire [4-1:0] node38505;
	wire [4-1:0] node38506;
	wire [4-1:0] node38508;
	wire [4-1:0] node38509;
	wire [4-1:0] node38512;
	wire [4-1:0] node38515;
	wire [4-1:0] node38516;
	wire [4-1:0] node38517;
	wire [4-1:0] node38521;
	wire [4-1:0] node38522;
	wire [4-1:0] node38525;
	wire [4-1:0] node38528;
	wire [4-1:0] node38529;
	wire [4-1:0] node38530;
	wire [4-1:0] node38531;
	wire [4-1:0] node38534;
	wire [4-1:0] node38537;
	wire [4-1:0] node38538;
	wire [4-1:0] node38541;
	wire [4-1:0] node38544;
	wire [4-1:0] node38545;
	wire [4-1:0] node38549;
	wire [4-1:0] node38550;
	wire [4-1:0] node38551;
	wire [4-1:0] node38552;
	wire [4-1:0] node38555;
	wire [4-1:0] node38558;
	wire [4-1:0] node38559;
	wire [4-1:0] node38561;
	wire [4-1:0] node38564;
	wire [4-1:0] node38565;
	wire [4-1:0] node38569;
	wire [4-1:0] node38570;
	wire [4-1:0] node38571;
	wire [4-1:0] node38574;
	wire [4-1:0] node38577;
	wire [4-1:0] node38578;
	wire [4-1:0] node38579;
	wire [4-1:0] node38582;
	wire [4-1:0] node38585;
	wire [4-1:0] node38586;
	wire [4-1:0] node38589;
	wire [4-1:0] node38591;
	wire [4-1:0] node38594;
	wire [4-1:0] node38595;
	wire [4-1:0] node38596;
	wire [4-1:0] node38597;
	wire [4-1:0] node38598;
	wire [4-1:0] node38601;
	wire [4-1:0] node38604;
	wire [4-1:0] node38605;
	wire [4-1:0] node38608;
	wire [4-1:0] node38611;
	wire [4-1:0] node38612;
	wire [4-1:0] node38613;
	wire [4-1:0] node38615;
	wire [4-1:0] node38618;
	wire [4-1:0] node38619;
	wire [4-1:0] node38622;
	wire [4-1:0] node38625;
	wire [4-1:0] node38626;
	wire [4-1:0] node38627;
	wire [4-1:0] node38632;
	wire [4-1:0] node38633;
	wire [4-1:0] node38634;
	wire [4-1:0] node38635;
	wire [4-1:0] node38638;
	wire [4-1:0] node38641;
	wire [4-1:0] node38642;
	wire [4-1:0] node38645;
	wire [4-1:0] node38648;
	wire [4-1:0] node38649;
	wire [4-1:0] node38650;
	wire [4-1:0] node38654;
	wire [4-1:0] node38655;
	wire [4-1:0] node38658;
	wire [4-1:0] node38661;
	wire [4-1:0] node38662;
	wire [4-1:0] node38663;
	wire [4-1:0] node38664;
	wire [4-1:0] node38665;
	wire [4-1:0] node38666;
	wire [4-1:0] node38667;
	wire [4-1:0] node38671;
	wire [4-1:0] node38672;
	wire [4-1:0] node38675;
	wire [4-1:0] node38678;
	wire [4-1:0] node38679;
	wire [4-1:0] node38680;
	wire [4-1:0] node38682;
	wire [4-1:0] node38685;
	wire [4-1:0] node38687;
	wire [4-1:0] node38690;
	wire [4-1:0] node38691;
	wire [4-1:0] node38694;
	wire [4-1:0] node38697;
	wire [4-1:0] node38698;
	wire [4-1:0] node38699;
	wire [4-1:0] node38703;
	wire [4-1:0] node38704;
	wire [4-1:0] node38705;
	wire [4-1:0] node38708;
	wire [4-1:0] node38711;
	wire [4-1:0] node38712;
	wire [4-1:0] node38715;
	wire [4-1:0] node38718;
	wire [4-1:0] node38719;
	wire [4-1:0] node38720;
	wire [4-1:0] node38721;
	wire [4-1:0] node38722;
	wire [4-1:0] node38723;
	wire [4-1:0] node38726;
	wire [4-1:0] node38729;
	wire [4-1:0] node38730;
	wire [4-1:0] node38731;
	wire [4-1:0] node38734;
	wire [4-1:0] node38738;
	wire [4-1:0] node38739;
	wire [4-1:0] node38743;
	wire [4-1:0] node38744;
	wire [4-1:0] node38746;
	wire [4-1:0] node38749;
	wire [4-1:0] node38750;
	wire [4-1:0] node38752;
	wire [4-1:0] node38755;
	wire [4-1:0] node38757;
	wire [4-1:0] node38759;
	wire [4-1:0] node38762;
	wire [4-1:0] node38763;
	wire [4-1:0] node38764;
	wire [4-1:0] node38767;
	wire [4-1:0] node38770;
	wire [4-1:0] node38771;
	wire [4-1:0] node38772;
	wire [4-1:0] node38776;
	wire [4-1:0] node38777;
	wire [4-1:0] node38778;
	wire [4-1:0] node38781;
	wire [4-1:0] node38784;
	wire [4-1:0] node38786;
	wire [4-1:0] node38789;
	wire [4-1:0] node38790;
	wire [4-1:0] node38791;
	wire [4-1:0] node38792;
	wire [4-1:0] node38793;
	wire [4-1:0] node38794;
	wire [4-1:0] node38796;
	wire [4-1:0] node38799;
	wire [4-1:0] node38801;
	wire [4-1:0] node38804;
	wire [4-1:0] node38807;
	wire [4-1:0] node38808;
	wire [4-1:0] node38810;
	wire [4-1:0] node38813;
	wire [4-1:0] node38814;
	wire [4-1:0] node38816;
	wire [4-1:0] node38819;
	wire [4-1:0] node38820;
	wire [4-1:0] node38824;
	wire [4-1:0] node38825;
	wire [4-1:0] node38826;
	wire [4-1:0] node38827;
	wire [4-1:0] node38829;
	wire [4-1:0] node38832;
	wire [4-1:0] node38833;
	wire [4-1:0] node38837;
	wire [4-1:0] node38839;
	wire [4-1:0] node38840;
	wire [4-1:0] node38844;
	wire [4-1:0] node38846;
	wire [4-1:0] node38848;
	wire [4-1:0] node38849;
	wire [4-1:0] node38851;
	wire [4-1:0] node38854;
	wire [4-1:0] node38855;
	wire [4-1:0] node38859;
	wire [4-1:0] node38860;
	wire [4-1:0] node38861;
	wire [4-1:0] node38862;
	wire [4-1:0] node38863;
	wire [4-1:0] node38865;
	wire [4-1:0] node38867;
	wire [4-1:0] node38870;
	wire [4-1:0] node38871;
	wire [4-1:0] node38875;
	wire [4-1:0] node38876;
	wire [4-1:0] node38878;
	wire [4-1:0] node38881;
	wire [4-1:0] node38883;
	wire [4-1:0] node38886;
	wire [4-1:0] node38887;
	wire [4-1:0] node38888;
	wire [4-1:0] node38891;
	wire [4-1:0] node38894;
	wire [4-1:0] node38896;
	wire [4-1:0] node38897;
	wire [4-1:0] node38900;
	wire [4-1:0] node38903;
	wire [4-1:0] node38904;
	wire [4-1:0] node38905;
	wire [4-1:0] node38906;
	wire [4-1:0] node38907;
	wire [4-1:0] node38910;
	wire [4-1:0] node38913;
	wire [4-1:0] node38914;
	wire [4-1:0] node38915;
	wire [4-1:0] node38920;
	wire [4-1:0] node38921;
	wire [4-1:0] node38922;
	wire [4-1:0] node38926;
	wire [4-1:0] node38927;
	wire [4-1:0] node38930;
	wire [4-1:0] node38933;
	wire [4-1:0] node38934;
	wire [4-1:0] node38935;
	wire [4-1:0] node38936;
	wire [4-1:0] node38937;
	wire [4-1:0] node38940;
	wire [4-1:0] node38944;
	wire [4-1:0] node38945;
	wire [4-1:0] node38946;
	wire [4-1:0] node38949;
	wire [4-1:0] node38953;
	wire [4-1:0] node38954;
	wire [4-1:0] node38955;
	wire [4-1:0] node38957;
	wire [4-1:0] node38960;
	wire [4-1:0] node38963;
	wire [4-1:0] node38964;
	wire [4-1:0] node38967;
	wire [4-1:0] node38970;
	wire [4-1:0] node38971;
	wire [4-1:0] node38972;
	wire [4-1:0] node38973;
	wire [4-1:0] node38974;
	wire [4-1:0] node38975;
	wire [4-1:0] node38976;
	wire [4-1:0] node38977;
	wire [4-1:0] node38978;
	wire [4-1:0] node38979;
	wire [4-1:0] node38980;
	wire [4-1:0] node38984;
	wire [4-1:0] node38985;
	wire [4-1:0] node38988;
	wire [4-1:0] node38991;
	wire [4-1:0] node38992;
	wire [4-1:0] node38994;
	wire [4-1:0] node38995;
	wire [4-1:0] node38998;
	wire [4-1:0] node39001;
	wire [4-1:0] node39002;
	wire [4-1:0] node39006;
	wire [4-1:0] node39007;
	wire [4-1:0] node39008;
	wire [4-1:0] node39009;
	wire [4-1:0] node39010;
	wire [4-1:0] node39015;
	wire [4-1:0] node39017;
	wire [4-1:0] node39018;
	wire [4-1:0] node39021;
	wire [4-1:0] node39024;
	wire [4-1:0] node39025;
	wire [4-1:0] node39026;
	wire [4-1:0] node39030;
	wire [4-1:0] node39031;
	wire [4-1:0] node39033;
	wire [4-1:0] node39035;
	wire [4-1:0] node39038;
	wire [4-1:0] node39040;
	wire [4-1:0] node39043;
	wire [4-1:0] node39044;
	wire [4-1:0] node39045;
	wire [4-1:0] node39046;
	wire [4-1:0] node39047;
	wire [4-1:0] node39050;
	wire [4-1:0] node39053;
	wire [4-1:0] node39054;
	wire [4-1:0] node39057;
	wire [4-1:0] node39060;
	wire [4-1:0] node39061;
	wire [4-1:0] node39062;
	wire [4-1:0] node39066;
	wire [4-1:0] node39067;
	wire [4-1:0] node39070;
	wire [4-1:0] node39073;
	wire [4-1:0] node39074;
	wire [4-1:0] node39075;
	wire [4-1:0] node39077;
	wire [4-1:0] node39078;
	wire [4-1:0] node39082;
	wire [4-1:0] node39084;
	wire [4-1:0] node39087;
	wire [4-1:0] node39088;
	wire [4-1:0] node39091;
	wire [4-1:0] node39094;
	wire [4-1:0] node39095;
	wire [4-1:0] node39096;
	wire [4-1:0] node39097;
	wire [4-1:0] node39098;
	wire [4-1:0] node39100;
	wire [4-1:0] node39103;
	wire [4-1:0] node39105;
	wire [4-1:0] node39108;
	wire [4-1:0] node39109;
	wire [4-1:0] node39110;
	wire [4-1:0] node39113;
	wire [4-1:0] node39116;
	wire [4-1:0] node39117;
	wire [4-1:0] node39119;
	wire [4-1:0] node39122;
	wire [4-1:0] node39125;
	wire [4-1:0] node39126;
	wire [4-1:0] node39127;
	wire [4-1:0] node39128;
	wire [4-1:0] node39131;
	wire [4-1:0] node39134;
	wire [4-1:0] node39135;
	wire [4-1:0] node39138;
	wire [4-1:0] node39141;
	wire [4-1:0] node39142;
	wire [4-1:0] node39143;
	wire [4-1:0] node39145;
	wire [4-1:0] node39146;
	wire [4-1:0] node39149;
	wire [4-1:0] node39152;
	wire [4-1:0] node39153;
	wire [4-1:0] node39157;
	wire [4-1:0] node39158;
	wire [4-1:0] node39159;
	wire [4-1:0] node39160;
	wire [4-1:0] node39163;
	wire [4-1:0] node39168;
	wire [4-1:0] node39169;
	wire [4-1:0] node39170;
	wire [4-1:0] node39171;
	wire [4-1:0] node39172;
	wire [4-1:0] node39176;
	wire [4-1:0] node39177;
	wire [4-1:0] node39181;
	wire [4-1:0] node39182;
	wire [4-1:0] node39185;
	wire [4-1:0] node39188;
	wire [4-1:0] node39189;
	wire [4-1:0] node39191;
	wire [4-1:0] node39192;
	wire [4-1:0] node39193;
	wire [4-1:0] node39196;
	wire [4-1:0] node39200;
	wire [4-1:0] node39201;
	wire [4-1:0] node39202;
	wire [4-1:0] node39205;
	wire [4-1:0] node39208;
	wire [4-1:0] node39210;
	wire [4-1:0] node39211;
	wire [4-1:0] node39214;
	wire [4-1:0] node39217;
	wire [4-1:0] node39218;
	wire [4-1:0] node39219;
	wire [4-1:0] node39220;
	wire [4-1:0] node39221;
	wire [4-1:0] node39222;
	wire [4-1:0] node39223;
	wire [4-1:0] node39226;
	wire [4-1:0] node39229;
	wire [4-1:0] node39230;
	wire [4-1:0] node39232;
	wire [4-1:0] node39235;
	wire [4-1:0] node39238;
	wire [4-1:0] node39239;
	wire [4-1:0] node39240;
	wire [4-1:0] node39243;
	wire [4-1:0] node39246;
	wire [4-1:0] node39247;
	wire [4-1:0] node39251;
	wire [4-1:0] node39252;
	wire [4-1:0] node39253;
	wire [4-1:0] node39254;
	wire [4-1:0] node39257;
	wire [4-1:0] node39260;
	wire [4-1:0] node39261;
	wire [4-1:0] node39262;
	wire [4-1:0] node39267;
	wire [4-1:0] node39268;
	wire [4-1:0] node39269;
	wire [4-1:0] node39270;
	wire [4-1:0] node39272;
	wire [4-1:0] node39275;
	wire [4-1:0] node39276;
	wire [4-1:0] node39281;
	wire [4-1:0] node39282;
	wire [4-1:0] node39285;
	wire [4-1:0] node39288;
	wire [4-1:0] node39289;
	wire [4-1:0] node39290;
	wire [4-1:0] node39291;
	wire [4-1:0] node39292;
	wire [4-1:0] node39293;
	wire [4-1:0] node39298;
	wire [4-1:0] node39299;
	wire [4-1:0] node39302;
	wire [4-1:0] node39305;
	wire [4-1:0] node39306;
	wire [4-1:0] node39307;
	wire [4-1:0] node39309;
	wire [4-1:0] node39310;
	wire [4-1:0] node39313;
	wire [4-1:0] node39316;
	wire [4-1:0] node39317;
	wire [4-1:0] node39318;
	wire [4-1:0] node39321;
	wire [4-1:0] node39325;
	wire [4-1:0] node39326;
	wire [4-1:0] node39328;
	wire [4-1:0] node39332;
	wire [4-1:0] node39333;
	wire [4-1:0] node39334;
	wire [4-1:0] node39335;
	wire [4-1:0] node39338;
	wire [4-1:0] node39341;
	wire [4-1:0] node39342;
	wire [4-1:0] node39343;
	wire [4-1:0] node39345;
	wire [4-1:0] node39349;
	wire [4-1:0] node39350;
	wire [4-1:0] node39354;
	wire [4-1:0] node39355;
	wire [4-1:0] node39356;
	wire [4-1:0] node39357;
	wire [4-1:0] node39360;
	wire [4-1:0] node39364;
	wire [4-1:0] node39365;
	wire [4-1:0] node39366;
	wire [4-1:0] node39369;
	wire [4-1:0] node39373;
	wire [4-1:0] node39374;
	wire [4-1:0] node39375;
	wire [4-1:0] node39376;
	wire [4-1:0] node39377;
	wire [4-1:0] node39378;
	wire [4-1:0] node39379;
	wire [4-1:0] node39382;
	wire [4-1:0] node39385;
	wire [4-1:0] node39386;
	wire [4-1:0] node39389;
	wire [4-1:0] node39392;
	wire [4-1:0] node39393;
	wire [4-1:0] node39394;
	wire [4-1:0] node39397;
	wire [4-1:0] node39400;
	wire [4-1:0] node39401;
	wire [4-1:0] node39405;
	wire [4-1:0] node39406;
	wire [4-1:0] node39408;
	wire [4-1:0] node39409;
	wire [4-1:0] node39412;
	wire [4-1:0] node39415;
	wire [4-1:0] node39416;
	wire [4-1:0] node39419;
	wire [4-1:0] node39422;
	wire [4-1:0] node39423;
	wire [4-1:0] node39424;
	wire [4-1:0] node39425;
	wire [4-1:0] node39427;
	wire [4-1:0] node39430;
	wire [4-1:0] node39431;
	wire [4-1:0] node39434;
	wire [4-1:0] node39437;
	wire [4-1:0] node39438;
	wire [4-1:0] node39440;
	wire [4-1:0] node39442;
	wire [4-1:0] node39445;
	wire [4-1:0] node39447;
	wire [4-1:0] node39448;
	wire [4-1:0] node39452;
	wire [4-1:0] node39453;
	wire [4-1:0] node39456;
	wire [4-1:0] node39458;
	wire [4-1:0] node39459;
	wire [4-1:0] node39463;
	wire [4-1:0] node39464;
	wire [4-1:0] node39465;
	wire [4-1:0] node39466;
	wire [4-1:0] node39467;
	wire [4-1:0] node39468;
	wire [4-1:0] node39469;
	wire [4-1:0] node39474;
	wire [4-1:0] node39475;
	wire [4-1:0] node39478;
	wire [4-1:0] node39481;
	wire [4-1:0] node39482;
	wire [4-1:0] node39486;
	wire [4-1:0] node39487;
	wire [4-1:0] node39490;
	wire [4-1:0] node39493;
	wire [4-1:0] node39494;
	wire [4-1:0] node39495;
	wire [4-1:0] node39496;
	wire [4-1:0] node39498;
	wire [4-1:0] node39501;
	wire [4-1:0] node39502;
	wire [4-1:0] node39506;
	wire [4-1:0] node39507;
	wire [4-1:0] node39508;
	wire [4-1:0] node39511;
	wire [4-1:0] node39514;
	wire [4-1:0] node39515;
	wire [4-1:0] node39519;
	wire [4-1:0] node39520;
	wire [4-1:0] node39521;
	wire [4-1:0] node39522;
	wire [4-1:0] node39526;
	wire [4-1:0] node39527;
	wire [4-1:0] node39531;
	wire [4-1:0] node39532;
	wire [4-1:0] node39535;
	wire [4-1:0] node39538;
	wire [4-1:0] node39539;
	wire [4-1:0] node39540;
	wire [4-1:0] node39541;
	wire [4-1:0] node39542;
	wire [4-1:0] node39543;
	wire [4-1:0] node39544;
	wire [4-1:0] node39545;
	wire [4-1:0] node39546;
	wire [4-1:0] node39547;
	wire [4-1:0] node39551;
	wire [4-1:0] node39554;
	wire [4-1:0] node39556;
	wire [4-1:0] node39559;
	wire [4-1:0] node39560;
	wire [4-1:0] node39561;
	wire [4-1:0] node39562;
	wire [4-1:0] node39565;
	wire [4-1:0] node39569;
	wire [4-1:0] node39570;
	wire [4-1:0] node39572;
	wire [4-1:0] node39576;
	wire [4-1:0] node39577;
	wire [4-1:0] node39578;
	wire [4-1:0] node39579;
	wire [4-1:0] node39583;
	wire [4-1:0] node39586;
	wire [4-1:0] node39587;
	wire [4-1:0] node39590;
	wire [4-1:0] node39593;
	wire [4-1:0] node39594;
	wire [4-1:0] node39595;
	wire [4-1:0] node39596;
	wire [4-1:0] node39600;
	wire [4-1:0] node39601;
	wire [4-1:0] node39603;
	wire [4-1:0] node39607;
	wire [4-1:0] node39608;
	wire [4-1:0] node39609;
	wire [4-1:0] node39610;
	wire [4-1:0] node39613;
	wire [4-1:0] node39616;
	wire [4-1:0] node39617;
	wire [4-1:0] node39621;
	wire [4-1:0] node39622;
	wire [4-1:0] node39625;
	wire [4-1:0] node39628;
	wire [4-1:0] node39629;
	wire [4-1:0] node39630;
	wire [4-1:0] node39631;
	wire [4-1:0] node39632;
	wire [4-1:0] node39635;
	wire [4-1:0] node39637;
	wire [4-1:0] node39640;
	wire [4-1:0] node39641;
	wire [4-1:0] node39642;
	wire [4-1:0] node39643;
	wire [4-1:0] node39648;
	wire [4-1:0] node39650;
	wire [4-1:0] node39652;
	wire [4-1:0] node39655;
	wire [4-1:0] node39656;
	wire [4-1:0] node39657;
	wire [4-1:0] node39658;
	wire [4-1:0] node39660;
	wire [4-1:0] node39663;
	wire [4-1:0] node39664;
	wire [4-1:0] node39668;
	wire [4-1:0] node39669;
	wire [4-1:0] node39670;
	wire [4-1:0] node39674;
	wire [4-1:0] node39676;
	wire [4-1:0] node39679;
	wire [4-1:0] node39680;
	wire [4-1:0] node39681;
	wire [4-1:0] node39683;
	wire [4-1:0] node39686;
	wire [4-1:0] node39689;
	wire [4-1:0] node39690;
	wire [4-1:0] node39694;
	wire [4-1:0] node39695;
	wire [4-1:0] node39696;
	wire [4-1:0] node39697;
	wire [4-1:0] node39699;
	wire [4-1:0] node39700;
	wire [4-1:0] node39703;
	wire [4-1:0] node39706;
	wire [4-1:0] node39708;
	wire [4-1:0] node39711;
	wire [4-1:0] node39712;
	wire [4-1:0] node39715;
	wire [4-1:0] node39716;
	wire [4-1:0] node39720;
	wire [4-1:0] node39721;
	wire [4-1:0] node39723;
	wire [4-1:0] node39724;
	wire [4-1:0] node39726;
	wire [4-1:0] node39729;
	wire [4-1:0] node39730;
	wire [4-1:0] node39733;
	wire [4-1:0] node39736;
	wire [4-1:0] node39737;
	wire [4-1:0] node39738;
	wire [4-1:0] node39739;
	wire [4-1:0] node39744;
	wire [4-1:0] node39746;
	wire [4-1:0] node39748;
	wire [4-1:0] node39751;
	wire [4-1:0] node39752;
	wire [4-1:0] node39753;
	wire [4-1:0] node39754;
	wire [4-1:0] node39755;
	wire [4-1:0] node39756;
	wire [4-1:0] node39759;
	wire [4-1:0] node39762;
	wire [4-1:0] node39763;
	wire [4-1:0] node39764;
	wire [4-1:0] node39767;
	wire [4-1:0] node39770;
	wire [4-1:0] node39771;
	wire [4-1:0] node39774;
	wire [4-1:0] node39775;
	wire [4-1:0] node39779;
	wire [4-1:0] node39780;
	wire [4-1:0] node39783;
	wire [4-1:0] node39786;
	wire [4-1:0] node39787;
	wire [4-1:0] node39788;
	wire [4-1:0] node39789;
	wire [4-1:0] node39790;
	wire [4-1:0] node39794;
	wire [4-1:0] node39795;
	wire [4-1:0] node39799;
	wire [4-1:0] node39800;
	wire [4-1:0] node39804;
	wire [4-1:0] node39805;
	wire [4-1:0] node39806;
	wire [4-1:0] node39808;
	wire [4-1:0] node39811;
	wire [4-1:0] node39812;
	wire [4-1:0] node39816;
	wire [4-1:0] node39817;
	wire [4-1:0] node39818;
	wire [4-1:0] node39819;
	wire [4-1:0] node39822;
	wire [4-1:0] node39827;
	wire [4-1:0] node39828;
	wire [4-1:0] node39829;
	wire [4-1:0] node39830;
	wire [4-1:0] node39832;
	wire [4-1:0] node39835;
	wire [4-1:0] node39838;
	wire [4-1:0] node39839;
	wire [4-1:0] node39840;
	wire [4-1:0] node39842;
	wire [4-1:0] node39844;
	wire [4-1:0] node39847;
	wire [4-1:0] node39848;
	wire [4-1:0] node39849;
	wire [4-1:0] node39854;
	wire [4-1:0] node39855;
	wire [4-1:0] node39858;
	wire [4-1:0] node39861;
	wire [4-1:0] node39862;
	wire [4-1:0] node39863;
	wire [4-1:0] node39864;
	wire [4-1:0] node39866;
	wire [4-1:0] node39869;
	wire [4-1:0] node39870;
	wire [4-1:0] node39874;
	wire [4-1:0] node39876;
	wire [4-1:0] node39879;
	wire [4-1:0] node39880;
	wire [4-1:0] node39881;
	wire [4-1:0] node39883;
	wire [4-1:0] node39886;
	wire [4-1:0] node39888;
	wire [4-1:0] node39889;
	wire [4-1:0] node39893;
	wire [4-1:0] node39894;
	wire [4-1:0] node39895;
	wire [4-1:0] node39898;
	wire [4-1:0] node39902;
	wire [4-1:0] node39903;
	wire [4-1:0] node39904;
	wire [4-1:0] node39905;
	wire [4-1:0] node39906;
	wire [4-1:0] node39907;
	wire [4-1:0] node39910;
	wire [4-1:0] node39911;
	wire [4-1:0] node39915;
	wire [4-1:0] node39916;
	wire [4-1:0] node39917;
	wire [4-1:0] node39920;
	wire [4-1:0] node39923;
	wire [4-1:0] node39924;
	wire [4-1:0] node39927;
	wire [4-1:0] node39930;
	wire [4-1:0] node39931;
	wire [4-1:0] node39932;
	wire [4-1:0] node39933;
	wire [4-1:0] node39934;
	wire [4-1:0] node39937;
	wire [4-1:0] node39940;
	wire [4-1:0] node39941;
	wire [4-1:0] node39945;
	wire [4-1:0] node39947;
	wire [4-1:0] node39949;
	wire [4-1:0] node39952;
	wire [4-1:0] node39954;
	wire [4-1:0] node39955;
	wire [4-1:0] node39958;
	wire [4-1:0] node39961;
	wire [4-1:0] node39962;
	wire [4-1:0] node39963;
	wire [4-1:0] node39964;
	wire [4-1:0] node39966;
	wire [4-1:0] node39967;
	wire [4-1:0] node39971;
	wire [4-1:0] node39972;
	wire [4-1:0] node39973;
	wire [4-1:0] node39974;
	wire [4-1:0] node39977;
	wire [4-1:0] node39980;
	wire [4-1:0] node39981;
	wire [4-1:0] node39985;
	wire [4-1:0] node39987;
	wire [4-1:0] node39989;
	wire [4-1:0] node39992;
	wire [4-1:0] node39993;
	wire [4-1:0] node39994;
	wire [4-1:0] node39997;
	wire [4-1:0] node40001;
	wire [4-1:0] node40002;
	wire [4-1:0] node40003;
	wire [4-1:0] node40004;
	wire [4-1:0] node40005;
	wire [4-1:0] node40006;
	wire [4-1:0] node40011;
	wire [4-1:0] node40013;
	wire [4-1:0] node40014;
	wire [4-1:0] node40018;
	wire [4-1:0] node40020;
	wire [4-1:0] node40022;
	wire [4-1:0] node40023;
	wire [4-1:0] node40027;
	wire [4-1:0] node40028;
	wire [4-1:0] node40029;
	wire [4-1:0] node40030;
	wire [4-1:0] node40033;
	wire [4-1:0] node40036;
	wire [4-1:0] node40038;
	wire [4-1:0] node40039;
	wire [4-1:0] node40043;
	wire [4-1:0] node40044;
	wire [4-1:0] node40045;
	wire [4-1:0] node40048;
	wire [4-1:0] node40052;
	wire [4-1:0] node40053;
	wire [4-1:0] node40054;
	wire [4-1:0] node40055;
	wire [4-1:0] node40056;
	wire [4-1:0] node40058;
	wire [4-1:0] node40059;
	wire [4-1:0] node40060;
	wire [4-1:0] node40064;
	wire [4-1:0] node40067;
	wire [4-1:0] node40068;
	wire [4-1:0] node40072;
	wire [4-1:0] node40073;
	wire [4-1:0] node40074;
	wire [4-1:0] node40075;
	wire [4-1:0] node40077;
	wire [4-1:0] node40080;
	wire [4-1:0] node40082;
	wire [4-1:0] node40085;
	wire [4-1:0] node40086;
	wire [4-1:0] node40090;
	wire [4-1:0] node40092;
	wire [4-1:0] node40094;
	wire [4-1:0] node40097;
	wire [4-1:0] node40098;
	wire [4-1:0] node40099;
	wire [4-1:0] node40100;
	wire [4-1:0] node40101;
	wire [4-1:0] node40105;
	wire [4-1:0] node40106;
	wire [4-1:0] node40110;
	wire [4-1:0] node40111;
	wire [4-1:0] node40113;
	wire [4-1:0] node40115;
	wire [4-1:0] node40118;
	wire [4-1:0] node40119;
	wire [4-1:0] node40120;
	wire [4-1:0] node40123;
	wire [4-1:0] node40127;
	wire [4-1:0] node40128;
	wire [4-1:0] node40131;
	wire [4-1:0] node40132;
	wire [4-1:0] node40133;
	wire [4-1:0] node40137;
	wire [4-1:0] node40138;
	wire [4-1:0] node40142;
	wire [4-1:0] node40143;
	wire [4-1:0] node40144;
	wire [4-1:0] node40145;
	wire [4-1:0] node40147;
	wire [4-1:0] node40148;
	wire [4-1:0] node40151;
	wire [4-1:0] node40154;
	wire [4-1:0] node40155;
	wire [4-1:0] node40156;
	wire [4-1:0] node40159;
	wire [4-1:0] node40162;
	wire [4-1:0] node40163;
	wire [4-1:0] node40166;
	wire [4-1:0] node40169;
	wire [4-1:0] node40170;
	wire [4-1:0] node40171;
	wire [4-1:0] node40172;
	wire [4-1:0] node40177;
	wire [4-1:0] node40178;
	wire [4-1:0] node40181;
	wire [4-1:0] node40182;
	wire [4-1:0] node40186;
	wire [4-1:0] node40187;
	wire [4-1:0] node40188;
	wire [4-1:0] node40189;
	wire [4-1:0] node40191;
	wire [4-1:0] node40192;
	wire [4-1:0] node40195;
	wire [4-1:0] node40198;
	wire [4-1:0] node40200;
	wire [4-1:0] node40203;
	wire [4-1:0] node40204;
	wire [4-1:0] node40206;
	wire [4-1:0] node40208;
	wire [4-1:0] node40212;
	wire [4-1:0] node40213;
	wire [4-1:0] node40214;
	wire [4-1:0] node40218;
	wire [4-1:0] node40220;
	wire [4-1:0] node40221;
	wire [4-1:0] node40222;
	wire [4-1:0] node40225;
	wire [4-1:0] node40229;
	wire [4-1:0] node40230;
	wire [4-1:0] node40231;
	wire [4-1:0] node40232;
	wire [4-1:0] node40233;
	wire [4-1:0] node40234;
	wire [4-1:0] node40235;
	wire [4-1:0] node40236;
	wire [4-1:0] node40238;
	wire [4-1:0] node40239;
	wire [4-1:0] node40241;
	wire [4-1:0] node40245;
	wire [4-1:0] node40246;
	wire [4-1:0] node40247;
	wire [4-1:0] node40251;
	wire [4-1:0] node40252;
	wire [4-1:0] node40255;
	wire [4-1:0] node40258;
	wire [4-1:0] node40259;
	wire [4-1:0] node40260;
	wire [4-1:0] node40261;
	wire [4-1:0] node40262;
	wire [4-1:0] node40265;
	wire [4-1:0] node40269;
	wire [4-1:0] node40272;
	wire [4-1:0] node40273;
	wire [4-1:0] node40274;
	wire [4-1:0] node40278;
	wire [4-1:0] node40279;
	wire [4-1:0] node40283;
	wire [4-1:0] node40284;
	wire [4-1:0] node40285;
	wire [4-1:0] node40286;
	wire [4-1:0] node40290;
	wire [4-1:0] node40293;
	wire [4-1:0] node40294;
	wire [4-1:0] node40295;
	wire [4-1:0] node40296;
	wire [4-1:0] node40300;
	wire [4-1:0] node40303;
	wire [4-1:0] node40304;
	wire [4-1:0] node40305;
	wire [4-1:0] node40309;
	wire [4-1:0] node40310;
	wire [4-1:0] node40313;
	wire [4-1:0] node40314;
	wire [4-1:0] node40318;
	wire [4-1:0] node40319;
	wire [4-1:0] node40320;
	wire [4-1:0] node40321;
	wire [4-1:0] node40322;
	wire [4-1:0] node40326;
	wire [4-1:0] node40327;
	wire [4-1:0] node40331;
	wire [4-1:0] node40332;
	wire [4-1:0] node40333;
	wire [4-1:0] node40337;
	wire [4-1:0] node40338;
	wire [4-1:0] node40342;
	wire [4-1:0] node40343;
	wire [4-1:0] node40345;
	wire [4-1:0] node40348;
	wire [4-1:0] node40350;
	wire [4-1:0] node40351;
	wire [4-1:0] node40355;
	wire [4-1:0] node40356;
	wire [4-1:0] node40357;
	wire [4-1:0] node40358;
	wire [4-1:0] node40359;
	wire [4-1:0] node40360;
	wire [4-1:0] node40363;
	wire [4-1:0] node40366;
	wire [4-1:0] node40367;
	wire [4-1:0] node40370;
	wire [4-1:0] node40373;
	wire [4-1:0] node40374;
	wire [4-1:0] node40375;
	wire [4-1:0] node40376;
	wire [4-1:0] node40379;
	wire [4-1:0] node40382;
	wire [4-1:0] node40383;
	wire [4-1:0] node40387;
	wire [4-1:0] node40388;
	wire [4-1:0] node40391;
	wire [4-1:0] node40394;
	wire [4-1:0] node40395;
	wire [4-1:0] node40396;
	wire [4-1:0] node40398;
	wire [4-1:0] node40400;
	wire [4-1:0] node40401;
	wire [4-1:0] node40404;
	wire [4-1:0] node40407;
	wire [4-1:0] node40410;
	wire [4-1:0] node40411;
	wire [4-1:0] node40412;
	wire [4-1:0] node40414;
	wire [4-1:0] node40418;
	wire [4-1:0] node40419;
	wire [4-1:0] node40421;
	wire [4-1:0] node40422;
	wire [4-1:0] node40427;
	wire [4-1:0] node40428;
	wire [4-1:0] node40429;
	wire [4-1:0] node40430;
	wire [4-1:0] node40431;
	wire [4-1:0] node40433;
	wire [4-1:0] node40436;
	wire [4-1:0] node40437;
	wire [4-1:0] node40440;
	wire [4-1:0] node40443;
	wire [4-1:0] node40444;
	wire [4-1:0] node40445;
	wire [4-1:0] node40448;
	wire [4-1:0] node40452;
	wire [4-1:0] node40453;
	wire [4-1:0] node40454;
	wire [4-1:0] node40455;
	wire [4-1:0] node40458;
	wire [4-1:0] node40461;
	wire [4-1:0] node40462;
	wire [4-1:0] node40465;
	wire [4-1:0] node40468;
	wire [4-1:0] node40469;
	wire [4-1:0] node40470;
	wire [4-1:0] node40473;
	wire [4-1:0] node40477;
	wire [4-1:0] node40478;
	wire [4-1:0] node40479;
	wire [4-1:0] node40481;
	wire [4-1:0] node40482;
	wire [4-1:0] node40486;
	wire [4-1:0] node40487;
	wire [4-1:0] node40489;
	wire [4-1:0] node40493;
	wire [4-1:0] node40494;
	wire [4-1:0] node40495;
	wire [4-1:0] node40498;
	wire [4-1:0] node40501;
	wire [4-1:0] node40502;
	wire [4-1:0] node40504;
	wire [4-1:0] node40507;
	wire [4-1:0] node40508;
	wire [4-1:0] node40511;
	wire [4-1:0] node40514;
	wire [4-1:0] node40515;
	wire [4-1:0] node40516;
	wire [4-1:0] node40517;
	wire [4-1:0] node40518;
	wire [4-1:0] node40519;
	wire [4-1:0] node40520;
	wire [4-1:0] node40523;
	wire [4-1:0] node40526;
	wire [4-1:0] node40529;
	wire [4-1:0] node40530;
	wire [4-1:0] node40531;
	wire [4-1:0] node40532;
	wire [4-1:0] node40533;
	wire [4-1:0] node40537;
	wire [4-1:0] node40538;
	wire [4-1:0] node40541;
	wire [4-1:0] node40545;
	wire [4-1:0] node40547;
	wire [4-1:0] node40549;
	wire [4-1:0] node40552;
	wire [4-1:0] node40553;
	wire [4-1:0] node40554;
	wire [4-1:0] node40555;
	wire [4-1:0] node40558;
	wire [4-1:0] node40561;
	wire [4-1:0] node40562;
	wire [4-1:0] node40564;
	wire [4-1:0] node40565;
	wire [4-1:0] node40570;
	wire [4-1:0] node40571;
	wire [4-1:0] node40573;
	wire [4-1:0] node40574;
	wire [4-1:0] node40577;
	wire [4-1:0] node40580;
	wire [4-1:0] node40581;
	wire [4-1:0] node40584;
	wire [4-1:0] node40587;
	wire [4-1:0] node40588;
	wire [4-1:0] node40589;
	wire [4-1:0] node40590;
	wire [4-1:0] node40591;
	wire [4-1:0] node40595;
	wire [4-1:0] node40597;
	wire [4-1:0] node40598;
	wire [4-1:0] node40601;
	wire [4-1:0] node40604;
	wire [4-1:0] node40605;
	wire [4-1:0] node40606;
	wire [4-1:0] node40607;
	wire [4-1:0] node40610;
	wire [4-1:0] node40614;
	wire [4-1:0] node40615;
	wire [4-1:0] node40616;
	wire [4-1:0] node40621;
	wire [4-1:0] node40622;
	wire [4-1:0] node40623;
	wire [4-1:0] node40625;
	wire [4-1:0] node40627;
	wire [4-1:0] node40630;
	wire [4-1:0] node40632;
	wire [4-1:0] node40633;
	wire [4-1:0] node40636;
	wire [4-1:0] node40639;
	wire [4-1:0] node40640;
	wire [4-1:0] node40641;
	wire [4-1:0] node40642;
	wire [4-1:0] node40643;
	wire [4-1:0] node40646;
	wire [4-1:0] node40650;
	wire [4-1:0] node40651;
	wire [4-1:0] node40655;
	wire [4-1:0] node40657;
	wire [4-1:0] node40660;
	wire [4-1:0] node40661;
	wire [4-1:0] node40662;
	wire [4-1:0] node40663;
	wire [4-1:0] node40664;
	wire [4-1:0] node40665;
	wire [4-1:0] node40666;
	wire [4-1:0] node40667;
	wire [4-1:0] node40670;
	wire [4-1:0] node40673;
	wire [4-1:0] node40674;
	wire [4-1:0] node40677;
	wire [4-1:0] node40681;
	wire [4-1:0] node40682;
	wire [4-1:0] node40685;
	wire [4-1:0] node40688;
	wire [4-1:0] node40689;
	wire [4-1:0] node40690;
	wire [4-1:0] node40692;
	wire [4-1:0] node40694;
	wire [4-1:0] node40697;
	wire [4-1:0] node40698;
	wire [4-1:0] node40701;
	wire [4-1:0] node40704;
	wire [4-1:0] node40705;
	wire [4-1:0] node40708;
	wire [4-1:0] node40709;
	wire [4-1:0] node40712;
	wire [4-1:0] node40715;
	wire [4-1:0] node40716;
	wire [4-1:0] node40717;
	wire [4-1:0] node40718;
	wire [4-1:0] node40721;
	wire [4-1:0] node40724;
	wire [4-1:0] node40725;
	wire [4-1:0] node40726;
	wire [4-1:0] node40727;
	wire [4-1:0] node40730;
	wire [4-1:0] node40733;
	wire [4-1:0] node40735;
	wire [4-1:0] node40739;
	wire [4-1:0] node40740;
	wire [4-1:0] node40741;
	wire [4-1:0] node40744;
	wire [4-1:0] node40747;
	wire [4-1:0] node40748;
	wire [4-1:0] node40749;
	wire [4-1:0] node40751;
	wire [4-1:0] node40754;
	wire [4-1:0] node40755;
	wire [4-1:0] node40759;
	wire [4-1:0] node40760;
	wire [4-1:0] node40764;
	wire [4-1:0] node40765;
	wire [4-1:0] node40766;
	wire [4-1:0] node40767;
	wire [4-1:0] node40769;
	wire [4-1:0] node40770;
	wire [4-1:0] node40774;
	wire [4-1:0] node40777;
	wire [4-1:0] node40778;
	wire [4-1:0] node40779;
	wire [4-1:0] node40782;
	wire [4-1:0] node40784;
	wire [4-1:0] node40787;
	wire [4-1:0] node40788;
	wire [4-1:0] node40792;
	wire [4-1:0] node40793;
	wire [4-1:0] node40794;
	wire [4-1:0] node40795;
	wire [4-1:0] node40796;
	wire [4-1:0] node40800;
	wire [4-1:0] node40801;
	wire [4-1:0] node40805;
	wire [4-1:0] node40806;
	wire [4-1:0] node40809;
	wire [4-1:0] node40812;
	wire [4-1:0] node40813;
	wire [4-1:0] node40814;
	wire [4-1:0] node40815;
	wire [4-1:0] node40819;
	wire [4-1:0] node40822;
	wire [4-1:0] node40823;
	wire [4-1:0] node40824;
	wire [4-1:0] node40828;
	wire [4-1:0] node40829;
	wire [4-1:0] node40830;
	wire [4-1:0] node40833;
	wire [4-1:0] node40837;
	wire [4-1:0] node40838;
	wire [4-1:0] node40839;
	wire [4-1:0] node40840;
	wire [4-1:0] node40841;
	wire [4-1:0] node40842;
	wire [4-1:0] node40843;
	wire [4-1:0] node40844;
	wire [4-1:0] node40846;
	wire [4-1:0] node40848;
	wire [4-1:0] node40852;
	wire [4-1:0] node40854;
	wire [4-1:0] node40855;
	wire [4-1:0] node40856;
	wire [4-1:0] node40859;
	wire [4-1:0] node40863;
	wire [4-1:0] node40864;
	wire [4-1:0] node40865;
	wire [4-1:0] node40866;
	wire [4-1:0] node40869;
	wire [4-1:0] node40873;
	wire [4-1:0] node40874;
	wire [4-1:0] node40877;
	wire [4-1:0] node40880;
	wire [4-1:0] node40881;
	wire [4-1:0] node40882;
	wire [4-1:0] node40883;
	wire [4-1:0] node40884;
	wire [4-1:0] node40885;
	wire [4-1:0] node40888;
	wire [4-1:0] node40893;
	wire [4-1:0] node40895;
	wire [4-1:0] node40896;
	wire [4-1:0] node40898;
	wire [4-1:0] node40902;
	wire [4-1:0] node40903;
	wire [4-1:0] node40904;
	wire [4-1:0] node40905;
	wire [4-1:0] node40906;
	wire [4-1:0] node40910;
	wire [4-1:0] node40912;
	wire [4-1:0] node40916;
	wire [4-1:0] node40918;
	wire [4-1:0] node40921;
	wire [4-1:0] node40922;
	wire [4-1:0] node40923;
	wire [4-1:0] node40924;
	wire [4-1:0] node40925;
	wire [4-1:0] node40926;
	wire [4-1:0] node40929;
	wire [4-1:0] node40930;
	wire [4-1:0] node40934;
	wire [4-1:0] node40936;
	wire [4-1:0] node40938;
	wire [4-1:0] node40941;
	wire [4-1:0] node40942;
	wire [4-1:0] node40946;
	wire [4-1:0] node40947;
	wire [4-1:0] node40948;
	wire [4-1:0] node40949;
	wire [4-1:0] node40952;
	wire [4-1:0] node40954;
	wire [4-1:0] node40957;
	wire [4-1:0] node40959;
	wire [4-1:0] node40962;
	wire [4-1:0] node40964;
	wire [4-1:0] node40965;
	wire [4-1:0] node40967;
	wire [4-1:0] node40970;
	wire [4-1:0] node40973;
	wire [4-1:0] node40974;
	wire [4-1:0] node40975;
	wire [4-1:0] node40977;
	wire [4-1:0] node40979;
	wire [4-1:0] node40980;
	wire [4-1:0] node40983;
	wire [4-1:0] node40986;
	wire [4-1:0] node40987;
	wire [4-1:0] node40988;
	wire [4-1:0] node40990;
	wire [4-1:0] node40995;
	wire [4-1:0] node40996;
	wire [4-1:0] node40997;
	wire [4-1:0] node40998;
	wire [4-1:0] node40999;
	wire [4-1:0] node41002;
	wire [4-1:0] node41005;
	wire [4-1:0] node41006;
	wire [4-1:0] node41010;
	wire [4-1:0] node41011;
	wire [4-1:0] node41015;
	wire [4-1:0] node41016;
	wire [4-1:0] node41019;
	wire [4-1:0] node41022;
	wire [4-1:0] node41023;
	wire [4-1:0] node41024;
	wire [4-1:0] node41025;
	wire [4-1:0] node41026;
	wire [4-1:0] node41027;
	wire [4-1:0] node41028;
	wire [4-1:0] node41033;
	wire [4-1:0] node41035;
	wire [4-1:0] node41037;
	wire [4-1:0] node41038;
	wire [4-1:0] node41041;
	wire [4-1:0] node41044;
	wire [4-1:0] node41045;
	wire [4-1:0] node41046;
	wire [4-1:0] node41050;
	wire [4-1:0] node41052;
	wire [4-1:0] node41055;
	wire [4-1:0] node41056;
	wire [4-1:0] node41057;
	wire [4-1:0] node41058;
	wire [4-1:0] node41060;
	wire [4-1:0] node41062;
	wire [4-1:0] node41065;
	wire [4-1:0] node41066;
	wire [4-1:0] node41067;
	wire [4-1:0] node41070;
	wire [4-1:0] node41074;
	wire [4-1:0] node41075;
	wire [4-1:0] node41076;
	wire [4-1:0] node41079;
	wire [4-1:0] node41080;
	wire [4-1:0] node41085;
	wire [4-1:0] node41086;
	wire [4-1:0] node41087;
	wire [4-1:0] node41090;
	wire [4-1:0] node41093;
	wire [4-1:0] node41094;
	wire [4-1:0] node41097;
	wire [4-1:0] node41100;
	wire [4-1:0] node41101;
	wire [4-1:0] node41102;
	wire [4-1:0] node41103;
	wire [4-1:0] node41105;
	wire [4-1:0] node41107;
	wire [4-1:0] node41108;
	wire [4-1:0] node41111;
	wire [4-1:0] node41114;
	wire [4-1:0] node41116;
	wire [4-1:0] node41118;
	wire [4-1:0] node41119;
	wire [4-1:0] node41122;
	wire [4-1:0] node41125;
	wire [4-1:0] node41126;
	wire [4-1:0] node41127;
	wire [4-1:0] node41130;
	wire [4-1:0] node41133;
	wire [4-1:0] node41135;
	wire [4-1:0] node41138;
	wire [4-1:0] node41139;
	wire [4-1:0] node41140;
	wire [4-1:0] node41141;
	wire [4-1:0] node41145;
	wire [4-1:0] node41147;
	wire [4-1:0] node41148;
	wire [4-1:0] node41152;
	wire [4-1:0] node41153;
	wire [4-1:0] node41154;
	wire [4-1:0] node41157;
	wire [4-1:0] node41160;
	wire [4-1:0] node41161;
	wire [4-1:0] node41163;
	wire [4-1:0] node41165;
	wire [4-1:0] node41168;
	wire [4-1:0] node41169;
	wire [4-1:0] node41173;
	wire [4-1:0] node41174;
	wire [4-1:0] node41175;
	wire [4-1:0] node41176;
	wire [4-1:0] node41177;
	wire [4-1:0] node41178;
	wire [4-1:0] node41181;
	wire [4-1:0] node41182;
	wire [4-1:0] node41184;
	wire [4-1:0] node41187;
	wire [4-1:0] node41189;
	wire [4-1:0] node41192;
	wire [4-1:0] node41193;
	wire [4-1:0] node41194;
	wire [4-1:0] node41197;
	wire [4-1:0] node41200;
	wire [4-1:0] node41201;
	wire [4-1:0] node41205;
	wire [4-1:0] node41206;
	wire [4-1:0] node41207;
	wire [4-1:0] node41208;
	wire [4-1:0] node41210;
	wire [4-1:0] node41213;
	wire [4-1:0] node41214;
	wire [4-1:0] node41217;
	wire [4-1:0] node41220;
	wire [4-1:0] node41222;
	wire [4-1:0] node41223;
	wire [4-1:0] node41226;
	wire [4-1:0] node41229;
	wire [4-1:0] node41230;
	wire [4-1:0] node41231;
	wire [4-1:0] node41234;
	wire [4-1:0] node41237;
	wire [4-1:0] node41239;
	wire [4-1:0] node41242;
	wire [4-1:0] node41243;
	wire [4-1:0] node41244;
	wire [4-1:0] node41245;
	wire [4-1:0] node41246;
	wire [4-1:0] node41247;
	wire [4-1:0] node41248;
	wire [4-1:0] node41251;
	wire [4-1:0] node41255;
	wire [4-1:0] node41256;
	wire [4-1:0] node41260;
	wire [4-1:0] node41261;
	wire [4-1:0] node41264;
	wire [4-1:0] node41266;
	wire [4-1:0] node41269;
	wire [4-1:0] node41270;
	wire [4-1:0] node41272;
	wire [4-1:0] node41273;
	wire [4-1:0] node41274;
	wire [4-1:0] node41278;
	wire [4-1:0] node41279;
	wire [4-1:0] node41283;
	wire [4-1:0] node41284;
	wire [4-1:0] node41285;
	wire [4-1:0] node41286;
	wire [4-1:0] node41289;
	wire [4-1:0] node41293;
	wire [4-1:0] node41295;
	wire [4-1:0] node41296;
	wire [4-1:0] node41299;
	wire [4-1:0] node41302;
	wire [4-1:0] node41303;
	wire [4-1:0] node41304;
	wire [4-1:0] node41305;
	wire [4-1:0] node41308;
	wire [4-1:0] node41309;
	wire [4-1:0] node41313;
	wire [4-1:0] node41314;
	wire [4-1:0] node41317;
	wire [4-1:0] node41319;
	wire [4-1:0] node41322;
	wire [4-1:0] node41323;
	wire [4-1:0] node41324;
	wire [4-1:0] node41325;
	wire [4-1:0] node41329;
	wire [4-1:0] node41331;
	wire [4-1:0] node41334;
	wire [4-1:0] node41335;
	wire [4-1:0] node41338;
	wire [4-1:0] node41341;
	wire [4-1:0] node41342;
	wire [4-1:0] node41343;
	wire [4-1:0] node41344;
	wire [4-1:0] node41345;
	wire [4-1:0] node41347;
	wire [4-1:0] node41349;
	wire [4-1:0] node41352;
	wire [4-1:0] node41354;
	wire [4-1:0] node41356;
	wire [4-1:0] node41359;
	wire [4-1:0] node41360;
	wire [4-1:0] node41361;
	wire [4-1:0] node41364;
	wire [4-1:0] node41367;
	wire [4-1:0] node41368;
	wire [4-1:0] node41369;
	wire [4-1:0] node41374;
	wire [4-1:0] node41375;
	wire [4-1:0] node41376;
	wire [4-1:0] node41377;
	wire [4-1:0] node41378;
	wire [4-1:0] node41382;
	wire [4-1:0] node41383;
	wire [4-1:0] node41386;
	wire [4-1:0] node41389;
	wire [4-1:0] node41391;
	wire [4-1:0] node41392;
	wire [4-1:0] node41395;
	wire [4-1:0] node41398;
	wire [4-1:0] node41399;
	wire [4-1:0] node41401;
	wire [4-1:0] node41404;
	wire [4-1:0] node41406;
	wire [4-1:0] node41409;
	wire [4-1:0] node41410;
	wire [4-1:0] node41411;
	wire [4-1:0] node41412;
	wire [4-1:0] node41413;
	wire [4-1:0] node41415;
	wire [4-1:0] node41418;
	wire [4-1:0] node41419;
	wire [4-1:0] node41423;
	wire [4-1:0] node41424;
	wire [4-1:0] node41426;
	wire [4-1:0] node41430;
	wire [4-1:0] node41431;
	wire [4-1:0] node41432;
	wire [4-1:0] node41433;
	wire [4-1:0] node41436;
	wire [4-1:0] node41439;
	wire [4-1:0] node41440;
	wire [4-1:0] node41443;
	wire [4-1:0] node41446;
	wire [4-1:0] node41447;
	wire [4-1:0] node41450;
	wire [4-1:0] node41453;
	wire [4-1:0] node41454;
	wire [4-1:0] node41455;
	wire [4-1:0] node41456;
	wire [4-1:0] node41458;
	wire [4-1:0] node41462;
	wire [4-1:0] node41464;
	wire [4-1:0] node41465;
	wire [4-1:0] node41469;
	wire [4-1:0] node41470;
	wire [4-1:0] node41471;
	wire [4-1:0] node41474;
	wire [4-1:0] node41475;
	wire [4-1:0] node41476;
	wire [4-1:0] node41479;
	wire [4-1:0] node41482;
	wire [4-1:0] node41483;
	wire [4-1:0] node41487;
	wire [4-1:0] node41489;
	wire [4-1:0] node41490;
	wire [4-1:0] node41493;
	wire [4-1:0] node41496;
	wire [4-1:0] node41497;
	wire [4-1:0] node41498;
	wire [4-1:0] node41499;
	wire [4-1:0] node41500;
	wire [4-1:0] node41501;
	wire [4-1:0] node41502;
	wire [4-1:0] node41503;
	wire [4-1:0] node41504;
	wire [4-1:0] node41506;
	wire [4-1:0] node41507;
	wire [4-1:0] node41508;
	wire [4-1:0] node41511;
	wire [4-1:0] node41515;
	wire [4-1:0] node41516;
	wire [4-1:0] node41519;
	wire [4-1:0] node41521;
	wire [4-1:0] node41524;
	wire [4-1:0] node41525;
	wire [4-1:0] node41526;
	wire [4-1:0] node41528;
	wire [4-1:0] node41529;
	wire [4-1:0] node41533;
	wire [4-1:0] node41535;
	wire [4-1:0] node41538;
	wire [4-1:0] node41539;
	wire [4-1:0] node41542;
	wire [4-1:0] node41545;
	wire [4-1:0] node41546;
	wire [4-1:0] node41547;
	wire [4-1:0] node41549;
	wire [4-1:0] node41550;
	wire [4-1:0] node41551;
	wire [4-1:0] node41554;
	wire [4-1:0] node41558;
	wire [4-1:0] node41559;
	wire [4-1:0] node41560;
	wire [4-1:0] node41563;
	wire [4-1:0] node41566;
	wire [4-1:0] node41567;
	wire [4-1:0] node41570;
	wire [4-1:0] node41573;
	wire [4-1:0] node41574;
	wire [4-1:0] node41576;
	wire [4-1:0] node41577;
	wire [4-1:0] node41578;
	wire [4-1:0] node41583;
	wire [4-1:0] node41584;
	wire [4-1:0] node41586;
	wire [4-1:0] node41589;
	wire [4-1:0] node41590;
	wire [4-1:0] node41594;
	wire [4-1:0] node41595;
	wire [4-1:0] node41596;
	wire [4-1:0] node41597;
	wire [4-1:0] node41598;
	wire [4-1:0] node41599;
	wire [4-1:0] node41601;
	wire [4-1:0] node41605;
	wire [4-1:0] node41606;
	wire [4-1:0] node41610;
	wire [4-1:0] node41611;
	wire [4-1:0] node41612;
	wire [4-1:0] node41615;
	wire [4-1:0] node41618;
	wire [4-1:0] node41619;
	wire [4-1:0] node41623;
	wire [4-1:0] node41624;
	wire [4-1:0] node41625;
	wire [4-1:0] node41627;
	wire [4-1:0] node41630;
	wire [4-1:0] node41633;
	wire [4-1:0] node41634;
	wire [4-1:0] node41635;
	wire [4-1:0] node41636;
	wire [4-1:0] node41639;
	wire [4-1:0] node41644;
	wire [4-1:0] node41645;
	wire [4-1:0] node41646;
	wire [4-1:0] node41647;
	wire [4-1:0] node41648;
	wire [4-1:0] node41649;
	wire [4-1:0] node41652;
	wire [4-1:0] node41656;
	wire [4-1:0] node41657;
	wire [4-1:0] node41661;
	wire [4-1:0] node41662;
	wire [4-1:0] node41664;
	wire [4-1:0] node41667;
	wire [4-1:0] node41668;
	wire [4-1:0] node41671;
	wire [4-1:0] node41674;
	wire [4-1:0] node41675;
	wire [4-1:0] node41676;
	wire [4-1:0] node41678;
	wire [4-1:0] node41681;
	wire [4-1:0] node41683;
	wire [4-1:0] node41686;
	wire [4-1:0] node41688;
	wire [4-1:0] node41689;
	wire [4-1:0] node41692;
	wire [4-1:0] node41695;
	wire [4-1:0] node41696;
	wire [4-1:0] node41697;
	wire [4-1:0] node41698;
	wire [4-1:0] node41699;
	wire [4-1:0] node41700;
	wire [4-1:0] node41702;
	wire [4-1:0] node41705;
	wire [4-1:0] node41706;
	wire [4-1:0] node41709;
	wire [4-1:0] node41712;
	wire [4-1:0] node41713;
	wire [4-1:0] node41714;
	wire [4-1:0] node41717;
	wire [4-1:0] node41721;
	wire [4-1:0] node41722;
	wire [4-1:0] node41723;
	wire [4-1:0] node41724;
	wire [4-1:0] node41727;
	wire [4-1:0] node41730;
	wire [4-1:0] node41731;
	wire [4-1:0] node41734;
	wire [4-1:0] node41737;
	wire [4-1:0] node41738;
	wire [4-1:0] node41739;
	wire [4-1:0] node41740;
	wire [4-1:0] node41744;
	wire [4-1:0] node41746;
	wire [4-1:0] node41749;
	wire [4-1:0] node41750;
	wire [4-1:0] node41754;
	wire [4-1:0] node41755;
	wire [4-1:0] node41756;
	wire [4-1:0] node41757;
	wire [4-1:0] node41758;
	wire [4-1:0] node41763;
	wire [4-1:0] node41765;
	wire [4-1:0] node41766;
	wire [4-1:0] node41770;
	wire [4-1:0] node41771;
	wire [4-1:0] node41772;
	wire [4-1:0] node41773;
	wire [4-1:0] node41776;
	wire [4-1:0] node41779;
	wire [4-1:0] node41781;
	wire [4-1:0] node41784;
	wire [4-1:0] node41785;
	wire [4-1:0] node41787;
	wire [4-1:0] node41790;
	wire [4-1:0] node41793;
	wire [4-1:0] node41794;
	wire [4-1:0] node41795;
	wire [4-1:0] node41796;
	wire [4-1:0] node41797;
	wire [4-1:0] node41798;
	wire [4-1:0] node41801;
	wire [4-1:0] node41805;
	wire [4-1:0] node41806;
	wire [4-1:0] node41807;
	wire [4-1:0] node41808;
	wire [4-1:0] node41812;
	wire [4-1:0] node41814;
	wire [4-1:0] node41817;
	wire [4-1:0] node41818;
	wire [4-1:0] node41822;
	wire [4-1:0] node41823;
	wire [4-1:0] node41824;
	wire [4-1:0] node41825;
	wire [4-1:0] node41829;
	wire [4-1:0] node41832;
	wire [4-1:0] node41833;
	wire [4-1:0] node41836;
	wire [4-1:0] node41839;
	wire [4-1:0] node41840;
	wire [4-1:0] node41841;
	wire [4-1:0] node41842;
	wire [4-1:0] node41844;
	wire [4-1:0] node41847;
	wire [4-1:0] node41849;
	wire [4-1:0] node41852;
	wire [4-1:0] node41853;
	wire [4-1:0] node41854;
	wire [4-1:0] node41856;
	wire [4-1:0] node41859;
	wire [4-1:0] node41861;
	wire [4-1:0] node41865;
	wire [4-1:0] node41866;
	wire [4-1:0] node41867;
	wire [4-1:0] node41869;
	wire [4-1:0] node41871;
	wire [4-1:0] node41875;
	wire [4-1:0] node41876;
	wire [4-1:0] node41878;
	wire [4-1:0] node41882;
	wire [4-1:0] node41883;
	wire [4-1:0] node41884;
	wire [4-1:0] node41885;
	wire [4-1:0] node41886;
	wire [4-1:0] node41887;
	wire [4-1:0] node41888;
	wire [4-1:0] node41889;
	wire [4-1:0] node41892;
	wire [4-1:0] node41896;
	wire [4-1:0] node41897;
	wire [4-1:0] node41898;
	wire [4-1:0] node41901;
	wire [4-1:0] node41902;
	wire [4-1:0] node41906;
	wire [4-1:0] node41907;
	wire [4-1:0] node41911;
	wire [4-1:0] node41912;
	wire [4-1:0] node41913;
	wire [4-1:0] node41914;
	wire [4-1:0] node41917;
	wire [4-1:0] node41918;
	wire [4-1:0] node41922;
	wire [4-1:0] node41923;
	wire [4-1:0] node41926;
	wire [4-1:0] node41929;
	wire [4-1:0] node41931;
	wire [4-1:0] node41932;
	wire [4-1:0] node41935;
	wire [4-1:0] node41938;
	wire [4-1:0] node41939;
	wire [4-1:0] node41940;
	wire [4-1:0] node41941;
	wire [4-1:0] node41942;
	wire [4-1:0] node41945;
	wire [4-1:0] node41948;
	wire [4-1:0] node41949;
	wire [4-1:0] node41952;
	wire [4-1:0] node41954;
	wire [4-1:0] node41957;
	wire [4-1:0] node41958;
	wire [4-1:0] node41959;
	wire [4-1:0] node41962;
	wire [4-1:0] node41965;
	wire [4-1:0] node41968;
	wire [4-1:0] node41969;
	wire [4-1:0] node41971;
	wire [4-1:0] node41972;
	wire [4-1:0] node41975;
	wire [4-1:0] node41978;
	wire [4-1:0] node41979;
	wire [4-1:0] node41980;
	wire [4-1:0] node41984;
	wire [4-1:0] node41985;
	wire [4-1:0] node41989;
	wire [4-1:0] node41990;
	wire [4-1:0] node41991;
	wire [4-1:0] node41992;
	wire [4-1:0] node41994;
	wire [4-1:0] node41995;
	wire [4-1:0] node41997;
	wire [4-1:0] node42000;
	wire [4-1:0] node42003;
	wire [4-1:0] node42006;
	wire [4-1:0] node42007;
	wire [4-1:0] node42008;
	wire [4-1:0] node42010;
	wire [4-1:0] node42013;
	wire [4-1:0] node42015;
	wire [4-1:0] node42018;
	wire [4-1:0] node42020;
	wire [4-1:0] node42022;
	wire [4-1:0] node42023;
	wire [4-1:0] node42027;
	wire [4-1:0] node42028;
	wire [4-1:0] node42029;
	wire [4-1:0] node42031;
	wire [4-1:0] node42032;
	wire [4-1:0] node42036;
	wire [4-1:0] node42037;
	wire [4-1:0] node42040;
	wire [4-1:0] node42042;
	wire [4-1:0] node42044;
	wire [4-1:0] node42047;
	wire [4-1:0] node42048;
	wire [4-1:0] node42049;
	wire [4-1:0] node42050;
	wire [4-1:0] node42054;
	wire [4-1:0] node42057;
	wire [4-1:0] node42058;
	wire [4-1:0] node42060;
	wire [4-1:0] node42062;
	wire [4-1:0] node42065;
	wire [4-1:0] node42067;
	wire [4-1:0] node42070;
	wire [4-1:0] node42071;
	wire [4-1:0] node42072;
	wire [4-1:0] node42073;
	wire [4-1:0] node42074;
	wire [4-1:0] node42076;
	wire [4-1:0] node42079;
	wire [4-1:0] node42080;
	wire [4-1:0] node42082;
	wire [4-1:0] node42085;
	wire [4-1:0] node42086;
	wire [4-1:0] node42090;
	wire [4-1:0] node42091;
	wire [4-1:0] node42092;
	wire [4-1:0] node42095;
	wire [4-1:0] node42098;
	wire [4-1:0] node42099;
	wire [4-1:0] node42103;
	wire [4-1:0] node42104;
	wire [4-1:0] node42105;
	wire [4-1:0] node42106;
	wire [4-1:0] node42107;
	wire [4-1:0] node42110;
	wire [4-1:0] node42113;
	wire [4-1:0] node42114;
	wire [4-1:0] node42117;
	wire [4-1:0] node42120;
	wire [4-1:0] node42122;
	wire [4-1:0] node42124;
	wire [4-1:0] node42127;
	wire [4-1:0] node42128;
	wire [4-1:0] node42129;
	wire [4-1:0] node42130;
	wire [4-1:0] node42133;
	wire [4-1:0] node42136;
	wire [4-1:0] node42137;
	wire [4-1:0] node42141;
	wire [4-1:0] node42142;
	wire [4-1:0] node42143;
	wire [4-1:0] node42147;
	wire [4-1:0] node42148;
	wire [4-1:0] node42152;
	wire [4-1:0] node42153;
	wire [4-1:0] node42154;
	wire [4-1:0] node42155;
	wire [4-1:0] node42156;
	wire [4-1:0] node42157;
	wire [4-1:0] node42161;
	wire [4-1:0] node42162;
	wire [4-1:0] node42163;
	wire [4-1:0] node42166;
	wire [4-1:0] node42169;
	wire [4-1:0] node42171;
	wire [4-1:0] node42174;
	wire [4-1:0] node42175;
	wire [4-1:0] node42177;
	wire [4-1:0] node42181;
	wire [4-1:0] node42182;
	wire [4-1:0] node42183;
	wire [4-1:0] node42185;
	wire [4-1:0] node42188;
	wire [4-1:0] node42189;
	wire [4-1:0] node42191;
	wire [4-1:0] node42195;
	wire [4-1:0] node42196;
	wire [4-1:0] node42199;
	wire [4-1:0] node42200;
	wire [4-1:0] node42204;
	wire [4-1:0] node42205;
	wire [4-1:0] node42206;
	wire [4-1:0] node42207;
	wire [4-1:0] node42208;
	wire [4-1:0] node42209;
	wire [4-1:0] node42212;
	wire [4-1:0] node42215;
	wire [4-1:0] node42217;
	wire [4-1:0] node42221;
	wire [4-1:0] node42222;
	wire [4-1:0] node42223;
	wire [4-1:0] node42226;
	wire [4-1:0] node42229;
	wire [4-1:0] node42230;
	wire [4-1:0] node42234;
	wire [4-1:0] node42235;
	wire [4-1:0] node42236;
	wire [4-1:0] node42237;
	wire [4-1:0] node42238;
	wire [4-1:0] node42244;
	wire [4-1:0] node42246;
	wire [4-1:0] node42247;
	wire [4-1:0] node42251;
	wire [4-1:0] node42252;
	wire [4-1:0] node42253;
	wire [4-1:0] node42254;
	wire [4-1:0] node42255;
	wire [4-1:0] node42256;
	wire [4-1:0] node42257;
	wire [4-1:0] node42259;
	wire [4-1:0] node42260;
	wire [4-1:0] node42263;
	wire [4-1:0] node42266;
	wire [4-1:0] node42267;
	wire [4-1:0] node42268;
	wire [4-1:0] node42272;
	wire [4-1:0] node42273;
	wire [4-1:0] node42277;
	wire [4-1:0] node42278;
	wire [4-1:0] node42279;
	wire [4-1:0] node42280;
	wire [4-1:0] node42285;
	wire [4-1:0] node42287;
	wire [4-1:0] node42290;
	wire [4-1:0] node42291;
	wire [4-1:0] node42292;
	wire [4-1:0] node42293;
	wire [4-1:0] node42295;
	wire [4-1:0] node42296;
	wire [4-1:0] node42301;
	wire [4-1:0] node42304;
	wire [4-1:0] node42305;
	wire [4-1:0] node42306;
	wire [4-1:0] node42307;
	wire [4-1:0] node42310;
	wire [4-1:0] node42313;
	wire [4-1:0] node42314;
	wire [4-1:0] node42318;
	wire [4-1:0] node42319;
	wire [4-1:0] node42322;
	wire [4-1:0] node42325;
	wire [4-1:0] node42326;
	wire [4-1:0] node42327;
	wire [4-1:0] node42328;
	wire [4-1:0] node42329;
	wire [4-1:0] node42330;
	wire [4-1:0] node42333;
	wire [4-1:0] node42336;
	wire [4-1:0] node42338;
	wire [4-1:0] node42341;
	wire [4-1:0] node42342;
	wire [4-1:0] node42343;
	wire [4-1:0] node42346;
	wire [4-1:0] node42350;
	wire [4-1:0] node42351;
	wire [4-1:0] node42352;
	wire [4-1:0] node42354;
	wire [4-1:0] node42357;
	wire [4-1:0] node42359;
	wire [4-1:0] node42362;
	wire [4-1:0] node42363;
	wire [4-1:0] node42366;
	wire [4-1:0] node42369;
	wire [4-1:0] node42370;
	wire [4-1:0] node42371;
	wire [4-1:0] node42372;
	wire [4-1:0] node42376;
	wire [4-1:0] node42377;
	wire [4-1:0] node42380;
	wire [4-1:0] node42381;
	wire [4-1:0] node42385;
	wire [4-1:0] node42386;
	wire [4-1:0] node42387;
	wire [4-1:0] node42390;
	wire [4-1:0] node42391;
	wire [4-1:0] node42393;
	wire [4-1:0] node42397;
	wire [4-1:0] node42398;
	wire [4-1:0] node42400;
	wire [4-1:0] node42403;
	wire [4-1:0] node42405;
	wire [4-1:0] node42408;
	wire [4-1:0] node42409;
	wire [4-1:0] node42410;
	wire [4-1:0] node42411;
	wire [4-1:0] node42412;
	wire [4-1:0] node42413;
	wire [4-1:0] node42415;
	wire [4-1:0] node42418;
	wire [4-1:0] node42420;
	wire [4-1:0] node42422;
	wire [4-1:0] node42425;
	wire [4-1:0] node42426;
	wire [4-1:0] node42428;
	wire [4-1:0] node42429;
	wire [4-1:0] node42432;
	wire [4-1:0] node42435;
	wire [4-1:0] node42437;
	wire [4-1:0] node42440;
	wire [4-1:0] node42441;
	wire [4-1:0] node42443;
	wire [4-1:0] node42444;
	wire [4-1:0] node42445;
	wire [4-1:0] node42449;
	wire [4-1:0] node42450;
	wire [4-1:0] node42454;
	wire [4-1:0] node42457;
	wire [4-1:0] node42458;
	wire [4-1:0] node42459;
	wire [4-1:0] node42460;
	wire [4-1:0] node42461;
	wire [4-1:0] node42465;
	wire [4-1:0] node42466;
	wire [4-1:0] node42469;
	wire [4-1:0] node42472;
	wire [4-1:0] node42473;
	wire [4-1:0] node42474;
	wire [4-1:0] node42478;
	wire [4-1:0] node42481;
	wire [4-1:0] node42482;
	wire [4-1:0] node42483;
	wire [4-1:0] node42485;
	wire [4-1:0] node42488;
	wire [4-1:0] node42490;
	wire [4-1:0] node42491;
	wire [4-1:0] node42495;
	wire [4-1:0] node42498;
	wire [4-1:0] node42499;
	wire [4-1:0] node42500;
	wire [4-1:0] node42501;
	wire [4-1:0] node42502;
	wire [4-1:0] node42503;
	wire [4-1:0] node42506;
	wire [4-1:0] node42510;
	wire [4-1:0] node42512;
	wire [4-1:0] node42515;
	wire [4-1:0] node42516;
	wire [4-1:0] node42517;
	wire [4-1:0] node42521;
	wire [4-1:0] node42523;
	wire [4-1:0] node42525;
	wire [4-1:0] node42528;
	wire [4-1:0] node42529;
	wire [4-1:0] node42530;
	wire [4-1:0] node42531;
	wire [4-1:0] node42532;
	wire [4-1:0] node42533;
	wire [4-1:0] node42538;
	wire [4-1:0] node42540;
	wire [4-1:0] node42543;
	wire [4-1:0] node42544;
	wire [4-1:0] node42548;
	wire [4-1:0] node42549;
	wire [4-1:0] node42550;
	wire [4-1:0] node42551;
	wire [4-1:0] node42555;
	wire [4-1:0] node42556;
	wire [4-1:0] node42560;
	wire [4-1:0] node42561;
	wire [4-1:0] node42563;
	wire [4-1:0] node42566;
	wire [4-1:0] node42567;
	wire [4-1:0] node42568;
	wire [4-1:0] node42573;
	wire [4-1:0] node42574;
	wire [4-1:0] node42575;
	wire [4-1:0] node42576;
	wire [4-1:0] node42577;
	wire [4-1:0] node42578;
	wire [4-1:0] node42580;
	wire [4-1:0] node42581;
	wire [4-1:0] node42584;
	wire [4-1:0] node42587;
	wire [4-1:0] node42588;
	wire [4-1:0] node42589;
	wire [4-1:0] node42592;
	wire [4-1:0] node42596;
	wire [4-1:0] node42597;
	wire [4-1:0] node42598;
	wire [4-1:0] node42600;
	wire [4-1:0] node42603;
	wire [4-1:0] node42606;
	wire [4-1:0] node42607;
	wire [4-1:0] node42609;
	wire [4-1:0] node42612;
	wire [4-1:0] node42613;
	wire [4-1:0] node42617;
	wire [4-1:0] node42618;
	wire [4-1:0] node42619;
	wire [4-1:0] node42620;
	wire [4-1:0] node42621;
	wire [4-1:0] node42625;
	wire [4-1:0] node42626;
	wire [4-1:0] node42629;
	wire [4-1:0] node42632;
	wire [4-1:0] node42633;
	wire [4-1:0] node42636;
	wire [4-1:0] node42637;
	wire [4-1:0] node42640;
	wire [4-1:0] node42642;
	wire [4-1:0] node42645;
	wire [4-1:0] node42646;
	wire [4-1:0] node42647;
	wire [4-1:0] node42651;
	wire [4-1:0] node42652;
	wire [4-1:0] node42653;
	wire [4-1:0] node42654;
	wire [4-1:0] node42657;
	wire [4-1:0] node42661;
	wire [4-1:0] node42662;
	wire [4-1:0] node42666;
	wire [4-1:0] node42667;
	wire [4-1:0] node42668;
	wire [4-1:0] node42669;
	wire [4-1:0] node42670;
	wire [4-1:0] node42671;
	wire [4-1:0] node42676;
	wire [4-1:0] node42677;
	wire [4-1:0] node42680;
	wire [4-1:0] node42683;
	wire [4-1:0] node42684;
	wire [4-1:0] node42685;
	wire [4-1:0] node42686;
	wire [4-1:0] node42690;
	wire [4-1:0] node42693;
	wire [4-1:0] node42694;
	wire [4-1:0] node42695;
	wire [4-1:0] node42697;
	wire [4-1:0] node42700;
	wire [4-1:0] node42701;
	wire [4-1:0] node42705;
	wire [4-1:0] node42706;
	wire [4-1:0] node42709;
	wire [4-1:0] node42712;
	wire [4-1:0] node42713;
	wire [4-1:0] node42714;
	wire [4-1:0] node42715;
	wire [4-1:0] node42716;
	wire [4-1:0] node42720;
	wire [4-1:0] node42721;
	wire [4-1:0] node42725;
	wire [4-1:0] node42726;
	wire [4-1:0] node42727;
	wire [4-1:0] node42731;
	wire [4-1:0] node42733;
	wire [4-1:0] node42736;
	wire [4-1:0] node42737;
	wire [4-1:0] node42738;
	wire [4-1:0] node42741;
	wire [4-1:0] node42743;
	wire [4-1:0] node42746;
	wire [4-1:0] node42747;
	wire [4-1:0] node42748;
	wire [4-1:0] node42750;
	wire [4-1:0] node42753;
	wire [4-1:0] node42756;
	wire [4-1:0] node42758;
	wire [4-1:0] node42761;
	wire [4-1:0] node42762;
	wire [4-1:0] node42763;
	wire [4-1:0] node42764;
	wire [4-1:0] node42765;
	wire [4-1:0] node42766;
	wire [4-1:0] node42767;
	wire [4-1:0] node42770;
	wire [4-1:0] node42773;
	wire [4-1:0] node42775;
	wire [4-1:0] node42778;
	wire [4-1:0] node42779;
	wire [4-1:0] node42780;
	wire [4-1:0] node42783;
	wire [4-1:0] node42784;
	wire [4-1:0] node42787;
	wire [4-1:0] node42790;
	wire [4-1:0] node42791;
	wire [4-1:0] node42792;
	wire [4-1:0] node42796;
	wire [4-1:0] node42799;
	wire [4-1:0] node42800;
	wire [4-1:0] node42801;
	wire [4-1:0] node42804;
	wire [4-1:0] node42807;
	wire [4-1:0] node42808;
	wire [4-1:0] node42809;
	wire [4-1:0] node42813;
	wire [4-1:0] node42815;
	wire [4-1:0] node42818;
	wire [4-1:0] node42819;
	wire [4-1:0] node42820;
	wire [4-1:0] node42821;
	wire [4-1:0] node42822;
	wire [4-1:0] node42824;
	wire [4-1:0] node42828;
	wire [4-1:0] node42829;
	wire [4-1:0] node42832;
	wire [4-1:0] node42835;
	wire [4-1:0] node42836;
	wire [4-1:0] node42838;
	wire [4-1:0] node42839;
	wire [4-1:0] node42843;
	wire [4-1:0] node42844;
	wire [4-1:0] node42848;
	wire [4-1:0] node42849;
	wire [4-1:0] node42850;
	wire [4-1:0] node42851;
	wire [4-1:0] node42855;
	wire [4-1:0] node42856;
	wire [4-1:0] node42858;
	wire [4-1:0] node42862;
	wire [4-1:0] node42863;
	wire [4-1:0] node42867;
	wire [4-1:0] node42868;
	wire [4-1:0] node42869;
	wire [4-1:0] node42870;
	wire [4-1:0] node42871;
	wire [4-1:0] node42875;
	wire [4-1:0] node42876;
	wire [4-1:0] node42878;
	wire [4-1:0] node42881;
	wire [4-1:0] node42882;
	wire [4-1:0] node42885;
	wire [4-1:0] node42888;
	wire [4-1:0] node42889;
	wire [4-1:0] node42890;
	wire [4-1:0] node42892;
	wire [4-1:0] node42895;
	wire [4-1:0] node42896;
	wire [4-1:0] node42900;
	wire [4-1:0] node42901;
	wire [4-1:0] node42902;
	wire [4-1:0] node42903;
	wire [4-1:0] node42908;
	wire [4-1:0] node42909;
	wire [4-1:0] node42912;
	wire [4-1:0] node42915;
	wire [4-1:0] node42916;
	wire [4-1:0] node42917;
	wire [4-1:0] node42918;
	wire [4-1:0] node42921;
	wire [4-1:0] node42922;
	wire [4-1:0] node42924;
	wire [4-1:0] node42927;
	wire [4-1:0] node42929;
	wire [4-1:0] node42932;
	wire [4-1:0] node42933;
	wire [4-1:0] node42934;
	wire [4-1:0] node42937;
	wire [4-1:0] node42940;
	wire [4-1:0] node42942;
	wire [4-1:0] node42945;
	wire [4-1:0] node42946;
	wire [4-1:0] node42947;
	wire [4-1:0] node42950;
	wire [4-1:0] node42951;
	wire [4-1:0] node42954;
	wire [4-1:0] node42957;
	wire [4-1:0] node42958;
	wire [4-1:0] node42959;
	wire [4-1:0] node42961;
	wire [4-1:0] node42965;
	wire [4-1:0] node42966;
	wire [4-1:0] node42968;
	wire [4-1:0] node42972;
	wire [4-1:0] node42973;
	wire [4-1:0] node42974;
	wire [4-1:0] node42975;
	wire [4-1:0] node42976;
	wire [4-1:0] node42977;
	wire [4-1:0] node42978;
	wire [4-1:0] node42979;
	wire [4-1:0] node42980;
	wire [4-1:0] node42981;
	wire [4-1:0] node42985;
	wire [4-1:0] node42988;
	wire [4-1:0] node42989;
	wire [4-1:0] node42990;
	wire [4-1:0] node42991;
	wire [4-1:0] node42994;
	wire [4-1:0] node42997;
	wire [4-1:0] node42999;
	wire [4-1:0] node43002;
	wire [4-1:0] node43003;
	wire [4-1:0] node43005;
	wire [4-1:0] node43009;
	wire [4-1:0] node43010;
	wire [4-1:0] node43013;
	wire [4-1:0] node43014;
	wire [4-1:0] node43015;
	wire [4-1:0] node43017;
	wire [4-1:0] node43020;
	wire [4-1:0] node43021;
	wire [4-1:0] node43025;
	wire [4-1:0] node43026;
	wire [4-1:0] node43030;
	wire [4-1:0] node43031;
	wire [4-1:0] node43032;
	wire [4-1:0] node43033;
	wire [4-1:0] node43034;
	wire [4-1:0] node43037;
	wire [4-1:0] node43040;
	wire [4-1:0] node43041;
	wire [4-1:0] node43045;
	wire [4-1:0] node43046;
	wire [4-1:0] node43050;
	wire [4-1:0] node43051;
	wire [4-1:0] node43054;
	wire [4-1:0] node43055;
	wire [4-1:0] node43057;
	wire [4-1:0] node43060;
	wire [4-1:0] node43061;
	wire [4-1:0] node43064;
	wire [4-1:0] node43067;
	wire [4-1:0] node43068;
	wire [4-1:0] node43069;
	wire [4-1:0] node43070;
	wire [4-1:0] node43071;
	wire [4-1:0] node43072;
	wire [4-1:0] node43074;
	wire [4-1:0] node43078;
	wire [4-1:0] node43079;
	wire [4-1:0] node43083;
	wire [4-1:0] node43084;
	wire [4-1:0] node43085;
	wire [4-1:0] node43088;
	wire [4-1:0] node43091;
	wire [4-1:0] node43093;
	wire [4-1:0] node43096;
	wire [4-1:0] node43097;
	wire [4-1:0] node43099;
	wire [4-1:0] node43101;
	wire [4-1:0] node43102;
	wire [4-1:0] node43105;
	wire [4-1:0] node43108;
	wire [4-1:0] node43109;
	wire [4-1:0] node43113;
	wire [4-1:0] node43114;
	wire [4-1:0] node43115;
	wire [4-1:0] node43116;
	wire [4-1:0] node43117;
	wire [4-1:0] node43118;
	wire [4-1:0] node43121;
	wire [4-1:0] node43125;
	wire [4-1:0] node43127;
	wire [4-1:0] node43130;
	wire [4-1:0] node43131;
	wire [4-1:0] node43132;
	wire [4-1:0] node43135;
	wire [4-1:0] node43139;
	wire [4-1:0] node43140;
	wire [4-1:0] node43141;
	wire [4-1:0] node43142;
	wire [4-1:0] node43143;
	wire [4-1:0] node43146;
	wire [4-1:0] node43151;
	wire [4-1:0] node43153;
	wire [4-1:0] node43156;
	wire [4-1:0] node43157;
	wire [4-1:0] node43158;
	wire [4-1:0] node43159;
	wire [4-1:0] node43160;
	wire [4-1:0] node43161;
	wire [4-1:0] node43162;
	wire [4-1:0] node43165;
	wire [4-1:0] node43168;
	wire [4-1:0] node43169;
	wire [4-1:0] node43171;
	wire [4-1:0] node43175;
	wire [4-1:0] node43176;
	wire [4-1:0] node43177;
	wire [4-1:0] node43179;
	wire [4-1:0] node43182;
	wire [4-1:0] node43183;
	wire [4-1:0] node43187;
	wire [4-1:0] node43188;
	wire [4-1:0] node43191;
	wire [4-1:0] node43194;
	wire [4-1:0] node43195;
	wire [4-1:0] node43196;
	wire [4-1:0] node43198;
	wire [4-1:0] node43199;
	wire [4-1:0] node43203;
	wire [4-1:0] node43205;
	wire [4-1:0] node43208;
	wire [4-1:0] node43209;
	wire [4-1:0] node43210;
	wire [4-1:0] node43212;
	wire [4-1:0] node43215;
	wire [4-1:0] node43216;
	wire [4-1:0] node43220;
	wire [4-1:0] node43221;
	wire [4-1:0] node43223;
	wire [4-1:0] node43227;
	wire [4-1:0] node43228;
	wire [4-1:0] node43229;
	wire [4-1:0] node43230;
	wire [4-1:0] node43231;
	wire [4-1:0] node43235;
	wire [4-1:0] node43237;
	wire [4-1:0] node43240;
	wire [4-1:0] node43241;
	wire [4-1:0] node43245;
	wire [4-1:0] node43246;
	wire [4-1:0] node43247;
	wire [4-1:0] node43248;
	wire [4-1:0] node43250;
	wire [4-1:0] node43254;
	wire [4-1:0] node43256;
	wire [4-1:0] node43259;
	wire [4-1:0] node43260;
	wire [4-1:0] node43262;
	wire [4-1:0] node43265;
	wire [4-1:0] node43266;
	wire [4-1:0] node43268;
	wire [4-1:0] node43272;
	wire [4-1:0] node43273;
	wire [4-1:0] node43274;
	wire [4-1:0] node43275;
	wire [4-1:0] node43277;
	wire [4-1:0] node43280;
	wire [4-1:0] node43281;
	wire [4-1:0] node43284;
	wire [4-1:0] node43287;
	wire [4-1:0] node43288;
	wire [4-1:0] node43291;
	wire [4-1:0] node43294;
	wire [4-1:0] node43295;
	wire [4-1:0] node43296;
	wire [4-1:0] node43297;
	wire [4-1:0] node43298;
	wire [4-1:0] node43299;
	wire [4-1:0] node43302;
	wire [4-1:0] node43305;
	wire [4-1:0] node43307;
	wire [4-1:0] node43310;
	wire [4-1:0] node43312;
	wire [4-1:0] node43315;
	wire [4-1:0] node43317;
	wire [4-1:0] node43319;
	wire [4-1:0] node43322;
	wire [4-1:0] node43323;
	wire [4-1:0] node43324;
	wire [4-1:0] node43327;
	wire [4-1:0] node43330;
	wire [4-1:0] node43331;
	wire [4-1:0] node43333;
	wire [4-1:0] node43336;
	wire [4-1:0] node43337;
	wire [4-1:0] node43340;
	wire [4-1:0] node43343;
	wire [4-1:0] node43344;
	wire [4-1:0] node43345;
	wire [4-1:0] node43346;
	wire [4-1:0] node43347;
	wire [4-1:0] node43348;
	wire [4-1:0] node43349;
	wire [4-1:0] node43350;
	wire [4-1:0] node43353;
	wire [4-1:0] node43354;
	wire [4-1:0] node43359;
	wire [4-1:0] node43360;
	wire [4-1:0] node43362;
	wire [4-1:0] node43365;
	wire [4-1:0] node43367;
	wire [4-1:0] node43370;
	wire [4-1:0] node43371;
	wire [4-1:0] node43372;
	wire [4-1:0] node43373;
	wire [4-1:0] node43374;
	wire [4-1:0] node43380;
	wire [4-1:0] node43381;
	wire [4-1:0] node43383;
	wire [4-1:0] node43386;
	wire [4-1:0] node43387;
	wire [4-1:0] node43390;
	wire [4-1:0] node43393;
	wire [4-1:0] node43394;
	wire [4-1:0] node43395;
	wire [4-1:0] node43396;
	wire [4-1:0] node43398;
	wire [4-1:0] node43399;
	wire [4-1:0] node43402;
	wire [4-1:0] node43405;
	wire [4-1:0] node43407;
	wire [4-1:0] node43410;
	wire [4-1:0] node43413;
	wire [4-1:0] node43414;
	wire [4-1:0] node43415;
	wire [4-1:0] node43416;
	wire [4-1:0] node43418;
	wire [4-1:0] node43421;
	wire [4-1:0] node43424;
	wire [4-1:0] node43425;
	wire [4-1:0] node43428;
	wire [4-1:0] node43431;
	wire [4-1:0] node43433;
	wire [4-1:0] node43434;
	wire [4-1:0] node43438;
	wire [4-1:0] node43439;
	wire [4-1:0] node43440;
	wire [4-1:0] node43441;
	wire [4-1:0] node43442;
	wire [4-1:0] node43443;
	wire [4-1:0] node43447;
	wire [4-1:0] node43450;
	wire [4-1:0] node43451;
	wire [4-1:0] node43452;
	wire [4-1:0] node43453;
	wire [4-1:0] node43458;
	wire [4-1:0] node43459;
	wire [4-1:0] node43463;
	wire [4-1:0] node43464;
	wire [4-1:0] node43465;
	wire [4-1:0] node43468;
	wire [4-1:0] node43471;
	wire [4-1:0] node43472;
	wire [4-1:0] node43474;
	wire [4-1:0] node43477;
	wire [4-1:0] node43478;
	wire [4-1:0] node43481;
	wire [4-1:0] node43484;
	wire [4-1:0] node43485;
	wire [4-1:0] node43486;
	wire [4-1:0] node43489;
	wire [4-1:0] node43492;
	wire [4-1:0] node43493;
	wire [4-1:0] node43494;
	wire [4-1:0] node43498;
	wire [4-1:0] node43499;
	wire [4-1:0] node43501;
	wire [4-1:0] node43504;
	wire [4-1:0] node43505;
	wire [4-1:0] node43508;
	wire [4-1:0] node43511;
	wire [4-1:0] node43512;
	wire [4-1:0] node43513;
	wire [4-1:0] node43514;
	wire [4-1:0] node43515;
	wire [4-1:0] node43516;
	wire [4-1:0] node43519;
	wire [4-1:0] node43522;
	wire [4-1:0] node43523;
	wire [4-1:0] node43524;
	wire [4-1:0] node43527;
	wire [4-1:0] node43529;
	wire [4-1:0] node43532;
	wire [4-1:0] node43533;
	wire [4-1:0] node43536;
	wire [4-1:0] node43539;
	wire [4-1:0] node43540;
	wire [4-1:0] node43541;
	wire [4-1:0] node43544;
	wire [4-1:0] node43545;
	wire [4-1:0] node43546;
	wire [4-1:0] node43551;
	wire [4-1:0] node43552;
	wire [4-1:0] node43555;
	wire [4-1:0] node43558;
	wire [4-1:0] node43559;
	wire [4-1:0] node43560;
	wire [4-1:0] node43561;
	wire [4-1:0] node43562;
	wire [4-1:0] node43567;
	wire [4-1:0] node43568;
	wire [4-1:0] node43569;
	wire [4-1:0] node43572;
	wire [4-1:0] node43575;
	wire [4-1:0] node43576;
	wire [4-1:0] node43577;
	wire [4-1:0] node43582;
	wire [4-1:0] node43583;
	wire [4-1:0] node43585;
	wire [4-1:0] node43586;
	wire [4-1:0] node43587;
	wire [4-1:0] node43591;
	wire [4-1:0] node43592;
	wire [4-1:0] node43596;
	wire [4-1:0] node43597;
	wire [4-1:0] node43598;
	wire [4-1:0] node43601;
	wire [4-1:0] node43605;
	wire [4-1:0] node43606;
	wire [4-1:0] node43607;
	wire [4-1:0] node43608;
	wire [4-1:0] node43610;
	wire [4-1:0] node43611;
	wire [4-1:0] node43612;
	wire [4-1:0] node43617;
	wire [4-1:0] node43619;
	wire [4-1:0] node43622;
	wire [4-1:0] node43623;
	wire [4-1:0] node43625;
	wire [4-1:0] node43628;
	wire [4-1:0] node43629;
	wire [4-1:0] node43633;
	wire [4-1:0] node43634;
	wire [4-1:0] node43635;
	wire [4-1:0] node43638;
	wire [4-1:0] node43641;
	wire [4-1:0] node43642;
	wire [4-1:0] node43643;
	wire [4-1:0] node43646;
	wire [4-1:0] node43649;
	wire [4-1:0] node43651;
	wire [4-1:0] node43652;
	wire [4-1:0] node43656;
	wire [4-1:0] node43657;
	wire [4-1:0] node43658;
	wire [4-1:0] node43659;
	wire [4-1:0] node43660;
	wire [4-1:0] node43661;
	wire [4-1:0] node43662;
	wire [4-1:0] node43663;
	wire [4-1:0] node43665;
	wire [4-1:0] node43668;
	wire [4-1:0] node43669;
	wire [4-1:0] node43672;
	wire [4-1:0] node43675;
	wire [4-1:0] node43676;
	wire [4-1:0] node43678;
	wire [4-1:0] node43681;
	wire [4-1:0] node43683;
	wire [4-1:0] node43686;
	wire [4-1:0] node43687;
	wire [4-1:0] node43688;
	wire [4-1:0] node43691;
	wire [4-1:0] node43693;
	wire [4-1:0] node43696;
	wire [4-1:0] node43698;
	wire [4-1:0] node43699;
	wire [4-1:0] node43702;
	wire [4-1:0] node43705;
	wire [4-1:0] node43706;
	wire [4-1:0] node43707;
	wire [4-1:0] node43708;
	wire [4-1:0] node43711;
	wire [4-1:0] node43714;
	wire [4-1:0] node43716;
	wire [4-1:0] node43717;
	wire [4-1:0] node43720;
	wire [4-1:0] node43723;
	wire [4-1:0] node43724;
	wire [4-1:0] node43726;
	wire [4-1:0] node43727;
	wire [4-1:0] node43730;
	wire [4-1:0] node43733;
	wire [4-1:0] node43734;
	wire [4-1:0] node43736;
	wire [4-1:0] node43739;
	wire [4-1:0] node43740;
	wire [4-1:0] node43741;
	wire [4-1:0] node43744;
	wire [4-1:0] node43747;
	wire [4-1:0] node43748;
	wire [4-1:0] node43752;
	wire [4-1:0] node43753;
	wire [4-1:0] node43754;
	wire [4-1:0] node43755;
	wire [4-1:0] node43756;
	wire [4-1:0] node43759;
	wire [4-1:0] node43760;
	wire [4-1:0] node43762;
	wire [4-1:0] node43766;
	wire [4-1:0] node43767;
	wire [4-1:0] node43768;
	wire [4-1:0] node43770;
	wire [4-1:0] node43773;
	wire [4-1:0] node43776;
	wire [4-1:0] node43778;
	wire [4-1:0] node43781;
	wire [4-1:0] node43783;
	wire [4-1:0] node43784;
	wire [4-1:0] node43786;
	wire [4-1:0] node43788;
	wire [4-1:0] node43791;
	wire [4-1:0] node43793;
	wire [4-1:0] node43796;
	wire [4-1:0] node43797;
	wire [4-1:0] node43798;
	wire [4-1:0] node43800;
	wire [4-1:0] node43802;
	wire [4-1:0] node43805;
	wire [4-1:0] node43806;
	wire [4-1:0] node43808;
	wire [4-1:0] node43809;
	wire [4-1:0] node43813;
	wire [4-1:0] node43816;
	wire [4-1:0] node43817;
	wire [4-1:0] node43818;
	wire [4-1:0] node43820;
	wire [4-1:0] node43822;
	wire [4-1:0] node43825;
	wire [4-1:0] node43828;
	wire [4-1:0] node43829;
	wire [4-1:0] node43830;
	wire [4-1:0] node43834;
	wire [4-1:0] node43836;
	wire [4-1:0] node43839;
	wire [4-1:0] node43840;
	wire [4-1:0] node43841;
	wire [4-1:0] node43842;
	wire [4-1:0] node43843;
	wire [4-1:0] node43844;
	wire [4-1:0] node43847;
	wire [4-1:0] node43850;
	wire [4-1:0] node43852;
	wire [4-1:0] node43853;
	wire [4-1:0] node43855;
	wire [4-1:0] node43858;
	wire [4-1:0] node43861;
	wire [4-1:0] node43862;
	wire [4-1:0] node43863;
	wire [4-1:0] node43865;
	wire [4-1:0] node43868;
	wire [4-1:0] node43869;
	wire [4-1:0] node43871;
	wire [4-1:0] node43874;
	wire [4-1:0] node43877;
	wire [4-1:0] node43878;
	wire [4-1:0] node43881;
	wire [4-1:0] node43882;
	wire [4-1:0] node43885;
	wire [4-1:0] node43888;
	wire [4-1:0] node43889;
	wire [4-1:0] node43890;
	wire [4-1:0] node43891;
	wire [4-1:0] node43894;
	wire [4-1:0] node43897;
	wire [4-1:0] node43898;
	wire [4-1:0] node43900;
	wire [4-1:0] node43903;
	wire [4-1:0] node43905;
	wire [4-1:0] node43908;
	wire [4-1:0] node43909;
	wire [4-1:0] node43910;
	wire [4-1:0] node43911;
	wire [4-1:0] node43914;
	wire [4-1:0] node43918;
	wire [4-1:0] node43919;
	wire [4-1:0] node43920;
	wire [4-1:0] node43923;
	wire [4-1:0] node43926;
	wire [4-1:0] node43928;
	wire [4-1:0] node43929;
	wire [4-1:0] node43932;
	wire [4-1:0] node43935;
	wire [4-1:0] node43936;
	wire [4-1:0] node43937;
	wire [4-1:0] node43938;
	wire [4-1:0] node43939;
	wire [4-1:0] node43940;
	wire [4-1:0] node43943;
	wire [4-1:0] node43946;
	wire [4-1:0] node43947;
	wire [4-1:0] node43950;
	wire [4-1:0] node43953;
	wire [4-1:0] node43954;
	wire [4-1:0] node43956;
	wire [4-1:0] node43958;
	wire [4-1:0] node43961;
	wire [4-1:0] node43963;
	wire [4-1:0] node43966;
	wire [4-1:0] node43967;
	wire [4-1:0] node43969;
	wire [4-1:0] node43971;
	wire [4-1:0] node43974;
	wire [4-1:0] node43975;
	wire [4-1:0] node43977;
	wire [4-1:0] node43980;
	wire [4-1:0] node43982;
	wire [4-1:0] node43985;
	wire [4-1:0] node43986;
	wire [4-1:0] node43987;
	wire [4-1:0] node43990;
	wire [4-1:0] node43993;
	wire [4-1:0] node43994;
	wire [4-1:0] node43995;
	wire [4-1:0] node43996;
	wire [4-1:0] node44000;
	wire [4-1:0] node44002;
	wire [4-1:0] node44005;
	wire [4-1:0] node44006;
	wire [4-1:0] node44007;
	wire [4-1:0] node44008;
	wire [4-1:0] node44013;
	wire [4-1:0] node44015;
	wire [4-1:0] node44018;
	wire [4-1:0] node44019;
	wire [4-1:0] node44020;
	wire [4-1:0] node44021;
	wire [4-1:0] node44022;
	wire [4-1:0] node44023;
	wire [4-1:0] node44024;
	wire [4-1:0] node44025;
	wire [4-1:0] node44028;
	wire [4-1:0] node44031;
	wire [4-1:0] node44032;
	wire [4-1:0] node44035;
	wire [4-1:0] node44038;
	wire [4-1:0] node44039;
	wire [4-1:0] node44040;
	wire [4-1:0] node44044;
	wire [4-1:0] node44046;
	wire [4-1:0] node44049;
	wire [4-1:0] node44050;
	wire [4-1:0] node44051;
	wire [4-1:0] node44052;
	wire [4-1:0] node44055;
	wire [4-1:0] node44058;
	wire [4-1:0] node44059;
	wire [4-1:0] node44062;
	wire [4-1:0] node44065;
	wire [4-1:0] node44066;
	wire [4-1:0] node44067;
	wire [4-1:0] node44070;
	wire [4-1:0] node44071;
	wire [4-1:0] node44074;
	wire [4-1:0] node44078;
	wire [4-1:0] node44079;
	wire [4-1:0] node44080;
	wire [4-1:0] node44081;
	wire [4-1:0] node44083;
	wire [4-1:0] node44086;
	wire [4-1:0] node44089;
	wire [4-1:0] node44090;
	wire [4-1:0] node44094;
	wire [4-1:0] node44095;
	wire [4-1:0] node44096;
	wire [4-1:0] node44099;
	wire [4-1:0] node44102;
	wire [4-1:0] node44105;
	wire [4-1:0] node44106;
	wire [4-1:0] node44107;
	wire [4-1:0] node44108;
	wire [4-1:0] node44109;
	wire [4-1:0] node44113;
	wire [4-1:0] node44114;
	wire [4-1:0] node44118;
	wire [4-1:0] node44119;
	wire [4-1:0] node44120;
	wire [4-1:0] node44123;
	wire [4-1:0] node44126;
	wire [4-1:0] node44127;
	wire [4-1:0] node44128;
	wire [4-1:0] node44131;
	wire [4-1:0] node44135;
	wire [4-1:0] node44136;
	wire [4-1:0] node44137;
	wire [4-1:0] node44138;
	wire [4-1:0] node44141;
	wire [4-1:0] node44144;
	wire [4-1:0] node44146;
	wire [4-1:0] node44149;
	wire [4-1:0] node44150;
	wire [4-1:0] node44151;
	wire [4-1:0] node44154;
	wire [4-1:0] node44157;
	wire [4-1:0] node44158;
	wire [4-1:0] node44160;
	wire [4-1:0] node44164;
	wire [4-1:0] node44165;
	wire [4-1:0] node44166;
	wire [4-1:0] node44167;
	wire [4-1:0] node44168;
	wire [4-1:0] node44170;
	wire [4-1:0] node44173;
	wire [4-1:0] node44174;
	wire [4-1:0] node44175;
	wire [4-1:0] node44178;
	wire [4-1:0] node44181;
	wire [4-1:0] node44182;
	wire [4-1:0] node44185;
	wire [4-1:0] node44188;
	wire [4-1:0] node44189;
	wire [4-1:0] node44190;
	wire [4-1:0] node44191;
	wire [4-1:0] node44195;
	wire [4-1:0] node44197;
	wire [4-1:0] node44198;
	wire [4-1:0] node44202;
	wire [4-1:0] node44203;
	wire [4-1:0] node44204;
	wire [4-1:0] node44206;
	wire [4-1:0] node44209;
	wire [4-1:0] node44210;
	wire [4-1:0] node44213;
	wire [4-1:0] node44216;
	wire [4-1:0] node44217;
	wire [4-1:0] node44220;
	wire [4-1:0] node44223;
	wire [4-1:0] node44224;
	wire [4-1:0] node44225;
	wire [4-1:0] node44226;
	wire [4-1:0] node44229;
	wire [4-1:0] node44232;
	wire [4-1:0] node44235;
	wire [4-1:0] node44236;
	wire [4-1:0] node44237;
	wire [4-1:0] node44239;
	wire [4-1:0] node44242;
	wire [4-1:0] node44243;
	wire [4-1:0] node44244;
	wire [4-1:0] node44249;
	wire [4-1:0] node44250;
	wire [4-1:0] node44252;
	wire [4-1:0] node44254;
	wire [4-1:0] node44257;
	wire [4-1:0] node44258;
	wire [4-1:0] node44262;
	wire [4-1:0] node44263;
	wire [4-1:0] node44264;
	wire [4-1:0] node44265;
	wire [4-1:0] node44266;
	wire [4-1:0] node44268;
	wire [4-1:0] node44270;
	wire [4-1:0] node44273;
	wire [4-1:0] node44276;
	wire [4-1:0] node44277;
	wire [4-1:0] node44279;
	wire [4-1:0] node44282;
	wire [4-1:0] node44285;
	wire [4-1:0] node44286;
	wire [4-1:0] node44287;
	wire [4-1:0] node44289;
	wire [4-1:0] node44292;
	wire [4-1:0] node44293;
	wire [4-1:0] node44296;
	wire [4-1:0] node44299;
	wire [4-1:0] node44300;
	wire [4-1:0] node44304;
	wire [4-1:0] node44305;
	wire [4-1:0] node44306;
	wire [4-1:0] node44307;
	wire [4-1:0] node44308;
	wire [4-1:0] node44311;
	wire [4-1:0] node44314;
	wire [4-1:0] node44316;
	wire [4-1:0] node44319;
	wire [4-1:0] node44320;
	wire [4-1:0] node44323;
	wire [4-1:0] node44326;
	wire [4-1:0] node44327;
	wire [4-1:0] node44328;
	wire [4-1:0] node44331;
	wire [4-1:0] node44334;
	wire [4-1:0] node44335;
	wire [4-1:0] node44338;

	assign outp = (inp[14]) ? node24864 : node1;
		assign node1 = (inp[11]) ? node12493 : node2;
			assign node2 = (inp[5]) ? node6078 : node3;
				assign node3 = (inp[7]) ? node2999 : node4;
					assign node4 = (inp[6]) ? node1542 : node5;
						assign node5 = (inp[1]) ? node779 : node6;
							assign node6 = (inp[13]) ? node386 : node7;
								assign node7 = (inp[9]) ? node155 : node8;
									assign node8 = (inp[4]) ? node92 : node9;
										assign node9 = (inp[12]) ? node47 : node10;
											assign node10 = (inp[8]) ? node28 : node11;
												assign node11 = (inp[2]) ? node21 : node12;
													assign node12 = (inp[10]) ? node14 : 4'b1101;
														assign node14 = (inp[0]) ? node18 : node15;
															assign node15 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node18 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node21 = (inp[15]) ? node25 : node22;
														assign node22 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node25 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node28 = (inp[2]) ? node40 : node29;
													assign node29 = (inp[3]) ? node35 : node30;
														assign node30 = (inp[0]) ? node32 : 4'b1100;
															assign node32 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node35 = (inp[15]) ? node37 : 4'b1110;
															assign node37 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node40 = (inp[0]) ? node44 : node41;
														assign node41 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node44 = (inp[15]) ? 4'b1111 : 4'b1101;
											assign node47 = (inp[10]) ? node73 : node48;
												assign node48 = (inp[15]) ? node60 : node49;
													assign node49 = (inp[0]) ? node55 : node50;
														assign node50 = (inp[2]) ? 4'b1110 : node51;
															assign node51 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node55 = (inp[2]) ? node57 : 4'b1100;
															assign node57 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node60 = (inp[0]) ? 4'b1110 : node61;
														assign node61 = (inp[3]) ? node67 : node62;
															assign node62 = (inp[8]) ? node64 : 4'b1101;
																assign node64 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node67 = (inp[2]) ? node69 : 4'b1100;
																assign node69 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node73 = (inp[0]) ? node85 : node74;
													assign node74 = (inp[15]) ? node78 : node75;
														assign node75 = (inp[3]) ? 4'b1011 : 4'b1010;
														assign node78 = (inp[8]) ? node82 : node79;
															assign node79 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node82 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node85 = (inp[15]) ? node89 : node86;
														assign node86 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node89 = (inp[2]) ? 4'b1010 : 4'b1011;
										assign node92 = (inp[12]) ? node124 : node93;
											assign node93 = (inp[15]) ? node109 : node94;
												assign node94 = (inp[0]) ? node102 : node95;
													assign node95 = (inp[2]) ? node99 : node96;
														assign node96 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node99 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node102 = (inp[2]) ? node106 : node103;
														assign node103 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node106 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node109 = (inp[0]) ? node119 : node110;
													assign node110 = (inp[3]) ? node114 : node111;
														assign node111 = (inp[10]) ? 4'b1000 : 4'b1001;
														assign node114 = (inp[2]) ? 4'b1001 : node115;
															assign node115 = (inp[10]) ? 4'b1001 : 4'b1000;
													assign node119 = (inp[2]) ? node121 : 4'b1011;
														assign node121 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node124 = (inp[10]) ? node144 : node125;
												assign node125 = (inp[15]) ? node139 : node126;
													assign node126 = (inp[0]) ? node134 : node127;
														assign node127 = (inp[8]) ? node131 : node128;
															assign node128 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node131 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node134 = (inp[3]) ? node136 : 4'b1001;
															assign node136 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node139 = (inp[3]) ? node141 : 4'b1000;
														assign node141 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node144 = (inp[8]) ? node148 : node145;
													assign node145 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node148 = (inp[2]) ? node150 : 4'b1100;
														assign node150 = (inp[0]) ? 4'b1101 : node151;
															assign node151 = (inp[3]) ? 4'b1111 : 4'b1101;
									assign node155 = (inp[4]) ? node275 : node156;
										assign node156 = (inp[12]) ? node214 : node157;
											assign node157 = (inp[3]) ? node181 : node158;
												assign node158 = (inp[0]) ? node168 : node159;
													assign node159 = (inp[15]) ? 4'b1000 : node160;
														assign node160 = (inp[2]) ? node164 : node161;
															assign node161 = (inp[8]) ? 4'b1010 : 4'b1011;
															assign node164 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node168 = (inp[15]) ? node172 : node169;
														assign node169 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node172 = (inp[10]) ? node174 : 4'b1011;
															assign node174 = (inp[2]) ? node178 : node175;
																assign node175 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node178 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node181 = (inp[8]) ? node197 : node182;
													assign node182 = (inp[2]) ? node190 : node183;
														assign node183 = (inp[10]) ? node187 : node184;
															assign node184 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node187 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node190 = (inp[15]) ? node194 : node191;
															assign node191 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node194 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node197 = (inp[2]) ? node205 : node198;
														assign node198 = (inp[10]) ? 4'b1000 : node199;
															assign node199 = (inp[0]) ? node201 : 4'b1010;
																assign node201 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node205 = (inp[10]) ? 4'b1011 : node206;
															assign node206 = (inp[15]) ? node210 : node207;
																assign node207 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node210 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node214 = (inp[10]) ? node240 : node215;
												assign node215 = (inp[15]) ? node227 : node216;
													assign node216 = (inp[0]) ? node222 : node217;
														assign node217 = (inp[3]) ? 4'b1010 : node218;
															assign node218 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node222 = (inp[2]) ? node224 : 4'b1000;
															assign node224 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node227 = (inp[0]) ? node235 : node228;
														assign node228 = (inp[3]) ? node230 : 4'b1001;
															assign node230 = (inp[8]) ? 4'b1000 : node231;
																assign node231 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node235 = (inp[8]) ? 4'b1010 : node236;
															assign node236 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node240 = (inp[15]) ? node256 : node241;
													assign node241 = (inp[3]) ? node249 : node242;
														assign node242 = (inp[0]) ? 4'b1101 : node243;
															assign node243 = (inp[8]) ? node245 : 4'b1111;
																assign node245 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node249 = (inp[0]) ? node251 : 4'b1101;
															assign node251 = (inp[2]) ? 4'b1110 : node252;
																assign node252 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node256 = (inp[8]) ? node264 : node257;
														assign node257 = (inp[3]) ? node261 : node258;
															assign node258 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node261 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node264 = (inp[2]) ? node270 : node265;
															assign node265 = (inp[3]) ? 4'b1100 : node266;
																assign node266 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node270 = (inp[3]) ? node272 : 4'b1101;
																assign node272 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node275 = (inp[10]) ? node329 : node276;
											assign node276 = (inp[2]) ? node306 : node277;
												assign node277 = (inp[8]) ? node287 : node278;
													assign node278 = (inp[15]) ? 4'b1111 : node279;
														assign node279 = (inp[0]) ? node283 : node280;
															assign node280 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node283 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node287 = (inp[3]) ? node301 : node288;
														assign node288 = (inp[12]) ? node296 : node289;
															assign node289 = (inp[0]) ? node293 : node290;
																assign node290 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node293 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node296 = (inp[15]) ? node298 : 4'b1110;
																assign node298 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node301 = (inp[15]) ? node303 : 4'b1100;
															assign node303 = (inp[12]) ? 4'b1100 : 4'b1110;
												assign node306 = (inp[8]) ? node326 : node307;
													assign node307 = (inp[15]) ? node319 : node308;
														assign node308 = (inp[12]) ? node314 : node309;
															assign node309 = (inp[3]) ? node311 : 4'b1100;
																assign node311 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node314 = (inp[0]) ? 4'b1100 : node315;
																assign node315 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node319 = (inp[3]) ? node323 : node320;
															assign node320 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node323 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node326 = (inp[12]) ? 4'b1111 : 4'b1101;
											assign node329 = (inp[12]) ? node357 : node330;
												assign node330 = (inp[0]) ? node350 : node331;
													assign node331 = (inp[15]) ? node343 : node332;
														assign node332 = (inp[3]) ? node340 : node333;
															assign node333 = (inp[8]) ? node337 : node334;
																assign node334 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node337 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node340 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node343 = (inp[3]) ? node345 : 4'b1101;
															assign node345 = (inp[8]) ? node347 : 4'b1111;
																assign node347 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node350 = (inp[8]) ? node354 : node351;
														assign node351 = (inp[2]) ? 4'b1110 : 4'b1101;
														assign node354 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node357 = (inp[2]) ? node367 : node358;
													assign node358 = (inp[8]) ? 4'b1000 : node359;
														assign node359 = (inp[0]) ? node363 : node360;
															assign node360 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node363 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node367 = (inp[8]) ? node379 : node368;
														assign node368 = (inp[15]) ? node374 : node369;
															assign node369 = (inp[3]) ? 4'b1000 : node370;
																assign node370 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node374 = (inp[0]) ? node376 : 4'b1010;
																assign node376 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node379 = (inp[15]) ? node381 : 4'b1011;
															assign node381 = (inp[0]) ? node383 : 4'b1011;
																assign node383 = (inp[3]) ? 4'b1001 : 4'b1011;
								assign node386 = (inp[2]) ? node610 : node387;
									assign node387 = (inp[8]) ? node507 : node388;
										assign node388 = (inp[10]) ? node452 : node389;
											assign node389 = (inp[15]) ? node423 : node390;
												assign node390 = (inp[0]) ? node400 : node391;
													assign node391 = (inp[9]) ? node395 : node392;
														assign node392 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node395 = (inp[3]) ? 4'b1101 : node396;
															assign node396 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node400 = (inp[12]) ? node412 : node401;
														assign node401 = (inp[3]) ? node409 : node402;
															assign node402 = (inp[4]) ? node406 : node403;
																assign node403 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node406 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node409 = (inp[9]) ? 4'b1111 : 4'b1101;
														assign node412 = (inp[3]) ? node418 : node413;
															assign node413 = (inp[9]) ? 4'b1101 : node414;
																assign node414 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node418 = (inp[9]) ? 4'b1001 : node419;
																assign node419 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node423 = (inp[0]) ? node433 : node424;
													assign node424 = (inp[9]) ? node428 : node425;
														assign node425 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node428 = (inp[4]) ? node430 : 4'b1001;
															assign node430 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node433 = (inp[3]) ? node447 : node434;
														assign node434 = (inp[12]) ? node440 : node435;
															assign node435 = (inp[9]) ? 4'b1011 : node436;
																assign node436 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node440 = (inp[9]) ? node444 : node441;
																assign node441 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node444 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node447 = (inp[4]) ? 4'b1101 : node448;
															assign node448 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node452 = (inp[4]) ? node478 : node453;
												assign node453 = (inp[15]) ? node469 : node454;
													assign node454 = (inp[0]) ? node460 : node455;
														assign node455 = (inp[9]) ? node457 : 4'b1111;
															assign node457 = (inp[3]) ? 4'b1011 : 4'b1111;
														assign node460 = (inp[9]) ? node464 : node461;
															assign node461 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node464 = (inp[12]) ? node466 : 4'b1001;
																assign node466 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node469 = (inp[0]) ? 4'b1011 : node470;
														assign node470 = (inp[3]) ? node472 : 4'b1001;
															assign node472 = (inp[12]) ? 4'b1111 : node473;
																assign node473 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node478 = (inp[15]) ? node494 : node479;
													assign node479 = (inp[3]) ? node489 : node480;
														assign node480 = (inp[0]) ? 4'b1101 : node481;
															assign node481 = (inp[12]) ? node485 : node482;
																assign node482 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node485 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node489 = (inp[12]) ? node491 : 4'b1011;
															assign node491 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node494 = (inp[0]) ? node498 : node495;
														assign node495 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node498 = (inp[3]) ? node500 : 4'b1111;
															assign node500 = (inp[9]) ? node504 : node501;
																assign node501 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node504 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node507 = (inp[12]) ? node551 : node508;
											assign node508 = (inp[15]) ? node528 : node509;
												assign node509 = (inp[0]) ? node513 : node510;
													assign node510 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node513 = (inp[10]) ? node521 : node514;
														assign node514 = (inp[4]) ? node518 : node515;
															assign node515 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node518 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node521 = (inp[3]) ? 4'b1110 : node522;
															assign node522 = (inp[4]) ? 4'b1100 : node523;
																assign node523 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node528 = (inp[0]) ? node542 : node529;
													assign node529 = (inp[3]) ? node537 : node530;
														assign node530 = (inp[9]) ? node534 : node531;
															assign node531 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node534 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node537 = (inp[9]) ? node539 : 4'b1000;
															assign node539 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node542 = (inp[4]) ? node546 : node543;
														assign node543 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node546 = (inp[3]) ? 4'b1100 : node547;
															assign node547 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node551 = (inp[4]) ? node579 : node552;
												assign node552 = (inp[3]) ? node564 : node553;
													assign node553 = (inp[15]) ? node561 : node554;
														assign node554 = (inp[9]) ? node558 : node555;
															assign node555 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node558 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node561 = (inp[10]) ? 4'b1110 : 4'b1100;
													assign node564 = (inp[15]) ? node568 : node565;
														assign node565 = (inp[0]) ? 4'b1110 : 4'b1010;
														assign node568 = (inp[10]) ? node572 : node569;
															assign node569 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node572 = (inp[9]) ? node576 : node573;
																assign node573 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node576 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node579 = (inp[0]) ? node599 : node580;
													assign node580 = (inp[3]) ? node590 : node581;
														assign node581 = (inp[15]) ? 4'b1000 : node582;
															assign node582 = (inp[10]) ? node586 : node583;
																assign node583 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node586 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node590 = (inp[15]) ? node592 : 4'b1100;
															assign node592 = (inp[9]) ? node596 : node593;
																assign node593 = (inp[10]) ? 4'b1110 : 4'b1000;
																assign node596 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node599 = (inp[10]) ? node603 : node600;
														assign node600 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node603 = (inp[9]) ? node605 : 4'b1110;
															assign node605 = (inp[3]) ? node607 : 4'b1010;
																assign node607 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node610 = (inp[8]) ? node696 : node611;
										assign node611 = (inp[3]) ? node653 : node612;
											assign node612 = (inp[9]) ? node636 : node613;
												assign node613 = (inp[4]) ? node625 : node614;
													assign node614 = (inp[10]) ? node620 : node615;
														assign node615 = (inp[12]) ? node617 : 4'b1100;
															assign node617 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node620 = (inp[12]) ? 4'b1010 : node621;
															assign node621 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node625 = (inp[12]) ? node631 : node626;
														assign node626 = (inp[15]) ? node628 : 4'b1010;
															assign node628 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node631 = (inp[10]) ? 4'b1100 : node632;
															assign node632 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node636 = (inp[15]) ? node644 : node637;
													assign node637 = (inp[0]) ? 4'b1000 : node638;
														assign node638 = (inp[10]) ? 4'b1010 : node639;
															assign node639 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node644 = (inp[0]) ? node646 : 4'b1000;
														assign node646 = (inp[12]) ? node648 : 4'b1010;
															assign node648 = (inp[10]) ? 4'b1110 : node649;
																assign node649 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node653 = (inp[0]) ? node675 : node654;
												assign node654 = (inp[4]) ? node666 : node655;
													assign node655 = (inp[10]) ? node659 : node656;
														assign node656 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node659 = (inp[12]) ? node663 : node660;
															assign node660 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node663 = (inp[15]) ? 4'b1000 : 4'b1100;
													assign node666 = (inp[9]) ? node672 : node667;
														assign node667 = (inp[10]) ? node669 : 4'b1010;
															assign node669 = (inp[12]) ? 4'b1100 : 4'b1010;
														assign node672 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node675 = (inp[15]) ? node687 : node676;
													assign node676 = (inp[10]) ? node678 : 4'b1000;
														assign node678 = (inp[4]) ? 4'b1110 : node679;
															assign node679 = (inp[12]) ? node683 : node680;
																assign node680 = (inp[9]) ? 4'b1000 : 4'b1100;
																assign node683 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node687 = (inp[4]) ? node691 : node688;
														assign node688 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node691 = (inp[9]) ? node693 : 4'b1010;
															assign node693 = (inp[10]) ? 4'b1000 : 4'b1100;
										assign node696 = (inp[9]) ? node746 : node697;
											assign node697 = (inp[4]) ? node721 : node698;
												assign node698 = (inp[12]) ? node712 : node699;
													assign node699 = (inp[3]) ? node707 : node700;
														assign node700 = (inp[15]) ? node704 : node701;
															assign node701 = (inp[10]) ? 4'b0111 : 4'b0101;
															assign node704 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node707 = (inp[10]) ? 4'b0101 : node708;
															assign node708 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node712 = (inp[10]) ? node714 : 4'b0111;
														assign node714 = (inp[15]) ? node718 : node715;
															assign node715 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node718 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node721 = (inp[12]) ? node735 : node722;
													assign node722 = (inp[3]) ? node730 : node723;
														assign node723 = (inp[15]) ? node727 : node724;
															assign node724 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node727 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node730 = (inp[15]) ? node732 : 4'b0011;
															assign node732 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node735 = (inp[10]) ? node743 : node736;
														assign node736 = (inp[3]) ? node740 : node737;
															assign node737 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node740 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node743 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node746 = (inp[4]) ? node760 : node747;
												assign node747 = (inp[12]) ? node753 : node748;
													assign node748 = (inp[15]) ? 4'b0011 : node749;
														assign node749 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node753 = (inp[10]) ? node755 : 4'b0001;
														assign node755 = (inp[0]) ? node757 : 4'b0111;
															assign node757 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node760 = (inp[3]) ? node770 : node761;
													assign node761 = (inp[10]) ? node765 : node762;
														assign node762 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node765 = (inp[0]) ? node767 : 4'b0001;
															assign node767 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node770 = (inp[12]) ? node776 : node771;
														assign node771 = (inp[15]) ? node773 : 4'b0111;
															assign node773 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node776 = (inp[15]) ? 4'b0111 : 4'b0101;
							assign node779 = (inp[13]) ? node1157 : node780;
								assign node780 = (inp[2]) ? node974 : node781;
									assign node781 = (inp[8]) ? node877 : node782;
										assign node782 = (inp[10]) ? node816 : node783;
											assign node783 = (inp[15]) ? node791 : node784;
												assign node784 = (inp[0]) ? 4'b1001 : node785;
													assign node785 = (inp[9]) ? 4'b1011 : node786;
														assign node786 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node791 = (inp[0]) ? node799 : node792;
													assign node792 = (inp[4]) ? node796 : node793;
														assign node793 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node796 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node799 = (inp[12]) ? node811 : node800;
														assign node800 = (inp[3]) ? node808 : node801;
															assign node801 = (inp[9]) ? node805 : node802;
																assign node802 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node805 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node808 = (inp[9]) ? 4'b1101 : 4'b1111;
														assign node811 = (inp[4]) ? 4'b1011 : node812;
															assign node812 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node816 = (inp[0]) ? node840 : node817;
												assign node817 = (inp[15]) ? node827 : node818;
													assign node818 = (inp[9]) ? 4'b1011 : node819;
														assign node819 = (inp[4]) ? node823 : node820;
															assign node820 = (inp[3]) ? 4'b1011 : 4'b1111;
															assign node823 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node827 = (inp[4]) ? node837 : node828;
														assign node828 = (inp[3]) ? node830 : 4'b1101;
															assign node830 = (inp[12]) ? node834 : node831;
																assign node831 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node834 = (inp[9]) ? 4'b1111 : 4'b1001;
														assign node837 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node840 = (inp[15]) ? node860 : node841;
													assign node841 = (inp[3]) ? node851 : node842;
														assign node842 = (inp[4]) ? node844 : 4'b1101;
															assign node844 = (inp[12]) ? node848 : node845;
																assign node845 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node848 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node851 = (inp[12]) ? 4'b1011 : node852;
															assign node852 = (inp[9]) ? node856 : node853;
																assign node853 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node856 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node860 = (inp[9]) ? node866 : node861;
														assign node861 = (inp[3]) ? 4'b1011 : node862;
															assign node862 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node866 = (inp[3]) ? node872 : node867;
															assign node867 = (inp[4]) ? node869 : 4'b1011;
																assign node869 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node872 = (inp[12]) ? 4'b1101 : node873;
																assign node873 = (inp[4]) ? 4'b1101 : 4'b1011;
										assign node877 = (inp[0]) ? node927 : node878;
											assign node878 = (inp[15]) ? node908 : node879;
												assign node879 = (inp[12]) ? node895 : node880;
													assign node880 = (inp[3]) ? node890 : node881;
														assign node881 = (inp[10]) ? node887 : node882;
															assign node882 = (inp[9]) ? 4'b1110 : node883;
																assign node883 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node887 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node890 = (inp[4]) ? 4'b1010 : node891;
															assign node891 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node895 = (inp[3]) ? node905 : node896;
														assign node896 = (inp[4]) ? node898 : 4'b1110;
															assign node898 = (inp[10]) ? node902 : node899;
																assign node899 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node902 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node905 = (inp[10]) ? 4'b1100 : 4'b1110;
												assign node908 = (inp[3]) ? node918 : node909;
													assign node909 = (inp[10]) ? 4'b1100 : node910;
														assign node910 = (inp[4]) ? node914 : node911;
															assign node911 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node914 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node918 = (inp[9]) ? node924 : node919;
														assign node919 = (inp[4]) ? 4'b1000 : node920;
															assign node920 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node924 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node927 = (inp[15]) ? node953 : node928;
												assign node928 = (inp[12]) ? node938 : node929;
													assign node929 = (inp[10]) ? 4'b1000 : node930;
														assign node930 = (inp[3]) ? 4'b1000 : node931;
															assign node931 = (inp[9]) ? 4'b1100 : node932;
																assign node932 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node938 = (inp[3]) ? node946 : node939;
														assign node939 = (inp[9]) ? 4'b1000 : node940;
															assign node940 = (inp[4]) ? node942 : 4'b1100;
																assign node942 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node946 = (inp[4]) ? 4'b1110 : node947;
															assign node947 = (inp[9]) ? 4'b1000 : node948;
																assign node948 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node953 = (inp[3]) ? node963 : node954;
													assign node954 = (inp[10]) ? 4'b1010 : node955;
														assign node955 = (inp[4]) ? node959 : node956;
															assign node956 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node959 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node963 = (inp[10]) ? node965 : 4'b1010;
														assign node965 = (inp[4]) ? node969 : node966;
															assign node966 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node969 = (inp[9]) ? node971 : 4'b1100;
																assign node971 = (inp[12]) ? 4'b1000 : 4'b1100;
									assign node974 = (inp[8]) ? node1070 : node975;
										assign node975 = (inp[12]) ? node1021 : node976;
											assign node976 = (inp[9]) ? node990 : node977;
												assign node977 = (inp[4]) ? node983 : node978;
													assign node978 = (inp[0]) ? 4'b1110 : node979;
														assign node979 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node983 = (inp[3]) ? node985 : 4'b1010;
														assign node985 = (inp[10]) ? 4'b1010 : node986;
															assign node986 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node990 = (inp[4]) ? node1004 : node991;
													assign node991 = (inp[10]) ? node997 : node992;
														assign node992 = (inp[15]) ? 4'b1000 : node993;
															assign node993 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node997 = (inp[15]) ? node1001 : node998;
															assign node998 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node1001 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node1004 = (inp[10]) ? node1014 : node1005;
														assign node1005 = (inp[15]) ? 4'b1100 : node1006;
															assign node1006 = (inp[0]) ? node1010 : node1007;
																assign node1007 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node1010 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node1014 = (inp[0]) ? 4'b1110 : node1015;
															assign node1015 = (inp[3]) ? 4'b1110 : node1016;
																assign node1016 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node1021 = (inp[3]) ? node1045 : node1022;
												assign node1022 = (inp[10]) ? node1034 : node1023;
													assign node1023 = (inp[0]) ? node1031 : node1024;
														assign node1024 = (inp[15]) ? node1026 : 4'b1010;
															assign node1026 = (inp[9]) ? 4'b1000 : node1027;
																assign node1027 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node1031 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node1034 = (inp[4]) ? node1040 : node1035;
														assign node1035 = (inp[0]) ? 4'b1000 : node1036;
															assign node1036 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node1040 = (inp[0]) ? node1042 : 4'b1110;
															assign node1042 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node1045 = (inp[0]) ? node1059 : node1046;
													assign node1046 = (inp[9]) ? node1052 : node1047;
														assign node1047 = (inp[10]) ? node1049 : 4'b1110;
															assign node1049 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node1052 = (inp[10]) ? node1056 : node1053;
															assign node1053 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node1056 = (inp[15]) ? 4'b1110 : 4'b1000;
													assign node1059 = (inp[9]) ? node1067 : node1060;
														assign node1060 = (inp[15]) ? 4'b1100 : node1061;
															assign node1061 = (inp[10]) ? 4'b1000 : node1062;
																assign node1062 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node1067 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node1070 = (inp[12]) ? node1110 : node1071;
											assign node1071 = (inp[9]) ? node1091 : node1072;
												assign node1072 = (inp[4]) ? node1076 : node1073;
													assign node1073 = (inp[10]) ? 4'b0111 : 4'b0101;
													assign node1076 = (inp[3]) ? node1082 : node1077;
														assign node1077 = (inp[0]) ? node1079 : 4'b0011;
															assign node1079 = (inp[10]) ? 4'b0001 : 4'b0011;
														assign node1082 = (inp[10]) ? 4'b0011 : node1083;
															assign node1083 = (inp[15]) ? node1087 : node1084;
																assign node1084 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node1087 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node1091 = (inp[4]) ? node1099 : node1092;
													assign node1092 = (inp[10]) ? 4'b0001 : node1093;
														assign node1093 = (inp[0]) ? 4'b0011 : node1094;
															assign node1094 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node1099 = (inp[0]) ? node1101 : 4'b0111;
														assign node1101 = (inp[10]) ? node1105 : node1102;
															assign node1102 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node1105 = (inp[15]) ? node1107 : 4'b0111;
																assign node1107 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node1110 = (inp[9]) ? node1126 : node1111;
												assign node1111 = (inp[0]) ? node1117 : node1112;
													assign node1112 = (inp[15]) ? 4'b0101 : node1113;
														assign node1113 = (inp[4]) ? 4'b0101 : 4'b0111;
													assign node1117 = (inp[4]) ? node1119 : 4'b0101;
														assign node1119 = (inp[10]) ? node1121 : 4'b0011;
															assign node1121 = (inp[15]) ? node1123 : 4'b0111;
																assign node1123 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node1126 = (inp[3]) ? node1138 : node1127;
													assign node1127 = (inp[0]) ? node1133 : node1128;
														assign node1128 = (inp[10]) ? node1130 : 4'b0001;
															assign node1130 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node1133 = (inp[15]) ? 4'b0011 : node1134;
															assign node1134 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node1138 = (inp[10]) ? node1152 : node1139;
														assign node1139 = (inp[4]) ? node1145 : node1140;
															assign node1140 = (inp[15]) ? node1142 : 4'b0001;
																assign node1142 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node1145 = (inp[0]) ? node1149 : node1146;
																assign node1146 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node1149 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node1152 = (inp[4]) ? node1154 : 4'b0111;
															assign node1154 = (inp[15]) ? 4'b0011 : 4'b0001;
								assign node1157 = (inp[12]) ? node1325 : node1158;
									assign node1158 = (inp[9]) ? node1236 : node1159;
										assign node1159 = (inp[4]) ? node1207 : node1160;
											assign node1160 = (inp[8]) ? node1188 : node1161;
												assign node1161 = (inp[2]) ? node1171 : node1162;
													assign node1162 = (inp[3]) ? 4'b0111 : node1163;
														assign node1163 = (inp[10]) ? node1165 : 4'b0101;
															assign node1165 = (inp[15]) ? node1167 : 4'b0111;
																assign node1167 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node1171 = (inp[3]) ? node1183 : node1172;
														assign node1172 = (inp[10]) ? node1178 : node1173;
															assign node1173 = (inp[0]) ? node1175 : 4'b0110;
																assign node1175 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node1178 = (inp[0]) ? 4'b0100 : node1179;
																assign node1179 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node1183 = (inp[10]) ? node1185 : 4'b0100;
															assign node1185 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node1188 = (inp[2]) ? node1200 : node1189;
													assign node1189 = (inp[10]) ? node1195 : node1190;
														assign node1190 = (inp[0]) ? 4'b0110 : node1191;
															assign node1191 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node1195 = (inp[3]) ? 4'b0100 : node1196;
															assign node1196 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node1200 = (inp[15]) ? node1204 : node1201;
														assign node1201 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node1204 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node1207 = (inp[0]) ? node1221 : node1208;
												assign node1208 = (inp[15]) ? node1216 : node1209;
													assign node1209 = (inp[8]) ? node1213 : node1210;
														assign node1210 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node1213 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node1216 = (inp[2]) ? node1218 : 4'b0001;
														assign node1218 = (inp[8]) ? 4'b0001 : 4'b0000;
												assign node1221 = (inp[15]) ? node1229 : node1222;
													assign node1222 = (inp[2]) ? node1226 : node1223;
														assign node1223 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node1226 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node1229 = (inp[8]) ? node1233 : node1230;
														assign node1230 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node1233 = (inp[2]) ? 4'b0011 : 4'b0010;
										assign node1236 = (inp[4]) ? node1264 : node1237;
											assign node1237 = (inp[2]) ? node1253 : node1238;
												assign node1238 = (inp[8]) ? node1246 : node1239;
													assign node1239 = (inp[3]) ? node1241 : 4'b0001;
														assign node1241 = (inp[15]) ? node1243 : 4'b0011;
															assign node1243 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node1246 = (inp[15]) ? node1250 : node1247;
														assign node1247 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node1250 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node1253 = (inp[8]) ? 4'b0011 : node1254;
													assign node1254 = (inp[10]) ? 4'b0010 : node1255;
														assign node1255 = (inp[3]) ? node1257 : 4'b0000;
															assign node1257 = (inp[15]) ? node1259 : 4'b0010;
																assign node1259 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node1264 = (inp[3]) ? node1292 : node1265;
												assign node1265 = (inp[2]) ? node1275 : node1266;
													assign node1266 = (inp[8]) ? 4'b0110 : node1267;
														assign node1267 = (inp[0]) ? node1271 : node1268;
															assign node1268 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node1271 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node1275 = (inp[8]) ? node1285 : node1276;
														assign node1276 = (inp[10]) ? node1278 : 4'b0100;
															assign node1278 = (inp[0]) ? node1282 : node1279;
																assign node1279 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node1282 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node1285 = (inp[0]) ? node1289 : node1286;
															assign node1286 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node1289 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node1292 = (inp[0]) ? node1312 : node1293;
													assign node1293 = (inp[15]) ? node1305 : node1294;
														assign node1294 = (inp[10]) ? node1300 : node1295;
															assign node1295 = (inp[8]) ? 4'b0100 : node1296;
																assign node1296 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node1300 = (inp[8]) ? node1302 : 4'b0101;
																assign node1302 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node1305 = (inp[2]) ? node1309 : node1306;
															assign node1306 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node1309 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node1312 = (inp[15]) ? node1318 : node1313;
														assign node1313 = (inp[2]) ? 4'b0111 : node1314;
															assign node1314 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node1318 = (inp[8]) ? node1322 : node1319;
															assign node1319 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node1322 = (inp[2]) ? 4'b0101 : 4'b0100;
									assign node1325 = (inp[4]) ? node1443 : node1326;
										assign node1326 = (inp[3]) ? node1392 : node1327;
											assign node1327 = (inp[8]) ? node1359 : node1328;
												assign node1328 = (inp[2]) ? node1346 : node1329;
													assign node1329 = (inp[9]) ? node1337 : node1330;
														assign node1330 = (inp[10]) ? 4'b0001 : node1331;
															assign node1331 = (inp[0]) ? 4'b0101 : node1332;
																assign node1332 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node1337 = (inp[10]) ? 4'b0101 : node1338;
															assign node1338 = (inp[0]) ? node1342 : node1339;
																assign node1339 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node1342 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node1346 = (inp[9]) ? node1356 : node1347;
														assign node1347 = (inp[10]) ? node1353 : node1348;
															assign node1348 = (inp[15]) ? 4'b0110 : node1349;
																assign node1349 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node1353 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node1356 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node1359 = (inp[2]) ? node1381 : node1360;
													assign node1360 = (inp[9]) ? node1372 : node1361;
														assign node1361 = (inp[10]) ? node1367 : node1362;
															assign node1362 = (inp[0]) ? node1364 : 4'b0100;
																assign node1364 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node1367 = (inp[15]) ? 4'b0000 : node1368;
																assign node1368 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node1372 = (inp[10]) ? node1374 : 4'b0010;
															assign node1374 = (inp[0]) ? node1378 : node1375;
																assign node1375 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node1378 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node1381 = (inp[0]) ? node1385 : node1382;
														assign node1382 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node1385 = (inp[15]) ? node1387 : 4'b0101;
															assign node1387 = (inp[10]) ? node1389 : 4'b0011;
																assign node1389 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node1392 = (inp[9]) ? node1412 : node1393;
												assign node1393 = (inp[10]) ? node1397 : node1394;
													assign node1394 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node1397 = (inp[8]) ? node1401 : node1398;
														assign node1398 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node1401 = (inp[2]) ? node1407 : node1402;
															assign node1402 = (inp[0]) ? 4'b0010 : node1403;
																assign node1403 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node1407 = (inp[0]) ? node1409 : 4'b0001;
																assign node1409 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node1412 = (inp[10]) ? node1424 : node1413;
													assign node1413 = (inp[8]) ? node1417 : node1414;
														assign node1414 = (inp[2]) ? 4'b0010 : 4'b0001;
														assign node1417 = (inp[2]) ? 4'b0001 : node1418;
															assign node1418 = (inp[0]) ? node1420 : 4'b0000;
																assign node1420 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node1424 = (inp[8]) ? node1432 : node1425;
														assign node1425 = (inp[2]) ? node1427 : 4'b0111;
															assign node1427 = (inp[15]) ? 4'b0110 : node1428;
																assign node1428 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node1432 = (inp[2]) ? node1438 : node1433;
															assign node1433 = (inp[0]) ? node1435 : 4'b0100;
																assign node1435 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node1438 = (inp[15]) ? node1440 : 4'b0101;
																assign node1440 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node1443 = (inp[0]) ? node1487 : node1444;
											assign node1444 = (inp[15]) ? node1464 : node1445;
												assign node1445 = (inp[3]) ? node1451 : node1446;
													assign node1446 = (inp[9]) ? 4'b0111 : node1447;
														assign node1447 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node1451 = (inp[8]) ? node1461 : node1452;
														assign node1452 = (inp[2]) ? node1454 : 4'b0001;
															assign node1454 = (inp[9]) ? node1458 : node1455;
																assign node1455 = (inp[10]) ? 4'b0100 : 4'b0010;
																assign node1458 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node1461 = (inp[10]) ? 4'b0100 : 4'b0101;
												assign node1464 = (inp[3]) ? node1478 : node1465;
													assign node1465 = (inp[8]) ? node1475 : node1466;
														assign node1466 = (inp[2]) ? node1472 : node1467;
															assign node1467 = (inp[10]) ? 4'b0101 : node1468;
																assign node1468 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node1472 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node1475 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node1478 = (inp[10]) ? node1482 : node1479;
														assign node1479 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node1482 = (inp[9]) ? 4'b0011 : node1483;
															assign node1483 = (inp[8]) ? 4'b0111 : 4'b0110;
											assign node1487 = (inp[8]) ? node1513 : node1488;
												assign node1488 = (inp[2]) ? node1504 : node1489;
													assign node1489 = (inp[10]) ? node1495 : node1490;
														assign node1490 = (inp[3]) ? 4'b0101 : node1491;
															assign node1491 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node1495 = (inp[9]) ? 4'b0011 : node1496;
															assign node1496 = (inp[3]) ? node1500 : node1497;
																assign node1497 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node1500 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node1504 = (inp[9]) ? node1510 : node1505;
														assign node1505 = (inp[10]) ? 4'b0100 : node1506;
															assign node1506 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node1510 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node1513 = (inp[2]) ? node1533 : node1514;
													assign node1514 = (inp[15]) ? node1526 : node1515;
														assign node1515 = (inp[3]) ? node1521 : node1516;
															assign node1516 = (inp[9]) ? 4'b0000 : node1517;
																assign node1517 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node1521 = (inp[9]) ? node1523 : 4'b0000;
																assign node1523 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node1526 = (inp[3]) ? 4'b0100 : node1527;
															assign node1527 = (inp[9]) ? 4'b0010 : node1528;
																assign node1528 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node1533 = (inp[15]) ? node1535 : 4'b0001;
														assign node1535 = (inp[10]) ? node1539 : node1536;
															assign node1536 = (inp[3]) ? 4'b0011 : 4'b0111;
															assign node1539 = (inp[9]) ? 4'b0001 : 4'b0101;
						assign node1542 = (inp[1]) ? node2226 : node1543;
							assign node1543 = (inp[2]) ? node1875 : node1544;
								assign node1544 = (inp[8]) ? node1696 : node1545;
									assign node1545 = (inp[15]) ? node1619 : node1546;
										assign node1546 = (inp[0]) ? node1574 : node1547;
											assign node1547 = (inp[9]) ? node1559 : node1548;
												assign node1548 = (inp[4]) ? node1554 : node1549;
													assign node1549 = (inp[10]) ? node1551 : 4'b0111;
														assign node1551 = (inp[13]) ? 4'b0111 : 4'b0011;
													assign node1554 = (inp[10]) ? node1556 : 4'b0011;
														assign node1556 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node1559 = (inp[4]) ? node1565 : node1560;
													assign node1560 = (inp[12]) ? node1562 : 4'b0011;
														assign node1562 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node1565 = (inp[3]) ? node1571 : node1566;
														assign node1566 = (inp[12]) ? node1568 : 4'b0111;
															assign node1568 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node1571 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node1574 = (inp[3]) ? node1608 : node1575;
												assign node1575 = (inp[12]) ? node1601 : node1576;
													assign node1576 = (inp[10]) ? node1592 : node1577;
														assign node1577 = (inp[13]) ? node1585 : node1578;
															assign node1578 = (inp[4]) ? node1582 : node1579;
																assign node1579 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node1582 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node1585 = (inp[4]) ? node1589 : node1586;
																assign node1586 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node1589 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node1592 = (inp[13]) ? node1598 : node1593;
															assign node1593 = (inp[4]) ? node1595 : 4'b0001;
																assign node1595 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node1598 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node1601 = (inp[13]) ? node1603 : 4'b0101;
														assign node1603 = (inp[9]) ? node1605 : 4'b0001;
															assign node1605 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node1608 = (inp[4]) ? node1612 : node1609;
													assign node1609 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node1612 = (inp[9]) ? node1614 : 4'b0001;
														assign node1614 = (inp[12]) ? node1616 : 4'b0111;
															assign node1616 = (inp[10]) ? 4'b0011 : 4'b0111;
										assign node1619 = (inp[0]) ? node1659 : node1620;
											assign node1620 = (inp[3]) ? node1638 : node1621;
												assign node1621 = (inp[9]) ? node1631 : node1622;
													assign node1622 = (inp[12]) ? node1626 : node1623;
														assign node1623 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node1626 = (inp[10]) ? node1628 : 4'b0001;
															assign node1628 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node1631 = (inp[4]) ? node1633 : 4'b0001;
														assign node1633 = (inp[12]) ? node1635 : 4'b0101;
															assign node1635 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node1638 = (inp[10]) ? node1644 : node1639;
													assign node1639 = (inp[9]) ? 4'b0001 : node1640;
														assign node1640 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node1644 = (inp[4]) ? node1652 : node1645;
														assign node1645 = (inp[13]) ? 4'b0001 : node1646;
															assign node1646 = (inp[9]) ? 4'b0111 : node1647;
																assign node1647 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node1652 = (inp[12]) ? node1656 : node1653;
															assign node1653 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node1656 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node1659 = (inp[3]) ? node1679 : node1660;
												assign node1660 = (inp[12]) ? node1666 : node1661;
													assign node1661 = (inp[4]) ? 4'b0011 : node1662;
														assign node1662 = (inp[13]) ? 4'b0011 : 4'b0111;
													assign node1666 = (inp[13]) ? node1674 : node1667;
														assign node1667 = (inp[9]) ? node1669 : 4'b0011;
															assign node1669 = (inp[10]) ? 4'b0011 : node1670;
																assign node1670 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node1674 = (inp[10]) ? 4'b0111 : node1675;
															assign node1675 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node1679 = (inp[9]) ? node1689 : node1680;
													assign node1680 = (inp[13]) ? node1682 : 4'b0011;
														assign node1682 = (inp[4]) ? node1686 : node1683;
															assign node1683 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node1686 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node1689 = (inp[4]) ? 4'b0101 : node1690;
														assign node1690 = (inp[10]) ? node1692 : 4'b0011;
															assign node1692 = (inp[12]) ? 4'b0101 : 4'b0011;
									assign node1696 = (inp[4]) ? node1790 : node1697;
										assign node1697 = (inp[9]) ? node1749 : node1698;
											assign node1698 = (inp[12]) ? node1724 : node1699;
												assign node1699 = (inp[3]) ? node1711 : node1700;
													assign node1700 = (inp[10]) ? node1702 : 4'b0110;
														assign node1702 = (inp[13]) ? node1704 : 4'b0110;
															assign node1704 = (inp[15]) ? node1708 : node1705;
																assign node1705 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node1708 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node1711 = (inp[13]) ? node1719 : node1712;
														assign node1712 = (inp[15]) ? node1716 : node1713;
															assign node1713 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node1716 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node1719 = (inp[15]) ? node1721 : 4'b0100;
															assign node1721 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node1724 = (inp[10]) ? node1736 : node1725;
													assign node1725 = (inp[13]) ? node1729 : node1726;
														assign node1726 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node1729 = (inp[3]) ? node1731 : 4'b0100;
															assign node1731 = (inp[15]) ? node1733 : 4'b0100;
																assign node1733 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node1736 = (inp[3]) ? node1744 : node1737;
														assign node1737 = (inp[15]) ? node1741 : node1738;
															assign node1738 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node1741 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node1744 = (inp[15]) ? node1746 : 4'b0000;
															assign node1746 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node1749 = (inp[12]) ? node1771 : node1750;
												assign node1750 = (inp[3]) ? node1766 : node1751;
													assign node1751 = (inp[10]) ? node1759 : node1752;
														assign node1752 = (inp[13]) ? node1754 : 4'b0010;
															assign node1754 = (inp[0]) ? node1756 : 4'b0000;
																assign node1756 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node1759 = (inp[15]) ? node1763 : node1760;
															assign node1760 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node1763 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node1766 = (inp[0]) ? node1768 : 4'b0000;
														assign node1768 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node1771 = (inp[10]) ? node1781 : node1772;
													assign node1772 = (inp[13]) ? 4'b0010 : node1773;
														assign node1773 = (inp[15]) ? node1777 : node1774;
															assign node1774 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node1777 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node1781 = (inp[3]) ? 4'b0110 : node1782;
														assign node1782 = (inp[13]) ? 4'b0100 : node1783;
															assign node1783 = (inp[15]) ? 4'b0110 : node1784;
																assign node1784 = (inp[0]) ? 4'b0100 : 4'b0110;
										assign node1790 = (inp[9]) ? node1830 : node1791;
											assign node1791 = (inp[12]) ? node1799 : node1792;
												assign node1792 = (inp[15]) ? node1796 : node1793;
													assign node1793 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node1796 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node1799 = (inp[10]) ? node1811 : node1800;
													assign node1800 = (inp[3]) ? node1802 : 4'b0000;
														assign node1802 = (inp[13]) ? node1806 : node1803;
															assign node1803 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node1806 = (inp[15]) ? node1808 : 4'b0000;
																assign node1808 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node1811 = (inp[3]) ? node1823 : node1812;
														assign node1812 = (inp[13]) ? node1818 : node1813;
															assign node1813 = (inp[15]) ? node1815 : 4'b0100;
																assign node1815 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node1818 = (inp[0]) ? node1820 : 4'b0110;
																assign node1820 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node1823 = (inp[13]) ? node1825 : 4'b0110;
															assign node1825 = (inp[15]) ? 4'b0110 : node1826;
																assign node1826 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node1830 = (inp[12]) ? node1852 : node1831;
												assign node1831 = (inp[0]) ? node1845 : node1832;
													assign node1832 = (inp[13]) ? node1840 : node1833;
														assign node1833 = (inp[15]) ? node1837 : node1834;
															assign node1834 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node1837 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node1840 = (inp[10]) ? 4'b0110 : node1841;
															assign node1841 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node1845 = (inp[3]) ? node1849 : node1846;
														assign node1846 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node1849 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node1852 = (inp[10]) ? node1862 : node1853;
													assign node1853 = (inp[15]) ? node1855 : 4'b0100;
														assign node1855 = (inp[13]) ? node1857 : 4'b0110;
															assign node1857 = (inp[0]) ? node1859 : 4'b0110;
																assign node1859 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node1862 = (inp[0]) ? node1868 : node1863;
														assign node1863 = (inp[15]) ? 4'b0000 : node1864;
															assign node1864 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node1868 = (inp[13]) ? node1870 : 4'b0010;
															assign node1870 = (inp[3]) ? 4'b0010 : node1871;
																assign node1871 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node1875 = (inp[8]) ? node2023 : node1876;
									assign node1876 = (inp[15]) ? node1950 : node1877;
										assign node1877 = (inp[0]) ? node1917 : node1878;
											assign node1878 = (inp[3]) ? node1898 : node1879;
												assign node1879 = (inp[9]) ? node1891 : node1880;
													assign node1880 = (inp[4]) ? node1886 : node1881;
														assign node1881 = (inp[10]) ? node1883 : 4'b0110;
															assign node1883 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node1886 = (inp[10]) ? node1888 : 4'b0010;
															assign node1888 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node1891 = (inp[4]) ? 4'b0110 : node1892;
														assign node1892 = (inp[13]) ? 4'b0010 : node1893;
															assign node1893 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node1898 = (inp[4]) ? node1906 : node1899;
													assign node1899 = (inp[9]) ? 4'b0010 : node1900;
														assign node1900 = (inp[12]) ? node1902 : 4'b0110;
															assign node1902 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node1906 = (inp[9]) ? node1912 : node1907;
														assign node1907 = (inp[13]) ? 4'b0010 : node1908;
															assign node1908 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node1912 = (inp[10]) ? node1914 : 4'b0100;
															assign node1914 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node1917 = (inp[3]) ? node1933 : node1918;
												assign node1918 = (inp[4]) ? node1924 : node1919;
													assign node1919 = (inp[9]) ? node1921 : 4'b0100;
														assign node1921 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node1924 = (inp[12]) ? node1926 : 4'b0000;
														assign node1926 = (inp[9]) ? node1930 : node1927;
															assign node1927 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node1930 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node1933 = (inp[12]) ? node1941 : node1934;
													assign node1934 = (inp[9]) ? node1938 : node1935;
														assign node1935 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node1938 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node1941 = (inp[9]) ? node1947 : node1942;
														assign node1942 = (inp[13]) ? node1944 : 4'b0000;
															assign node1944 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node1947 = (inp[13]) ? 4'b0010 : 4'b0110;
										assign node1950 = (inp[0]) ? node1992 : node1951;
											assign node1951 = (inp[3]) ? node1973 : node1952;
												assign node1952 = (inp[4]) ? node1964 : node1953;
													assign node1953 = (inp[12]) ? node1957 : node1954;
														assign node1954 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node1957 = (inp[9]) ? node1961 : node1958;
															assign node1958 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node1961 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node1964 = (inp[12]) ? node1968 : node1965;
														assign node1965 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node1968 = (inp[10]) ? node1970 : 4'b0100;
															assign node1970 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node1973 = (inp[4]) ? node1987 : node1974;
													assign node1974 = (inp[9]) ? node1982 : node1975;
														assign node1975 = (inp[13]) ? node1977 : 4'b0100;
															assign node1977 = (inp[10]) ? node1979 : 4'b0100;
																assign node1979 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node1982 = (inp[13]) ? node1984 : 4'b0000;
															assign node1984 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node1987 = (inp[9]) ? node1989 : 4'b0000;
														assign node1989 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node1992 = (inp[3]) ? node2008 : node1993;
												assign node1993 = (inp[12]) ? node2001 : node1994;
													assign node1994 = (inp[4]) ? node1998 : node1995;
														assign node1995 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node1998 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node2001 = (inp[10]) ? 4'b0110 : node2002;
														assign node2002 = (inp[13]) ? node2004 : 4'b0110;
															assign node2004 = (inp[9]) ? 4'b0110 : 4'b0010;
												assign node2008 = (inp[13]) ? node2016 : node2009;
													assign node2009 = (inp[4]) ? 4'b0100 : node2010;
														assign node2010 = (inp[12]) ? 4'b0100 : node2011;
															assign node2011 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node2016 = (inp[9]) ? node2018 : 4'b0010;
														assign node2018 = (inp[4]) ? node2020 : 4'b0010;
															assign node2020 = (inp[12]) ? 4'b0000 : 4'b0100;
									assign node2023 = (inp[13]) ? node2127 : node2024;
										assign node2024 = (inp[12]) ? node2076 : node2025;
											assign node2025 = (inp[3]) ? node2043 : node2026;
												assign node2026 = (inp[9]) ? node2036 : node2027;
													assign node2027 = (inp[4]) ? node2033 : node2028;
														assign node2028 = (inp[0]) ? 4'b0111 : node2029;
															assign node2029 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node2033 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node2036 = (inp[4]) ? node2038 : 4'b0001;
														assign node2038 = (inp[15]) ? node2040 : 4'b0101;
															assign node2040 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node2043 = (inp[15]) ? node2065 : node2044;
													assign node2044 = (inp[0]) ? node2054 : node2045;
														assign node2045 = (inp[10]) ? node2049 : node2046;
															assign node2046 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node2049 = (inp[9]) ? 4'b0011 : node2050;
																assign node2050 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node2054 = (inp[10]) ? node2060 : node2055;
															assign node2055 = (inp[4]) ? node2057 : 4'b0001;
																assign node2057 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node2060 = (inp[9]) ? 4'b0001 : node2061;
																assign node2061 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node2065 = (inp[0]) ? node2073 : node2066;
														assign node2066 = (inp[10]) ? 4'b0001 : node2067;
															assign node2067 = (inp[9]) ? 4'b0001 : node2068;
																assign node2068 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node2073 = (inp[4]) ? 4'b0101 : 4'b0011;
											assign node2076 = (inp[0]) ? node2100 : node2077;
												assign node2077 = (inp[15]) ? node2085 : node2078;
													assign node2078 = (inp[10]) ? node2082 : node2079;
														assign node2079 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node2082 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node2085 = (inp[3]) ? node2093 : node2086;
														assign node2086 = (inp[9]) ? 4'b0101 : node2087;
															assign node2087 = (inp[4]) ? 4'b0101 : node2088;
																assign node2088 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node2093 = (inp[4]) ? 4'b0011 : node2094;
															assign node2094 = (inp[10]) ? 4'b0001 : node2095;
																assign node2095 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node2100 = (inp[4]) ? node2112 : node2101;
													assign node2101 = (inp[9]) ? node2105 : node2102;
														assign node2102 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node2105 = (inp[10]) ? node2109 : node2106;
															assign node2106 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node2109 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node2112 = (inp[15]) ? node2120 : node2113;
														assign node2113 = (inp[9]) ? node2115 : 4'b0001;
															assign node2115 = (inp[3]) ? 4'b0111 : node2116;
																assign node2116 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node2120 = (inp[9]) ? node2124 : node2121;
															assign node2121 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node2124 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node2127 = (inp[10]) ? node2181 : node2128;
											assign node2128 = (inp[12]) ? node2160 : node2129;
												assign node2129 = (inp[4]) ? node2141 : node2130;
													assign node2130 = (inp[9]) ? node2134 : node2131;
														assign node2131 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node2134 = (inp[0]) ? node2138 : node2135;
															assign node2135 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node2138 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node2141 = (inp[9]) ? node2149 : node2142;
														assign node2142 = (inp[0]) ? node2146 : node2143;
															assign node2143 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node2146 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node2149 = (inp[3]) ? node2155 : node2150;
															assign node2150 = (inp[0]) ? node2152 : 4'b1111;
																assign node2152 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node2155 = (inp[15]) ? 4'b1101 : node2156;
																assign node2156 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node2160 = (inp[0]) ? node2174 : node2161;
													assign node2161 = (inp[3]) ? node2165 : node2162;
														assign node2162 = (inp[15]) ? 4'b1101 : 4'b1011;
														assign node2165 = (inp[15]) ? node2171 : node2166;
															assign node2166 = (inp[9]) ? node2168 : 4'b1011;
																assign node2168 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node2171 = (inp[9]) ? 4'b1011 : 4'b1001;
													assign node2174 = (inp[9]) ? node2178 : node2175;
														assign node2175 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node2178 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node2181 = (inp[0]) ? node2209 : node2182;
												assign node2182 = (inp[3]) ? node2200 : node2183;
													assign node2183 = (inp[15]) ? node2191 : node2184;
														assign node2184 = (inp[9]) ? node2188 : node2185;
															assign node2185 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node2188 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node2191 = (inp[12]) ? node2193 : 4'b1001;
															assign node2193 = (inp[4]) ? node2197 : node2194;
																assign node2194 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node2197 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node2200 = (inp[15]) ? 4'b1111 : node2201;
														assign node2201 = (inp[4]) ? node2205 : node2202;
															assign node2202 = (inp[12]) ? 4'b1011 : 4'b1101;
															assign node2205 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node2209 = (inp[4]) ? node2219 : node2210;
													assign node2210 = (inp[9]) ? node2214 : node2211;
														assign node2211 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node2214 = (inp[3]) ? node2216 : 4'b1111;
															assign node2216 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node2219 = (inp[9]) ? 4'b1011 : node2220;
														assign node2220 = (inp[3]) ? 4'b1111 : node2221;
															assign node2221 = (inp[15]) ? 4'b1111 : 4'b1101;
							assign node2226 = (inp[13]) ? node2600 : node2227;
								assign node2227 = (inp[8]) ? node2417 : node2228;
									assign node2228 = (inp[2]) ? node2304 : node2229;
										assign node2229 = (inp[0]) ? node2263 : node2230;
											assign node2230 = (inp[15]) ? node2246 : node2231;
												assign node2231 = (inp[4]) ? node2241 : node2232;
													assign node2232 = (inp[12]) ? node2234 : 4'b0011;
														assign node2234 = (inp[10]) ? node2238 : node2235;
															assign node2235 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node2238 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node2241 = (inp[9]) ? node2243 : 4'b0011;
														assign node2243 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node2246 = (inp[9]) ? node2258 : node2247;
													assign node2247 = (inp[4]) ? node2253 : node2248;
														assign node2248 = (inp[12]) ? node2250 : 4'b0101;
															assign node2250 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node2253 = (inp[12]) ? node2255 : 4'b0001;
															assign node2255 = (inp[3]) ? 4'b0001 : 4'b0101;
													assign node2258 = (inp[4]) ? node2260 : 4'b0001;
														assign node2260 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node2263 = (inp[15]) ? node2283 : node2264;
												assign node2264 = (inp[9]) ? node2270 : node2265;
													assign node2265 = (inp[4]) ? 4'b0001 : node2266;
														assign node2266 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node2270 = (inp[3]) ? node2276 : node2271;
														assign node2271 = (inp[4]) ? 4'b0101 : node2272;
															assign node2272 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node2276 = (inp[10]) ? node2278 : 4'b0111;
															assign node2278 = (inp[4]) ? node2280 : 4'b0111;
																assign node2280 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node2283 = (inp[9]) ? node2297 : node2284;
													assign node2284 = (inp[4]) ? node2290 : node2285;
														assign node2285 = (inp[10]) ? node2287 : 4'b0111;
															assign node2287 = (inp[3]) ? 4'b0111 : 4'b0011;
														assign node2290 = (inp[12]) ? node2292 : 4'b0011;
															assign node2292 = (inp[10]) ? node2294 : 4'b0011;
																assign node2294 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node2297 = (inp[4]) ? node2299 : 4'b0011;
														assign node2299 = (inp[12]) ? node2301 : 4'b0101;
															assign node2301 = (inp[3]) ? 4'b0001 : 4'b0011;
										assign node2304 = (inp[0]) ? node2354 : node2305;
											assign node2305 = (inp[15]) ? node2325 : node2306;
												assign node2306 = (inp[12]) ? node2316 : node2307;
													assign node2307 = (inp[4]) ? node2311 : node2308;
														assign node2308 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node2311 = (inp[9]) ? node2313 : 4'b0010;
															assign node2313 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node2316 = (inp[9]) ? 4'b0010 : node2317;
														assign node2317 = (inp[10]) ? node2321 : node2318;
															assign node2318 = (inp[3]) ? 4'b0010 : 4'b0110;
															assign node2321 = (inp[3]) ? 4'b0100 : 4'b0010;
												assign node2325 = (inp[10]) ? node2339 : node2326;
													assign node2326 = (inp[12]) ? node2332 : node2327;
														assign node2327 = (inp[4]) ? 4'b0000 : node2328;
															assign node2328 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node2332 = (inp[3]) ? 4'b0000 : node2333;
															assign node2333 = (inp[9]) ? node2335 : 4'b0000;
																assign node2335 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node2339 = (inp[3]) ? node2351 : node2340;
														assign node2340 = (inp[4]) ? node2346 : node2341;
															assign node2341 = (inp[12]) ? node2343 : 4'b0000;
																assign node2343 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node2346 = (inp[9]) ? node2348 : 4'b0100;
																assign node2348 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node2351 = (inp[9]) ? 4'b0110 : 4'b0000;
											assign node2354 = (inp[15]) ? node2380 : node2355;
												assign node2355 = (inp[3]) ? node2365 : node2356;
													assign node2356 = (inp[10]) ? node2358 : 4'b0000;
														assign node2358 = (inp[4]) ? 4'b0100 : node2359;
															assign node2359 = (inp[12]) ? node2361 : 4'b0000;
																assign node2361 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node2365 = (inp[4]) ? node2373 : node2366;
														assign node2366 = (inp[12]) ? node2370 : node2367;
															assign node2367 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node2370 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node2373 = (inp[9]) ? node2377 : node2374;
															assign node2374 = (inp[12]) ? 4'b0110 : 4'b0000;
															assign node2377 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node2380 = (inp[3]) ? node2400 : node2381;
													assign node2381 = (inp[12]) ? node2393 : node2382;
														assign node2382 = (inp[10]) ? node2388 : node2383;
															assign node2383 = (inp[4]) ? node2385 : 4'b0010;
																assign node2385 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node2388 = (inp[4]) ? node2390 : 4'b0110;
																assign node2390 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node2393 = (inp[10]) ? node2395 : 4'b0110;
															assign node2395 = (inp[9]) ? 4'b0010 : node2396;
																assign node2396 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node2400 = (inp[9]) ? node2410 : node2401;
														assign node2401 = (inp[4]) ? node2405 : node2402;
															assign node2402 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node2405 = (inp[12]) ? node2407 : 4'b0010;
																assign node2407 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node2410 = (inp[4]) ? node2412 : 4'b0010;
															assign node2412 = (inp[12]) ? node2414 : 4'b0100;
																assign node2414 = (inp[10]) ? 4'b0000 : 4'b0100;
									assign node2417 = (inp[2]) ? node2503 : node2418;
										assign node2418 = (inp[4]) ? node2456 : node2419;
											assign node2419 = (inp[15]) ? node2439 : node2420;
												assign node2420 = (inp[0]) ? node2432 : node2421;
													assign node2421 = (inp[10]) ? node2423 : 4'b0010;
														assign node2423 = (inp[3]) ? node2429 : node2424;
															assign node2424 = (inp[9]) ? node2426 : 4'b0110;
																assign node2426 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node2429 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node2432 = (inp[9]) ? node2434 : 4'b0100;
														assign node2434 = (inp[10]) ? node2436 : 4'b0000;
															assign node2436 = (inp[12]) ? 4'b0110 : 4'b0000;
												assign node2439 = (inp[0]) ? node2447 : node2440;
													assign node2440 = (inp[9]) ? node2442 : 4'b0100;
														assign node2442 = (inp[12]) ? node2444 : 4'b0000;
															assign node2444 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node2447 = (inp[9]) ? node2453 : node2448;
														assign node2448 = (inp[12]) ? node2450 : 4'b0110;
															assign node2450 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node2453 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node2456 = (inp[9]) ? node2482 : node2457;
												assign node2457 = (inp[12]) ? node2471 : node2458;
													assign node2458 = (inp[10]) ? node2466 : node2459;
														assign node2459 = (inp[3]) ? node2461 : 4'b0000;
															assign node2461 = (inp[15]) ? 4'b0010 : node2462;
																assign node2462 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node2466 = (inp[15]) ? node2468 : 4'b0010;
															assign node2468 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node2471 = (inp[10]) ? node2475 : node2472;
														assign node2472 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node2475 = (inp[15]) ? 4'b0110 : node2476;
															assign node2476 = (inp[3]) ? 4'b0100 : node2477;
																assign node2477 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node2482 = (inp[10]) ? node2492 : node2483;
													assign node2483 = (inp[3]) ? node2485 : 4'b0100;
														assign node2485 = (inp[15]) ? node2489 : node2486;
															assign node2486 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node2489 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node2492 = (inp[12]) ? node2496 : node2493;
														assign node2493 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node2496 = (inp[0]) ? node2498 : 4'b0000;
															assign node2498 = (inp[15]) ? node2500 : 4'b0010;
																assign node2500 = (inp[3]) ? 4'b0000 : 4'b0010;
										assign node2503 = (inp[0]) ? node2557 : node2504;
											assign node2504 = (inp[15]) ? node2524 : node2505;
												assign node2505 = (inp[3]) ? node2515 : node2506;
													assign node2506 = (inp[10]) ? node2510 : node2507;
														assign node2507 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node2510 = (inp[4]) ? 4'b1011 : node2511;
															assign node2511 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node2515 = (inp[10]) ? node2517 : 4'b1011;
														assign node2517 = (inp[9]) ? node2521 : node2518;
															assign node2518 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node2521 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node2524 = (inp[12]) ? node2550 : node2525;
													assign node2525 = (inp[3]) ? node2537 : node2526;
														assign node2526 = (inp[10]) ? node2532 : node2527;
															assign node2527 = (inp[4]) ? 4'b1101 : node2528;
																assign node2528 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node2532 = (inp[4]) ? 4'b1001 : node2533;
																assign node2533 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node2537 = (inp[10]) ? node2545 : node2538;
															assign node2538 = (inp[4]) ? node2542 : node2539;
																assign node2539 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node2542 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node2545 = (inp[9]) ? node2547 : 4'b1111;
																assign node2547 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node2550 = (inp[10]) ? 4'b1001 : node2551;
														assign node2551 = (inp[9]) ? 4'b1001 : node2552;
															assign node2552 = (inp[3]) ? 4'b1001 : 4'b1101;
											assign node2557 = (inp[15]) ? node2581 : node2558;
												assign node2558 = (inp[3]) ? node2568 : node2559;
													assign node2559 = (inp[9]) ? node2561 : 4'b1101;
														assign node2561 = (inp[12]) ? 4'b1001 : node2562;
															assign node2562 = (inp[4]) ? node2564 : 4'b1001;
																assign node2564 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node2568 = (inp[12]) ? node2576 : node2569;
														assign node2569 = (inp[9]) ? node2571 : 4'b1001;
															assign node2571 = (inp[4]) ? node2573 : 4'b1001;
																assign node2573 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node2576 = (inp[9]) ? node2578 : 4'b1111;
															assign node2578 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node2581 = (inp[3]) ? node2595 : node2582;
													assign node2582 = (inp[12]) ? node2590 : node2583;
														assign node2583 = (inp[10]) ? 4'b1011 : node2584;
															assign node2584 = (inp[4]) ? node2586 : 4'b1011;
																assign node2586 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node2590 = (inp[9]) ? node2592 : 4'b1111;
															assign node2592 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node2595 = (inp[10]) ? 4'b1001 : node2596;
														assign node2596 = (inp[9]) ? 4'b1101 : 4'b1111;
								assign node2600 = (inp[2]) ? node2816 : node2601;
									assign node2601 = (inp[8]) ? node2737 : node2602;
										assign node2602 = (inp[12]) ? node2670 : node2603;
											assign node2603 = (inp[4]) ? node2629 : node2604;
												assign node2604 = (inp[10]) ? node2612 : node2605;
													assign node2605 = (inp[9]) ? node2607 : 4'b1101;
														assign node2607 = (inp[15]) ? 4'b1001 : node2608;
															assign node2608 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node2612 = (inp[9]) ? node2620 : node2613;
														assign node2613 = (inp[15]) ? node2617 : node2614;
															assign node2614 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node2617 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node2620 = (inp[0]) ? 4'b1111 : node2621;
															assign node2621 = (inp[15]) ? node2625 : node2622;
																assign node2622 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node2625 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node2629 = (inp[3]) ? node2645 : node2630;
													assign node2630 = (inp[15]) ? node2638 : node2631;
														assign node2631 = (inp[10]) ? node2635 : node2632;
															assign node2632 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node2635 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node2638 = (inp[0]) ? node2640 : 4'b1001;
															assign node2640 = (inp[9]) ? 4'b1011 : node2641;
																assign node2641 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node2645 = (inp[15]) ? node2661 : node2646;
														assign node2646 = (inp[0]) ? node2654 : node2647;
															assign node2647 = (inp[9]) ? node2651 : node2648;
																assign node2648 = (inp[10]) ? 4'b1101 : 4'b1011;
																assign node2651 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node2654 = (inp[9]) ? node2658 : node2655;
																assign node2655 = (inp[10]) ? 4'b1111 : 4'b1001;
																assign node2658 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node2661 = (inp[0]) ? node2667 : node2662;
															assign node2662 = (inp[9]) ? 4'b1111 : node2663;
																assign node2663 = (inp[10]) ? 4'b1111 : 4'b1001;
															assign node2667 = (inp[9]) ? 4'b1001 : 4'b1101;
											assign node2670 = (inp[10]) ? node2712 : node2671;
												assign node2671 = (inp[3]) ? node2687 : node2672;
													assign node2672 = (inp[4]) ? node2680 : node2673;
														assign node2673 = (inp[9]) ? node2675 : 4'b1011;
															assign node2675 = (inp[15]) ? 4'b1111 : node2676;
																assign node2676 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node2680 = (inp[0]) ? node2684 : node2681;
															assign node2681 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node2684 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node2687 = (inp[9]) ? node2701 : node2688;
														assign node2688 = (inp[4]) ? node2696 : node2689;
															assign node2689 = (inp[15]) ? node2693 : node2690;
																assign node2690 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node2693 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node2696 = (inp[0]) ? node2698 : 4'b1101;
																assign node2698 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node2701 = (inp[4]) ? node2709 : node2702;
															assign node2702 = (inp[0]) ? node2706 : node2703;
																assign node2703 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node2706 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node2709 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node2712 = (inp[9]) ? node2726 : node2713;
													assign node2713 = (inp[4]) ? node2717 : node2714;
														assign node2714 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node2717 = (inp[0]) ? 4'b1101 : node2718;
															assign node2718 = (inp[3]) ? node2722 : node2719;
																assign node2719 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node2722 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node2726 = (inp[4]) ? node2730 : node2727;
														assign node2727 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node2730 = (inp[0]) ? 4'b1011 : node2731;
															assign node2731 = (inp[15]) ? 4'b1001 : node2732;
																assign node2732 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node2737 = (inp[12]) ? node2771 : node2738;
											assign node2738 = (inp[4]) ? node2760 : node2739;
												assign node2739 = (inp[0]) ? node2753 : node2740;
													assign node2740 = (inp[15]) ? node2750 : node2741;
														assign node2741 = (inp[9]) ? node2745 : node2742;
															assign node2742 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node2745 = (inp[10]) ? node2747 : 4'b1010;
																assign node2747 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node2750 = (inp[3]) ? 4'b1000 : 4'b1100;
													assign node2753 = (inp[15]) ? node2755 : 4'b1000;
														assign node2755 = (inp[9]) ? 4'b1010 : node2756;
															assign node2756 = (inp[10]) ? 4'b1010 : 4'b1110;
												assign node2760 = (inp[15]) ? 4'b1000 : node2761;
													assign node2761 = (inp[10]) ? node2765 : node2762;
														assign node2762 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node2765 = (inp[0]) ? 4'b1110 : node2766;
															assign node2766 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node2771 = (inp[0]) ? node2793 : node2772;
												assign node2772 = (inp[3]) ? node2780 : node2773;
													assign node2773 = (inp[15]) ? node2775 : 4'b1010;
														assign node2775 = (inp[10]) ? 4'b1000 : node2776;
															assign node2776 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node2780 = (inp[15]) ? node2786 : node2781;
														assign node2781 = (inp[4]) ? node2783 : 4'b1100;
															assign node2783 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node2786 = (inp[9]) ? node2790 : node2787;
															assign node2787 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node2790 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node2793 = (inp[10]) ? node2809 : node2794;
													assign node2794 = (inp[9]) ? node2806 : node2795;
														assign node2795 = (inp[4]) ? node2799 : node2796;
															assign node2796 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node2799 = (inp[15]) ? node2803 : node2800;
																assign node2800 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node2803 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node2806 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node2809 = (inp[4]) ? node2813 : node2810;
														assign node2810 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node2813 = (inp[15]) ? 4'b1110 : 4'b1100;
									assign node2816 = (inp[8]) ? node2910 : node2817;
										assign node2817 = (inp[15]) ? node2877 : node2818;
											assign node2818 = (inp[0]) ? node2844 : node2819;
												assign node2819 = (inp[3]) ? node2835 : node2820;
													assign node2820 = (inp[10]) ? node2828 : node2821;
														assign node2821 = (inp[12]) ? 4'b1110 : node2822;
															assign node2822 = (inp[4]) ? 4'b1010 : node2823;
																assign node2823 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node2828 = (inp[12]) ? 4'b1010 : node2829;
															assign node2829 = (inp[9]) ? 4'b1110 : node2830;
																assign node2830 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node2835 = (inp[9]) ? node2841 : node2836;
														assign node2836 = (inp[4]) ? 4'b1100 : node2837;
															assign node2837 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node2841 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node2844 = (inp[3]) ? node2856 : node2845;
													assign node2845 = (inp[4]) ? node2847 : 4'b1000;
														assign node2847 = (inp[10]) ? 4'b1000 : node2848;
															assign node2848 = (inp[12]) ? node2852 : node2849;
																assign node2849 = (inp[9]) ? 4'b1100 : 4'b1000;
																assign node2852 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node2856 = (inp[4]) ? node2866 : node2857;
														assign node2857 = (inp[9]) ? node2863 : node2858;
															assign node2858 = (inp[12]) ? 4'b1000 : node2859;
																assign node2859 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node2863 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node2866 = (inp[9]) ? node2872 : node2867;
															assign node2867 = (inp[12]) ? 4'b1110 : node2868;
																assign node2868 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node2872 = (inp[10]) ? 4'b1010 : node2873;
																assign node2873 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node2877 = (inp[0]) ? node2895 : node2878;
												assign node2878 = (inp[3]) ? node2888 : node2879;
													assign node2879 = (inp[10]) ? node2881 : 4'b1100;
														assign node2881 = (inp[12]) ? 4'b1000 : node2882;
															assign node2882 = (inp[4]) ? node2884 : 4'b1100;
																assign node2884 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node2888 = (inp[4]) ? 4'b1110 : node2889;
														assign node2889 = (inp[12]) ? 4'b1110 : node2890;
															assign node2890 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node2895 = (inp[3]) ? node2903 : node2896;
													assign node2896 = (inp[12]) ? node2898 : 4'b1110;
														assign node2898 = (inp[9]) ? 4'b1010 : node2899;
															assign node2899 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node2903 = (inp[4]) ? node2907 : node2904;
														assign node2904 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node2907 = (inp[9]) ? 4'b1000 : 4'b1100;
										assign node2910 = (inp[4]) ? node2956 : node2911;
											assign node2911 = (inp[9]) ? node2933 : node2912;
												assign node2912 = (inp[12]) ? node2922 : node2913;
													assign node2913 = (inp[10]) ? node2919 : node2914;
														assign node2914 = (inp[15]) ? 4'b1111 : node2915;
															assign node2915 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node2919 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node2922 = (inp[3]) ? node2928 : node2923;
														assign node2923 = (inp[0]) ? node2925 : 4'b1001;
															assign node2925 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node2928 = (inp[10]) ? 4'b1011 : node2929;
															assign node2929 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node2933 = (inp[10]) ? node2945 : node2934;
													assign node2934 = (inp[12]) ? node2942 : node2935;
														assign node2935 = (inp[0]) ? node2939 : node2936;
															assign node2936 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node2939 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node2942 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node2945 = (inp[3]) ? node2951 : node2946;
														assign node2946 = (inp[15]) ? node2948 : 4'b1111;
															assign node2948 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node2951 = (inp[15]) ? node2953 : 4'b1101;
															assign node2953 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node2956 = (inp[9]) ? node2978 : node2957;
												assign node2957 = (inp[12]) ? node2965 : node2958;
													assign node2958 = (inp[10]) ? node2960 : 4'b1001;
														assign node2960 = (inp[0]) ? node2962 : 4'b1101;
															assign node2962 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node2965 = (inp[0]) ? node2973 : node2966;
														assign node2966 = (inp[15]) ? node2970 : node2967;
															assign node2967 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node2970 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node2973 = (inp[3]) ? 4'b1101 : node2974;
															assign node2974 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node2978 = (inp[12]) ? node2994 : node2979;
													assign node2979 = (inp[10]) ? node2987 : node2980;
														assign node2980 = (inp[3]) ? node2982 : 4'b1101;
															assign node2982 = (inp[0]) ? node2984 : 4'b1111;
																assign node2984 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node2987 = (inp[15]) ? node2991 : node2988;
															assign node2988 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node2991 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node2994 = (inp[15]) ? node2996 : 4'b1001;
														assign node2996 = (inp[3]) ? 4'b1001 : 4'b1011;
					assign node2999 = (inp[6]) ? node4523 : node3000;
						assign node3000 = (inp[1]) ? node3818 : node3001;
							assign node3001 = (inp[13]) ? node3443 : node3002;
								assign node3002 = (inp[0]) ? node3216 : node3003;
									assign node3003 = (inp[15]) ? node3113 : node3004;
										assign node3004 = (inp[3]) ? node3058 : node3005;
											assign node3005 = (inp[12]) ? node3029 : node3006;
												assign node3006 = (inp[10]) ? node3020 : node3007;
													assign node3007 = (inp[4]) ? node3015 : node3008;
														assign node3008 = (inp[9]) ? 4'b1011 : node3009;
															assign node3009 = (inp[8]) ? 4'b1111 : node3010;
																assign node3010 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node3015 = (inp[8]) ? 4'b1110 : node3016;
															assign node3016 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node3020 = (inp[4]) ? node3024 : node3021;
														assign node3021 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node3024 = (inp[2]) ? node3026 : 4'b1011;
															assign node3026 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node3029 = (inp[8]) ? node3047 : node3030;
													assign node3030 = (inp[2]) ? node3032 : 4'b1010;
														assign node3032 = (inp[9]) ? node3040 : node3033;
															assign node3033 = (inp[10]) ? node3037 : node3034;
																assign node3034 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node3037 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node3040 = (inp[4]) ? node3044 : node3041;
																assign node3041 = (inp[10]) ? 4'b1111 : 4'b1011;
																assign node3044 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node3047 = (inp[2]) ? node3053 : node3048;
														assign node3048 = (inp[4]) ? node3050 : 4'b1111;
															assign node3050 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node3053 = (inp[10]) ? node3055 : 4'b1110;
															assign node3055 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node3058 = (inp[9]) ? node3090 : node3059;
												assign node3059 = (inp[4]) ? node3073 : node3060;
													assign node3060 = (inp[10]) ? node3066 : node3061;
														assign node3061 = (inp[8]) ? 4'b1110 : node3062;
															assign node3062 = (inp[12]) ? 4'b1111 : 4'b1110;
														assign node3066 = (inp[12]) ? node3068 : 4'b1110;
															assign node3068 = (inp[2]) ? 4'b1010 : node3069;
																assign node3069 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node3073 = (inp[10]) ? node3083 : node3074;
														assign node3074 = (inp[12]) ? node3078 : node3075;
															assign node3075 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node3078 = (inp[8]) ? 4'b1010 : node3079;
																assign node3079 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node3083 = (inp[12]) ? node3087 : node3084;
															assign node3084 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node3087 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node3090 = (inp[4]) ? node3100 : node3091;
													assign node3091 = (inp[12]) ? node3097 : node3092;
														assign node3092 = (inp[2]) ? 4'b1010 : node3093;
															assign node3093 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node3097 = (inp[8]) ? 4'b1011 : 4'b1101;
													assign node3100 = (inp[12]) ? node3110 : node3101;
														assign node3101 = (inp[10]) ? node3107 : node3102;
															assign node3102 = (inp[8]) ? node3104 : 4'b1101;
																assign node3104 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node3107 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node3110 = (inp[10]) ? 4'b1001 : 4'b1101;
										assign node3113 = (inp[3]) ? node3177 : node3114;
											assign node3114 = (inp[4]) ? node3148 : node3115;
												assign node3115 = (inp[9]) ? node3127 : node3116;
													assign node3116 = (inp[12]) ? node3124 : node3117;
														assign node3117 = (inp[10]) ? node3119 : 4'b1101;
															assign node3119 = (inp[2]) ? node3121 : 4'b1100;
																assign node3121 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node3124 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node3127 = (inp[12]) ? node3137 : node3128;
														assign node3128 = (inp[10]) ? node3130 : 4'b1000;
															assign node3130 = (inp[8]) ? node3134 : node3131;
																assign node3131 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node3134 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node3137 = (inp[10]) ? node3143 : node3138;
															assign node3138 = (inp[2]) ? node3140 : 4'b1001;
																assign node3140 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node3143 = (inp[2]) ? node3145 : 4'b1100;
																assign node3145 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node3148 = (inp[9]) ? node3160 : node3149;
													assign node3149 = (inp[10]) ? node3155 : node3150;
														assign node3150 = (inp[8]) ? node3152 : 4'b1001;
															assign node3152 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node3155 = (inp[12]) ? node3157 : 4'b1000;
															assign node3157 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node3160 = (inp[10]) ? node3168 : node3161;
														assign node3161 = (inp[2]) ? node3165 : node3162;
															assign node3162 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node3165 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node3168 = (inp[12]) ? node3170 : 4'b1101;
															assign node3170 = (inp[8]) ? node3174 : node3171;
																assign node3171 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node3174 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node3177 = (inp[9]) ? node3191 : node3178;
												assign node3178 = (inp[8]) ? node3184 : node3179;
													assign node3179 = (inp[2]) ? 4'b1001 : node3180;
														assign node3180 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node3184 = (inp[2]) ? node3188 : node3185;
														assign node3185 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node3188 = (inp[4]) ? 4'b1110 : 4'b1100;
												assign node3191 = (inp[4]) ? node3203 : node3192;
													assign node3192 = (inp[8]) ? node3196 : node3193;
														assign node3193 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node3196 = (inp[2]) ? 4'b1000 : node3197;
															assign node3197 = (inp[12]) ? node3199 : 4'b1001;
																assign node3199 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node3203 = (inp[12]) ? node3209 : node3204;
														assign node3204 = (inp[2]) ? 4'b1110 : node3205;
															assign node3205 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node3209 = (inp[10]) ? node3211 : 4'b1110;
															assign node3211 = (inp[2]) ? node3213 : 4'b1011;
																assign node3213 = (inp[8]) ? 4'b1010 : 4'b1011;
									assign node3216 = (inp[15]) ? node3316 : node3217;
										assign node3217 = (inp[3]) ? node3259 : node3218;
											assign node3218 = (inp[10]) ? node3236 : node3219;
												assign node3219 = (inp[4]) ? node3227 : node3220;
													assign node3220 = (inp[9]) ? 4'b1001 : node3221;
														assign node3221 = (inp[12]) ? node3223 : 4'b1101;
															assign node3223 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node3227 = (inp[9]) ? node3229 : 4'b1000;
														assign node3229 = (inp[8]) ? node3233 : node3230;
															assign node3230 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node3233 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node3236 = (inp[4]) ? node3248 : node3237;
													assign node3237 = (inp[9]) ? node3243 : node3238;
														assign node3238 = (inp[12]) ? 4'b1001 : node3239;
															assign node3239 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node3243 = (inp[12]) ? 4'b1100 : node3244;
															assign node3244 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node3248 = (inp[2]) ? node3252 : node3249;
														assign node3249 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node3252 = (inp[8]) ? node3256 : node3253;
															assign node3253 = (inp[12]) ? 4'b1101 : 4'b1001;
															assign node3256 = (inp[12]) ? 4'b1100 : 4'b1000;
											assign node3259 = (inp[9]) ? node3285 : node3260;
												assign node3260 = (inp[4]) ? node3272 : node3261;
													assign node3261 = (inp[2]) ? node3267 : node3262;
														assign node3262 = (inp[10]) ? node3264 : 4'b1100;
															assign node3264 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node3267 = (inp[8]) ? 4'b1100 : node3268;
															assign node3268 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node3272 = (inp[10]) ? node3280 : node3273;
														assign node3273 = (inp[8]) ? node3277 : node3274;
															assign node3274 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node3277 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node3280 = (inp[12]) ? 4'b1111 : node3281;
															assign node3281 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node3285 = (inp[4]) ? node3301 : node3286;
													assign node3286 = (inp[10]) ? node3294 : node3287;
														assign node3287 = (inp[2]) ? node3291 : node3288;
															assign node3288 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node3291 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node3294 = (inp[12]) ? node3296 : 4'b1001;
															assign node3296 = (inp[8]) ? 4'b1111 : node3297;
																assign node3297 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node3301 = (inp[12]) ? node3309 : node3302;
														assign node3302 = (inp[2]) ? node3306 : node3303;
															assign node3303 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node3306 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node3309 = (inp[10]) ? node3311 : 4'b1110;
															assign node3311 = (inp[8]) ? 4'b1011 : node3312;
																assign node3312 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node3316 = (inp[3]) ? node3378 : node3317;
											assign node3317 = (inp[2]) ? node3353 : node3318;
												assign node3318 = (inp[8]) ? node3340 : node3319;
													assign node3319 = (inp[12]) ? node3333 : node3320;
														assign node3320 = (inp[10]) ? node3328 : node3321;
															assign node3321 = (inp[4]) ? node3325 : node3322;
																assign node3322 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node3325 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node3328 = (inp[9]) ? 4'b1110 : node3329;
																assign node3329 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node3333 = (inp[10]) ? node3335 : 4'b1110;
															assign node3335 = (inp[9]) ? node3337 : 4'b1110;
																assign node3337 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node3340 = (inp[10]) ? node3346 : node3341;
														assign node3341 = (inp[4]) ? 4'b1011 : node3342;
															assign node3342 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node3346 = (inp[9]) ? node3348 : 4'b1111;
															assign node3348 = (inp[12]) ? 4'b1111 : node3349;
																assign node3349 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node3353 = (inp[8]) ? node3369 : node3354;
													assign node3354 = (inp[12]) ? node3362 : node3355;
														assign node3355 = (inp[4]) ? node3359 : node3356;
															assign node3356 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node3359 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node3362 = (inp[4]) ? 4'b1011 : node3363;
															assign node3363 = (inp[10]) ? node3365 : 4'b1011;
																assign node3365 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node3369 = (inp[12]) ? 4'b1010 : node3370;
														assign node3370 = (inp[9]) ? node3374 : node3371;
															assign node3371 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node3374 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node3378 = (inp[4]) ? node3416 : node3379;
												assign node3379 = (inp[9]) ? node3405 : node3380;
													assign node3380 = (inp[10]) ? node3390 : node3381;
														assign node3381 = (inp[12]) ? node3383 : 4'b1110;
															assign node3383 = (inp[8]) ? node3387 : node3384;
																assign node3384 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node3387 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node3390 = (inp[12]) ? node3398 : node3391;
															assign node3391 = (inp[8]) ? node3395 : node3392;
																assign node3392 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node3395 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node3398 = (inp[8]) ? node3402 : node3399;
																assign node3399 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node3402 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node3405 = (inp[12]) ? node3411 : node3406;
														assign node3406 = (inp[2]) ? 4'b1011 : node3407;
															assign node3407 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node3411 = (inp[10]) ? node3413 : 4'b1010;
															assign node3413 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node3416 = (inp[9]) ? node3430 : node3417;
													assign node3417 = (inp[12]) ? node3423 : node3418;
														assign node3418 = (inp[2]) ? node3420 : 4'b1011;
															assign node3420 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node3423 = (inp[10]) ? node3425 : 4'b1011;
															assign node3425 = (inp[8]) ? node3427 : 4'b1101;
																assign node3427 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node3430 = (inp[12]) ? node3440 : node3431;
														assign node3431 = (inp[10]) ? 4'b1101 : node3432;
															assign node3432 = (inp[2]) ? node3436 : node3433;
																assign node3433 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node3436 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node3440 = (inp[2]) ? 4'b1101 : 4'b1000;
								assign node3443 = (inp[2]) ? node3641 : node3444;
									assign node3444 = (inp[8]) ? node3548 : node3445;
										assign node3445 = (inp[10]) ? node3481 : node3446;
											assign node3446 = (inp[4]) ? node3464 : node3447;
												assign node3447 = (inp[9]) ? node3455 : node3448;
													assign node3448 = (inp[15]) ? node3452 : node3449;
														assign node3449 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node3452 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node3455 = (inp[12]) ? 4'b1000 : node3456;
														assign node3456 = (inp[15]) ? node3460 : node3457;
															assign node3457 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node3460 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node3464 = (inp[9]) ? node3470 : node3465;
													assign node3465 = (inp[12]) ? node3467 : 4'b1000;
														assign node3467 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node3470 = (inp[3]) ? node3478 : node3471;
														assign node3471 = (inp[15]) ? node3475 : node3472;
															assign node3472 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node3475 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node3478 = (inp[12]) ? 4'b1110 : 4'b1100;
											assign node3481 = (inp[0]) ? node3511 : node3482;
												assign node3482 = (inp[15]) ? node3504 : node3483;
													assign node3483 = (inp[3]) ? node3495 : node3484;
														assign node3484 = (inp[9]) ? node3490 : node3485;
															assign node3485 = (inp[12]) ? node3487 : 4'b1110;
																assign node3487 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node3490 = (inp[12]) ? node3492 : 4'b1010;
																assign node3492 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node3495 = (inp[4]) ? 4'b1100 : node3496;
															assign node3496 = (inp[12]) ? node3500 : node3497;
																assign node3497 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node3500 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node3504 = (inp[4]) ? node3508 : node3505;
														assign node3505 = (inp[3]) ? 4'b1100 : 4'b1000;
														assign node3508 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node3511 = (inp[15]) ? node3523 : node3512;
													assign node3512 = (inp[3]) ? node3514 : 4'b1000;
														assign node3514 = (inp[12]) ? node3518 : node3515;
															assign node3515 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node3518 = (inp[9]) ? node3520 : 4'b1110;
																assign node3520 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node3523 = (inp[3]) ? node3539 : node3524;
														assign node3524 = (inp[4]) ? node3532 : node3525;
															assign node3525 = (inp[12]) ? node3529 : node3526;
																assign node3526 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node3529 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node3532 = (inp[12]) ? node3536 : node3533;
																assign node3533 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node3536 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node3539 = (inp[4]) ? node3545 : node3540;
															assign node3540 = (inp[12]) ? 4'b1010 : node3541;
																assign node3541 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node3545 = (inp[12]) ? 4'b1100 : 4'b1010;
										assign node3548 = (inp[9]) ? node3590 : node3549;
											assign node3549 = (inp[4]) ? node3567 : node3550;
												assign node3550 = (inp[12]) ? node3558 : node3551;
													assign node3551 = (inp[15]) ? node3555 : node3552;
														assign node3552 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node3555 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node3558 = (inp[10]) ? node3564 : node3559;
														assign node3559 = (inp[0]) ? node3561 : 4'b0101;
															assign node3561 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node3564 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node3567 = (inp[10]) ? node3585 : node3568;
													assign node3568 = (inp[3]) ? node3580 : node3569;
														assign node3569 = (inp[12]) ? node3575 : node3570;
															assign node3570 = (inp[0]) ? 4'b0001 : node3571;
																assign node3571 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node3575 = (inp[15]) ? node3577 : 4'b0011;
																assign node3577 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node3580 = (inp[0]) ? node3582 : 4'b0011;
															assign node3582 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node3585 = (inp[12]) ? 4'b0111 : node3586;
														assign node3586 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node3590 = (inp[4]) ? node3618 : node3591;
												assign node3591 = (inp[12]) ? node3603 : node3592;
													assign node3592 = (inp[3]) ? node3598 : node3593;
														assign node3593 = (inp[15]) ? node3595 : 4'b0011;
															assign node3595 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node3598 = (inp[0]) ? 4'b0001 : node3599;
															assign node3599 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node3603 = (inp[10]) ? node3611 : node3604;
														assign node3604 = (inp[3]) ? node3606 : 4'b0001;
															assign node3606 = (inp[15]) ? node3608 : 4'b0001;
																assign node3608 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node3611 = (inp[0]) ? 4'b0111 : node3612;
															assign node3612 = (inp[15]) ? 4'b0101 : node3613;
																assign node3613 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node3618 = (inp[15]) ? node3632 : node3619;
													assign node3619 = (inp[12]) ? node3627 : node3620;
														assign node3620 = (inp[0]) ? node3624 : node3621;
															assign node3621 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node3624 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node3627 = (inp[10]) ? node3629 : 4'b0101;
															assign node3629 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node3632 = (inp[10]) ? 4'b0111 : node3633;
														assign node3633 = (inp[12]) ? node3637 : node3634;
															assign node3634 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node3637 = (inp[3]) ? 4'b0101 : 4'b0111;
									assign node3641 = (inp[8]) ? node3739 : node3642;
										assign node3642 = (inp[12]) ? node3680 : node3643;
											assign node3643 = (inp[0]) ? node3661 : node3644;
												assign node3644 = (inp[15]) ? node3652 : node3645;
													assign node3645 = (inp[3]) ? node3647 : 4'b0111;
														assign node3647 = (inp[4]) ? 4'b0101 : node3648;
															assign node3648 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node3652 = (inp[3]) ? 4'b0101 : node3653;
														assign node3653 = (inp[9]) ? node3657 : node3654;
															assign node3654 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node3657 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node3661 = (inp[15]) ? node3671 : node3662;
													assign node3662 = (inp[4]) ? node3666 : node3663;
														assign node3663 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node3666 = (inp[9]) ? node3668 : 4'b0001;
															assign node3668 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node3671 = (inp[9]) ? node3675 : node3672;
														assign node3672 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node3675 = (inp[4]) ? node3677 : 4'b0011;
															assign node3677 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node3680 = (inp[0]) ? node3704 : node3681;
												assign node3681 = (inp[15]) ? node3695 : node3682;
													assign node3682 = (inp[4]) ? node3688 : node3683;
														assign node3683 = (inp[3]) ? 4'b0011 : node3684;
															assign node3684 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node3688 = (inp[3]) ? 4'b0101 : node3689;
															assign node3689 = (inp[9]) ? 4'b0111 : node3690;
																assign node3690 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node3695 = (inp[4]) ? node3701 : node3696;
														assign node3696 = (inp[9]) ? node3698 : 4'b0101;
															assign node3698 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node3701 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node3704 = (inp[15]) ? node3718 : node3705;
													assign node3705 = (inp[3]) ? node3715 : node3706;
														assign node3706 = (inp[9]) ? 4'b0101 : node3707;
															assign node3707 = (inp[10]) ? node3711 : node3708;
																assign node3708 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node3711 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node3715 = (inp[10]) ? 4'b0111 : 4'b0101;
													assign node3718 = (inp[3]) ? node3730 : node3719;
														assign node3719 = (inp[4]) ? node3725 : node3720;
															assign node3720 = (inp[9]) ? node3722 : 4'b0111;
																assign node3722 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node3725 = (inp[9]) ? node3727 : 4'b0011;
																assign node3727 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node3730 = (inp[10]) ? 4'b0101 : node3731;
															assign node3731 = (inp[9]) ? node3735 : node3732;
																assign node3732 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node3735 = (inp[4]) ? 4'b0101 : 4'b0011;
										assign node3739 = (inp[15]) ? node3789 : node3740;
											assign node3740 = (inp[0]) ? node3766 : node3741;
												assign node3741 = (inp[4]) ? node3753 : node3742;
													assign node3742 = (inp[9]) ? node3748 : node3743;
														assign node3743 = (inp[12]) ? node3745 : 4'b0110;
															assign node3745 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node3748 = (inp[3]) ? 4'b0010 : node3749;
															assign node3749 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node3753 = (inp[9]) ? node3759 : node3754;
														assign node3754 = (inp[10]) ? node3756 : 4'b0010;
															assign node3756 = (inp[3]) ? 4'b0100 : 4'b0010;
														assign node3759 = (inp[3]) ? 4'b0100 : node3760;
															assign node3760 = (inp[12]) ? node3762 : 4'b0110;
																assign node3762 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node3766 = (inp[3]) ? node3782 : node3767;
													assign node3767 = (inp[10]) ? node3773 : node3768;
														assign node3768 = (inp[9]) ? node3770 : 4'b0000;
															assign node3770 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node3773 = (inp[4]) ? node3775 : 4'b0100;
															assign node3775 = (inp[12]) ? node3779 : node3776;
																assign node3776 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node3779 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node3782 = (inp[12]) ? 4'b0110 : node3783;
														assign node3783 = (inp[9]) ? 4'b0110 : node3784;
															assign node3784 = (inp[4]) ? 4'b0000 : 4'b0100;
											assign node3789 = (inp[0]) ? node3807 : node3790;
												assign node3790 = (inp[9]) ? node3800 : node3791;
													assign node3791 = (inp[4]) ? node3795 : node3792;
														assign node3792 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node3795 = (inp[10]) ? node3797 : 4'b0000;
															assign node3797 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node3800 = (inp[4]) ? 4'b0110 : node3801;
														assign node3801 = (inp[10]) ? node3803 : 4'b0000;
															assign node3803 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node3807 = (inp[12]) ? node3809 : 4'b0010;
													assign node3809 = (inp[4]) ? 4'b0100 : node3810;
														assign node3810 = (inp[3]) ? node3812 : 4'b0110;
															assign node3812 = (inp[10]) ? node3814 : 4'b0010;
																assign node3814 = (inp[9]) ? 4'b0100 : 4'b0010;
							assign node3818 = (inp[13]) ? node4178 : node3819;
								assign node3819 = (inp[2]) ? node4005 : node3820;
									assign node3820 = (inp[8]) ? node3902 : node3821;
										assign node3821 = (inp[9]) ? node3855 : node3822;
											assign node3822 = (inp[4]) ? node3836 : node3823;
												assign node3823 = (inp[10]) ? node3831 : node3824;
													assign node3824 = (inp[0]) ? node3828 : node3825;
														assign node3825 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node3828 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node3831 = (inp[12]) ? 4'b1000 : node3832;
														assign node3832 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node3836 = (inp[10]) ? node3842 : node3837;
													assign node3837 = (inp[15]) ? 4'b1000 : node3838;
														assign node3838 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node3842 = (inp[12]) ? node3848 : node3843;
														assign node3843 = (inp[15]) ? node3845 : 4'b1000;
															assign node3845 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node3848 = (inp[0]) ? 4'b1110 : node3849;
															assign node3849 = (inp[15]) ? 4'b1110 : node3850;
																assign node3850 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node3855 = (inp[4]) ? node3877 : node3856;
												assign node3856 = (inp[12]) ? node3868 : node3857;
													assign node3857 = (inp[3]) ? node3859 : 4'b1010;
														assign node3859 = (inp[10]) ? node3863 : node3860;
															assign node3860 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node3863 = (inp[0]) ? 4'b1010 : node3864;
																assign node3864 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node3868 = (inp[10]) ? node3874 : node3869;
														assign node3869 = (inp[15]) ? 4'b1000 : node3870;
															assign node3870 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node3874 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node3877 = (inp[12]) ? node3889 : node3878;
													assign node3878 = (inp[3]) ? node3884 : node3879;
														assign node3879 = (inp[10]) ? node3881 : 4'b1100;
															assign node3881 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node3884 = (inp[0]) ? 4'b1110 : node3885;
															assign node3885 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node3889 = (inp[10]) ? node3897 : node3890;
														assign node3890 = (inp[0]) ? node3892 : 4'b1110;
															assign node3892 = (inp[3]) ? 4'b1110 : node3893;
																assign node3893 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node3897 = (inp[15]) ? 4'b1000 : node3898;
															assign node3898 = (inp[0]) ? 4'b1010 : 4'b1000;
										assign node3902 = (inp[10]) ? node3944 : node3903;
											assign node3903 = (inp[4]) ? node3927 : node3904;
												assign node3904 = (inp[9]) ? node3914 : node3905;
													assign node3905 = (inp[12]) ? 4'b0101 : node3906;
														assign node3906 = (inp[3]) ? node3908 : 4'b0111;
															assign node3908 = (inp[0]) ? 4'b0101 : node3909;
																assign node3909 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node3914 = (inp[3]) ? node3922 : node3915;
														assign node3915 = (inp[15]) ? node3919 : node3916;
															assign node3916 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node3919 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node3922 = (inp[15]) ? node3924 : 4'b0001;
															assign node3924 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node3927 = (inp[9]) ? node3935 : node3928;
													assign node3928 = (inp[0]) ? node3932 : node3929;
														assign node3929 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node3932 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node3935 = (inp[12]) ? 4'b0111 : node3936;
														assign node3936 = (inp[0]) ? 4'b0101 : node3937;
															assign node3937 = (inp[15]) ? node3939 : 4'b0111;
																assign node3939 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node3944 = (inp[0]) ? node3984 : node3945;
												assign node3945 = (inp[15]) ? node3969 : node3946;
													assign node3946 = (inp[3]) ? node3956 : node3947;
														assign node3947 = (inp[12]) ? node3949 : 4'b0111;
															assign node3949 = (inp[9]) ? node3953 : node3950;
																assign node3950 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node3953 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node3956 = (inp[9]) ? node3964 : node3957;
															assign node3957 = (inp[4]) ? node3961 : node3958;
																assign node3958 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node3961 = (inp[12]) ? 4'b0101 : 4'b0011;
															assign node3964 = (inp[4]) ? node3966 : 4'b0101;
																assign node3966 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node3969 = (inp[4]) ? node3979 : node3970;
														assign node3970 = (inp[3]) ? node3976 : node3971;
															assign node3971 = (inp[12]) ? 4'b0101 : node3972;
																assign node3972 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node3976 = (inp[9]) ? 4'b0111 : 4'b0101;
														assign node3979 = (inp[9]) ? node3981 : 4'b0001;
															assign node3981 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node3984 = (inp[3]) ? node3992 : node3985;
													assign node3985 = (inp[12]) ? node3987 : 4'b0101;
														assign node3987 = (inp[4]) ? node3989 : 4'b0001;
															assign node3989 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node3992 = (inp[12]) ? node4002 : node3993;
														assign node3993 = (inp[15]) ? node3999 : node3994;
															assign node3994 = (inp[9]) ? 4'b0111 : node3995;
																assign node3995 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node3999 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node4002 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node4005 = (inp[8]) ? node4099 : node4006;
										assign node4006 = (inp[15]) ? node4042 : node4007;
											assign node4007 = (inp[0]) ? node4025 : node4008;
												assign node4008 = (inp[9]) ? node4014 : node4009;
													assign node4009 = (inp[4]) ? 4'b0011 : node4010;
														assign node4010 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node4014 = (inp[12]) ? node4016 : 4'b0101;
														assign node4016 = (inp[4]) ? node4022 : node4017;
															assign node4017 = (inp[10]) ? node4019 : 4'b0011;
																assign node4019 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node4022 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node4025 = (inp[3]) ? node4031 : node4026;
													assign node4026 = (inp[4]) ? 4'b0101 : node4027;
														assign node4027 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node4031 = (inp[4]) ? node4037 : node4032;
														assign node4032 = (inp[9]) ? 4'b0001 : node4033;
															assign node4033 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node4037 = (inp[12]) ? node4039 : 4'b0001;
															assign node4039 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node4042 = (inp[0]) ? node4072 : node4043;
												assign node4043 = (inp[3]) ? node4057 : node4044;
													assign node4044 = (inp[10]) ? 4'b0101 : node4045;
														assign node4045 = (inp[12]) ? node4051 : node4046;
															assign node4046 = (inp[9]) ? 4'b0101 : node4047;
																assign node4047 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node4051 = (inp[4]) ? 4'b0001 : node4052;
																assign node4052 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node4057 = (inp[4]) ? node4067 : node4058;
														assign node4058 = (inp[9]) ? node4064 : node4059;
															assign node4059 = (inp[12]) ? node4061 : 4'b0101;
																assign node4061 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node4064 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node4067 = (inp[9]) ? 4'b0111 : node4068;
															assign node4068 = (inp[12]) ? 4'b0111 : 4'b0001;
												assign node4072 = (inp[3]) ? node4086 : node4073;
													assign node4073 = (inp[9]) ? node4081 : node4074;
														assign node4074 = (inp[4]) ? node4076 : 4'b0111;
															assign node4076 = (inp[10]) ? node4078 : 4'b0011;
																assign node4078 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node4081 = (inp[12]) ? node4083 : 4'b0011;
															assign node4083 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node4086 = (inp[4]) ? node4090 : node4087;
														assign node4087 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node4090 = (inp[12]) ? node4092 : 4'b0101;
															assign node4092 = (inp[10]) ? node4096 : node4093;
																assign node4093 = (inp[9]) ? 4'b0101 : 4'b0011;
																assign node4096 = (inp[9]) ? 4'b0001 : 4'b0101;
										assign node4099 = (inp[12]) ? node4139 : node4100;
											assign node4100 = (inp[15]) ? node4124 : node4101;
												assign node4101 = (inp[0]) ? node4109 : node4102;
													assign node4102 = (inp[4]) ? node4104 : 4'b0010;
														assign node4104 = (inp[10]) ? 4'b0100 : node4105;
															assign node4105 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node4109 = (inp[3]) ? node4119 : node4110;
														assign node4110 = (inp[10]) ? node4112 : 4'b0100;
															assign node4112 = (inp[4]) ? node4116 : node4113;
																assign node4113 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node4116 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node4119 = (inp[9]) ? 4'b0000 : node4120;
															assign node4120 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node4124 = (inp[0]) ? node4132 : node4125;
													assign node4125 = (inp[4]) ? node4129 : node4126;
														assign node4126 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node4129 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node4132 = (inp[4]) ? node4136 : node4133;
														assign node4133 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node4136 = (inp[9]) ? 4'b0100 : 4'b0010;
											assign node4139 = (inp[9]) ? node4161 : node4140;
												assign node4140 = (inp[3]) ? node4148 : node4141;
													assign node4141 = (inp[10]) ? 4'b0010 : node4142;
														assign node4142 = (inp[4]) ? node4144 : 4'b0100;
															assign node4144 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node4148 = (inp[4]) ? node4152 : node4149;
														assign node4149 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node4152 = (inp[10]) ? node4158 : node4153;
															assign node4153 = (inp[0]) ? node4155 : 4'b0000;
																assign node4155 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node4158 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node4161 = (inp[10]) ? node4173 : node4162;
													assign node4162 = (inp[4]) ? node4164 : 4'b0010;
														assign node4164 = (inp[3]) ? node4166 : 4'b0110;
															assign node4166 = (inp[15]) ? node4170 : node4167;
																assign node4167 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node4170 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node4173 = (inp[3]) ? node4175 : 4'b0100;
														assign node4175 = (inp[0]) ? 4'b0100 : 4'b0110;
								assign node4178 = (inp[2]) ? node4366 : node4179;
									assign node4179 = (inp[8]) ? node4277 : node4180;
										assign node4180 = (inp[10]) ? node4222 : node4181;
											assign node4181 = (inp[0]) ? node4203 : node4182;
												assign node4182 = (inp[15]) ? node4196 : node4183;
													assign node4183 = (inp[12]) ? node4191 : node4184;
														assign node4184 = (inp[9]) ? node4188 : node4185;
															assign node4185 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node4188 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node4191 = (inp[9]) ? node4193 : 4'b0010;
															assign node4193 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node4196 = (inp[3]) ? node4198 : 4'b0000;
														assign node4198 = (inp[4]) ? 4'b0110 : node4199;
															assign node4199 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node4203 = (inp[15]) ? node4219 : node4204;
													assign node4204 = (inp[3]) ? node4212 : node4205;
														assign node4205 = (inp[4]) ? node4209 : node4206;
															assign node4206 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node4209 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node4212 = (inp[9]) ? node4216 : node4213;
															assign node4213 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node4216 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node4219 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node4222 = (inp[3]) ? node4244 : node4223;
												assign node4223 = (inp[9]) ? node4233 : node4224;
													assign node4224 = (inp[12]) ? node4228 : node4225;
														assign node4225 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node4228 = (inp[0]) ? node4230 : 4'b0000;
															assign node4230 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node4233 = (inp[12]) ? node4241 : node4234;
														assign node4234 = (inp[4]) ? 4'b0100 : node4235;
															assign node4235 = (inp[0]) ? node4237 : 4'b0010;
																assign node4237 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node4241 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node4244 = (inp[4]) ? node4262 : node4245;
													assign node4245 = (inp[12]) ? node4253 : node4246;
														assign node4246 = (inp[9]) ? 4'b0000 : node4247;
															assign node4247 = (inp[0]) ? node4249 : 4'b0100;
																assign node4249 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node4253 = (inp[9]) ? node4259 : node4254;
															assign node4254 = (inp[0]) ? node4256 : 4'b0000;
																assign node4256 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node4259 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node4262 = (inp[12]) ? node4274 : node4263;
														assign node4263 = (inp[9]) ? node4269 : node4264;
															assign node4264 = (inp[0]) ? node4266 : 4'b0010;
																assign node4266 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node4269 = (inp[15]) ? node4271 : 4'b0100;
																assign node4271 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node4274 = (inp[9]) ? 4'b0010 : 4'b0110;
										assign node4277 = (inp[15]) ? node4321 : node4278;
											assign node4278 = (inp[0]) ? node4298 : node4279;
												assign node4279 = (inp[9]) ? node4287 : node4280;
													assign node4280 = (inp[4]) ? 4'b0011 : node4281;
														assign node4281 = (inp[10]) ? node4283 : 4'b0111;
															assign node4283 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node4287 = (inp[4]) ? node4293 : node4288;
														assign node4288 = (inp[12]) ? node4290 : 4'b0011;
															assign node4290 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node4293 = (inp[3]) ? 4'b0101 : node4294;
															assign node4294 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node4298 = (inp[4]) ? node4306 : node4299;
													assign node4299 = (inp[9]) ? 4'b0001 : node4300;
														assign node4300 = (inp[10]) ? node4302 : 4'b0101;
															assign node4302 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node4306 = (inp[3]) ? node4312 : node4307;
														assign node4307 = (inp[12]) ? 4'b0101 : node4308;
															assign node4308 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node4312 = (inp[12]) ? node4314 : 4'b0001;
															assign node4314 = (inp[9]) ? node4318 : node4315;
																assign node4315 = (inp[10]) ? 4'b0111 : 4'b0001;
																assign node4318 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node4321 = (inp[0]) ? node4343 : node4322;
												assign node4322 = (inp[3]) ? node4336 : node4323;
													assign node4323 = (inp[9]) ? node4331 : node4324;
														assign node4324 = (inp[4]) ? node4328 : node4325;
															assign node4325 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node4328 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node4331 = (inp[10]) ? 4'b0001 : node4332;
															assign node4332 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node4336 = (inp[9]) ? node4340 : node4337;
														assign node4337 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node4340 = (inp[4]) ? 4'b0111 : 4'b0001;
												assign node4343 = (inp[3]) ? node4353 : node4344;
													assign node4344 = (inp[9]) ? node4350 : node4345;
														assign node4345 = (inp[4]) ? 4'b0011 : node4346;
															assign node4346 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node4350 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node4353 = (inp[4]) ? node4357 : node4354;
														assign node4354 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node4357 = (inp[9]) ? node4361 : node4358;
															assign node4358 = (inp[12]) ? 4'b0101 : 4'b0011;
															assign node4361 = (inp[10]) ? node4363 : 4'b0101;
																assign node4363 = (inp[12]) ? 4'b0001 : 4'b0101;
									assign node4366 = (inp[8]) ? node4442 : node4367;
										assign node4367 = (inp[15]) ? node4409 : node4368;
											assign node4368 = (inp[0]) ? node4386 : node4369;
												assign node4369 = (inp[4]) ? node4375 : node4370;
													assign node4370 = (inp[9]) ? node4372 : 4'b0111;
														assign node4372 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node4375 = (inp[3]) ? node4381 : node4376;
														assign node4376 = (inp[12]) ? 4'b0011 : node4377;
															assign node4377 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node4381 = (inp[9]) ? 4'b0101 : node4382;
															assign node4382 = (inp[12]) ? 4'b0101 : 4'b0011;
												assign node4386 = (inp[3]) ? node4394 : node4387;
													assign node4387 = (inp[10]) ? 4'b0101 : node4388;
														assign node4388 = (inp[9]) ? node4390 : 4'b0101;
															assign node4390 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node4394 = (inp[9]) ? node4404 : node4395;
														assign node4395 = (inp[4]) ? node4401 : node4396;
															assign node4396 = (inp[10]) ? node4398 : 4'b0101;
																assign node4398 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node4401 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node4404 = (inp[10]) ? node4406 : 4'b0111;
															assign node4406 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node4409 = (inp[0]) ? node4425 : node4410;
												assign node4410 = (inp[3]) ? node4418 : node4411;
													assign node4411 = (inp[12]) ? 4'b0001 : node4412;
														assign node4412 = (inp[4]) ? 4'b0101 : node4413;
															assign node4413 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node4418 = (inp[9]) ? node4420 : 4'b0001;
														assign node4420 = (inp[10]) ? 4'b0111 : node4421;
															assign node4421 = (inp[4]) ? 4'b0111 : 4'b0001;
												assign node4425 = (inp[4]) ? node4433 : node4426;
													assign node4426 = (inp[9]) ? 4'b0011 : node4427;
														assign node4427 = (inp[10]) ? node4429 : 4'b0111;
															assign node4429 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node4433 = (inp[10]) ? node4439 : node4434;
														assign node4434 = (inp[9]) ? node4436 : 4'b0011;
															assign node4436 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node4439 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node4442 = (inp[10]) ? node4482 : node4443;
											assign node4443 = (inp[0]) ? node4467 : node4444;
												assign node4444 = (inp[15]) ? node4452 : node4445;
													assign node4445 = (inp[4]) ? node4449 : node4446;
														assign node4446 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node4449 = (inp[3]) ? 4'b0100 : 4'b0010;
													assign node4452 = (inp[12]) ? node4458 : node4453;
														assign node4453 = (inp[9]) ? 4'b0000 : node4454;
															assign node4454 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node4458 = (inp[3]) ? node4464 : node4459;
															assign node4459 = (inp[4]) ? 4'b0100 : node4460;
																assign node4460 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node4464 = (inp[9]) ? 4'b0110 : 4'b0000;
												assign node4467 = (inp[15]) ? node4475 : node4468;
													assign node4468 = (inp[4]) ? node4470 : 4'b0000;
														assign node4470 = (inp[9]) ? node4472 : 4'b0000;
															assign node4472 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node4475 = (inp[9]) ? node4477 : 4'b0010;
														assign node4477 = (inp[4]) ? node4479 : 4'b0010;
															assign node4479 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node4482 = (inp[9]) ? node4506 : node4483;
												assign node4483 = (inp[15]) ? node4495 : node4484;
													assign node4484 = (inp[0]) ? node4490 : node4485;
														assign node4485 = (inp[4]) ? 4'b0100 : node4486;
															assign node4486 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node4490 = (inp[12]) ? node4492 : 4'b0100;
															assign node4492 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node4495 = (inp[0]) ? node4501 : node4496;
														assign node4496 = (inp[12]) ? node4498 : 4'b0100;
															assign node4498 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node4501 = (inp[12]) ? node4503 : 4'b0110;
															assign node4503 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node4506 = (inp[4]) ? node4520 : node4507;
													assign node4507 = (inp[12]) ? node4513 : node4508;
														assign node4508 = (inp[3]) ? node4510 : 4'b0010;
															assign node4510 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node4513 = (inp[15]) ? node4515 : 4'b0110;
															assign node4515 = (inp[3]) ? 4'b0110 : node4516;
																assign node4516 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node4520 = (inp[12]) ? 4'b0010 : 4'b0110;
						assign node4523 = (inp[13]) ? node5301 : node4524;
							assign node4524 = (inp[1]) ? node4932 : node4525;
								assign node4525 = (inp[12]) ? node4699 : node4526;
									assign node4526 = (inp[8]) ? node4618 : node4527;
										assign node4527 = (inp[2]) ? node4567 : node4528;
											assign node4528 = (inp[4]) ? node4544 : node4529;
												assign node4529 = (inp[9]) ? node4537 : node4530;
													assign node4530 = (inp[15]) ? node4534 : node4531;
														assign node4531 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node4534 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node4537 = (inp[3]) ? node4539 : 4'b0010;
														assign node4539 = (inp[0]) ? 4'b0000 : node4540;
															assign node4540 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node4544 = (inp[9]) ? node4560 : node4545;
													assign node4545 = (inp[10]) ? node4551 : node4546;
														assign node4546 = (inp[15]) ? 4'b0010 : node4547;
															assign node4547 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node4551 = (inp[3]) ? node4553 : 4'b0000;
															assign node4553 = (inp[15]) ? node4557 : node4554;
																assign node4554 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node4557 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node4560 = (inp[0]) ? node4564 : node4561;
														assign node4561 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node4564 = (inp[10]) ? 4'b0110 : 4'b0100;
											assign node4567 = (inp[3]) ? node4593 : node4568;
												assign node4568 = (inp[4]) ? node4582 : node4569;
													assign node4569 = (inp[9]) ? node4577 : node4570;
														assign node4570 = (inp[15]) ? node4574 : node4571;
															assign node4571 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node4574 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node4577 = (inp[0]) ? 4'b0001 : node4578;
															assign node4578 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node4582 = (inp[9]) ? node4590 : node4583;
														assign node4583 = (inp[0]) ? node4587 : node4584;
															assign node4584 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node4587 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node4590 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node4593 = (inp[9]) ? node4603 : node4594;
													assign node4594 = (inp[4]) ? 4'b0011 : node4595;
														assign node4595 = (inp[0]) ? node4599 : node4596;
															assign node4596 = (inp[10]) ? 4'b0111 : 4'b0101;
															assign node4599 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node4603 = (inp[4]) ? node4613 : node4604;
														assign node4604 = (inp[10]) ? 4'b0001 : node4605;
															assign node4605 = (inp[0]) ? node4609 : node4606;
																assign node4606 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node4609 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node4613 = (inp[0]) ? node4615 : 4'b0101;
															assign node4615 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node4618 = (inp[2]) ? node4664 : node4619;
											assign node4619 = (inp[3]) ? node4639 : node4620;
												assign node4620 = (inp[0]) ? node4632 : node4621;
													assign node4621 = (inp[15]) ? node4625 : node4622;
														assign node4622 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node4625 = (inp[9]) ? node4629 : node4626;
															assign node4626 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node4629 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node4632 = (inp[15]) ? node4634 : 4'b0001;
														assign node4634 = (inp[4]) ? 4'b0111 : node4635;
															assign node4635 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node4639 = (inp[9]) ? node4651 : node4640;
													assign node4640 = (inp[4]) ? node4644 : node4641;
														assign node4641 = (inp[10]) ? 4'b0111 : 4'b0101;
														assign node4644 = (inp[0]) ? node4648 : node4645;
															assign node4645 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node4648 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node4651 = (inp[4]) ? 4'b0101 : node4652;
														assign node4652 = (inp[10]) ? node4658 : node4653;
															assign node4653 = (inp[15]) ? 4'b0001 : node4654;
																assign node4654 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node4658 = (inp[0]) ? node4660 : 4'b0001;
																assign node4660 = (inp[15]) ? 4'b0011 : 4'b0001;
											assign node4664 = (inp[9]) ? node4680 : node4665;
												assign node4665 = (inp[4]) ? node4673 : node4666;
													assign node4666 = (inp[15]) ? node4670 : node4667;
														assign node4667 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node4670 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node4673 = (inp[15]) ? node4677 : node4674;
														assign node4674 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node4677 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node4680 = (inp[4]) ? node4686 : node4681;
													assign node4681 = (inp[15]) ? node4683 : 4'b0010;
														assign node4683 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node4686 = (inp[0]) ? node4692 : node4687;
														assign node4687 = (inp[3]) ? node4689 : 4'b0100;
															assign node4689 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node4692 = (inp[3]) ? node4696 : node4693;
															assign node4693 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node4696 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node4699 = (inp[3]) ? node4833 : node4700;
										assign node4700 = (inp[8]) ? node4766 : node4701;
											assign node4701 = (inp[2]) ? node4735 : node4702;
												assign node4702 = (inp[10]) ? node4718 : node4703;
													assign node4703 = (inp[15]) ? node4713 : node4704;
														assign node4704 = (inp[0]) ? node4706 : 4'b0010;
															assign node4706 = (inp[4]) ? node4710 : node4707;
																assign node4707 = (inp[9]) ? 4'b0000 : 4'b0100;
																assign node4710 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node4713 = (inp[4]) ? node4715 : 4'b0100;
															assign node4715 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node4718 = (inp[4]) ? node4730 : node4719;
														assign node4719 = (inp[9]) ? node4727 : node4720;
															assign node4720 = (inp[0]) ? node4724 : node4721;
																assign node4721 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node4724 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node4727 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node4730 = (inp[9]) ? 4'b0000 : node4731;
															assign node4731 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node4735 = (inp[15]) ? node4753 : node4736;
													assign node4736 = (inp[0]) ? node4744 : node4737;
														assign node4737 = (inp[9]) ? 4'b0111 : node4738;
															assign node4738 = (inp[10]) ? 4'b0011 : node4739;
																assign node4739 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node4744 = (inp[4]) ? 4'b0001 : node4745;
															assign node4745 = (inp[9]) ? node4749 : node4746;
																assign node4746 = (inp[10]) ? 4'b0001 : 4'b0101;
																assign node4749 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node4753 = (inp[0]) ? node4759 : node4754;
														assign node4754 = (inp[4]) ? node4756 : 4'b0101;
															assign node4756 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node4759 = (inp[9]) ? 4'b0111 : node4760;
															assign node4760 = (inp[4]) ? 4'b0111 : node4761;
																assign node4761 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node4766 = (inp[2]) ? node4806 : node4767;
												assign node4767 = (inp[15]) ? node4785 : node4768;
													assign node4768 = (inp[0]) ? 4'b0101 : node4769;
														assign node4769 = (inp[10]) ? node4777 : node4770;
															assign node4770 = (inp[9]) ? node4774 : node4771;
																assign node4771 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node4774 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node4777 = (inp[9]) ? node4781 : node4778;
																assign node4778 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node4781 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node4785 = (inp[0]) ? node4799 : node4786;
														assign node4786 = (inp[9]) ? node4794 : node4787;
															assign node4787 = (inp[4]) ? node4791 : node4788;
																assign node4788 = (inp[10]) ? 4'b0001 : 4'b0101;
																assign node4791 = (inp[10]) ? 4'b0101 : 4'b0001;
															assign node4794 = (inp[4]) ? 4'b0101 : node4795;
																assign node4795 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node4799 = (inp[9]) ? 4'b0111 : node4800;
															assign node4800 = (inp[10]) ? 4'b0011 : node4801;
																assign node4801 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node4806 = (inp[10]) ? node4822 : node4807;
													assign node4807 = (inp[4]) ? node4819 : node4808;
														assign node4808 = (inp[9]) ? node4816 : node4809;
															assign node4809 = (inp[0]) ? node4813 : node4810;
																assign node4810 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node4813 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node4816 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node4819 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node4822 = (inp[15]) ? 4'b0000 : node4823;
														assign node4823 = (inp[0]) ? node4829 : node4824;
															assign node4824 = (inp[9]) ? 4'b0110 : node4825;
																assign node4825 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node4829 = (inp[4]) ? 4'b0100 : 4'b0000;
										assign node4833 = (inp[8]) ? node4883 : node4834;
											assign node4834 = (inp[2]) ? node4864 : node4835;
												assign node4835 = (inp[15]) ? node4851 : node4836;
													assign node4836 = (inp[0]) ? node4848 : node4837;
														assign node4837 = (inp[9]) ? node4843 : node4838;
															assign node4838 = (inp[10]) ? node4840 : 4'b0010;
																assign node4840 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node4843 = (inp[4]) ? node4845 : 4'b0100;
																assign node4845 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node4848 = (inp[10]) ? 4'b0010 : 4'b0000;
													assign node4851 = (inp[0]) ? node4859 : node4852;
														assign node4852 = (inp[9]) ? node4854 : 4'b0110;
															assign node4854 = (inp[10]) ? node4856 : 4'b0110;
																assign node4856 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node4859 = (inp[9]) ? 4'b0100 : node4860;
															assign node4860 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node4864 = (inp[4]) ? node4876 : node4865;
													assign node4865 = (inp[15]) ? node4867 : 4'b0111;
														assign node4867 = (inp[0]) ? node4873 : node4868;
															assign node4868 = (inp[10]) ? node4870 : 4'b0001;
																assign node4870 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node4873 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node4876 = (inp[15]) ? 4'b0111 : node4877;
														assign node4877 = (inp[9]) ? 4'b0111 : node4878;
															assign node4878 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node4883 = (inp[2]) ? node4911 : node4884;
												assign node4884 = (inp[9]) ? node4896 : node4885;
													assign node4885 = (inp[10]) ? node4889 : node4886;
														assign node4886 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node4889 = (inp[4]) ? node4893 : node4890;
															assign node4890 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node4893 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node4896 = (inp[15]) ? node4902 : node4897;
														assign node4897 = (inp[4]) ? 4'b0011 : node4898;
															assign node4898 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node4902 = (inp[4]) ? node4906 : node4903;
															assign node4903 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node4906 = (inp[10]) ? 4'b0011 : node4907;
																assign node4907 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node4911 = (inp[0]) ? node4923 : node4912;
													assign node4912 = (inp[4]) ? node4914 : 4'b0100;
														assign node4914 = (inp[15]) ? 4'b0000 : node4915;
															assign node4915 = (inp[9]) ? node4919 : node4916;
																assign node4916 = (inp[10]) ? 4'b0100 : 4'b0010;
																assign node4919 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node4923 = (inp[4]) ? node4929 : node4924;
														assign node4924 = (inp[10]) ? node4926 : 4'b0010;
															assign node4926 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node4929 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node4932 = (inp[8]) ? node5108 : node4933;
									assign node4933 = (inp[2]) ? node5021 : node4934;
										assign node4934 = (inp[0]) ? node4972 : node4935;
											assign node4935 = (inp[15]) ? node4959 : node4936;
												assign node4936 = (inp[9]) ? node4950 : node4937;
													assign node4937 = (inp[3]) ? node4947 : node4938;
														assign node4938 = (inp[12]) ? node4940 : 4'b0110;
															assign node4940 = (inp[4]) ? node4944 : node4941;
																assign node4941 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node4944 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node4947 = (inp[4]) ? 4'b0100 : 4'b0110;
													assign node4950 = (inp[4]) ? node4952 : 4'b0010;
														assign node4952 = (inp[3]) ? 4'b0100 : node4953;
															assign node4953 = (inp[10]) ? node4955 : 4'b0110;
																assign node4955 = (inp[12]) ? 4'b0010 : 4'b0110;
												assign node4959 = (inp[9]) ? node4965 : node4960;
													assign node4960 = (inp[10]) ? 4'b0000 : node4961;
														assign node4961 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node4965 = (inp[4]) ? node4969 : node4966;
														assign node4966 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node4969 = (inp[12]) ? 4'b0100 : 4'b0110;
											assign node4972 = (inp[15]) ? node4990 : node4973;
												assign node4973 = (inp[3]) ? 4'b0000 : node4974;
													assign node4974 = (inp[4]) ? node4982 : node4975;
														assign node4975 = (inp[9]) ? 4'b0000 : node4976;
															assign node4976 = (inp[10]) ? node4978 : 4'b0100;
																assign node4978 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node4982 = (inp[9]) ? 4'b0100 : node4983;
															assign node4983 = (inp[12]) ? node4985 : 4'b0000;
																assign node4985 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node4990 = (inp[3]) ? node5004 : node4991;
													assign node4991 = (inp[12]) ? node4993 : 4'b0110;
														assign node4993 = (inp[4]) ? node4999 : node4994;
															assign node4994 = (inp[10]) ? 4'b0110 : node4995;
																assign node4995 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node4999 = (inp[10]) ? 4'b0010 : node5000;
																assign node5000 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node5004 = (inp[12]) ? node5010 : node5005;
														assign node5005 = (inp[10]) ? 4'b0010 : node5006;
															assign node5006 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node5010 = (inp[10]) ? node5016 : node5011;
															assign node5011 = (inp[9]) ? 4'b0100 : node5012;
																assign node5012 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node5016 = (inp[4]) ? node5018 : 4'b0100;
																assign node5018 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node5021 = (inp[10]) ? node5073 : node5022;
											assign node5022 = (inp[9]) ? node5044 : node5023;
												assign node5023 = (inp[3]) ? node5035 : node5024;
													assign node5024 = (inp[15]) ? node5032 : node5025;
														assign node5025 = (inp[0]) ? node5027 : 4'b1011;
															assign node5027 = (inp[12]) ? 4'b1101 : node5028;
																assign node5028 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node5032 = (inp[0]) ? 4'b1011 : 4'b1101;
													assign node5035 = (inp[4]) ? node5039 : node5036;
														assign node5036 = (inp[0]) ? 4'b1001 : 4'b1101;
														assign node5039 = (inp[15]) ? node5041 : 4'b1111;
															assign node5041 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node5044 = (inp[3]) ? node5056 : node5045;
													assign node5045 = (inp[4]) ? node5047 : 4'b1011;
														assign node5047 = (inp[12]) ? node5051 : node5048;
															assign node5048 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node5051 = (inp[0]) ? 4'b1001 : node5052;
																assign node5052 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node5056 = (inp[4]) ? node5070 : node5057;
														assign node5057 = (inp[12]) ? node5065 : node5058;
															assign node5058 = (inp[0]) ? node5062 : node5059;
																assign node5059 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node5062 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node5065 = (inp[15]) ? 4'b1111 : node5066;
																assign node5066 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node5070 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node5073 = (inp[9]) ? node5093 : node5074;
												assign node5074 = (inp[4]) ? node5076 : 4'b1011;
													assign node5076 = (inp[15]) ? node5084 : node5077;
														assign node5077 = (inp[12]) ? node5079 : 4'b1101;
															assign node5079 = (inp[0]) ? 4'b1111 : node5080;
																assign node5080 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node5084 = (inp[12]) ? node5086 : 4'b1111;
															assign node5086 = (inp[0]) ? node5090 : node5087;
																assign node5087 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node5090 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node5093 = (inp[4]) ? node5105 : node5094;
													assign node5094 = (inp[3]) ? node5100 : node5095;
														assign node5095 = (inp[0]) ? node5097 : 4'b1101;
															assign node5097 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node5100 = (inp[0]) ? node5102 : 4'b1111;
															assign node5102 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node5105 = (inp[15]) ? 4'b1011 : 4'b1001;
									assign node5108 = (inp[2]) ? node5218 : node5109;
										assign node5109 = (inp[15]) ? node5159 : node5110;
											assign node5110 = (inp[0]) ? node5142 : node5111;
												assign node5111 = (inp[3]) ? node5127 : node5112;
													assign node5112 = (inp[10]) ? node5122 : node5113;
														assign node5113 = (inp[9]) ? node5115 : 4'b1011;
															assign node5115 = (inp[12]) ? node5119 : node5116;
																assign node5116 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node5119 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node5122 = (inp[9]) ? 4'b1011 : node5123;
															assign node5123 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node5127 = (inp[12]) ? node5135 : node5128;
														assign node5128 = (inp[4]) ? 4'b1011 : node5129;
															assign node5129 = (inp[10]) ? 4'b1011 : node5130;
																assign node5130 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node5135 = (inp[9]) ? node5139 : node5136;
															assign node5136 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node5139 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node5142 = (inp[3]) ? node5144 : 4'b1101;
													assign node5144 = (inp[4]) ? node5152 : node5145;
														assign node5145 = (inp[12]) ? 4'b1111 : node5146;
															assign node5146 = (inp[9]) ? node5148 : 4'b1001;
																assign node5148 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node5152 = (inp[9]) ? node5154 : 4'b1111;
															assign node5154 = (inp[12]) ? 4'b1011 : node5155;
																assign node5155 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node5159 = (inp[0]) ? node5181 : node5160;
												assign node5160 = (inp[3]) ? node5172 : node5161;
													assign node5161 = (inp[4]) ? node5169 : node5162;
														assign node5162 = (inp[9]) ? node5164 : 4'b1001;
															assign node5164 = (inp[12]) ? 4'b1101 : node5165;
																assign node5165 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node5169 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node5172 = (inp[10]) ? node5178 : node5173;
														assign node5173 = (inp[9]) ? 4'b1111 : node5174;
															assign node5174 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node5178 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node5181 = (inp[3]) ? node5199 : node5182;
													assign node5182 = (inp[12]) ? node5192 : node5183;
														assign node5183 = (inp[4]) ? node5185 : 4'b1111;
															assign node5185 = (inp[10]) ? node5189 : node5186;
																assign node5186 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node5189 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node5192 = (inp[4]) ? node5196 : node5193;
															assign node5193 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node5196 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node5199 = (inp[9]) ? node5209 : node5200;
														assign node5200 = (inp[12]) ? 4'b1011 : node5201;
															assign node5201 = (inp[10]) ? node5205 : node5202;
																assign node5202 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node5205 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node5209 = (inp[4]) ? node5213 : node5210;
															assign node5210 = (inp[10]) ? 4'b1101 : 4'b1011;
															assign node5213 = (inp[10]) ? 4'b1001 : node5214;
																assign node5214 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node5218 = (inp[0]) ? node5248 : node5219;
											assign node5219 = (inp[15]) ? node5237 : node5220;
												assign node5220 = (inp[4]) ? node5226 : node5221;
													assign node5221 = (inp[9]) ? node5223 : 4'b1010;
														assign node5223 = (inp[3]) ? 4'b1010 : 4'b1110;
													assign node5226 = (inp[3]) ? node5232 : node5227;
														assign node5227 = (inp[9]) ? 4'b1010 : node5228;
															assign node5228 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node5232 = (inp[12]) ? node5234 : 4'b1010;
															assign node5234 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node5237 = (inp[3]) ? node5245 : node5238;
													assign node5238 = (inp[4]) ? 4'b1000 : node5239;
														assign node5239 = (inp[10]) ? node5241 : 4'b1100;
															assign node5241 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node5245 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node5248 = (inp[15]) ? node5280 : node5249;
												assign node5249 = (inp[3]) ? node5269 : node5250;
													assign node5250 = (inp[12]) ? node5262 : node5251;
														assign node5251 = (inp[4]) ? node5257 : node5252;
															assign node5252 = (inp[10]) ? node5254 : 4'b1000;
																assign node5254 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node5257 = (inp[10]) ? node5259 : 4'b1100;
																assign node5259 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node5262 = (inp[10]) ? 4'b1100 : node5263;
															assign node5263 = (inp[9]) ? node5265 : 4'b1100;
																assign node5265 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node5269 = (inp[4]) ? node5275 : node5270;
														assign node5270 = (inp[10]) ? node5272 : 4'b1000;
															assign node5272 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node5275 = (inp[9]) ? node5277 : 4'b1110;
															assign node5277 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node5280 = (inp[3]) ? node5294 : node5281;
													assign node5281 = (inp[4]) ? node5291 : node5282;
														assign node5282 = (inp[10]) ? node5288 : node5283;
															assign node5283 = (inp[12]) ? 4'b1110 : node5284;
																assign node5284 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node5288 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node5291 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node5294 = (inp[10]) ? node5298 : node5295;
														assign node5295 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node5298 = (inp[4]) ? 4'b1000 : 4'b1100;
							assign node5301 = (inp[1]) ? node5649 : node5302;
								assign node5302 = (inp[8]) ? node5464 : node5303;
									assign node5303 = (inp[2]) ? node5381 : node5304;
										assign node5304 = (inp[9]) ? node5352 : node5305;
											assign node5305 = (inp[4]) ? node5331 : node5306;
												assign node5306 = (inp[10]) ? node5314 : node5307;
													assign node5307 = (inp[15]) ? node5311 : node5308;
														assign node5308 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node5311 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node5314 = (inp[12]) ? node5322 : node5315;
														assign node5315 = (inp[15]) ? node5319 : node5316;
															assign node5316 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node5319 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node5322 = (inp[3]) ? node5326 : node5323;
															assign node5323 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node5326 = (inp[0]) ? 4'b0010 : node5327;
																assign node5327 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node5331 = (inp[12]) ? node5341 : node5332;
													assign node5332 = (inp[3]) ? node5334 : 4'b0000;
														assign node5334 = (inp[0]) ? node5338 : node5335;
															assign node5335 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node5338 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node5341 = (inp[10]) ? node5347 : node5342;
														assign node5342 = (inp[15]) ? 4'b0010 : node5343;
															assign node5343 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node5347 = (inp[15]) ? node5349 : 4'b0110;
															assign node5349 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node5352 = (inp[4]) ? node5366 : node5353;
												assign node5353 = (inp[12]) ? node5355 : 4'b0000;
													assign node5355 = (inp[10]) ? node5361 : node5356;
														assign node5356 = (inp[15]) ? 4'b0000 : node5357;
															assign node5357 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node5361 = (inp[0]) ? 4'b0110 : node5362;
															assign node5362 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node5366 = (inp[3]) ? node5372 : node5367;
													assign node5367 = (inp[0]) ? node5369 : 4'b0000;
														assign node5369 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node5372 = (inp[12]) ? node5378 : node5373;
														assign node5373 = (inp[0]) ? node5375 : 4'b0100;
															assign node5375 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node5378 = (inp[10]) ? 4'b0000 : 4'b0100;
										assign node5381 = (inp[0]) ? node5415 : node5382;
											assign node5382 = (inp[15]) ? node5400 : node5383;
												assign node5383 = (inp[3]) ? node5387 : node5384;
													assign node5384 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node5387 = (inp[9]) ? node5393 : node5388;
														assign node5388 = (inp[4]) ? 4'b1101 : node5389;
															assign node5389 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node5393 = (inp[4]) ? node5395 : 4'b1101;
															assign node5395 = (inp[12]) ? 4'b1001 : node5396;
																assign node5396 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node5400 = (inp[3]) ? node5408 : node5401;
													assign node5401 = (inp[10]) ? node5403 : 4'b1001;
														assign node5403 = (inp[4]) ? node5405 : 4'b1101;
															assign node5405 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node5408 = (inp[4]) ? node5410 : 4'b1001;
														assign node5410 = (inp[12]) ? node5412 : 4'b1111;
															assign node5412 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node5415 = (inp[12]) ? node5445 : node5416;
												assign node5416 = (inp[15]) ? node5430 : node5417;
													assign node5417 = (inp[3]) ? node5423 : node5418;
														assign node5418 = (inp[4]) ? 4'b1001 : node5419;
															assign node5419 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node5423 = (inp[4]) ? node5425 : 4'b1001;
															assign node5425 = (inp[10]) ? node5427 : 4'b1111;
																assign node5427 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node5430 = (inp[3]) ? node5442 : node5431;
														assign node5431 = (inp[4]) ? node5437 : node5432;
															assign node5432 = (inp[10]) ? node5434 : 4'b1111;
																assign node5434 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node5437 = (inp[10]) ? node5439 : 4'b1011;
																assign node5439 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node5442 = (inp[4]) ? 4'b1101 : 4'b1011;
												assign node5445 = (inp[3]) ? node5453 : node5446;
													assign node5446 = (inp[15]) ? 4'b1111 : node5447;
														assign node5447 = (inp[4]) ? 4'b1101 : node5448;
															assign node5448 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node5453 = (inp[15]) ? node5459 : node5454;
														assign node5454 = (inp[9]) ? node5456 : 4'b1111;
															assign node5456 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node5459 = (inp[4]) ? node5461 : 4'b1011;
															assign node5461 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node5464 = (inp[2]) ? node5548 : node5465;
										assign node5465 = (inp[9]) ? node5515 : node5466;
											assign node5466 = (inp[4]) ? node5494 : node5467;
												assign node5467 = (inp[10]) ? node5479 : node5468;
													assign node5468 = (inp[12]) ? node5474 : node5469;
														assign node5469 = (inp[0]) ? 4'b1111 : node5470;
															assign node5470 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node5474 = (inp[0]) ? node5476 : 4'b1011;
															assign node5476 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node5479 = (inp[3]) ? node5485 : node5480;
														assign node5480 = (inp[12]) ? 4'b1011 : node5481;
															assign node5481 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5485 = (inp[12]) ? 4'b1001 : node5486;
															assign node5486 = (inp[0]) ? node5490 : node5487;
																assign node5487 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node5490 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node5494 = (inp[10]) ? node5500 : node5495;
													assign node5495 = (inp[12]) ? 4'b1111 : node5496;
														assign node5496 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node5500 = (inp[15]) ? node5510 : node5501;
														assign node5501 = (inp[12]) ? 4'b1111 : node5502;
															assign node5502 = (inp[0]) ? node5506 : node5503;
																assign node5503 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node5506 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node5510 = (inp[3]) ? node5512 : 4'b1111;
															assign node5512 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node5515 = (inp[4]) ? node5533 : node5516;
												assign node5516 = (inp[12]) ? node5524 : node5517;
													assign node5517 = (inp[10]) ? 4'b1101 : node5518;
														assign node5518 = (inp[15]) ? 4'b1011 : node5519;
															assign node5519 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node5524 = (inp[3]) ? node5530 : node5525;
														assign node5525 = (inp[0]) ? 4'b1101 : node5526;
															assign node5526 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node5530 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node5533 = (inp[3]) ? node5539 : node5534;
													assign node5534 = (inp[0]) ? 4'b1001 : node5535;
														assign node5535 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node5539 = (inp[0]) ? node5545 : node5540;
														assign node5540 = (inp[15]) ? 4'b1011 : node5541;
															assign node5541 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node5545 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node5548 = (inp[9]) ? node5590 : node5549;
											assign node5549 = (inp[4]) ? node5571 : node5550;
												assign node5550 = (inp[12]) ? node5558 : node5551;
													assign node5551 = (inp[10]) ? node5555 : node5552;
														assign node5552 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node5555 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node5558 = (inp[3]) ? node5566 : node5559;
														assign node5559 = (inp[10]) ? node5563 : node5560;
															assign node5560 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node5563 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node5566 = (inp[0]) ? node5568 : 4'b1010;
															assign node5568 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node5571 = (inp[10]) ? node5581 : node5572;
													assign node5572 = (inp[12]) ? 4'b1110 : node5573;
														assign node5573 = (inp[15]) ? node5577 : node5574;
															assign node5574 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node5577 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node5581 = (inp[0]) ? node5583 : 4'b1110;
														assign node5583 = (inp[3]) ? node5587 : node5584;
															assign node5584 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node5587 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node5590 = (inp[4]) ? node5620 : node5591;
												assign node5591 = (inp[12]) ? node5607 : node5592;
													assign node5592 = (inp[10]) ? node5598 : node5593;
														assign node5593 = (inp[3]) ? node5595 : 4'b1000;
															assign node5595 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node5598 = (inp[15]) ? node5600 : 4'b1110;
															assign node5600 = (inp[3]) ? node5604 : node5601;
																assign node5601 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node5604 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node5607 = (inp[0]) ? node5613 : node5608;
														assign node5608 = (inp[15]) ? node5610 : 4'b1110;
															assign node5610 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node5613 = (inp[15]) ? node5617 : node5614;
															assign node5614 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node5617 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node5620 = (inp[10]) ? node5636 : node5621;
													assign node5621 = (inp[12]) ? node5633 : node5622;
														assign node5622 = (inp[15]) ? node5628 : node5623;
															assign node5623 = (inp[0]) ? 4'b1100 : node5624;
																assign node5624 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node5628 = (inp[3]) ? 4'b1110 : node5629;
																assign node5629 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node5633 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node5636 = (inp[3]) ? node5642 : node5637;
														assign node5637 = (inp[0]) ? node5639 : 4'b1010;
															assign node5639 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node5642 = (inp[0]) ? node5646 : node5643;
															assign node5643 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node5646 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node5649 = (inp[12]) ? node5879 : node5650;
									assign node5650 = (inp[0]) ? node5760 : node5651;
										assign node5651 = (inp[15]) ? node5719 : node5652;
											assign node5652 = (inp[3]) ? node5690 : node5653;
												assign node5653 = (inp[10]) ? node5677 : node5654;
													assign node5654 = (inp[9]) ? node5664 : node5655;
														assign node5655 = (inp[4]) ? 4'b1011 : node5656;
															assign node5656 = (inp[2]) ? node5660 : node5657;
																assign node5657 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node5660 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node5664 = (inp[4]) ? node5672 : node5665;
															assign node5665 = (inp[8]) ? node5669 : node5666;
																assign node5666 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node5669 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node5672 = (inp[8]) ? 4'b1111 : node5673;
																assign node5673 = (inp[2]) ? 4'b1111 : 4'b1110;
													assign node5677 = (inp[4]) ? node5687 : node5678;
														assign node5678 = (inp[9]) ? node5680 : 4'b1011;
															assign node5680 = (inp[2]) ? node5684 : node5681;
																assign node5681 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node5684 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node5687 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node5690 = (inp[9]) ? node5706 : node5691;
													assign node5691 = (inp[10]) ? node5701 : node5692;
														assign node5692 = (inp[4]) ? node5694 : 4'b1111;
															assign node5694 = (inp[8]) ? node5698 : node5695;
																assign node5695 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node5698 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node5701 = (inp[4]) ? node5703 : 4'b1011;
															assign node5703 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node5706 = (inp[10]) ? node5714 : node5707;
														assign node5707 = (inp[4]) ? node5711 : node5708;
															assign node5708 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node5711 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node5714 = (inp[8]) ? 4'b1100 : node5715;
															assign node5715 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node5719 = (inp[3]) ? node5735 : node5720;
												assign node5720 = (inp[4]) ? node5730 : node5721;
													assign node5721 = (inp[9]) ? node5723 : 4'b1101;
														assign node5723 = (inp[10]) ? 4'b1101 : node5724;
															assign node5724 = (inp[2]) ? 4'b1001 : node5725;
																assign node5725 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node5730 = (inp[10]) ? 4'b1100 : node5731;
														assign node5731 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node5735 = (inp[9]) ? node5747 : node5736;
													assign node5736 = (inp[4]) ? node5744 : node5737;
														assign node5737 = (inp[10]) ? node5741 : node5738;
															assign node5738 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node5741 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node5744 = (inp[10]) ? 4'b1111 : 4'b1000;
													assign node5747 = (inp[10]) ? node5751 : node5748;
														assign node5748 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node5751 = (inp[4]) ? node5755 : node5752;
															assign node5752 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node5755 = (inp[8]) ? 4'b1010 : node5756;
																assign node5756 = (inp[2]) ? 4'b1011 : 4'b1010;
										assign node5760 = (inp[15]) ? node5824 : node5761;
											assign node5761 = (inp[3]) ? node5787 : node5762;
												assign node5762 = (inp[2]) ? node5774 : node5763;
													assign node5763 = (inp[8]) ? 4'b1001 : node5764;
														assign node5764 = (inp[10]) ? node5766 : 4'b1000;
															assign node5766 = (inp[9]) ? node5770 : node5767;
																assign node5767 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node5770 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node5774 = (inp[8]) ? node5782 : node5775;
														assign node5775 = (inp[4]) ? node5777 : 4'b1101;
															assign node5777 = (inp[10]) ? node5779 : 4'b1101;
																assign node5779 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node5782 = (inp[4]) ? node5784 : 4'b1100;
															assign node5784 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node5787 = (inp[4]) ? node5803 : node5788;
													assign node5788 = (inp[10]) ? node5798 : node5789;
														assign node5789 = (inp[9]) ? node5793 : node5790;
															assign node5790 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node5793 = (inp[2]) ? node5795 : 4'b1001;
																assign node5795 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node5798 = (inp[9]) ? 4'b1110 : node5799;
															assign node5799 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node5803 = (inp[9]) ? node5813 : node5804;
														assign node5804 = (inp[10]) ? node5808 : node5805;
															assign node5805 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node5808 = (inp[2]) ? node5810 : 4'b1111;
																assign node5810 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node5813 = (inp[10]) ? node5821 : node5814;
															assign node5814 = (inp[2]) ? node5818 : node5815;
																assign node5815 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node5818 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node5821 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node5824 = (inp[3]) ? node5844 : node5825;
												assign node5825 = (inp[8]) ? node5835 : node5826;
													assign node5826 = (inp[2]) ? node5830 : node5827;
														assign node5827 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node5830 = (inp[9]) ? node5832 : 4'b1111;
															assign node5832 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node5835 = (inp[2]) ? 4'b1010 : node5836;
														assign node5836 = (inp[4]) ? node5838 : 4'b1011;
															assign node5838 = (inp[9]) ? node5840 : 4'b1111;
																assign node5840 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node5844 = (inp[10]) ? node5862 : node5845;
													assign node5845 = (inp[8]) ? node5859 : node5846;
														assign node5846 = (inp[2]) ? node5854 : node5847;
															assign node5847 = (inp[4]) ? node5851 : node5848;
																assign node5848 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node5851 = (inp[9]) ? 4'b1100 : 4'b1010;
															assign node5854 = (inp[4]) ? 4'b1011 : node5855;
																assign node5855 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node5859 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node5862 = (inp[4]) ? node5868 : node5863;
														assign node5863 = (inp[9]) ? 4'b1100 : node5864;
															assign node5864 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node5868 = (inp[9]) ? node5876 : node5869;
															assign node5869 = (inp[8]) ? node5873 : node5870;
																assign node5870 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node5873 = (inp[2]) ? 4'b1100 : 4'b1101;
															assign node5876 = (inp[8]) ? 4'b1001 : 4'b1000;
									assign node5879 = (inp[4]) ? node5985 : node5880;
										assign node5880 = (inp[9]) ? node5932 : node5881;
											assign node5881 = (inp[2]) ? node5905 : node5882;
												assign node5882 = (inp[8]) ? node5888 : node5883;
													assign node5883 = (inp[0]) ? 4'b1010 : node5884;
														assign node5884 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node5888 = (inp[10]) ? node5898 : node5889;
														assign node5889 = (inp[3]) ? node5891 : 4'b1011;
															assign node5891 = (inp[15]) ? node5895 : node5892;
																assign node5892 = (inp[0]) ? 4'b1001 : 4'b1011;
																assign node5895 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node5898 = (inp[15]) ? node5902 : node5899;
															assign node5899 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node5902 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node5905 = (inp[8]) ? node5921 : node5906;
													assign node5906 = (inp[3]) ? node5914 : node5907;
														assign node5907 = (inp[0]) ? node5911 : node5908;
															assign node5908 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node5911 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node5914 = (inp[15]) ? node5918 : node5915;
															assign node5915 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node5918 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node5921 = (inp[3]) ? 4'b1000 : node5922;
														assign node5922 = (inp[10]) ? node5924 : 4'b1000;
															assign node5924 = (inp[0]) ? node5928 : node5925;
																assign node5925 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node5928 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node5932 = (inp[0]) ? node5960 : node5933;
												assign node5933 = (inp[2]) ? node5949 : node5934;
													assign node5934 = (inp[8]) ? node5942 : node5935;
														assign node5935 = (inp[10]) ? node5937 : 4'b1100;
															assign node5937 = (inp[15]) ? 4'b1110 : node5938;
																assign node5938 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node5942 = (inp[15]) ? node5946 : node5943;
															assign node5943 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node5946 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node5949 = (inp[8]) ? node5955 : node5950;
														assign node5950 = (inp[3]) ? node5952 : 4'b1111;
															assign node5952 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node5955 = (inp[15]) ? node5957 : 4'b1110;
															assign node5957 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node5960 = (inp[10]) ? node5968 : node5961;
													assign node5961 = (inp[8]) ? node5963 : 4'b1101;
														assign node5963 = (inp[3]) ? node5965 : 4'b1111;
															assign node5965 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node5968 = (inp[8]) ? node5978 : node5969;
														assign node5969 = (inp[2]) ? node5973 : node5970;
															assign node5970 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node5973 = (inp[15]) ? 4'b1111 : node5974;
																assign node5974 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node5978 = (inp[2]) ? 4'b1100 : node5979;
															assign node5979 = (inp[15]) ? 4'b1101 : node5980;
																assign node5980 = (inp[3]) ? 4'b1111 : 4'b1101;
										assign node5985 = (inp[9]) ? node6033 : node5986;
											assign node5986 = (inp[10]) ? node6014 : node5987;
												assign node5987 = (inp[15]) ? node5993 : node5988;
													assign node5988 = (inp[0]) ? 4'b1101 : node5989;
														assign node5989 = (inp[8]) ? 4'b1101 : 4'b1110;
													assign node5993 = (inp[2]) ? node6005 : node5994;
														assign node5994 = (inp[8]) ? node5998 : node5995;
															assign node5995 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node5998 = (inp[0]) ? node6002 : node5999;
																assign node5999 = (inp[3]) ? 4'b1111 : 4'b1101;
																assign node6002 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node6005 = (inp[8]) ? node6009 : node6006;
															assign node6006 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node6009 = (inp[3]) ? 4'b1100 : node6010;
																assign node6010 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node6014 = (inp[15]) ? node6024 : node6015;
													assign node6015 = (inp[8]) ? node6017 : 4'b1111;
														assign node6017 = (inp[2]) ? node6019 : 4'b1111;
															assign node6019 = (inp[0]) ? node6021 : 4'b1100;
																assign node6021 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node6024 = (inp[8]) ? node6030 : node6025;
														assign node6025 = (inp[2]) ? node6027 : 4'b1100;
															assign node6027 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node6030 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node6033 = (inp[15]) ? node6057 : node6034;
												assign node6034 = (inp[3]) ? node6050 : node6035;
													assign node6035 = (inp[0]) ? node6041 : node6036;
														assign node6036 = (inp[8]) ? node6038 : 4'b1010;
															assign node6038 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node6041 = (inp[10]) ? node6047 : node6042;
															assign node6042 = (inp[8]) ? node6044 : 4'b1001;
																assign node6044 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node6047 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node6050 = (inp[0]) ? node6052 : 4'b1000;
														assign node6052 = (inp[2]) ? node6054 : 4'b1010;
															assign node6054 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node6057 = (inp[10]) ? node6067 : node6058;
													assign node6058 = (inp[2]) ? node6064 : node6059;
														assign node6059 = (inp[8]) ? node6061 : 4'b1000;
															assign node6061 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node6064 = (inp[8]) ? 4'b1000 : 4'b1011;
													assign node6067 = (inp[8]) ? node6075 : node6068;
														assign node6068 = (inp[2]) ? 4'b1001 : node6069;
															assign node6069 = (inp[0]) ? 4'b1000 : node6070;
																assign node6070 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node6075 = (inp[2]) ? 4'b1000 : 4'b1001;
				assign node6078 = (inp[13]) ? node9232 : node6079;
					assign node6079 = (inp[6]) ? node7701 : node6080;
						assign node6080 = (inp[1]) ? node6910 : node6081;
							assign node6081 = (inp[12]) ? node6477 : node6082;
								assign node6082 = (inp[0]) ? node6286 : node6083;
									assign node6083 = (inp[15]) ? node6201 : node6084;
										assign node6084 = (inp[3]) ? node6134 : node6085;
											assign node6085 = (inp[4]) ? node6115 : node6086;
												assign node6086 = (inp[9]) ? node6100 : node6087;
													assign node6087 = (inp[10]) ? node6095 : node6088;
														assign node6088 = (inp[7]) ? node6090 : 4'b1110;
															assign node6090 = (inp[8]) ? 4'b1111 : node6091;
																assign node6091 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node6095 = (inp[2]) ? 4'b1110 : node6096;
															assign node6096 = (inp[7]) ? 4'b1110 : 4'b1111;
													assign node6100 = (inp[7]) ? node6110 : node6101;
														assign node6101 = (inp[10]) ? 4'b1011 : node6102;
															assign node6102 = (inp[8]) ? node6106 : node6103;
																assign node6103 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node6106 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node6110 = (inp[8]) ? node6112 : 4'b1010;
															assign node6112 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node6115 = (inp[9]) ? node6125 : node6116;
													assign node6116 = (inp[8]) ? 4'b1011 : node6117;
														assign node6117 = (inp[10]) ? 4'b1010 : node6118;
															assign node6118 = (inp[7]) ? node6120 : 4'b1011;
																assign node6120 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node6125 = (inp[8]) ? 4'b1100 : node6126;
														assign node6126 = (inp[10]) ? node6128 : 4'b1100;
															assign node6128 = (inp[7]) ? 4'b1101 : node6129;
																assign node6129 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node6134 = (inp[2]) ? node6168 : node6135;
												assign node6135 = (inp[10]) ? node6151 : node6136;
													assign node6136 = (inp[7]) ? node6144 : node6137;
														assign node6137 = (inp[8]) ? node6139 : 4'b1101;
															assign node6139 = (inp[4]) ? node6141 : 4'b1000;
																assign node6141 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node6144 = (inp[8]) ? 4'b1101 : node6145;
															assign node6145 = (inp[4]) ? 4'b1100 : node6146;
																assign node6146 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node6151 = (inp[9]) ? node6161 : node6152;
														assign node6152 = (inp[4]) ? node6158 : node6153;
															assign node6153 = (inp[7]) ? 4'b1101 : node6154;
																assign node6154 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node6158 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node6161 = (inp[4]) ? 4'b1101 : node6162;
															assign node6162 = (inp[8]) ? 4'b1001 : node6163;
																assign node6163 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node6168 = (inp[4]) ? node6182 : node6169;
													assign node6169 = (inp[9]) ? node6177 : node6170;
														assign node6170 = (inp[10]) ? 4'b1101 : node6171;
															assign node6171 = (inp[7]) ? 4'b1101 : node6172;
																assign node6172 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node6177 = (inp[8]) ? 4'b1001 : node6178;
															assign node6178 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node6182 = (inp[9]) ? node6196 : node6183;
														assign node6183 = (inp[10]) ? node6191 : node6184;
															assign node6184 = (inp[8]) ? node6188 : node6185;
																assign node6185 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node6188 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node6191 = (inp[8]) ? node6193 : 4'b1001;
																assign node6193 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node6196 = (inp[8]) ? node6198 : 4'b1100;
															assign node6198 = (inp[7]) ? 4'b1100 : 4'b1101;
										assign node6201 = (inp[3]) ? node6265 : node6202;
											assign node6202 = (inp[9]) ? node6232 : node6203;
												assign node6203 = (inp[4]) ? node6211 : node6204;
													assign node6204 = (inp[7]) ? 4'b1101 : node6205;
														assign node6205 = (inp[2]) ? node6207 : 4'b1100;
															assign node6207 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node6211 = (inp[10]) ? node6221 : node6212;
														assign node6212 = (inp[7]) ? node6214 : 4'b1000;
															assign node6214 = (inp[8]) ? node6218 : node6215;
																assign node6215 = (inp[2]) ? 4'b1001 : 4'b1000;
																assign node6218 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node6221 = (inp[7]) ? node6227 : node6222;
															assign node6222 = (inp[8]) ? node6224 : 4'b1001;
																assign node6224 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node6227 = (inp[2]) ? 4'b1000 : node6228;
																assign node6228 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node6232 = (inp[4]) ? node6252 : node6233;
													assign node6233 = (inp[7]) ? node6241 : node6234;
														assign node6234 = (inp[10]) ? node6238 : node6235;
															assign node6235 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node6238 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node6241 = (inp[10]) ? node6247 : node6242;
															assign node6242 = (inp[2]) ? 4'b1000 : node6243;
																assign node6243 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node6247 = (inp[2]) ? node6249 : 4'b1000;
																assign node6249 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node6252 = (inp[2]) ? node6258 : node6253;
														assign node6253 = (inp[10]) ? 4'b1111 : node6254;
															assign node6254 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node6258 = (inp[10]) ? node6260 : 4'b1111;
															assign node6260 = (inp[8]) ? node6262 : 4'b1110;
																assign node6262 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node6265 = (inp[9]) ? node6277 : node6266;
												assign node6266 = (inp[4]) ? node6268 : 4'b1110;
													assign node6268 = (inp[2]) ? node6270 : 4'b1010;
														assign node6270 = (inp[8]) ? node6274 : node6271;
															assign node6271 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node6274 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node6277 = (inp[4]) ? node6283 : node6278;
													assign node6278 = (inp[8]) ? 4'b1011 : node6279;
														assign node6279 = (inp[10]) ? 4'b1011 : 4'b1010;
													assign node6283 = (inp[8]) ? 4'b1110 : 4'b1111;
									assign node6286 = (inp[2]) ? node6384 : node6287;
										assign node6287 = (inp[3]) ? node6343 : node6288;
											assign node6288 = (inp[15]) ? node6320 : node6289;
												assign node6289 = (inp[4]) ? node6307 : node6290;
													assign node6290 = (inp[9]) ? node6294 : node6291;
														assign node6291 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node6294 = (inp[10]) ? node6302 : node6295;
															assign node6295 = (inp[8]) ? node6299 : node6296;
																assign node6296 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node6299 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node6302 = (inp[7]) ? 4'b1000 : node6303;
																assign node6303 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node6307 = (inp[9]) ? node6315 : node6308;
														assign node6308 = (inp[7]) ? node6312 : node6309;
															assign node6309 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node6312 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node6315 = (inp[7]) ? 4'b1110 : node6316;
															assign node6316 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node6320 = (inp[4]) ? node6330 : node6321;
													assign node6321 = (inp[9]) ? node6325 : node6322;
														assign node6322 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node6325 = (inp[8]) ? node6327 : 4'b1011;
															assign node6327 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node6330 = (inp[9]) ? node6338 : node6331;
														assign node6331 = (inp[10]) ? node6333 : 4'b1011;
															assign node6333 = (inp[8]) ? node6335 : 4'b1010;
																assign node6335 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node6338 = (inp[8]) ? node6340 : 4'b1101;
															assign node6340 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node6343 = (inp[15]) ? node6369 : node6344;
												assign node6344 = (inp[10]) ? node6350 : node6345;
													assign node6345 = (inp[8]) ? 4'b1011 : node6346;
														assign node6346 = (inp[7]) ? 4'b1110 : 4'b1011;
													assign node6350 = (inp[8]) ? node6360 : node6351;
														assign node6351 = (inp[7]) ? 4'b1010 : node6352;
															assign node6352 = (inp[9]) ? node6356 : node6353;
																assign node6353 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node6356 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node6360 = (inp[7]) ? node6362 : 4'b1110;
															assign node6362 = (inp[4]) ? node6366 : node6363;
																assign node6363 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node6366 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node6369 = (inp[4]) ? node6373 : node6370;
													assign node6370 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node6373 = (inp[9]) ? node6377 : node6374;
														assign node6374 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node6377 = (inp[10]) ? 4'b1101 : node6378;
															assign node6378 = (inp[8]) ? node6380 : 4'b1100;
																assign node6380 = (inp[7]) ? 4'b1101 : 4'b1100;
										assign node6384 = (inp[7]) ? node6430 : node6385;
											assign node6385 = (inp[8]) ? node6411 : node6386;
												assign node6386 = (inp[9]) ? node6400 : node6387;
													assign node6387 = (inp[4]) ? node6393 : node6388;
														assign node6388 = (inp[15]) ? 4'b1110 : node6389;
															assign node6389 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node6393 = (inp[3]) ? node6397 : node6394;
															assign node6394 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node6397 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node6400 = (inp[4]) ? node6408 : node6401;
														assign node6401 = (inp[15]) ? node6405 : node6402;
															assign node6402 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node6405 = (inp[10]) ? 4'b1000 : 4'b1010;
														assign node6408 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node6411 = (inp[3]) ? node6425 : node6412;
													assign node6412 = (inp[15]) ? node6422 : node6413;
														assign node6413 = (inp[10]) ? node6417 : node6414;
															assign node6414 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node6417 = (inp[9]) ? 4'b1001 : node6418;
																assign node6418 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node6422 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node6425 = (inp[4]) ? node6427 : 4'b1011;
														assign node6427 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node6430 = (inp[8]) ? node6450 : node6431;
												assign node6431 = (inp[3]) ? node6441 : node6432;
													assign node6432 = (inp[15]) ? node6434 : 4'b1001;
														assign node6434 = (inp[9]) ? node6438 : node6435;
															assign node6435 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node6438 = (inp[4]) ? 4'b1101 : 4'b1011;
													assign node6441 = (inp[15]) ? node6443 : 4'b1011;
														assign node6443 = (inp[10]) ? node6445 : 4'b1101;
															assign node6445 = (inp[9]) ? 4'b1001 : node6446;
																assign node6446 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node6450 = (inp[10]) ? node6466 : node6451;
													assign node6451 = (inp[3]) ? node6461 : node6452;
														assign node6452 = (inp[15]) ? node6456 : node6453;
															assign node6453 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node6456 = (inp[4]) ? node6458 : 4'b1010;
																assign node6458 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node6461 = (inp[9]) ? 4'b1100 : node6462;
															assign node6462 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node6466 = (inp[4]) ? node6472 : node6467;
														assign node6467 = (inp[9]) ? node6469 : 4'b1100;
															assign node6469 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node6472 = (inp[9]) ? node6474 : 4'b1010;
															assign node6474 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node6477 = (inp[7]) ? node6669 : node6478;
									assign node6478 = (inp[10]) ? node6566 : node6479;
										assign node6479 = (inp[4]) ? node6517 : node6480;
											assign node6480 = (inp[9]) ? node6498 : node6481;
												assign node6481 = (inp[8]) ? node6489 : node6482;
													assign node6482 = (inp[2]) ? 4'b1110 : node6483;
														assign node6483 = (inp[15]) ? 4'b1111 : node6484;
															assign node6484 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node6489 = (inp[2]) ? 4'b1111 : node6490;
														assign node6490 = (inp[15]) ? 4'b1110 : node6491;
															assign node6491 = (inp[3]) ? node6493 : 4'b1110;
																assign node6493 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node6498 = (inp[0]) ? node6506 : node6499;
													assign node6499 = (inp[2]) ? node6503 : node6500;
														assign node6500 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node6503 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node6506 = (inp[3]) ? node6512 : node6507;
														assign node6507 = (inp[2]) ? 4'b1001 : node6508;
															assign node6508 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node6512 = (inp[15]) ? 4'b1001 : node6513;
															assign node6513 = (inp[8]) ? 4'b1011 : 4'b1010;
											assign node6517 = (inp[9]) ? node6537 : node6518;
												assign node6518 = (inp[8]) ? node6530 : node6519;
													assign node6519 = (inp[2]) ? node6523 : node6520;
														assign node6520 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node6523 = (inp[15]) ? node6525 : 4'b1010;
															assign node6525 = (inp[0]) ? node6527 : 4'b1000;
																assign node6527 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node6530 = (inp[15]) ? node6532 : 4'b1001;
														assign node6532 = (inp[0]) ? node6534 : 4'b1001;
															assign node6534 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node6537 = (inp[0]) ? node6551 : node6538;
													assign node6538 = (inp[15]) ? node6542 : node6539;
														assign node6539 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node6542 = (inp[3]) ? node6546 : node6543;
															assign node6543 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node6546 = (inp[2]) ? 4'b1111 : node6547;
																assign node6547 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node6551 = (inp[15]) ? node6561 : node6552;
														assign node6552 = (inp[3]) ? node6554 : 4'b1110;
															assign node6554 = (inp[8]) ? node6558 : node6555;
																assign node6555 = (inp[2]) ? 4'b1110 : 4'b1111;
																assign node6558 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node6561 = (inp[2]) ? 4'b1100 : node6562;
															assign node6562 = (inp[8]) ? 4'b1100 : 4'b1101;
										assign node6566 = (inp[0]) ? node6616 : node6567;
											assign node6567 = (inp[15]) ? node6587 : node6568;
												assign node6568 = (inp[3]) ? node6576 : node6569;
													assign node6569 = (inp[9]) ? node6573 : node6570;
														assign node6570 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node6573 = (inp[2]) ? 4'b1101 : 4'b1001;
													assign node6576 = (inp[2]) ? node6584 : node6577;
														assign node6577 = (inp[8]) ? 4'b1100 : node6578;
															assign node6578 = (inp[4]) ? node6580 : 4'b1001;
																assign node6580 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node6584 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node6587 = (inp[9]) ? node6601 : node6588;
													assign node6588 = (inp[4]) ? node6598 : node6589;
														assign node6589 = (inp[3]) ? node6593 : node6590;
															assign node6590 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node6593 = (inp[8]) ? node6595 : 4'b1010;
																assign node6595 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node6598 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node6601 = (inp[4]) ? node6611 : node6602;
														assign node6602 = (inp[3]) ? node6606 : node6603;
															assign node6603 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node6606 = (inp[2]) ? 4'b1111 : node6607;
																assign node6607 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node6611 = (inp[8]) ? 4'b1011 : node6612;
															assign node6612 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node6616 = (inp[15]) ? node6638 : node6617;
												assign node6617 = (inp[4]) ? node6629 : node6618;
													assign node6618 = (inp[9]) ? 4'b1111 : node6619;
														assign node6619 = (inp[3]) ? node6625 : node6620;
															assign node6620 = (inp[8]) ? 4'b1001 : node6621;
																assign node6621 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node6625 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node6629 = (inp[9]) ? node6635 : node6630;
														assign node6630 = (inp[3]) ? 4'b1110 : node6631;
															assign node6631 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node6635 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node6638 = (inp[4]) ? node6656 : node6639;
													assign node6639 = (inp[3]) ? node6649 : node6640;
														assign node6640 = (inp[9]) ? 4'b1100 : node6641;
															assign node6641 = (inp[2]) ? node6645 : node6642;
																assign node6642 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node6645 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node6649 = (inp[2]) ? node6653 : node6650;
															assign node6650 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node6653 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node6656 = (inp[9]) ? node6662 : node6657;
														assign node6657 = (inp[8]) ? 4'b1100 : node6658;
															assign node6658 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node6662 = (inp[2]) ? node6666 : node6663;
															assign node6663 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node6666 = (inp[8]) ? 4'b1001 : 4'b1000;
									assign node6669 = (inp[3]) ? node6799 : node6670;
										assign node6670 = (inp[15]) ? node6732 : node6671;
											assign node6671 = (inp[2]) ? node6705 : node6672;
												assign node6672 = (inp[8]) ? node6694 : node6673;
													assign node6673 = (inp[10]) ? node6679 : node6674;
														assign node6674 = (inp[4]) ? 4'b1110 : node6675;
															assign node6675 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node6679 = (inp[0]) ? node6687 : node6680;
															assign node6680 = (inp[4]) ? node6684 : node6681;
																assign node6681 = (inp[9]) ? 4'b1100 : 4'b1010;
																assign node6684 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node6687 = (inp[9]) ? node6691 : node6688;
																assign node6688 = (inp[4]) ? 4'b1110 : 4'b1000;
																assign node6691 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node6694 = (inp[9]) ? 4'b1111 : node6695;
														assign node6695 = (inp[0]) ? node6701 : node6696;
															assign node6696 = (inp[4]) ? 4'b1101 : node6697;
																assign node6697 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node6701 = (inp[4]) ? 4'b1111 : 4'b1101;
												assign node6705 = (inp[8]) ? node6715 : node6706;
													assign node6706 = (inp[9]) ? node6708 : 4'b1011;
														assign node6708 = (inp[0]) ? 4'b1111 : node6709;
															assign node6709 = (inp[4]) ? node6711 : 4'b1101;
																assign node6711 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node6715 = (inp[10]) ? node6721 : node6716;
														assign node6716 = (inp[0]) ? 4'b1000 : node6717;
															assign node6717 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node6721 = (inp[9]) ? node6729 : node6722;
															assign node6722 = (inp[4]) ? node6726 : node6723;
																assign node6723 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node6726 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node6729 = (inp[4]) ? 4'b1010 : 4'b1110;
											assign node6732 = (inp[10]) ? node6768 : node6733;
												assign node6733 = (inp[0]) ? node6751 : node6734;
													assign node6734 = (inp[9]) ? node6744 : node6735;
														assign node6735 = (inp[4]) ? node6741 : node6736;
															assign node6736 = (inp[8]) ? 4'b1100 : node6737;
																assign node6737 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node6741 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node6744 = (inp[4]) ? 4'b1111 : node6745;
															assign node6745 = (inp[8]) ? node6747 : 4'b1001;
																assign node6747 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node6751 = (inp[9]) ? node6763 : node6752;
														assign node6752 = (inp[4]) ? node6758 : node6753;
															assign node6753 = (inp[8]) ? 4'b1111 : node6754;
																assign node6754 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node6758 = (inp[8]) ? node6760 : 4'b1011;
																assign node6760 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node6763 = (inp[4]) ? 4'b1101 : node6764;
															assign node6764 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node6768 = (inp[0]) ? node6786 : node6769;
													assign node6769 = (inp[4]) ? node6779 : node6770;
														assign node6770 = (inp[9]) ? node6776 : node6771;
															assign node6771 = (inp[2]) ? 4'b1001 : node6772;
																assign node6772 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node6776 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node6779 = (inp[9]) ? 4'b1010 : node6780;
															assign node6780 = (inp[8]) ? node6782 : 4'b1111;
																assign node6782 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node6786 = (inp[4]) ? node6794 : node6787;
														assign node6787 = (inp[9]) ? node6789 : 4'b1010;
															assign node6789 = (inp[8]) ? node6791 : 4'b1100;
																assign node6791 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node6794 = (inp[8]) ? 4'b1100 : node6795;
															assign node6795 = (inp[2]) ? 4'b1101 : 4'b1100;
										assign node6799 = (inp[9]) ? node6849 : node6800;
											assign node6800 = (inp[15]) ? node6828 : node6801;
												assign node6801 = (inp[0]) ? node6813 : node6802;
													assign node6802 = (inp[2]) ? node6808 : node6803;
														assign node6803 = (inp[8]) ? node6805 : 4'b1100;
															assign node6805 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node6808 = (inp[8]) ? 4'b1000 : node6809;
															assign node6809 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node6813 = (inp[2]) ? node6823 : node6814;
														assign node6814 = (inp[8]) ? node6820 : node6815;
															assign node6815 = (inp[10]) ? 4'b1010 : node6816;
																assign node6816 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node6820 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node6823 = (inp[10]) ? 4'b1111 : node6824;
															assign node6824 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node6828 = (inp[0]) ? node6832 : node6829;
													assign node6829 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node6832 = (inp[4]) ? node6840 : node6833;
														assign node6833 = (inp[10]) ? 4'b1000 : node6834;
															assign node6834 = (inp[8]) ? 4'b1100 : node6835;
																assign node6835 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node6840 = (inp[10]) ? 4'b1100 : node6841;
															assign node6841 = (inp[2]) ? node6845 : node6842;
																assign node6842 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node6845 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node6849 = (inp[2]) ? node6875 : node6850;
												assign node6850 = (inp[8]) ? node6862 : node6851;
													assign node6851 = (inp[15]) ? node6859 : node6852;
														assign node6852 = (inp[0]) ? node6854 : 4'b1000;
															assign node6854 = (inp[10]) ? 4'b1010 : node6855;
																assign node6855 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node6859 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node6862 = (inp[15]) ? node6868 : node6863;
														assign node6863 = (inp[10]) ? node6865 : 4'b1101;
															assign node6865 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node6868 = (inp[4]) ? node6872 : node6869;
															assign node6869 = (inp[10]) ? 4'b1111 : 4'b1011;
															assign node6872 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node6875 = (inp[8]) ? node6895 : node6876;
													assign node6876 = (inp[10]) ? node6888 : node6877;
														assign node6877 = (inp[4]) ? node6881 : node6878;
															assign node6878 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node6881 = (inp[15]) ? node6885 : node6882;
																assign node6882 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node6885 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node6888 = (inp[4]) ? 4'b1011 : node6889;
															assign node6889 = (inp[15]) ? node6891 : 4'b1111;
																assign node6891 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node6895 = (inp[0]) ? node6903 : node6896;
														assign node6896 = (inp[15]) ? node6898 : 4'b1000;
															assign node6898 = (inp[4]) ? 4'b1110 : node6899;
																assign node6899 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node6903 = (inp[15]) ? node6905 : 4'b1010;
															assign node6905 = (inp[4]) ? 4'b1000 : node6906;
																assign node6906 = (inp[10]) ? 4'b1100 : 4'b1000;
							assign node6910 = (inp[7]) ? node7298 : node6911;
								assign node6911 = (inp[2]) ? node7117 : node6912;
									assign node6912 = (inp[8]) ? node7016 : node6913;
										assign node6913 = (inp[9]) ? node6969 : node6914;
											assign node6914 = (inp[4]) ? node6940 : node6915;
												assign node6915 = (inp[10]) ? node6927 : node6916;
													assign node6916 = (inp[0]) ? node6922 : node6917;
														assign node6917 = (inp[3]) ? node6919 : 4'b1111;
															assign node6919 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node6922 = (inp[3]) ? node6924 : 4'b1101;
															assign node6924 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node6927 = (inp[12]) ? node6935 : node6928;
														assign node6928 = (inp[3]) ? node6930 : 4'b1111;
															assign node6930 = (inp[0]) ? node6932 : 4'b1111;
																assign node6932 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node6935 = (inp[3]) ? node6937 : 4'b1011;
															assign node6937 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node6940 = (inp[12]) ? node6954 : node6941;
													assign node6941 = (inp[15]) ? node6949 : node6942;
														assign node6942 = (inp[3]) ? node6946 : node6943;
															assign node6943 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node6946 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node6949 = (inp[0]) ? 4'b1001 : node6950;
															assign node6950 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node6954 = (inp[10]) ? node6964 : node6955;
														assign node6955 = (inp[3]) ? node6957 : 4'b1011;
															assign node6957 = (inp[0]) ? node6961 : node6958;
																assign node6958 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node6961 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node6964 = (inp[3]) ? node6966 : 4'b1111;
															assign node6966 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node6969 = (inp[4]) ? node6995 : node6970;
												assign node6970 = (inp[10]) ? node6978 : node6971;
													assign node6971 = (inp[3]) ? 4'b1001 : node6972;
														assign node6972 = (inp[15]) ? node6974 : 4'b1001;
															assign node6974 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node6978 = (inp[12]) ? node6984 : node6979;
														assign node6979 = (inp[3]) ? node6981 : 4'b1001;
															assign node6981 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node6984 = (inp[3]) ? node6990 : node6985;
															assign node6985 = (inp[15]) ? node6987 : 4'b1101;
																assign node6987 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node6990 = (inp[15]) ? 4'b1111 : node6991;
																assign node6991 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node6995 = (inp[10]) ? node7003 : node6996;
													assign node6996 = (inp[0]) ? node7000 : node6997;
														assign node6997 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node7000 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node7003 = (inp[12]) ? node7007 : node7004;
														assign node7004 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node7007 = (inp[3]) ? node7009 : 4'b1001;
															assign node7009 = (inp[0]) ? node7013 : node7010;
																assign node7010 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node7013 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node7016 = (inp[10]) ? node7060 : node7017;
											assign node7017 = (inp[0]) ? node7037 : node7018;
												assign node7018 = (inp[12]) ? node7028 : node7019;
													assign node7019 = (inp[15]) ? node7025 : node7020;
														assign node7020 = (inp[9]) ? 4'b1100 : node7021;
															assign node7021 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node7025 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node7028 = (inp[15]) ? node7034 : node7029;
														assign node7029 = (inp[4]) ? node7031 : 4'b1110;
															assign node7031 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node7034 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node7037 = (inp[9]) ? node7045 : node7038;
													assign node7038 = (inp[4]) ? 4'b1010 : node7039;
														assign node7039 = (inp[12]) ? 4'b1110 : node7040;
															assign node7040 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node7045 = (inp[4]) ? node7057 : node7046;
														assign node7046 = (inp[12]) ? node7052 : node7047;
															assign node7047 = (inp[15]) ? 4'b1010 : node7048;
																assign node7048 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node7052 = (inp[3]) ? node7054 : 4'b1000;
																assign node7054 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node7057 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node7060 = (inp[4]) ? node7098 : node7061;
												assign node7061 = (inp[9]) ? node7083 : node7062;
													assign node7062 = (inp[12]) ? node7070 : node7063;
														assign node7063 = (inp[0]) ? 4'b1110 : node7064;
															assign node7064 = (inp[3]) ? node7066 : 4'b1100;
																assign node7066 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node7070 = (inp[15]) ? node7078 : node7071;
															assign node7071 = (inp[0]) ? node7075 : node7072;
																assign node7072 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node7075 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node7078 = (inp[3]) ? 4'b1010 : node7079;
																assign node7079 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node7083 = (inp[12]) ? node7091 : node7084;
														assign node7084 = (inp[3]) ? node7086 : 4'b1010;
															assign node7086 = (inp[15]) ? node7088 : 4'b1000;
																assign node7088 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node7091 = (inp[0]) ? node7095 : node7092;
															assign node7092 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node7095 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node7098 = (inp[9]) ? node7110 : node7099;
													assign node7099 = (inp[12]) ? node7105 : node7100;
														assign node7100 = (inp[0]) ? node7102 : 4'b1000;
															assign node7102 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node7105 = (inp[0]) ? node7107 : 4'b1100;
															assign node7107 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node7110 = (inp[12]) ? node7112 : 4'b1110;
														assign node7112 = (inp[15]) ? node7114 : 4'b1000;
															assign node7114 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node7117 = (inp[8]) ? node7215 : node7118;
										assign node7118 = (inp[0]) ? node7166 : node7119;
											assign node7119 = (inp[15]) ? node7139 : node7120;
												assign node7120 = (inp[3]) ? node7130 : node7121;
													assign node7121 = (inp[9]) ? node7125 : node7122;
														assign node7122 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node7125 = (inp[12]) ? node7127 : 4'b1100;
															assign node7127 = (inp[10]) ? 4'b1100 : 4'b1010;
													assign node7130 = (inp[4]) ? node7132 : 4'b1100;
														assign node7132 = (inp[10]) ? node7136 : node7133;
															assign node7133 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node7136 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node7139 = (inp[3]) ? node7157 : node7140;
													assign node7140 = (inp[9]) ? node7148 : node7141;
														assign node7141 = (inp[4]) ? node7143 : 4'b1100;
															assign node7143 = (inp[10]) ? node7145 : 4'b1000;
																assign node7145 = (inp[12]) ? 4'b1110 : 4'b1000;
														assign node7148 = (inp[4]) ? node7154 : node7149;
															assign node7149 = (inp[12]) ? node7151 : 4'b1000;
																assign node7151 = (inp[10]) ? 4'b1110 : 4'b1000;
															assign node7154 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node7157 = (inp[9]) ? node7161 : node7158;
														assign node7158 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node7161 = (inp[4]) ? 4'b1110 : node7162;
															assign node7162 = (inp[10]) ? 4'b1110 : 4'b1010;
											assign node7166 = (inp[15]) ? node7194 : node7167;
												assign node7167 = (inp[3]) ? node7185 : node7168;
													assign node7168 = (inp[10]) ? node7174 : node7169;
														assign node7169 = (inp[4]) ? 4'b1000 : node7170;
															assign node7170 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node7174 = (inp[12]) ? node7178 : node7175;
															assign node7175 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node7178 = (inp[4]) ? node7182 : node7179;
																assign node7179 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node7182 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node7185 = (inp[12]) ? node7191 : node7186;
														assign node7186 = (inp[4]) ? node7188 : 4'b1010;
															assign node7188 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node7191 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node7194 = (inp[3]) ? node7204 : node7195;
													assign node7195 = (inp[4]) ? node7197 : 4'b1010;
														assign node7197 = (inp[9]) ? 4'b1100 : node7198;
															assign node7198 = (inp[10]) ? node7200 : 4'b1010;
																assign node7200 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node7204 = (inp[4]) ? node7210 : node7205;
														assign node7205 = (inp[12]) ? 4'b1100 : node7206;
															assign node7206 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node7210 = (inp[9]) ? node7212 : 4'b1000;
															assign node7212 = (inp[10]) ? 4'b1000 : 4'b1100;
										assign node7215 = (inp[4]) ? node7259 : node7216;
											assign node7216 = (inp[9]) ? node7236 : node7217;
												assign node7217 = (inp[10]) ? node7231 : node7218;
													assign node7218 = (inp[0]) ? node7226 : node7219;
														assign node7219 = (inp[15]) ? node7223 : node7220;
															assign node7220 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node7223 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node7226 = (inp[15]) ? 4'b0111 : node7227;
															assign node7227 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node7231 = (inp[12]) ? 4'b0001 : node7232;
														assign node7232 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node7236 = (inp[10]) ? node7252 : node7237;
													assign node7237 = (inp[15]) ? node7247 : node7238;
														assign node7238 = (inp[12]) ? 4'b0001 : node7239;
															assign node7239 = (inp[3]) ? node7243 : node7240;
																assign node7240 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node7243 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node7247 = (inp[0]) ? node7249 : 4'b0011;
															assign node7249 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node7252 = (inp[12]) ? node7254 : 4'b0001;
														assign node7254 = (inp[0]) ? node7256 : 4'b0101;
															assign node7256 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node7259 = (inp[9]) ? node7289 : node7260;
												assign node7260 = (inp[12]) ? node7272 : node7261;
													assign node7261 = (inp[3]) ? node7267 : node7262;
														assign node7262 = (inp[15]) ? node7264 : 4'b0011;
															assign node7264 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node7267 = (inp[0]) ? node7269 : 4'b0001;
															assign node7269 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node7272 = (inp[10]) ? node7282 : node7273;
														assign node7273 = (inp[15]) ? node7275 : 4'b0001;
															assign node7275 = (inp[3]) ? node7279 : node7276;
																assign node7276 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node7279 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node7282 = (inp[15]) ? node7286 : node7283;
															assign node7283 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node7286 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node7289 = (inp[10]) ? node7295 : node7290;
													assign node7290 = (inp[15]) ? node7292 : 4'b0111;
														assign node7292 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node7295 = (inp[12]) ? 4'b0011 : 4'b0111;
								assign node7298 = (inp[8]) ? node7486 : node7299;
									assign node7299 = (inp[2]) ? node7407 : node7300;
										assign node7300 = (inp[10]) ? node7354 : node7301;
											assign node7301 = (inp[12]) ? node7327 : node7302;
												assign node7302 = (inp[15]) ? node7314 : node7303;
													assign node7303 = (inp[3]) ? node7309 : node7304;
														assign node7304 = (inp[0]) ? node7306 : 4'b1010;
															assign node7306 = (inp[4]) ? 4'b1110 : 4'b1100;
														assign node7309 = (inp[9]) ? 4'b1100 : node7310;
															assign node7310 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node7314 = (inp[9]) ? node7324 : node7315;
														assign node7315 = (inp[4]) ? node7317 : 4'b1100;
															assign node7317 = (inp[3]) ? node7321 : node7318;
																assign node7318 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node7321 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node7324 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node7327 = (inp[0]) ? node7341 : node7328;
													assign node7328 = (inp[9]) ? node7334 : node7329;
														assign node7329 = (inp[3]) ? 4'b1100 : node7330;
															assign node7330 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node7334 = (inp[4]) ? 4'b1110 : node7335;
															assign node7335 = (inp[15]) ? node7337 : 4'b1010;
																assign node7337 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node7341 = (inp[15]) ? node7349 : node7342;
														assign node7342 = (inp[4]) ? node7344 : 4'b1000;
															assign node7344 = (inp[9]) ? 4'b1110 : node7345;
																assign node7345 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node7349 = (inp[4]) ? node7351 : 4'b1110;
															assign node7351 = (inp[9]) ? 4'b1100 : 4'b1000;
											assign node7354 = (inp[9]) ? node7374 : node7355;
												assign node7355 = (inp[12]) ? node7363 : node7356;
													assign node7356 = (inp[15]) ? node7358 : 4'b1110;
														assign node7358 = (inp[3]) ? 4'b1110 : node7359;
															assign node7359 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node7363 = (inp[4]) ? node7367 : node7364;
														assign node7364 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node7367 = (inp[3]) ? 4'b1100 : node7368;
															assign node7368 = (inp[15]) ? 4'b1110 : node7369;
																assign node7369 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node7374 = (inp[3]) ? node7396 : node7375;
													assign node7375 = (inp[15]) ? node7383 : node7376;
														assign node7376 = (inp[0]) ? node7378 : 4'b1010;
															assign node7378 = (inp[12]) ? node7380 : 4'b1110;
																assign node7380 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node7383 = (inp[0]) ? node7391 : node7384;
															assign node7384 = (inp[4]) ? node7388 : node7385;
																assign node7385 = (inp[12]) ? 4'b1110 : 4'b1000;
																assign node7388 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node7391 = (inp[4]) ? 4'b1100 : node7392;
																assign node7392 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node7396 = (inp[0]) ? node7402 : node7397;
														assign node7397 = (inp[4]) ? 4'b1000 : node7398;
															assign node7398 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node7402 = (inp[15]) ? 4'b1000 : node7403;
															assign node7403 = (inp[4]) ? 4'b1110 : 4'b1010;
										assign node7407 = (inp[4]) ? node7447 : node7408;
											assign node7408 = (inp[9]) ? node7426 : node7409;
												assign node7409 = (inp[12]) ? node7419 : node7410;
													assign node7410 = (inp[15]) ? node7412 : 4'b0101;
														assign node7412 = (inp[0]) ? node7416 : node7413;
															assign node7413 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node7416 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node7419 = (inp[10]) ? 4'b0011 : node7420;
														assign node7420 = (inp[15]) ? 4'b0111 : node7421;
															assign node7421 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node7426 = (inp[10]) ? node7440 : node7427;
													assign node7427 = (inp[0]) ? node7433 : node7428;
														assign node7428 = (inp[3]) ? node7430 : 4'b0001;
															assign node7430 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node7433 = (inp[3]) ? node7437 : node7434;
															assign node7434 = (inp[12]) ? 4'b0011 : 4'b0001;
															assign node7437 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node7440 = (inp[12]) ? node7442 : 4'b0011;
														assign node7442 = (inp[15]) ? 4'b0111 : node7443;
															assign node7443 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node7447 = (inp[9]) ? node7469 : node7448;
												assign node7448 = (inp[12]) ? node7462 : node7449;
													assign node7449 = (inp[3]) ? node7457 : node7450;
														assign node7450 = (inp[15]) ? node7454 : node7451;
															assign node7451 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node7454 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node7457 = (inp[0]) ? node7459 : 4'b0011;
															assign node7459 = (inp[10]) ? 4'b0011 : 4'b0001;
													assign node7462 = (inp[10]) ? 4'b0101 : node7463;
														assign node7463 = (inp[3]) ? 4'b0011 : node7464;
															assign node7464 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node7469 = (inp[12]) ? node7477 : node7470;
													assign node7470 = (inp[15]) ? node7474 : node7471;
														assign node7471 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node7474 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node7477 = (inp[10]) ? node7479 : 4'b0101;
														assign node7479 = (inp[15]) ? node7483 : node7480;
															assign node7480 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node7483 = (inp[0]) ? 4'b0001 : 4'b0011;
									assign node7486 = (inp[2]) ? node7606 : node7487;
										assign node7487 = (inp[10]) ? node7543 : node7488;
											assign node7488 = (inp[4]) ? node7522 : node7489;
												assign node7489 = (inp[9]) ? node7507 : node7490;
													assign node7490 = (inp[12]) ? node7500 : node7491;
														assign node7491 = (inp[0]) ? 4'b0101 : node7492;
															assign node7492 = (inp[15]) ? node7496 : node7493;
																assign node7493 = (inp[3]) ? 4'b0101 : 4'b0111;
																assign node7496 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node7500 = (inp[0]) ? node7502 : 4'b0101;
															assign node7502 = (inp[3]) ? node7504 : 4'b0111;
																assign node7504 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node7507 = (inp[15]) ? 4'b0001 : node7508;
														assign node7508 = (inp[12]) ? node7514 : node7509;
															assign node7509 = (inp[0]) ? node7511 : 4'b0001;
																assign node7511 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node7514 = (inp[3]) ? node7518 : node7515;
																assign node7515 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node7518 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node7522 = (inp[9]) ? node7534 : node7523;
													assign node7523 = (inp[3]) ? node7529 : node7524;
														assign node7524 = (inp[0]) ? 4'b0011 : node7525;
															assign node7525 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node7529 = (inp[15]) ? node7531 : 4'b0001;
															assign node7531 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node7534 = (inp[12]) ? node7536 : 4'b0111;
														assign node7536 = (inp[0]) ? node7540 : node7537;
															assign node7537 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node7540 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node7543 = (inp[3]) ? node7579 : node7544;
												assign node7544 = (inp[9]) ? node7562 : node7545;
													assign node7545 = (inp[4]) ? node7553 : node7546;
														assign node7546 = (inp[15]) ? node7550 : node7547;
															assign node7547 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node7550 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node7553 = (inp[12]) ? node7555 : 4'b0011;
															assign node7555 = (inp[15]) ? node7559 : node7556;
																assign node7556 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node7559 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node7562 = (inp[15]) ? node7574 : node7563;
														assign node7563 = (inp[12]) ? node7569 : node7564;
															assign node7564 = (inp[4]) ? 4'b0101 : node7565;
																assign node7565 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node7569 = (inp[4]) ? 4'b0011 : node7570;
																assign node7570 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node7574 = (inp[12]) ? node7576 : 4'b0111;
															assign node7576 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node7579 = (inp[0]) ? node7591 : node7580;
													assign node7580 = (inp[15]) ? node7588 : node7581;
														assign node7581 = (inp[4]) ? 4'b0001 : node7582;
															assign node7582 = (inp[12]) ? 4'b0101 : node7583;
																assign node7583 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node7588 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node7591 = (inp[15]) ? 4'b0101 : node7592;
														assign node7592 = (inp[12]) ? node7598 : node7593;
															assign node7593 = (inp[4]) ? 4'b0011 : node7594;
																assign node7594 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node7598 = (inp[4]) ? node7602 : node7599;
																assign node7599 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node7602 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node7606 = (inp[12]) ? node7640 : node7607;
											assign node7607 = (inp[15]) ? node7629 : node7608;
												assign node7608 = (inp[0]) ? node7622 : node7609;
													assign node7609 = (inp[3]) ? node7617 : node7610;
														assign node7610 = (inp[4]) ? node7614 : node7611;
															assign node7611 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node7614 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node7617 = (inp[4]) ? 4'b0000 : node7618;
															assign node7618 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node7622 = (inp[9]) ? 4'b0110 : node7623;
														assign node7623 = (inp[4]) ? node7625 : 4'b0110;
															assign node7625 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node7629 = (inp[4]) ? node7635 : node7630;
													assign node7630 = (inp[9]) ? 4'b0010 : node7631;
														assign node7631 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node7635 = (inp[9]) ? node7637 : 4'b0000;
														assign node7637 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node7640 = (inp[0]) ? node7676 : node7641;
												assign node7641 = (inp[15]) ? node7657 : node7642;
													assign node7642 = (inp[10]) ? node7648 : node7643;
														assign node7643 = (inp[3]) ? 4'b0000 : node7644;
															assign node7644 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node7648 = (inp[4]) ? node7654 : node7649;
															assign node7649 = (inp[9]) ? 4'b0100 : node7650;
																assign node7650 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node7654 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node7657 = (inp[3]) ? node7663 : node7658;
														assign node7658 = (inp[10]) ? 4'b0110 : node7659;
															assign node7659 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node7663 = (inp[10]) ? node7669 : node7664;
															assign node7664 = (inp[4]) ? 4'b0010 : node7665;
																assign node7665 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node7669 = (inp[4]) ? node7673 : node7670;
																assign node7670 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node7673 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node7676 = (inp[15]) ? node7686 : node7677;
													assign node7677 = (inp[3]) ? node7679 : 4'b0000;
														assign node7679 = (inp[10]) ? 4'b0010 : node7680;
															assign node7680 = (inp[4]) ? 4'b0010 : node7681;
																assign node7681 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node7686 = (inp[9]) ? node7694 : node7687;
														assign node7687 = (inp[3]) ? node7689 : 4'b0010;
															assign node7689 = (inp[10]) ? 4'b0000 : node7690;
																assign node7690 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node7694 = (inp[4]) ? node7698 : node7695;
															assign node7695 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node7698 = (inp[10]) ? 4'b0000 : 4'b0100;
						assign node7701 = (inp[1]) ? node8529 : node7702;
							assign node7702 = (inp[7]) ? node8114 : node7703;
								assign node7703 = (inp[2]) ? node7897 : node7704;
									assign node7704 = (inp[8]) ? node7804 : node7705;
										assign node7705 = (inp[0]) ? node7765 : node7706;
											assign node7706 = (inp[15]) ? node7734 : node7707;
												assign node7707 = (inp[3]) ? node7723 : node7708;
													assign node7708 = (inp[4]) ? node7716 : node7709;
														assign node7709 = (inp[9]) ? 4'b0011 : node7710;
															assign node7710 = (inp[12]) ? node7712 : 4'b0111;
																assign node7712 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node7716 = (inp[12]) ? node7718 : 4'b0101;
															assign node7718 = (inp[10]) ? node7720 : 4'b0011;
																assign node7720 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node7723 = (inp[4]) ? node7729 : node7724;
														assign node7724 = (inp[12]) ? node7726 : 4'b0101;
															assign node7726 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node7729 = (inp[9]) ? node7731 : 4'b0001;
															assign node7731 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node7734 = (inp[3]) ? node7748 : node7735;
													assign node7735 = (inp[9]) ? node7739 : node7736;
														assign node7736 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node7739 = (inp[10]) ? node7743 : node7740;
															assign node7740 = (inp[4]) ? 4'b0111 : 4'b0001;
															assign node7743 = (inp[4]) ? node7745 : 4'b0111;
																assign node7745 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node7748 = (inp[12]) ? node7756 : node7749;
														assign node7749 = (inp[10]) ? node7751 : 4'b0011;
															assign node7751 = (inp[9]) ? node7753 : 4'b0011;
																assign node7753 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node7756 = (inp[4]) ? node7758 : 4'b0111;
															assign node7758 = (inp[10]) ? node7762 : node7759;
																assign node7759 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node7762 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node7765 = (inp[15]) ? node7785 : node7766;
												assign node7766 = (inp[3]) ? node7776 : node7767;
													assign node7767 = (inp[12]) ? node7769 : 4'b0001;
														assign node7769 = (inp[9]) ? node7773 : node7770;
															assign node7770 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node7773 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node7776 = (inp[9]) ? node7782 : node7777;
														assign node7777 = (inp[4]) ? 4'b0011 : node7778;
															assign node7778 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node7782 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node7785 = (inp[3]) ? node7795 : node7786;
													assign node7786 = (inp[10]) ? node7790 : node7787;
														assign node7787 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node7790 = (inp[4]) ? 4'b0101 : node7791;
															assign node7791 = (inp[12]) ? 4'b0101 : 4'b0111;
													assign node7795 = (inp[10]) ? 4'b0001 : node7796;
														assign node7796 = (inp[9]) ? node7800 : node7797;
															assign node7797 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node7800 = (inp[4]) ? 4'b0101 : 4'b0001;
										assign node7804 = (inp[4]) ? node7850 : node7805;
											assign node7805 = (inp[9]) ? node7829 : node7806;
												assign node7806 = (inp[12]) ? node7820 : node7807;
													assign node7807 = (inp[3]) ? node7813 : node7808;
														assign node7808 = (inp[10]) ? node7810 : 4'b0100;
															assign node7810 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node7813 = (inp[0]) ? node7817 : node7814;
															assign node7814 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node7817 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node7820 = (inp[10]) ? node7826 : node7821;
														assign node7821 = (inp[0]) ? 4'b0110 : node7822;
															assign node7822 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node7826 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node7829 = (inp[10]) ? node7837 : node7830;
													assign node7830 = (inp[0]) ? node7832 : 4'b0010;
														assign node7832 = (inp[15]) ? 4'b0000 : node7833;
															assign node7833 = (inp[12]) ? 4'b0010 : 4'b0000;
													assign node7837 = (inp[12]) ? node7841 : node7838;
														assign node7838 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node7841 = (inp[3]) ? node7843 : 4'b0110;
															assign node7843 = (inp[15]) ? node7847 : node7844;
																assign node7844 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node7847 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node7850 = (inp[9]) ? node7870 : node7851;
												assign node7851 = (inp[12]) ? node7861 : node7852;
													assign node7852 = (inp[15]) ? node7858 : node7853;
														assign node7853 = (inp[3]) ? node7855 : 4'b0000;
															assign node7855 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node7858 = (inp[10]) ? 4'b0000 : 4'b0010;
													assign node7861 = (inp[10]) ? 4'b0110 : node7862;
														assign node7862 = (inp[0]) ? node7864 : 4'b0000;
															assign node7864 = (inp[15]) ? node7866 : 4'b0010;
																assign node7866 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node7870 = (inp[10]) ? node7884 : node7871;
													assign node7871 = (inp[12]) ? node7873 : 4'b0110;
														assign node7873 = (inp[3]) ? node7879 : node7874;
															assign node7874 = (inp[15]) ? 4'b0110 : node7875;
																assign node7875 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node7879 = (inp[0]) ? node7881 : 4'b0110;
																assign node7881 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node7884 = (inp[12]) ? node7892 : node7885;
														assign node7885 = (inp[0]) ? node7889 : node7886;
															assign node7886 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node7889 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node7892 = (inp[15]) ? 4'b0010 : node7893;
															assign node7893 = (inp[0]) ? 4'b0010 : 4'b0000;
									assign node7897 = (inp[8]) ? node8017 : node7898;
										assign node7898 = (inp[12]) ? node7958 : node7899;
											assign node7899 = (inp[4]) ? node7929 : node7900;
												assign node7900 = (inp[9]) ? node7914 : node7901;
													assign node7901 = (inp[15]) ? node7907 : node7902;
														assign node7902 = (inp[0]) ? node7904 : 4'b0100;
															assign node7904 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node7907 = (inp[0]) ? node7911 : node7908;
															assign node7908 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node7911 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node7914 = (inp[15]) ? node7922 : node7915;
														assign node7915 = (inp[10]) ? node7917 : 4'b0000;
															assign node7917 = (inp[0]) ? 4'b0000 : node7918;
																assign node7918 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node7922 = (inp[3]) ? node7926 : node7923;
															assign node7923 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node7926 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node7929 = (inp[9]) ? node7947 : node7930;
													assign node7930 = (inp[10]) ? node7942 : node7931;
														assign node7931 = (inp[3]) ? node7937 : node7932;
															assign node7932 = (inp[15]) ? node7934 : 4'b0010;
																assign node7934 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node7937 = (inp[0]) ? 4'b0000 : node7938;
																assign node7938 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node7942 = (inp[3]) ? 4'b0010 : node7943;
															assign node7943 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node7947 = (inp[3]) ? node7953 : node7948;
														assign node7948 = (inp[15]) ? 4'b0110 : node7949;
															assign node7949 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node7953 = (inp[0]) ? node7955 : 4'b0100;
															assign node7955 = (inp[10]) ? 4'b0110 : 4'b0100;
											assign node7958 = (inp[9]) ? node7984 : node7959;
												assign node7959 = (inp[10]) ? node7977 : node7960;
													assign node7960 = (inp[4]) ? node7964 : node7961;
														assign node7961 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node7964 = (inp[3]) ? node7972 : node7965;
															assign node7965 = (inp[15]) ? node7969 : node7966;
																assign node7966 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node7969 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node7972 = (inp[15]) ? node7974 : 4'b0010;
																assign node7974 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node7977 = (inp[4]) ? 4'b0110 : node7978;
														assign node7978 = (inp[0]) ? 4'b0010 : node7979;
															assign node7979 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node7984 = (inp[0]) ? node8006 : node7985;
													assign node7985 = (inp[15]) ? node7995 : node7986;
														assign node7986 = (inp[10]) ? node7992 : node7987;
															assign node7987 = (inp[3]) ? node7989 : 4'b0010;
																assign node7989 = (inp[4]) ? 4'b0100 : 4'b0000;
															assign node7992 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node7995 = (inp[3]) ? node8001 : node7996;
															assign node7996 = (inp[10]) ? node7998 : 4'b0000;
																assign node7998 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node8001 = (inp[10]) ? 4'b0110 : node8002;
																assign node8002 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node8006 = (inp[15]) ? node8014 : node8007;
														assign node8007 = (inp[3]) ? 4'b0010 : node8008;
															assign node8008 = (inp[4]) ? node8010 : 4'b0110;
																assign node8010 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node8014 = (inp[4]) ? 4'b0100 : 4'b0010;
										assign node8017 = (inp[12]) ? node8073 : node8018;
											assign node8018 = (inp[4]) ? node8046 : node8019;
												assign node8019 = (inp[9]) ? node8029 : node8020;
													assign node8020 = (inp[15]) ? node8022 : 4'b0111;
														assign node8022 = (inp[0]) ? node8026 : node8023;
															assign node8023 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node8026 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node8029 = (inp[10]) ? node8037 : node8030;
														assign node8030 = (inp[0]) ? 4'b0011 : node8031;
															assign node8031 = (inp[15]) ? node8033 : 4'b0011;
																assign node8033 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node8037 = (inp[15]) ? 4'b0011 : node8038;
															assign node8038 = (inp[3]) ? node8042 : node8039;
																assign node8039 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node8042 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node8046 = (inp[9]) ? node8068 : node8047;
													assign node8047 = (inp[15]) ? node8063 : node8048;
														assign node8048 = (inp[10]) ? node8056 : node8049;
															assign node8049 = (inp[0]) ? node8053 : node8050;
																assign node8050 = (inp[3]) ? 4'b0001 : 4'b0011;
																assign node8053 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node8056 = (inp[0]) ? node8060 : node8057;
																assign node8057 = (inp[3]) ? 4'b0001 : 4'b0011;
																assign node8060 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node8063 = (inp[3]) ? node8065 : 4'b0001;
															assign node8065 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node8068 = (inp[10]) ? 4'b0101 : node8069;
														assign node8069 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node8073 = (inp[4]) ? node8099 : node8074;
												assign node8074 = (inp[15]) ? node8088 : node8075;
													assign node8075 = (inp[9]) ? node8081 : node8076;
														assign node8076 = (inp[3]) ? 4'b0001 : node8077;
															assign node8077 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node8081 = (inp[10]) ? 4'b0101 : node8082;
															assign node8082 = (inp[0]) ? node8084 : 4'b0001;
																assign node8084 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node8088 = (inp[10]) ? node8096 : node8089;
														assign node8089 = (inp[9]) ? node8093 : node8090;
															assign node8090 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node8093 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node8096 = (inp[0]) ? 4'b0011 : 4'b0111;
												assign node8099 = (inp[15]) ? node8103 : node8100;
													assign node8100 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node8103 = (inp[0]) ? node8105 : 4'b0111;
														assign node8105 = (inp[3]) ? 4'b0001 : node8106;
															assign node8106 = (inp[9]) ? node8110 : node8107;
																assign node8107 = (inp[10]) ? 4'b0101 : 4'b0011;
																assign node8110 = (inp[10]) ? 4'b0001 : 4'b0101;
								assign node8114 = (inp[0]) ? node8320 : node8115;
									assign node8115 = (inp[15]) ? node8217 : node8116;
										assign node8116 = (inp[3]) ? node8174 : node8117;
											assign node8117 = (inp[4]) ? node8145 : node8118;
												assign node8118 = (inp[9]) ? node8136 : node8119;
													assign node8119 = (inp[12]) ? node8133 : node8120;
														assign node8120 = (inp[10]) ? node8126 : node8121;
															assign node8121 = (inp[2]) ? node8123 : 4'b0110;
																assign node8123 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node8126 = (inp[2]) ? node8130 : node8127;
																assign node8127 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node8130 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node8133 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node8136 = (inp[10]) ? node8142 : node8137;
														assign node8137 = (inp[8]) ? node8139 : 4'b0010;
															assign node8139 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node8142 = (inp[12]) ? 4'b0100 : 4'b0011;
												assign node8145 = (inp[9]) ? node8161 : node8146;
													assign node8146 = (inp[12]) ? node8154 : node8147;
														assign node8147 = (inp[10]) ? node8149 : 4'b0010;
															assign node8149 = (inp[2]) ? 4'b0011 : node8150;
																assign node8150 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node8154 = (inp[10]) ? node8156 : 4'b0010;
															assign node8156 = (inp[2]) ? 4'b0101 : node8157;
																assign node8157 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node8161 = (inp[10]) ? node8167 : node8162;
														assign node8162 = (inp[8]) ? node8164 : 4'b0100;
															assign node8164 = (inp[12]) ? 4'b0101 : 4'b0100;
														assign node8167 = (inp[12]) ? 4'b0001 : node8168;
															assign node8168 = (inp[2]) ? node8170 : 4'b0101;
																assign node8170 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node8174 = (inp[4]) ? node8186 : node8175;
												assign node8175 = (inp[9]) ? node8179 : node8176;
													assign node8176 = (inp[12]) ? 4'b0101 : 4'b0100;
													assign node8179 = (inp[8]) ? 4'b0000 : node8180;
														assign node8180 = (inp[2]) ? 4'b0101 : node8181;
															assign node8181 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node8186 = (inp[9]) ? node8204 : node8187;
													assign node8187 = (inp[12]) ? node8195 : node8188;
														assign node8188 = (inp[8]) ? node8192 : node8189;
															assign node8189 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node8192 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node8195 = (inp[10]) ? node8199 : node8196;
															assign node8196 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node8199 = (inp[8]) ? 4'b0100 : node8200;
																assign node8200 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node8204 = (inp[12]) ? node8212 : node8205;
														assign node8205 = (inp[10]) ? node8207 : 4'b0100;
															assign node8207 = (inp[2]) ? node8209 : 4'b0101;
																assign node8209 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node8212 = (inp[10]) ? node8214 : 4'b0100;
															assign node8214 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node8217 = (inp[3]) ? node8263 : node8218;
											assign node8218 = (inp[4]) ? node8238 : node8219;
												assign node8219 = (inp[9]) ? node8227 : node8220;
													assign node8220 = (inp[2]) ? node8224 : node8221;
														assign node8221 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node8224 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node8227 = (inp[10]) ? node8235 : node8228;
														assign node8228 = (inp[12]) ? node8232 : node8229;
															assign node8229 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node8232 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node8235 = (inp[12]) ? 4'b0111 : 4'b0001;
												assign node8238 = (inp[9]) ? node8252 : node8239;
													assign node8239 = (inp[10]) ? node8247 : node8240;
														assign node8240 = (inp[12]) ? node8244 : node8241;
															assign node8241 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node8244 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node8247 = (inp[12]) ? 4'b0110 : node8248;
															assign node8248 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node8252 = (inp[12]) ? node8254 : 4'b0110;
														assign node8254 = (inp[10]) ? node8260 : node8255;
															assign node8255 = (inp[8]) ? 4'b0111 : node8256;
																assign node8256 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node8260 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node8263 = (inp[9]) ? node8293 : node8264;
												assign node8264 = (inp[4]) ? node8278 : node8265;
													assign node8265 = (inp[10]) ? node8273 : node8266;
														assign node8266 = (inp[8]) ? node8270 : node8267;
															assign node8267 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node8270 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node8273 = (inp[12]) ? 4'b0010 : node8274;
															assign node8274 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node8278 = (inp[12]) ? node8286 : node8279;
														assign node8279 = (inp[2]) ? node8283 : node8280;
															assign node8280 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node8283 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node8286 = (inp[10]) ? node8288 : 4'b0010;
															assign node8288 = (inp[2]) ? node8290 : 4'b0110;
																assign node8290 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node8293 = (inp[4]) ? node8303 : node8294;
													assign node8294 = (inp[8]) ? node8300 : node8295;
														assign node8295 = (inp[2]) ? 4'b0011 : node8296;
															assign node8296 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node8300 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node8303 = (inp[12]) ? node8311 : node8304;
														assign node8304 = (inp[10]) ? node8306 : 4'b0110;
															assign node8306 = (inp[8]) ? 4'b0111 : node8307;
																assign node8307 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node8311 = (inp[10]) ? node8315 : node8312;
															assign node8312 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node8315 = (inp[8]) ? 4'b0011 : node8316;
																assign node8316 = (inp[2]) ? 4'b0011 : 4'b0010;
									assign node8320 = (inp[15]) ? node8414 : node8321;
										assign node8321 = (inp[3]) ? node8375 : node8322;
											assign node8322 = (inp[9]) ? node8356 : node8323;
												assign node8323 = (inp[4]) ? node8341 : node8324;
													assign node8324 = (inp[10]) ? node8330 : node8325;
														assign node8325 = (inp[8]) ? node8327 : 4'b0100;
															assign node8327 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node8330 = (inp[12]) ? node8334 : node8331;
															assign node8331 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node8334 = (inp[2]) ? node8338 : node8335;
																assign node8335 = (inp[8]) ? 4'b0001 : 4'b0000;
																assign node8338 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node8341 = (inp[10]) ? node8353 : node8342;
														assign node8342 = (inp[12]) ? node8348 : node8343;
															assign node8343 = (inp[8]) ? 4'b0000 : node8344;
																assign node8344 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node8348 = (inp[8]) ? 4'b0001 : node8349;
																assign node8349 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node8353 = (inp[8]) ? 4'b0001 : 4'b0110;
												assign node8356 = (inp[4]) ? node8364 : node8357;
													assign node8357 = (inp[10]) ? node8359 : 4'b0000;
														assign node8359 = (inp[12]) ? 4'b0111 : node8360;
															assign node8360 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node8364 = (inp[8]) ? node8368 : node8365;
														assign node8365 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node8368 = (inp[2]) ? 4'b0110 : node8369;
															assign node8369 = (inp[12]) ? node8371 : 4'b0111;
																assign node8371 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node8375 = (inp[4]) ? node8387 : node8376;
												assign node8376 = (inp[9]) ? node8382 : node8377;
													assign node8377 = (inp[10]) ? node8379 : 4'b0110;
														assign node8379 = (inp[12]) ? 4'b0011 : 4'b0110;
													assign node8382 = (inp[10]) ? node8384 : 4'b0010;
														assign node8384 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node8387 = (inp[9]) ? node8401 : node8388;
													assign node8388 = (inp[12]) ? node8394 : node8389;
														assign node8389 = (inp[8]) ? node8391 : 4'b0011;
															assign node8391 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node8394 = (inp[10]) ? node8396 : 4'b0010;
															assign node8396 = (inp[2]) ? node8398 : 4'b0110;
																assign node8398 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node8401 = (inp[10]) ? node8409 : node8402;
														assign node8402 = (inp[12]) ? 4'b0111 : node8403;
															assign node8403 = (inp[2]) ? 4'b0110 : node8404;
																assign node8404 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node8409 = (inp[12]) ? 4'b0010 : node8410;
															assign node8410 = (inp[8]) ? 4'b0110 : 4'b0111;
										assign node8414 = (inp[3]) ? node8466 : node8415;
											assign node8415 = (inp[9]) ? node8443 : node8416;
												assign node8416 = (inp[4]) ? node8428 : node8417;
													assign node8417 = (inp[8]) ? node8425 : node8418;
														assign node8418 = (inp[2]) ? node8420 : 4'b0110;
															assign node8420 = (inp[12]) ? node8422 : 4'b0111;
																assign node8422 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node8425 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node8428 = (inp[10]) ? node8436 : node8429;
														assign node8429 = (inp[8]) ? node8433 : node8430;
															assign node8430 = (inp[12]) ? 4'b0011 : 4'b0010;
															assign node8433 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node8436 = (inp[12]) ? node8440 : node8437;
															assign node8437 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node8440 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node8443 = (inp[4]) ? node8453 : node8444;
													assign node8444 = (inp[12]) ? node8448 : node8445;
														assign node8445 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node8448 = (inp[8]) ? node8450 : 4'b0101;
															assign node8450 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node8453 = (inp[10]) ? node8459 : node8454;
														assign node8454 = (inp[8]) ? node8456 : 4'b0100;
															assign node8456 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node8459 = (inp[12]) ? node8461 : 4'b0101;
															assign node8461 = (inp[2]) ? 4'b0001 : node8462;
																assign node8462 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node8466 = (inp[12]) ? node8500 : node8467;
												assign node8467 = (inp[8]) ? node8479 : node8468;
													assign node8468 = (inp[2]) ? node8476 : node8469;
														assign node8469 = (inp[4]) ? node8473 : node8470;
															assign node8470 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node8473 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node8476 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node8479 = (inp[2]) ? node8489 : node8480;
														assign node8480 = (inp[10]) ? node8482 : 4'b0001;
															assign node8482 = (inp[4]) ? node8486 : node8483;
																assign node8483 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node8486 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node8489 = (inp[10]) ? node8495 : node8490;
															assign node8490 = (inp[4]) ? 4'b0100 : node8491;
																assign node8491 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node8495 = (inp[4]) ? node8497 : 4'b0000;
																assign node8497 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node8500 = (inp[10]) ? node8520 : node8501;
													assign node8501 = (inp[2]) ? node8509 : node8502;
														assign node8502 = (inp[8]) ? 4'b0101 : node8503;
															assign node8503 = (inp[4]) ? node8505 : 4'b0100;
																assign node8505 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node8509 = (inp[8]) ? node8515 : node8510;
															assign node8510 = (inp[4]) ? 4'b0001 : node8511;
																assign node8511 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node8515 = (inp[9]) ? node8517 : 4'b0000;
																assign node8517 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node8520 = (inp[9]) ? node8526 : node8521;
														assign node8521 = (inp[2]) ? node8523 : 4'b0100;
															assign node8523 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node8526 = (inp[4]) ? 4'b0000 : 4'b0100;
							assign node8529 = (inp[7]) ? node8931 : node8530;
								assign node8530 = (inp[2]) ? node8748 : node8531;
									assign node8531 = (inp[8]) ? node8653 : node8532;
										assign node8532 = (inp[4]) ? node8598 : node8533;
											assign node8533 = (inp[9]) ? node8559 : node8534;
												assign node8534 = (inp[12]) ? node8546 : node8535;
													assign node8535 = (inp[0]) ? node8541 : node8536;
														assign node8536 = (inp[15]) ? node8538 : 4'b0111;
															assign node8538 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node8541 = (inp[3]) ? node8543 : 4'b0101;
															assign node8543 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node8546 = (inp[10]) ? node8554 : node8547;
														assign node8547 = (inp[0]) ? 4'b0111 : node8548;
															assign node8548 = (inp[3]) ? node8550 : 4'b0101;
																assign node8550 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node8554 = (inp[3]) ? node8556 : 4'b0011;
															assign node8556 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node8559 = (inp[12]) ? node8581 : node8560;
													assign node8560 = (inp[10]) ? node8568 : node8561;
														assign node8561 = (inp[3]) ? node8563 : 4'b0001;
															assign node8563 = (inp[0]) ? 4'b0001 : node8564;
																assign node8564 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node8568 = (inp[15]) ? node8574 : node8569;
															assign node8569 = (inp[3]) ? 4'b0011 : node8570;
																assign node8570 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node8574 = (inp[3]) ? node8578 : node8575;
																assign node8575 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node8578 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node8581 = (inp[10]) ? node8591 : node8582;
														assign node8582 = (inp[3]) ? 4'b0001 : node8583;
															assign node8583 = (inp[0]) ? node8587 : node8584;
																assign node8584 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node8587 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node8591 = (inp[0]) ? node8595 : node8592;
															assign node8592 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node8595 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node8598 = (inp[9]) ? node8636 : node8599;
												assign node8599 = (inp[12]) ? node8621 : node8600;
													assign node8600 = (inp[10]) ? node8608 : node8601;
														assign node8601 = (inp[0]) ? node8603 : 4'b0011;
															assign node8603 = (inp[3]) ? node8605 : 4'b0011;
																assign node8605 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node8608 = (inp[0]) ? node8616 : node8609;
															assign node8609 = (inp[15]) ? node8613 : node8610;
																assign node8610 = (inp[3]) ? 4'b0001 : 4'b0011;
																assign node8613 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node8616 = (inp[15]) ? 4'b0011 : node8617;
																assign node8617 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node8621 = (inp[10]) ? node8631 : node8622;
														assign node8622 = (inp[0]) ? node8624 : 4'b0001;
															assign node8624 = (inp[15]) ? node8628 : node8625;
																assign node8625 = (inp[3]) ? 4'b0011 : 4'b0001;
																assign node8628 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node8631 = (inp[3]) ? node8633 : 4'b0111;
															assign node8633 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node8636 = (inp[12]) ? node8644 : node8637;
													assign node8637 = (inp[0]) ? node8641 : node8638;
														assign node8638 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node8641 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node8644 = (inp[10]) ? node8646 : 4'b0101;
														assign node8646 = (inp[0]) ? node8650 : node8647;
															assign node8647 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node8650 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node8653 = (inp[15]) ? node8697 : node8654;
											assign node8654 = (inp[0]) ? node8672 : node8655;
												assign node8655 = (inp[3]) ? node8663 : node8656;
													assign node8656 = (inp[10]) ? node8658 : 4'b0010;
														assign node8658 = (inp[12]) ? 4'b0100 : node8659;
															assign node8659 = (inp[9]) ? 4'b0100 : 4'b0110;
													assign node8663 = (inp[4]) ? node8669 : node8664;
														assign node8664 = (inp[12]) ? 4'b0000 : node8665;
															assign node8665 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node8669 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node8672 = (inp[3]) ? node8684 : node8673;
													assign node8673 = (inp[4]) ? node8677 : node8674;
														assign node8674 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node8677 = (inp[10]) ? node8681 : node8678;
															assign node8678 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node8681 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node8684 = (inp[9]) ? node8692 : node8685;
														assign node8685 = (inp[4]) ? node8687 : 4'b0110;
															assign node8687 = (inp[10]) ? node8689 : 4'b0010;
																assign node8689 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node8692 = (inp[4]) ? 4'b0110 : node8693;
															assign node8693 = (inp[12]) ? 4'b0110 : 4'b0010;
											assign node8697 = (inp[0]) ? node8727 : node8698;
												assign node8698 = (inp[3]) ? node8712 : node8699;
													assign node8699 = (inp[9]) ? node8703 : node8700;
														assign node8700 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node8703 = (inp[12]) ? node8705 : 4'b0000;
															assign node8705 = (inp[10]) ? node8709 : node8706;
																assign node8706 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node8709 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node8712 = (inp[9]) ? node8718 : node8713;
														assign node8713 = (inp[4]) ? node8715 : 4'b0110;
															assign node8715 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node8718 = (inp[12]) ? node8720 : 4'b0010;
															assign node8720 = (inp[10]) ? node8724 : node8721;
																assign node8721 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node8724 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node8727 = (inp[3]) ? node8741 : node8728;
													assign node8728 = (inp[9]) ? node8738 : node8729;
														assign node8729 = (inp[4]) ? node8733 : node8730;
															assign node8730 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node8733 = (inp[12]) ? node8735 : 4'b0010;
																assign node8735 = (inp[10]) ? 4'b0100 : 4'b0010;
														assign node8738 = (inp[4]) ? 4'b0000 : 4'b0010;
													assign node8741 = (inp[4]) ? node8743 : 4'b0000;
														assign node8743 = (inp[12]) ? 4'b0100 : node8744;
															assign node8744 = (inp[9]) ? 4'b0100 : 4'b0000;
									assign node8748 = (inp[8]) ? node8848 : node8749;
										assign node8749 = (inp[12]) ? node8787 : node8750;
											assign node8750 = (inp[0]) ? node8768 : node8751;
												assign node8751 = (inp[4]) ? node8759 : node8752;
													assign node8752 = (inp[9]) ? node8754 : 4'b0100;
														assign node8754 = (inp[15]) ? 4'b0000 : node8755;
															assign node8755 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node8759 = (inp[9]) ? node8765 : node8760;
														assign node8760 = (inp[3]) ? 4'b0010 : node8761;
															assign node8761 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node8765 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node8768 = (inp[9]) ? node8780 : node8769;
													assign node8769 = (inp[4]) ? 4'b0010 : node8770;
														assign node8770 = (inp[10]) ? node8772 : 4'b0110;
															assign node8772 = (inp[3]) ? node8776 : node8773;
																assign node8773 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node8776 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node8780 = (inp[4]) ? node8784 : node8781;
														assign node8781 = (inp[10]) ? 4'b0000 : 4'b0010;
														assign node8784 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node8787 = (inp[0]) ? node8815 : node8788;
												assign node8788 = (inp[15]) ? node8798 : node8789;
													assign node8789 = (inp[3]) ? node8793 : node8790;
														assign node8790 = (inp[4]) ? 4'b0100 : 4'b0110;
														assign node8793 = (inp[10]) ? node8795 : 4'b0000;
															assign node8795 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node8798 = (inp[9]) ? node8808 : node8799;
														assign node8799 = (inp[3]) ? 4'b0110 : node8800;
															assign node8800 = (inp[10]) ? node8804 : node8801;
																assign node8801 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node8804 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node8808 = (inp[3]) ? 4'b0010 : node8809;
															assign node8809 = (inp[10]) ? node8811 : 4'b0110;
																assign node8811 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node8815 = (inp[15]) ? node8837 : node8816;
													assign node8816 = (inp[3]) ? node8830 : node8817;
														assign node8817 = (inp[4]) ? node8823 : node8818;
															assign node8818 = (inp[10]) ? node8820 : 4'b0000;
																assign node8820 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node8823 = (inp[10]) ? node8827 : node8824;
																assign node8824 = (inp[9]) ? 4'b0110 : 4'b0000;
																assign node8827 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node8830 = (inp[4]) ? node8834 : node8831;
															assign node8831 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node8834 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node8837 = (inp[3]) ? node8845 : node8838;
														assign node8838 = (inp[9]) ? node8840 : 4'b0010;
															assign node8840 = (inp[10]) ? node8842 : 4'b0010;
																assign node8842 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node8845 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node8848 = (inp[10]) ? node8894 : node8849;
											assign node8849 = (inp[15]) ? node8877 : node8850;
												assign node8850 = (inp[0]) ? node8862 : node8851;
													assign node8851 = (inp[4]) ? node8857 : node8852;
														assign node8852 = (inp[3]) ? node8854 : 4'b1011;
															assign node8854 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node8857 = (inp[12]) ? 4'b1101 : node8858;
															assign node8858 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node8862 = (inp[3]) ? node8868 : node8863;
														assign node8863 = (inp[9]) ? 4'b1111 : node8864;
															assign node8864 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node8868 = (inp[4]) ? node8870 : 4'b1011;
															assign node8870 = (inp[12]) ? node8874 : node8871;
																assign node8871 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node8874 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node8877 = (inp[0]) ? node8885 : node8878;
													assign node8878 = (inp[3]) ? node8882 : node8879;
														assign node8879 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node8882 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node8885 = (inp[12]) ? node8887 : 4'b1101;
														assign node8887 = (inp[9]) ? node8891 : node8888;
															assign node8888 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node8891 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node8894 = (inp[15]) ? node8912 : node8895;
												assign node8895 = (inp[0]) ? node8903 : node8896;
													assign node8896 = (inp[9]) ? node8900 : node8897;
														assign node8897 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node8900 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node8903 = (inp[3]) ? node8907 : node8904;
														assign node8904 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node8907 = (inp[9]) ? 4'b1111 : node8908;
															assign node8908 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node8912 = (inp[0]) ? node8922 : node8913;
													assign node8913 = (inp[3]) ? 4'b1011 : node8914;
														assign node8914 = (inp[4]) ? node8918 : node8915;
															assign node8915 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node8918 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node8922 = (inp[9]) ? node8928 : node8923;
														assign node8923 = (inp[4]) ? 4'b1101 : node8924;
															assign node8924 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node8928 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node8931 = (inp[8]) ? node9097 : node8932;
									assign node8932 = (inp[2]) ? node9018 : node8933;
										assign node8933 = (inp[4]) ? node8971 : node8934;
											assign node8934 = (inp[9]) ? node8952 : node8935;
												assign node8935 = (inp[12]) ? node8945 : node8936;
													assign node8936 = (inp[3]) ? node8940 : node8937;
														assign node8937 = (inp[10]) ? 4'b0100 : 4'b0110;
														assign node8940 = (inp[15]) ? 4'b0110 : node8941;
															assign node8941 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node8945 = (inp[10]) ? 4'b0000 : node8946;
														assign node8946 = (inp[15]) ? 4'b0100 : node8947;
															assign node8947 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node8952 = (inp[10]) ? node8964 : node8953;
													assign node8953 = (inp[15]) ? node8959 : node8954;
														assign node8954 = (inp[3]) ? 4'b0000 : node8955;
															assign node8955 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node8959 = (inp[12]) ? node8961 : 4'b0010;
															assign node8961 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node8964 = (inp[12]) ? node8966 : 4'b0000;
														assign node8966 = (inp[0]) ? node8968 : 4'b0110;
															assign node8968 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node8971 = (inp[9]) ? node8999 : node8972;
												assign node8972 = (inp[10]) ? node8984 : node8973;
													assign node8973 = (inp[0]) ? node8979 : node8974;
														assign node8974 = (inp[3]) ? 4'b0000 : node8975;
															assign node8975 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node8979 = (inp[3]) ? 4'b0010 : node8980;
															assign node8980 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node8984 = (inp[12]) ? node8990 : node8985;
														assign node8985 = (inp[0]) ? 4'b0010 : node8986;
															assign node8986 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node8990 = (inp[3]) ? 4'b0100 : node8991;
															assign node8991 = (inp[0]) ? node8995 : node8992;
																assign node8992 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node8995 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node8999 = (inp[12]) ? node9005 : node9000;
													assign node9000 = (inp[15]) ? node9002 : 4'b0110;
														assign node9002 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node9005 = (inp[10]) ? node9011 : node9006;
														assign node9006 = (inp[0]) ? 4'b0100 : node9007;
															assign node9007 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node9011 = (inp[3]) ? node9013 : 4'b0000;
															assign node9013 = (inp[15]) ? 4'b0010 : node9014;
																assign node9014 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node9018 = (inp[15]) ? node9060 : node9019;
											assign node9019 = (inp[0]) ? node9035 : node9020;
												assign node9020 = (inp[10]) ? 4'b1101 : node9021;
													assign node9021 = (inp[3]) ? 4'b1001 : node9022;
														assign node9022 = (inp[9]) ? node9028 : node9023;
															assign node9023 = (inp[4]) ? 4'b1011 : node9024;
																assign node9024 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node9028 = (inp[12]) ? 4'b1101 : node9029;
																assign node9029 = (inp[4]) ? 4'b1101 : 4'b1011;
												assign node9035 = (inp[3]) ? node9051 : node9036;
													assign node9036 = (inp[4]) ? node9044 : node9037;
														assign node9037 = (inp[12]) ? 4'b1001 : node9038;
															assign node9038 = (inp[10]) ? 4'b1111 : node9039;
																assign node9039 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node9044 = (inp[9]) ? node9048 : node9045;
															assign node9045 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node9048 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node9051 = (inp[4]) ? node9053 : 4'b1111;
														assign node9053 = (inp[9]) ? 4'b1011 : node9054;
															assign node9054 = (inp[12]) ? 4'b1111 : node9055;
																assign node9055 = (inp[10]) ? 4'b1111 : 4'b1011;
											assign node9060 = (inp[0]) ? node9072 : node9061;
												assign node9061 = (inp[4]) ? node9067 : node9062;
													assign node9062 = (inp[3]) ? node9064 : 4'b1001;
														assign node9064 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node9067 = (inp[9]) ? node9069 : 4'b1111;
														assign node9069 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node9072 = (inp[3]) ? node9082 : node9073;
													assign node9073 = (inp[4]) ? node9079 : node9074;
														assign node9074 = (inp[9]) ? node9076 : 4'b1011;
															assign node9076 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node9079 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node9082 = (inp[10]) ? node9092 : node9083;
														assign node9083 = (inp[9]) ? 4'b1001 : node9084;
															assign node9084 = (inp[12]) ? node9088 : node9085;
																assign node9085 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node9088 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node9092 = (inp[9]) ? node9094 : 4'b1001;
															assign node9094 = (inp[4]) ? 4'b1001 : 4'b1101;
									assign node9097 = (inp[2]) ? node9157 : node9098;
										assign node9098 = (inp[15]) ? node9134 : node9099;
											assign node9099 = (inp[0]) ? node9117 : node9100;
												assign node9100 = (inp[3]) ? node9112 : node9101;
													assign node9101 = (inp[10]) ? node9105 : node9102;
														assign node9102 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node9105 = (inp[12]) ? 4'b1101 : node9106;
															assign node9106 = (inp[4]) ? node9108 : 4'b1011;
																assign node9108 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node9112 = (inp[9]) ? node9114 : 4'b1001;
														assign node9114 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node9117 = (inp[12]) ? node9125 : node9118;
													assign node9118 = (inp[9]) ? 4'b1111 : node9119;
														assign node9119 = (inp[10]) ? 4'b1111 : node9120;
															assign node9120 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node9125 = (inp[4]) ? node9131 : node9126;
														assign node9126 = (inp[3]) ? node9128 : 4'b1001;
															assign node9128 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node9131 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node9134 = (inp[0]) ? node9148 : node9135;
												assign node9135 = (inp[3]) ? node9141 : node9136;
													assign node9136 = (inp[4]) ? 4'b1111 : node9137;
														assign node9137 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node9141 = (inp[4]) ? node9143 : 4'b1111;
														assign node9143 = (inp[9]) ? node9145 : 4'b1111;
															assign node9145 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node9148 = (inp[9]) ? node9152 : node9149;
													assign node9149 = (inp[4]) ? 4'b1101 : 4'b1011;
													assign node9152 = (inp[4]) ? node9154 : 4'b1101;
														assign node9154 = (inp[10]) ? 4'b1001 : 4'b1101;
										assign node9157 = (inp[4]) ? node9203 : node9158;
											assign node9158 = (inp[9]) ? node9178 : node9159;
												assign node9159 = (inp[10]) ? node9171 : node9160;
													assign node9160 = (inp[12]) ? node9168 : node9161;
														assign node9161 = (inp[3]) ? 4'b1100 : node9162;
															assign node9162 = (inp[0]) ? node9164 : 4'b1110;
																assign node9164 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node9168 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node9171 = (inp[3]) ? node9173 : 4'b1000;
														assign node9173 = (inp[12]) ? node9175 : 4'b1010;
															assign node9175 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node9178 = (inp[10]) ? node9194 : node9179;
													assign node9179 = (inp[12]) ? node9181 : 4'b1010;
														assign node9181 = (inp[3]) ? node9189 : node9182;
															assign node9182 = (inp[15]) ? node9186 : node9183;
																assign node9183 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node9186 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node9189 = (inp[15]) ? node9191 : 4'b1110;
																assign node9191 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node9194 = (inp[12]) ? 4'b1100 : node9195;
														assign node9195 = (inp[15]) ? node9199 : node9196;
															assign node9196 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node9199 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node9203 = (inp[0]) ? node9219 : node9204;
												assign node9204 = (inp[15]) ? 4'b1010 : node9205;
													assign node9205 = (inp[9]) ? node9213 : node9206;
														assign node9206 = (inp[10]) ? 4'b1100 : node9207;
															assign node9207 = (inp[12]) ? 4'b1100 : node9208;
																assign node9208 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node9213 = (inp[10]) ? 4'b1000 : node9214;
															assign node9214 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node9219 = (inp[15]) ? node9223 : node9220;
													assign node9220 = (inp[12]) ? 4'b1010 : 4'b1110;
													assign node9223 = (inp[10]) ? 4'b1100 : node9224;
														assign node9224 = (inp[12]) ? 4'b1100 : node9225;
															assign node9225 = (inp[9]) ? 4'b1100 : node9226;
																assign node9226 = (inp[3]) ? 4'b1000 : 4'b1010;
					assign node9232 = (inp[6]) ? node10858 : node9233;
						assign node9233 = (inp[1]) ? node10059 : node9234;
							assign node9234 = (inp[7]) ? node9654 : node9235;
								assign node9235 = (inp[2]) ? node9447 : node9236;
									assign node9236 = (inp[8]) ? node9336 : node9237;
										assign node9237 = (inp[15]) ? node9283 : node9238;
											assign node9238 = (inp[0]) ? node9256 : node9239;
												assign node9239 = (inp[3]) ? node9249 : node9240;
													assign node9240 = (inp[9]) ? node9244 : node9241;
														assign node9241 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node9244 = (inp[4]) ? node9246 : 4'b1011;
															assign node9246 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node9249 = (inp[4]) ? node9251 : 4'b1001;
														assign node9251 = (inp[12]) ? node9253 : 4'b1001;
															assign node9253 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node9256 = (inp[3]) ? node9268 : node9257;
													assign node9257 = (inp[9]) ? node9265 : node9258;
														assign node9258 = (inp[4]) ? 4'b1001 : node9259;
															assign node9259 = (inp[12]) ? node9261 : 4'b1101;
																assign node9261 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node9265 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node9268 = (inp[12]) ? node9276 : node9269;
														assign node9269 = (inp[4]) ? node9273 : node9270;
															assign node9270 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node9273 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node9276 = (inp[10]) ? 4'b1111 : node9277;
															assign node9277 = (inp[4]) ? node9279 : 4'b1111;
																assign node9279 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node9283 = (inp[0]) ? node9303 : node9284;
												assign node9284 = (inp[3]) ? node9292 : node9285;
													assign node9285 = (inp[9]) ? node9289 : node9286;
														assign node9286 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node9289 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node9292 = (inp[12]) ? node9294 : 4'b1111;
														assign node9294 = (inp[10]) ? 4'b1011 : node9295;
															assign node9295 = (inp[4]) ? node9299 : node9296;
																assign node9296 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node9299 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node9303 = (inp[3]) ? node9319 : node9304;
													assign node9304 = (inp[9]) ? node9312 : node9305;
														assign node9305 = (inp[4]) ? node9307 : 4'b1111;
															assign node9307 = (inp[12]) ? node9309 : 4'b1011;
																assign node9309 = (inp[10]) ? 4'b1101 : 4'b1011;
														assign node9312 = (inp[4]) ? 4'b1101 : node9313;
															assign node9313 = (inp[10]) ? node9315 : 4'b1011;
																assign node9315 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node9319 = (inp[12]) ? node9327 : node9320;
														assign node9320 = (inp[9]) ? node9324 : node9321;
															assign node9321 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node9324 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node9327 = (inp[9]) ? node9329 : 4'b1001;
															assign node9329 = (inp[4]) ? node9333 : node9330;
																assign node9330 = (inp[10]) ? 4'b1101 : 4'b1001;
																assign node9333 = (inp[10]) ? 4'b1001 : 4'b1101;
										assign node9336 = (inp[0]) ? node9392 : node9337;
											assign node9337 = (inp[15]) ? node9365 : node9338;
												assign node9338 = (inp[3]) ? node9350 : node9339;
													assign node9339 = (inp[9]) ? node9345 : node9340;
														assign node9340 = (inp[4]) ? 4'b1010 : node9341;
															assign node9341 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node9345 = (inp[4]) ? node9347 : 4'b1010;
															assign node9347 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node9350 = (inp[4]) ? node9358 : node9351;
														assign node9351 = (inp[9]) ? node9353 : 4'b1100;
															assign node9353 = (inp[10]) ? node9355 : 4'b1000;
																assign node9355 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node9358 = (inp[9]) ? node9360 : 4'b1000;
															assign node9360 = (inp[12]) ? node9362 : 4'b1100;
																assign node9362 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node9365 = (inp[3]) ? node9377 : node9366;
													assign node9366 = (inp[9]) ? node9374 : node9367;
														assign node9367 = (inp[4]) ? 4'b1000 : node9368;
															assign node9368 = (inp[10]) ? node9370 : 4'b1100;
																assign node9370 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node9374 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node9377 = (inp[12]) ? node9383 : node9378;
														assign node9378 = (inp[4]) ? node9380 : 4'b1110;
															assign node9380 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node9383 = (inp[9]) ? 4'b1010 : node9384;
															assign node9384 = (inp[10]) ? node9388 : node9385;
																assign node9385 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node9388 = (inp[4]) ? 4'b1110 : 4'b1010;
											assign node9392 = (inp[12]) ? node9420 : node9393;
												assign node9393 = (inp[3]) ? node9407 : node9394;
													assign node9394 = (inp[15]) ? node9400 : node9395;
														assign node9395 = (inp[9]) ? node9397 : 4'b1000;
															assign node9397 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node9400 = (inp[9]) ? node9404 : node9401;
															assign node9401 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node9404 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node9407 = (inp[15]) ? node9417 : node9408;
														assign node9408 = (inp[10]) ? node9414 : node9409;
															assign node9409 = (inp[9]) ? node9411 : 4'b1010;
																assign node9411 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node9414 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node9417 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node9420 = (inp[15]) ? node9436 : node9421;
													assign node9421 = (inp[3]) ? node9425 : node9422;
														assign node9422 = (inp[9]) ? 4'b1110 : 4'b1100;
														assign node9425 = (inp[9]) ? node9431 : node9426;
															assign node9426 = (inp[4]) ? node9428 : 4'b1110;
																assign node9428 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node9431 = (inp[10]) ? node9433 : 4'b1010;
																assign node9433 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node9436 = (inp[10]) ? node9440 : node9437;
														assign node9437 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node9440 = (inp[3]) ? 4'b1100 : node9441;
															assign node9441 = (inp[4]) ? node9443 : 4'b1010;
																assign node9443 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node9447 = (inp[8]) ? node9545 : node9448;
										assign node9448 = (inp[10]) ? node9488 : node9449;
											assign node9449 = (inp[9]) ? node9471 : node9450;
												assign node9450 = (inp[4]) ? node9466 : node9451;
													assign node9451 = (inp[0]) ? node9459 : node9452;
														assign node9452 = (inp[3]) ? node9456 : node9453;
															assign node9453 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node9456 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node9459 = (inp[15]) ? node9463 : node9460;
															assign node9460 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node9463 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node9466 = (inp[12]) ? 4'b1010 : node9467;
														assign node9467 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node9471 = (inp[4]) ? node9481 : node9472;
													assign node9472 = (inp[12]) ? node9474 : 4'b1010;
														assign node9474 = (inp[15]) ? node9476 : 4'b1000;
															assign node9476 = (inp[3]) ? 4'b1010 : node9477;
																assign node9477 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node9481 = (inp[12]) ? node9483 : 4'b1110;
														assign node9483 = (inp[0]) ? node9485 : 4'b1100;
															assign node9485 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node9488 = (inp[15]) ? node9520 : node9489;
												assign node9489 = (inp[0]) ? node9505 : node9490;
													assign node9490 = (inp[3]) ? node9496 : node9491;
														assign node9491 = (inp[9]) ? node9493 : 4'b1010;
															assign node9493 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node9496 = (inp[9]) ? 4'b1000 : node9497;
															assign node9497 = (inp[4]) ? node9501 : node9498;
																assign node9498 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node9501 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node9505 = (inp[3]) ? node9513 : node9506;
														assign node9506 = (inp[4]) ? node9508 : 4'b1000;
															assign node9508 = (inp[12]) ? node9510 : 4'b1000;
																assign node9510 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node9513 = (inp[9]) ? node9517 : node9514;
															assign node9514 = (inp[12]) ? 4'b1010 : 4'b1110;
															assign node9517 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node9520 = (inp[3]) ? node9542 : node9521;
													assign node9521 = (inp[12]) ? node9531 : node9522;
														assign node9522 = (inp[0]) ? node9526 : node9523;
															assign node9523 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node9526 = (inp[4]) ? 4'b1010 : node9527;
																assign node9527 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node9531 = (inp[0]) ? node9537 : node9532;
															assign node9532 = (inp[4]) ? 4'b1110 : node9533;
																assign node9533 = (inp[9]) ? 4'b1110 : 4'b1000;
															assign node9537 = (inp[9]) ? node9539 : 4'b1100;
																assign node9539 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node9542 = (inp[4]) ? 4'b1100 : 4'b1000;
										assign node9545 = (inp[12]) ? node9597 : node9546;
											assign node9546 = (inp[4]) ? node9578 : node9547;
												assign node9547 = (inp[9]) ? node9561 : node9548;
													assign node9548 = (inp[3]) ? node9554 : node9549;
														assign node9549 = (inp[10]) ? 4'b0111 : node9550;
															assign node9550 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node9554 = (inp[10]) ? node9558 : node9555;
															assign node9555 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node9558 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node9561 = (inp[10]) ? node9567 : node9562;
														assign node9562 = (inp[3]) ? 4'b0011 : node9563;
															assign node9563 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node9567 = (inp[0]) ? node9573 : node9568;
															assign node9568 = (inp[15]) ? node9570 : 4'b0001;
																assign node9570 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node9573 = (inp[15]) ? node9575 : 4'b0011;
																assign node9575 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node9578 = (inp[9]) ? 4'b0111 : node9579;
													assign node9579 = (inp[10]) ? node9587 : node9580;
														assign node9580 = (inp[15]) ? node9582 : 4'b0001;
															assign node9582 = (inp[0]) ? 4'b0001 : node9583;
																assign node9583 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node9587 = (inp[15]) ? node9589 : 4'b0011;
															assign node9589 = (inp[3]) ? node9593 : node9590;
																assign node9590 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node9593 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node9597 = (inp[0]) ? node9631 : node9598;
												assign node9598 = (inp[15]) ? node9618 : node9599;
													assign node9599 = (inp[3]) ? node9611 : node9600;
														assign node9600 = (inp[4]) ? node9608 : node9601;
															assign node9601 = (inp[9]) ? node9605 : node9602;
																assign node9602 = (inp[10]) ? 4'b0011 : 4'b0111;
																assign node9605 = (inp[10]) ? 4'b0101 : 4'b0011;
															assign node9608 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node9611 = (inp[10]) ? 4'b0001 : node9612;
															assign node9612 = (inp[4]) ? node9614 : 4'b0101;
																assign node9614 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node9618 = (inp[10]) ? node9626 : node9619;
														assign node9619 = (inp[3]) ? 4'b0011 : node9620;
															assign node9620 = (inp[4]) ? 4'b0001 : node9621;
																assign node9621 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node9626 = (inp[9]) ? 4'b0111 : node9627;
															assign node9627 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node9631 = (inp[15]) ? node9639 : node9632;
													assign node9632 = (inp[10]) ? node9634 : 4'b0111;
														assign node9634 = (inp[9]) ? node9636 : 4'b0111;
															assign node9636 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node9639 = (inp[3]) ? node9647 : node9640;
														assign node9640 = (inp[9]) ? 4'b0101 : node9641;
															assign node9641 = (inp[10]) ? 4'b0011 : node9642;
																assign node9642 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node9647 = (inp[4]) ? 4'b0101 : node9648;
															assign node9648 = (inp[9]) ? node9650 : 4'b0101;
																assign node9650 = (inp[10]) ? 4'b0101 : 4'b0001;
								assign node9654 = (inp[8]) ? node9860 : node9655;
									assign node9655 = (inp[2]) ? node9755 : node9656;
										assign node9656 = (inp[4]) ? node9712 : node9657;
											assign node9657 = (inp[9]) ? node9683 : node9658;
												assign node9658 = (inp[10]) ? node9668 : node9659;
													assign node9659 = (inp[3]) ? node9661 : 4'b1100;
														assign node9661 = (inp[12]) ? node9663 : 4'b1110;
															assign node9663 = (inp[0]) ? node9665 : 4'b1100;
																assign node9665 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node9668 = (inp[12]) ? node9672 : node9669;
														assign node9669 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node9672 = (inp[3]) ? node9678 : node9673;
															assign node9673 = (inp[15]) ? node9675 : 4'b1000;
																assign node9675 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node9678 = (inp[15]) ? node9680 : 4'b1010;
																assign node9680 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node9683 = (inp[12]) ? node9701 : node9684;
													assign node9684 = (inp[0]) ? node9692 : node9685;
														assign node9685 = (inp[15]) ? node9689 : node9686;
															assign node9686 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node9689 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node9692 = (inp[10]) ? 4'b1010 : node9693;
															assign node9693 = (inp[3]) ? node9697 : node9694;
																assign node9694 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node9697 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node9701 = (inp[10]) ? node9709 : node9702;
														assign node9702 = (inp[0]) ? node9704 : 4'b1000;
															assign node9704 = (inp[3]) ? 4'b1000 : node9705;
																assign node9705 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node9709 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node9712 = (inp[9]) ? node9732 : node9713;
												assign node9713 = (inp[12]) ? node9721 : node9714;
													assign node9714 = (inp[0]) ? 4'b1010 : node9715;
														assign node9715 = (inp[15]) ? node9717 : 4'b1000;
															assign node9717 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node9721 = (inp[10]) ? node9725 : node9722;
														assign node9722 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node9725 = (inp[3]) ? 4'b1100 : node9726;
															assign node9726 = (inp[15]) ? 4'b1110 : node9727;
																assign node9727 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node9732 = (inp[12]) ? node9740 : node9733;
													assign node9733 = (inp[3]) ? node9735 : 4'b1100;
														assign node9735 = (inp[15]) ? node9737 : 4'b1100;
															assign node9737 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node9740 = (inp[10]) ? node9746 : node9741;
														assign node9741 = (inp[15]) ? node9743 : 4'b1110;
															assign node9743 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node9746 = (inp[3]) ? 4'b1000 : node9747;
															assign node9747 = (inp[0]) ? node9751 : node9748;
																assign node9748 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node9751 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node9755 = (inp[10]) ? node9803 : node9756;
											assign node9756 = (inp[9]) ? node9780 : node9757;
												assign node9757 = (inp[4]) ? node9773 : node9758;
													assign node9758 = (inp[3]) ? node9766 : node9759;
														assign node9759 = (inp[15]) ? node9763 : node9760;
															assign node9760 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node9763 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node9766 = (inp[15]) ? node9770 : node9767;
															assign node9767 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node9770 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node9773 = (inp[15]) ? node9775 : 4'b0011;
														assign node9775 = (inp[0]) ? 4'b0001 : node9776;
															assign node9776 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node9780 = (inp[4]) ? node9796 : node9781;
													assign node9781 = (inp[12]) ? node9789 : node9782;
														assign node9782 = (inp[15]) ? 4'b0011 : node9783;
															assign node9783 = (inp[0]) ? node9785 : 4'b0011;
																assign node9785 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node9789 = (inp[0]) ? 4'b0001 : node9790;
															assign node9790 = (inp[15]) ? 4'b0011 : node9791;
																assign node9791 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node9796 = (inp[15]) ? node9800 : node9797;
														assign node9797 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node9800 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node9803 = (inp[4]) ? node9839 : node9804;
												assign node9804 = (inp[9]) ? node9820 : node9805;
													assign node9805 = (inp[12]) ? node9807 : 4'b0111;
														assign node9807 = (inp[15]) ? node9813 : node9808;
															assign node9808 = (inp[3]) ? node9810 : 4'b0011;
																assign node9810 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node9813 = (inp[3]) ? node9817 : node9814;
																assign node9814 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node9817 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node9820 = (inp[12]) ? node9832 : node9821;
														assign node9821 = (inp[0]) ? node9827 : node9822;
															assign node9822 = (inp[15]) ? node9824 : 4'b0011;
																assign node9824 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node9827 = (inp[3]) ? 4'b0001 : node9828;
																assign node9828 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node9832 = (inp[3]) ? 4'b0101 : node9833;
															assign node9833 = (inp[0]) ? 4'b0111 : node9834;
																assign node9834 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node9839 = (inp[12]) ? node9853 : node9840;
													assign node9840 = (inp[9]) ? node9850 : node9841;
														assign node9841 = (inp[3]) ? node9843 : 4'b0001;
															assign node9843 = (inp[0]) ? node9847 : node9844;
																assign node9844 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node9847 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node9850 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node9853 = (inp[9]) ? 4'b0011 : node9854;
														assign node9854 = (inp[0]) ? node9856 : 4'b0111;
															assign node9856 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node9860 = (inp[2]) ? node9960 : node9861;
										assign node9861 = (inp[0]) ? node9903 : node9862;
											assign node9862 = (inp[15]) ? node9884 : node9863;
												assign node9863 = (inp[3]) ? node9877 : node9864;
													assign node9864 = (inp[10]) ? node9870 : node9865;
														assign node9865 = (inp[9]) ? 4'b0011 : node9866;
															assign node9866 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node9870 = (inp[9]) ? node9872 : 4'b0011;
															assign node9872 = (inp[4]) ? 4'b0101 : node9873;
																assign node9873 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node9877 = (inp[12]) ? 4'b0001 : node9878;
														assign node9878 = (inp[10]) ? 4'b0101 : node9879;
															assign node9879 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node9884 = (inp[3]) ? node9890 : node9885;
													assign node9885 = (inp[4]) ? 4'b0111 : node9886;
														assign node9886 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node9890 = (inp[4]) ? node9894 : node9891;
														assign node9891 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node9894 = (inp[9]) ? node9898 : node9895;
															assign node9895 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node9898 = (inp[12]) ? node9900 : 4'b0111;
																assign node9900 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node9903 = (inp[15]) ? node9935 : node9904;
												assign node9904 = (inp[3]) ? node9920 : node9905;
													assign node9905 = (inp[12]) ? node9911 : node9906;
														assign node9906 = (inp[4]) ? 4'b0001 : node9907;
															assign node9907 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node9911 = (inp[4]) ? node9913 : 4'b0001;
															assign node9913 = (inp[10]) ? node9917 : node9914;
																assign node9914 = (inp[9]) ? 4'b0111 : 4'b0001;
																assign node9917 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node9920 = (inp[10]) ? node9928 : node9921;
														assign node9921 = (inp[4]) ? node9925 : node9922;
															assign node9922 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node9925 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node9928 = (inp[12]) ? 4'b0111 : node9929;
															assign node9929 = (inp[4]) ? node9931 : 4'b0111;
																assign node9931 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node9935 = (inp[3]) ? node9945 : node9936;
													assign node9936 = (inp[4]) ? node9940 : node9937;
														assign node9937 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node9940 = (inp[9]) ? 4'b0101 : node9941;
															assign node9941 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node9945 = (inp[9]) ? node9955 : node9946;
														assign node9946 = (inp[4]) ? node9950 : node9947;
															assign node9947 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node9950 = (inp[12]) ? node9952 : 4'b0001;
																assign node9952 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node9955 = (inp[10]) ? node9957 : 4'b0001;
															assign node9957 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node9960 = (inp[4]) ? node10006 : node9961;
											assign node9961 = (inp[9]) ? node9987 : node9962;
												assign node9962 = (inp[12]) ? node9976 : node9963;
													assign node9963 = (inp[0]) ? node9971 : node9964;
														assign node9964 = (inp[15]) ? node9968 : node9965;
															assign node9965 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node9968 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node9971 = (inp[3]) ? 4'b0100 : node9972;
															assign node9972 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node9976 = (inp[10]) ? node9978 : 4'b0100;
														assign node9978 = (inp[3]) ? node9980 : 4'b0010;
															assign node9980 = (inp[0]) ? node9984 : node9981;
																assign node9981 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node9984 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node9987 = (inp[10]) ? node9995 : node9988;
													assign node9988 = (inp[3]) ? node9990 : 4'b0000;
														assign node9990 = (inp[15]) ? node9992 : 4'b0010;
															assign node9992 = (inp[12]) ? 4'b0000 : 4'b0010;
													assign node9995 = (inp[12]) ? node10001 : node9996;
														assign node9996 = (inp[0]) ? 4'b0000 : node9997;
															assign node9997 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node10001 = (inp[15]) ? node10003 : 4'b0110;
															assign node10003 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node10006 = (inp[9]) ? node10038 : node10007;
												assign node10007 = (inp[12]) ? node10027 : node10008;
													assign node10008 = (inp[0]) ? node10014 : node10009;
														assign node10009 = (inp[15]) ? node10011 : 4'b0010;
															assign node10011 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node10014 = (inp[10]) ? node10020 : node10015;
															assign node10015 = (inp[15]) ? node10017 : 4'b0000;
																assign node10017 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node10020 = (inp[3]) ? node10024 : node10021;
																assign node10021 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node10024 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node10027 = (inp[10]) ? node10033 : node10028;
														assign node10028 = (inp[0]) ? node10030 : 4'b0010;
															assign node10030 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node10033 = (inp[15]) ? 4'b0110 : node10034;
															assign node10034 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node10038 = (inp[10]) ? node10048 : node10039;
													assign node10039 = (inp[12]) ? node10043 : node10040;
														assign node10040 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node10043 = (inp[15]) ? node10045 : 4'b0110;
															assign node10045 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node10048 = (inp[12]) ? node10054 : node10049;
														assign node10049 = (inp[15]) ? 4'b0110 : node10050;
															assign node10050 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node10054 = (inp[15]) ? 4'b0000 : node10055;
															assign node10055 = (inp[0]) ? 4'b0010 : 4'b0000;
							assign node10059 = (inp[2]) ? node10449 : node10060;
								assign node10060 = (inp[9]) ? node10246 : node10061;
									assign node10061 = (inp[4]) ? node10167 : node10062;
										assign node10062 = (inp[12]) ? node10112 : node10063;
											assign node10063 = (inp[15]) ? node10091 : node10064;
												assign node10064 = (inp[10]) ? node10078 : node10065;
													assign node10065 = (inp[3]) ? node10075 : node10066;
														assign node10066 = (inp[0]) ? 4'b0101 : node10067;
															assign node10067 = (inp[8]) ? node10071 : node10068;
																assign node10068 = (inp[7]) ? 4'b0110 : 4'b0111;
																assign node10071 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node10075 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node10078 = (inp[7]) ? node10086 : node10079;
														assign node10079 = (inp[3]) ? node10083 : node10080;
															assign node10080 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node10083 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node10086 = (inp[8]) ? 4'b0101 : node10087;
															assign node10087 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node10091 = (inp[0]) ? node10103 : node10092;
													assign node10092 = (inp[3]) ? node10094 : 4'b0101;
														assign node10094 = (inp[10]) ? node10098 : node10095;
															assign node10095 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node10098 = (inp[8]) ? 4'b0111 : node10099;
																assign node10099 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node10103 = (inp[3]) ? 4'b0101 : node10104;
														assign node10104 = (inp[8]) ? node10108 : node10105;
															assign node10105 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node10108 = (inp[7]) ? 4'b0111 : 4'b0110;
											assign node10112 = (inp[10]) ? node10138 : node10113;
												assign node10113 = (inp[0]) ? node10121 : node10114;
													assign node10114 = (inp[8]) ? node10118 : node10115;
														assign node10115 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node10118 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node10121 = (inp[7]) ? node10131 : node10122;
														assign node10122 = (inp[8]) ? node10128 : node10123;
															assign node10123 = (inp[15]) ? 4'b0111 : node10124;
																assign node10124 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node10128 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node10131 = (inp[8]) ? 4'b0111 : node10132;
															assign node10132 = (inp[15]) ? 4'b0110 : node10133;
																assign node10133 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node10138 = (inp[15]) ? node10152 : node10139;
													assign node10139 = (inp[0]) ? node10145 : node10140;
														assign node10140 = (inp[8]) ? node10142 : 4'b0001;
															assign node10142 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node10145 = (inp[3]) ? node10147 : 4'b0000;
															assign node10147 = (inp[7]) ? node10149 : 4'b0010;
																assign node10149 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node10152 = (inp[8]) ? node10156 : node10153;
														assign node10153 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node10156 = (inp[7]) ? node10162 : node10157;
															assign node10157 = (inp[3]) ? 4'b0010 : node10158;
																assign node10158 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node10162 = (inp[3]) ? node10164 : 4'b0011;
																assign node10164 = (inp[0]) ? 4'b0001 : 4'b0011;
										assign node10167 = (inp[10]) ? node10203 : node10168;
											assign node10168 = (inp[8]) ? node10186 : node10169;
												assign node10169 = (inp[7]) ? node10177 : node10170;
													assign node10170 = (inp[12]) ? 4'b0001 : node10171;
														assign node10171 = (inp[15]) ? 4'b0011 : node10172;
															assign node10172 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node10177 = (inp[0]) ? 4'b0000 : node10178;
														assign node10178 = (inp[15]) ? node10182 : node10179;
															assign node10179 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node10182 = (inp[12]) ? 4'b0010 : 4'b0000;
												assign node10186 = (inp[7]) ? node10198 : node10187;
													assign node10187 = (inp[0]) ? node10193 : node10188;
														assign node10188 = (inp[3]) ? 4'b0010 : node10189;
															assign node10189 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node10193 = (inp[3]) ? node10195 : 4'b0000;
															assign node10195 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node10198 = (inp[3]) ? 4'b0011 : node10199;
														assign node10199 = (inp[0]) ? 4'b0011 : 4'b0001;
											assign node10203 = (inp[12]) ? node10227 : node10204;
												assign node10204 = (inp[8]) ? node10216 : node10205;
													assign node10205 = (inp[7]) ? node10209 : node10206;
														assign node10206 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node10209 = (inp[15]) ? node10211 : 4'b0010;
															assign node10211 = (inp[0]) ? 4'b0000 : node10212;
																assign node10212 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node10216 = (inp[7]) ? node10218 : 4'b0010;
														assign node10218 = (inp[0]) ? node10220 : 4'b0011;
															assign node10220 = (inp[3]) ? node10224 : node10221;
																assign node10221 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node10224 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node10227 = (inp[8]) ? node10237 : node10228;
													assign node10228 = (inp[7]) ? 4'b0110 : node10229;
														assign node10229 = (inp[0]) ? node10233 : node10230;
															assign node10230 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node10233 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node10237 = (inp[7]) ? node10243 : node10238;
														assign node10238 = (inp[15]) ? node10240 : 4'b0110;
															assign node10240 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node10243 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node10246 = (inp[4]) ? node10354 : node10247;
										assign node10247 = (inp[12]) ? node10301 : node10248;
											assign node10248 = (inp[7]) ? node10268 : node10249;
												assign node10249 = (inp[8]) ? node10259 : node10250;
													assign node10250 = (inp[3]) ? node10252 : 4'b0011;
														assign node10252 = (inp[10]) ? node10254 : 4'b0001;
															assign node10254 = (inp[15]) ? node10256 : 4'b0011;
																assign node10256 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node10259 = (inp[3]) ? 4'b0010 : node10260;
														assign node10260 = (inp[0]) ? node10264 : node10261;
															assign node10261 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node10264 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node10268 = (inp[8]) ? node10280 : node10269;
													assign node10269 = (inp[0]) ? node10275 : node10270;
														assign node10270 = (inp[15]) ? 4'b0000 : node10271;
															assign node10271 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node10275 = (inp[3]) ? node10277 : 4'b0010;
															assign node10277 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node10280 = (inp[10]) ? node10288 : node10281;
														assign node10281 = (inp[3]) ? node10283 : 4'b0001;
															assign node10283 = (inp[15]) ? 4'b0001 : node10284;
																assign node10284 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node10288 = (inp[3]) ? node10296 : node10289;
															assign node10289 = (inp[0]) ? node10293 : node10290;
																assign node10290 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node10293 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node10296 = (inp[15]) ? node10298 : 4'b0011;
																assign node10298 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node10301 = (inp[10]) ? node10331 : node10302;
												assign node10302 = (inp[0]) ? node10316 : node10303;
													assign node10303 = (inp[8]) ? node10313 : node10304;
														assign node10304 = (inp[7]) ? node10306 : 4'b0011;
															assign node10306 = (inp[15]) ? node10310 : node10307;
																assign node10307 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node10310 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node10313 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node10316 = (inp[15]) ? node10320 : node10317;
														assign node10317 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node10320 = (inp[3]) ? node10326 : node10321;
															assign node10321 = (inp[7]) ? 4'b0010 : node10322;
																assign node10322 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node10326 = (inp[7]) ? 4'b0000 : node10327;
																assign node10327 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node10331 = (inp[0]) ? node10343 : node10332;
													assign node10332 = (inp[15]) ? node10340 : node10333;
														assign node10333 = (inp[3]) ? node10335 : 4'b0101;
															assign node10335 = (inp[8]) ? 4'b0100 : node10336;
																assign node10336 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node10340 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node10343 = (inp[15]) ? node10351 : node10344;
														assign node10344 = (inp[8]) ? node10348 : node10345;
															assign node10345 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node10348 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node10351 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node10354 = (inp[10]) ? node10400 : node10355;
											assign node10355 = (inp[7]) ? node10375 : node10356;
												assign node10356 = (inp[8]) ? node10362 : node10357;
													assign node10357 = (inp[3]) ? node10359 : 4'b0111;
														assign node10359 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node10362 = (inp[12]) ? node10370 : node10363;
														assign node10363 = (inp[15]) ? node10367 : node10364;
															assign node10364 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node10367 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node10370 = (inp[0]) ? 4'b0110 : node10371;
															assign node10371 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node10375 = (inp[8]) ? node10387 : node10376;
													assign node10376 = (inp[3]) ? node10382 : node10377;
														assign node10377 = (inp[15]) ? node10379 : 4'b0100;
															assign node10379 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node10382 = (inp[0]) ? 4'b0110 : node10383;
															assign node10383 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node10387 = (inp[3]) ? node10395 : node10388;
														assign node10388 = (inp[15]) ? node10392 : node10389;
															assign node10389 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node10392 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node10395 = (inp[0]) ? node10397 : 4'b0101;
															assign node10397 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node10400 = (inp[12]) ? node10418 : node10401;
												assign node10401 = (inp[15]) ? node10409 : node10402;
													assign node10402 = (inp[0]) ? node10404 : 4'b0100;
														assign node10404 = (inp[7]) ? node10406 : 4'b0111;
															assign node10406 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node10409 = (inp[0]) ? node10413 : node10410;
														assign node10410 = (inp[3]) ? 4'b0111 : 4'b0110;
														assign node10413 = (inp[8]) ? 4'b0100 : node10414;
															assign node10414 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node10418 = (inp[8]) ? node10434 : node10419;
													assign node10419 = (inp[7]) ? node10429 : node10420;
														assign node10420 = (inp[3]) ? node10422 : 4'b0001;
															assign node10422 = (inp[15]) ? node10426 : node10423;
																assign node10423 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node10426 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node10429 = (inp[0]) ? 4'b0000 : node10430;
															assign node10430 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node10434 = (inp[7]) ? node10442 : node10435;
														assign node10435 = (inp[15]) ? node10439 : node10436;
															assign node10436 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node10439 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node10442 = (inp[3]) ? 4'b0011 : node10443;
															assign node10443 = (inp[0]) ? 4'b0001 : node10444;
																assign node10444 = (inp[15]) ? 4'b0011 : 4'b0001;
								assign node10449 = (inp[10]) ? node10653 : node10450;
									assign node10450 = (inp[15]) ? node10552 : node10451;
										assign node10451 = (inp[7]) ? node10493 : node10452;
											assign node10452 = (inp[8]) ? node10482 : node10453;
												assign node10453 = (inp[12]) ? node10469 : node10454;
													assign node10454 = (inp[9]) ? node10464 : node10455;
														assign node10455 = (inp[4]) ? 4'b0000 : node10456;
															assign node10456 = (inp[0]) ? node10460 : node10457;
																assign node10457 = (inp[3]) ? 4'b0100 : 4'b0110;
																assign node10460 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node10464 = (inp[3]) ? node10466 : 4'b0110;
															assign node10466 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node10469 = (inp[9]) ? node10477 : node10470;
														assign node10470 = (inp[3]) ? node10474 : node10471;
															assign node10471 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node10474 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node10477 = (inp[4]) ? node10479 : 4'b0000;
															assign node10479 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node10482 = (inp[4]) ? 4'b0101 : node10483;
													assign node10483 = (inp[9]) ? node10485 : 4'b0111;
														assign node10485 = (inp[12]) ? 4'b0001 : node10486;
															assign node10486 = (inp[3]) ? 4'b0011 : node10487;
																assign node10487 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node10493 = (inp[8]) ? node10525 : node10494;
												assign node10494 = (inp[12]) ? node10510 : node10495;
													assign node10495 = (inp[9]) ? node10503 : node10496;
														assign node10496 = (inp[4]) ? node10498 : 4'b0101;
															assign node10498 = (inp[3]) ? node10500 : 4'b0001;
																assign node10500 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node10503 = (inp[4]) ? node10507 : node10504;
															assign node10504 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node10507 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node10510 = (inp[4]) ? node10518 : node10511;
														assign node10511 = (inp[9]) ? node10513 : 4'b0111;
															assign node10513 = (inp[0]) ? 4'b0011 : node10514;
																assign node10514 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node10518 = (inp[9]) ? node10522 : node10519;
															assign node10519 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node10522 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node10525 = (inp[12]) ? node10541 : node10526;
													assign node10526 = (inp[9]) ? node10530 : node10527;
														assign node10527 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node10530 = (inp[4]) ? node10538 : node10531;
															assign node10531 = (inp[3]) ? node10535 : node10532;
																assign node10532 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node10535 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node10538 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node10541 = (inp[4]) ? node10543 : 4'b0010;
														assign node10543 = (inp[9]) ? 4'b0100 : node10544;
															assign node10544 = (inp[0]) ? node10548 : node10545;
																assign node10545 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node10548 = (inp[3]) ? 4'b0010 : 4'b0000;
										assign node10552 = (inp[0]) ? node10606 : node10553;
											assign node10553 = (inp[3]) ? node10583 : node10554;
												assign node10554 = (inp[9]) ? node10574 : node10555;
													assign node10555 = (inp[4]) ? node10567 : node10556;
														assign node10556 = (inp[12]) ? node10562 : node10557;
															assign node10557 = (inp[8]) ? node10559 : 4'b0101;
																assign node10559 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node10562 = (inp[7]) ? 4'b0100 : node10563;
																assign node10563 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node10567 = (inp[8]) ? node10571 : node10568;
															assign node10568 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node10571 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node10574 = (inp[4]) ? node10578 : node10575;
														assign node10575 = (inp[12]) ? 4'b0000 : 4'b0001;
														assign node10578 = (inp[8]) ? 4'b0110 : node10579;
															assign node10579 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node10583 = (inp[7]) ? node10593 : node10584;
													assign node10584 = (inp[8]) ? node10588 : node10585;
														assign node10585 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node10588 = (inp[4]) ? node10590 : 4'b0011;
															assign node10590 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node10593 = (inp[8]) ? 4'b0110 : node10594;
														assign node10594 = (inp[12]) ? node10600 : node10595;
															assign node10595 = (inp[4]) ? 4'b0011 : node10596;
																assign node10596 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node10600 = (inp[4]) ? 4'b0111 : node10601;
																assign node10601 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node10606 = (inp[3]) ? node10628 : node10607;
												assign node10607 = (inp[9]) ? node10623 : node10608;
													assign node10608 = (inp[4]) ? node10614 : node10609;
														assign node10609 = (inp[8]) ? node10611 : 4'b0110;
															assign node10611 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node10614 = (inp[12]) ? 4'b0011 : node10615;
															assign node10615 = (inp[7]) ? node10619 : node10616;
																assign node10616 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node10619 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node10623 = (inp[4]) ? 4'b0100 : node10624;
														assign node10624 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node10628 = (inp[7]) ? node10640 : node10629;
													assign node10629 = (inp[8]) ? node10637 : node10630;
														assign node10630 = (inp[9]) ? node10634 : node10631;
															assign node10631 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node10634 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node10637 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node10640 = (inp[8]) ? node10648 : node10641;
														assign node10641 = (inp[9]) ? node10645 : node10642;
															assign node10642 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node10645 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node10648 = (inp[4]) ? node10650 : 4'b0100;
															assign node10650 = (inp[9]) ? 4'b0100 : 4'b0000;
									assign node10653 = (inp[4]) ? node10763 : node10654;
										assign node10654 = (inp[8]) ? node10714 : node10655;
											assign node10655 = (inp[7]) ? node10691 : node10656;
												assign node10656 = (inp[3]) ? node10674 : node10657;
													assign node10657 = (inp[15]) ? node10665 : node10658;
														assign node10658 = (inp[0]) ? 4'b0100 : node10659;
															assign node10659 = (inp[9]) ? node10661 : 4'b0010;
																assign node10661 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node10665 = (inp[0]) ? node10669 : node10666;
															assign node10666 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node10669 = (inp[9]) ? 4'b0010 : node10670;
																assign node10670 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node10674 = (inp[0]) ? node10686 : node10675;
														assign node10675 = (inp[15]) ? node10681 : node10676;
															assign node10676 = (inp[9]) ? node10678 : 4'b0000;
																assign node10678 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node10681 = (inp[12]) ? 4'b0010 : node10682;
																assign node10682 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node10686 = (inp[9]) ? node10688 : 4'b0000;
															assign node10688 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node10691 = (inp[0]) ? node10703 : node10692;
													assign node10692 = (inp[12]) ? node10700 : node10693;
														assign node10693 = (inp[9]) ? node10697 : node10694;
															assign node10694 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node10697 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node10700 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node10703 = (inp[9]) ? node10709 : node10704;
														assign node10704 = (inp[3]) ? node10706 : 4'b0001;
															assign node10706 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node10709 = (inp[15]) ? node10711 : 4'b0111;
															assign node10711 = (inp[3]) ? 4'b0001 : 4'b0101;
											assign node10714 = (inp[7]) ? node10736 : node10715;
												assign node10715 = (inp[3]) ? node10723 : node10716;
													assign node10716 = (inp[0]) ? 4'b0011 : node10717;
														assign node10717 = (inp[12]) ? 4'b0101 : node10718;
															assign node10718 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node10723 = (inp[0]) ? node10731 : node10724;
														assign node10724 = (inp[9]) ? node10728 : node10725;
															assign node10725 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node10728 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node10731 = (inp[12]) ? node10733 : 4'b0111;
															assign node10733 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node10736 = (inp[0]) ? node10750 : node10737;
													assign node10737 = (inp[15]) ? node10741 : node10738;
														assign node10738 = (inp[3]) ? 4'b0000 : 4'b0110;
														assign node10741 = (inp[9]) ? node10747 : node10742;
															assign node10742 = (inp[3]) ? node10744 : 4'b0000;
																assign node10744 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node10747 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node10750 = (inp[15]) ? node10760 : node10751;
														assign node10751 = (inp[3]) ? node10753 : 4'b0110;
															assign node10753 = (inp[9]) ? node10757 : node10754;
																assign node10754 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node10757 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node10760 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node10763 = (inp[15]) ? node10815 : node10764;
											assign node10764 = (inp[0]) ? node10788 : node10765;
												assign node10765 = (inp[12]) ? node10779 : node10766;
													assign node10766 = (inp[9]) ? node10772 : node10767;
														assign node10767 = (inp[3]) ? node10769 : 4'b0010;
															assign node10769 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node10772 = (inp[7]) ? node10776 : node10773;
															assign node10773 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node10776 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node10779 = (inp[9]) ? node10781 : 4'b0101;
														assign node10781 = (inp[8]) ? node10785 : node10782;
															assign node10782 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node10785 = (inp[7]) ? 4'b0000 : 4'b0001;
												assign node10788 = (inp[12]) ? node10800 : node10789;
													assign node10789 = (inp[9]) ? node10795 : node10790;
														assign node10790 = (inp[3]) ? 4'b0011 : node10791;
															assign node10791 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node10795 = (inp[8]) ? node10797 : 4'b0111;
															assign node10797 = (inp[7]) ? 4'b0110 : 4'b0111;
													assign node10800 = (inp[9]) ? node10810 : node10801;
														assign node10801 = (inp[3]) ? node10803 : 4'b0110;
															assign node10803 = (inp[7]) ? node10807 : node10804;
																assign node10804 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node10807 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node10810 = (inp[8]) ? 4'b0010 : node10811;
															assign node10811 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node10815 = (inp[0]) ? node10841 : node10816;
												assign node10816 = (inp[9]) ? node10830 : node10817;
													assign node10817 = (inp[12]) ? node10825 : node10818;
														assign node10818 = (inp[3]) ? 4'b0010 : node10819;
															assign node10819 = (inp[7]) ? 4'b0000 : node10820;
																assign node10820 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node10825 = (inp[7]) ? 4'b0111 : node10826;
															assign node10826 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node10830 = (inp[12]) ? node10836 : node10831;
														assign node10831 = (inp[7]) ? node10833 : 4'b0110;
															assign node10833 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node10836 = (inp[7]) ? node10838 : 4'b0010;
															assign node10838 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node10841 = (inp[9]) ? node10849 : node10842;
													assign node10842 = (inp[12]) ? node10846 : node10843;
														assign node10843 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node10846 = (inp[3]) ? 4'b0100 : 4'b0101;
													assign node10849 = (inp[12]) ? node10851 : 4'b0101;
														assign node10851 = (inp[7]) ? node10855 : node10852;
															assign node10852 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node10855 = (inp[8]) ? 4'b0000 : 4'b0001;
						assign node10858 = (inp[1]) ? node11624 : node10859;
							assign node10859 = (inp[2]) ? node11255 : node10860;
								assign node10860 = (inp[8]) ? node11066 : node10861;
									assign node10861 = (inp[7]) ? node10951 : node10862;
										assign node10862 = (inp[3]) ? node10896 : node10863;
											assign node10863 = (inp[9]) ? node10883 : node10864;
												assign node10864 = (inp[4]) ? node10872 : node10865;
													assign node10865 = (inp[10]) ? node10869 : node10866;
														assign node10866 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node10869 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node10872 = (inp[10]) ? node10874 : 4'b0011;
														assign node10874 = (inp[12]) ? 4'b0101 : node10875;
															assign node10875 = (inp[15]) ? node10879 : node10876;
																assign node10876 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node10879 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node10883 = (inp[15]) ? node10889 : node10884;
													assign node10884 = (inp[0]) ? 4'b0111 : node10885;
														assign node10885 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node10889 = (inp[0]) ? node10891 : 4'b0111;
														assign node10891 = (inp[4]) ? 4'b0101 : node10892;
															assign node10892 = (inp[12]) ? 4'b0101 : 4'b0011;
											assign node10896 = (inp[10]) ? node10920 : node10897;
												assign node10897 = (inp[9]) ? node10909 : node10898;
													assign node10898 = (inp[4]) ? node10904 : node10899;
														assign node10899 = (inp[0]) ? 4'b0111 : node10900;
															assign node10900 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node10904 = (inp[0]) ? node10906 : 4'b0011;
															assign node10906 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node10909 = (inp[4]) ? node10915 : node10910;
														assign node10910 = (inp[12]) ? node10912 : 4'b0001;
															assign node10912 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node10915 = (inp[15]) ? 4'b0101 : node10916;
															assign node10916 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node10920 = (inp[0]) ? node10938 : node10921;
													assign node10921 = (inp[15]) ? node10927 : node10922;
														assign node10922 = (inp[4]) ? node10924 : 4'b0001;
															assign node10924 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node10927 = (inp[4]) ? node10933 : node10928;
															assign node10928 = (inp[12]) ? 4'b0111 : node10929;
																assign node10929 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node10933 = (inp[12]) ? node10935 : 4'b0011;
																assign node10935 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node10938 = (inp[15]) ? node10944 : node10939;
														assign node10939 = (inp[9]) ? node10941 : 4'b0011;
															assign node10941 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node10944 = (inp[12]) ? node10946 : 4'b0001;
															assign node10946 = (inp[4]) ? node10948 : 4'b0001;
																assign node10948 = (inp[9]) ? 4'b0001 : 4'b0101;
										assign node10951 = (inp[15]) ? node11005 : node10952;
											assign node10952 = (inp[0]) ? node10978 : node10953;
												assign node10953 = (inp[3]) ? node10967 : node10954;
													assign node10954 = (inp[4]) ? node10958 : node10955;
														assign node10955 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node10958 = (inp[10]) ? node10962 : node10959;
															assign node10959 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node10962 = (inp[9]) ? node10964 : 4'b0100;
																assign node10964 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node10967 = (inp[4]) ? node10975 : node10968;
														assign node10968 = (inp[9]) ? node10970 : 4'b0100;
															assign node10970 = (inp[12]) ? node10972 : 4'b0000;
																assign node10972 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node10975 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node10978 = (inp[3]) ? node10996 : node10979;
													assign node10979 = (inp[4]) ? node10985 : node10980;
														assign node10980 = (inp[9]) ? 4'b0000 : node10981;
															assign node10981 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node10985 = (inp[9]) ? node10991 : node10986;
															assign node10986 = (inp[12]) ? node10988 : 4'b0000;
																assign node10988 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node10991 = (inp[10]) ? node10993 : 4'b0110;
																assign node10993 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node10996 = (inp[9]) ? node11000 : node10997;
														assign node10997 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node11000 = (inp[4]) ? 4'b0110 : node11001;
															assign node11001 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node11005 = (inp[0]) ? node11039 : node11006;
												assign node11006 = (inp[3]) ? node11018 : node11007;
													assign node11007 = (inp[9]) ? node11011 : node11008;
														assign node11008 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node11011 = (inp[12]) ? node11015 : node11012;
															assign node11012 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node11015 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node11018 = (inp[10]) ? node11024 : node11019;
														assign node11019 = (inp[12]) ? node11021 : 4'b0010;
															assign node11021 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node11024 = (inp[9]) ? node11032 : node11025;
															assign node11025 = (inp[4]) ? node11029 : node11026;
																assign node11026 = (inp[12]) ? 4'b0010 : 4'b0110;
																assign node11029 = (inp[12]) ? 4'b0110 : 4'b0010;
															assign node11032 = (inp[12]) ? node11036 : node11033;
																assign node11033 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node11036 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node11039 = (inp[3]) ? node11053 : node11040;
													assign node11040 = (inp[4]) ? node11044 : node11041;
														assign node11041 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node11044 = (inp[9]) ? node11050 : node11045;
															assign node11045 = (inp[12]) ? node11047 : 4'b0010;
																assign node11047 = (inp[10]) ? 4'b0100 : 4'b0010;
															assign node11050 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node11053 = (inp[12]) ? node11061 : node11054;
														assign node11054 = (inp[9]) ? node11058 : node11055;
															assign node11055 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node11058 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node11061 = (inp[9]) ? 4'b0000 : node11062;
															assign node11062 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node11066 = (inp[7]) ? node11164 : node11067;
										assign node11067 = (inp[9]) ? node11117 : node11068;
											assign node11068 = (inp[4]) ? node11090 : node11069;
												assign node11069 = (inp[12]) ? node11077 : node11070;
													assign node11070 = (inp[15]) ? 4'b0100 : node11071;
														assign node11071 = (inp[0]) ? 4'b0100 : node11072;
															assign node11072 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node11077 = (inp[10]) ? node11081 : node11078;
														assign node11078 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node11081 = (inp[3]) ? node11083 : 4'b0010;
															assign node11083 = (inp[0]) ? node11087 : node11084;
																assign node11084 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node11087 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node11090 = (inp[10]) ? node11104 : node11091;
													assign node11091 = (inp[3]) ? node11099 : node11092;
														assign node11092 = (inp[15]) ? node11096 : node11093;
															assign node11093 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node11096 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node11099 = (inp[0]) ? 4'b0010 : node11100;
															assign node11100 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node11104 = (inp[12]) ? node11112 : node11105;
														assign node11105 = (inp[0]) ? 4'b0000 : node11106;
															assign node11106 = (inp[3]) ? node11108 : 4'b0000;
																assign node11108 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node11112 = (inp[0]) ? node11114 : 4'b0110;
															assign node11114 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node11117 = (inp[4]) ? node11137 : node11118;
												assign node11118 = (inp[12]) ? node11124 : node11119;
													assign node11119 = (inp[10]) ? 4'b0010 : node11120;
														assign node11120 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node11124 = (inp[10]) ? node11126 : 4'b0000;
														assign node11126 = (inp[3]) ? node11132 : node11127;
															assign node11127 = (inp[0]) ? 4'b0100 : node11128;
																assign node11128 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node11132 = (inp[0]) ? 4'b0110 : node11133;
																assign node11133 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node11137 = (inp[10]) ? node11155 : node11138;
													assign node11138 = (inp[3]) ? node11146 : node11139;
														assign node11139 = (inp[0]) ? node11143 : node11140;
															assign node11140 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node11143 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node11146 = (inp[12]) ? 4'b0100 : node11147;
															assign node11147 = (inp[15]) ? node11151 : node11148;
																assign node11148 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node11151 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node11155 = (inp[12]) ? node11159 : node11156;
														assign node11156 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node11159 = (inp[0]) ? 4'b0000 : node11160;
															assign node11160 = (inp[15]) ? 4'b0010 : 4'b0000;
										assign node11164 = (inp[12]) ? node11210 : node11165;
											assign node11165 = (inp[3]) ? node11197 : node11166;
												assign node11166 = (inp[0]) ? node11186 : node11167;
													assign node11167 = (inp[15]) ? node11179 : node11168;
														assign node11168 = (inp[4]) ? node11174 : node11169;
															assign node11169 = (inp[9]) ? 4'b1011 : node11170;
																assign node11170 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node11174 = (inp[9]) ? node11176 : 4'b1011;
																assign node11176 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node11179 = (inp[4]) ? node11181 : 4'b1101;
															assign node11181 = (inp[10]) ? node11183 : 4'b1111;
																assign node11183 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node11186 = (inp[10]) ? node11192 : node11187;
														assign node11187 = (inp[9]) ? 4'b1111 : node11188;
															assign node11188 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node11192 = (inp[9]) ? node11194 : 4'b1101;
															assign node11194 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node11197 = (inp[0]) ? node11207 : node11198;
													assign node11198 = (inp[15]) ? node11204 : node11199;
														assign node11199 = (inp[4]) ? 4'b1001 : node11200;
															assign node11200 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node11204 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node11207 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node11210 = (inp[9]) ? node11230 : node11211;
												assign node11211 = (inp[4]) ? node11217 : node11212;
													assign node11212 = (inp[15]) ? 4'b1011 : node11213;
														assign node11213 = (inp[10]) ? 4'b1001 : 4'b1011;
													assign node11217 = (inp[10]) ? node11223 : node11218;
														assign node11218 = (inp[15]) ? node11220 : 4'b1101;
															assign node11220 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node11223 = (inp[0]) ? node11227 : node11224;
															assign node11224 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node11227 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node11230 = (inp[4]) ? node11242 : node11231;
													assign node11231 = (inp[3]) ? node11237 : node11232;
														assign node11232 = (inp[0]) ? node11234 : 4'b1101;
															assign node11234 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node11237 = (inp[15]) ? 4'b1111 : node11238;
															assign node11238 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node11242 = (inp[10]) ? node11248 : node11243;
														assign node11243 = (inp[15]) ? 4'b1011 : node11244;
															assign node11244 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node11248 = (inp[3]) ? node11252 : node11249;
															assign node11249 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node11252 = (inp[15]) ? 4'b1001 : 4'b1011;
								assign node11255 = (inp[7]) ? node11439 : node11256;
									assign node11256 = (inp[8]) ? node11342 : node11257;
										assign node11257 = (inp[15]) ? node11287 : node11258;
											assign node11258 = (inp[0]) ? node11276 : node11259;
												assign node11259 = (inp[3]) ? node11269 : node11260;
													assign node11260 = (inp[4]) ? node11264 : node11261;
														assign node11261 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node11264 = (inp[9]) ? 4'b0100 : node11265;
															assign node11265 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node11269 = (inp[12]) ? 4'b0100 : node11270;
														assign node11270 = (inp[10]) ? node11272 : 4'b0000;
															assign node11272 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node11276 = (inp[9]) ? node11282 : node11277;
													assign node11277 = (inp[3]) ? node11279 : 4'b0000;
														assign node11279 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node11282 = (inp[4]) ? 4'b0110 : node11283;
														assign node11283 = (inp[10]) ? 4'b0110 : 4'b0010;
											assign node11287 = (inp[0]) ? node11319 : node11288;
												assign node11288 = (inp[3]) ? node11304 : node11289;
													assign node11289 = (inp[10]) ? node11295 : node11290;
														assign node11290 = (inp[4]) ? node11292 : 4'b0000;
															assign node11292 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node11295 = (inp[9]) ? node11297 : 4'b0100;
															assign node11297 = (inp[12]) ? node11301 : node11298;
																assign node11298 = (inp[4]) ? 4'b0110 : 4'b0000;
																assign node11301 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node11304 = (inp[12]) ? node11310 : node11305;
														assign node11305 = (inp[9]) ? 4'b0110 : node11306;
															assign node11306 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node11310 = (inp[9]) ? 4'b0010 : node11311;
															assign node11311 = (inp[10]) ? node11315 : node11312;
																assign node11312 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node11315 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node11319 = (inp[3]) ? node11331 : node11320;
													assign node11320 = (inp[10]) ? node11328 : node11321;
														assign node11321 = (inp[4]) ? node11325 : node11322;
															assign node11322 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node11325 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node11328 = (inp[12]) ? 4'b0000 : 4'b0010;
													assign node11331 = (inp[9]) ? node11335 : node11332;
														assign node11332 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node11335 = (inp[4]) ? 4'b0100 : node11336;
															assign node11336 = (inp[12]) ? node11338 : 4'b0000;
																assign node11338 = (inp[10]) ? 4'b0100 : 4'b0000;
										assign node11342 = (inp[12]) ? node11394 : node11343;
											assign node11343 = (inp[9]) ? node11371 : node11344;
												assign node11344 = (inp[0]) ? node11354 : node11345;
													assign node11345 = (inp[15]) ? node11349 : node11346;
														assign node11346 = (inp[3]) ? 4'b1001 : 4'b1101;
														assign node11349 = (inp[3]) ? 4'b1111 : node11350;
															assign node11350 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node11354 = (inp[3]) ? node11368 : node11355;
														assign node11355 = (inp[15]) ? node11363 : node11356;
															assign node11356 = (inp[4]) ? node11360 : node11357;
																assign node11357 = (inp[10]) ? 4'b1001 : 4'b1101;
																assign node11360 = (inp[10]) ? 4'b1111 : 4'b1001;
															assign node11363 = (inp[10]) ? 4'b1011 : node11364;
																assign node11364 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node11368 = (inp[4]) ? 4'b1111 : 4'b1101;
												assign node11371 = (inp[0]) ? node11385 : node11372;
													assign node11372 = (inp[4]) ? node11380 : node11373;
														assign node11373 = (inp[10]) ? 4'b1111 : node11374;
															assign node11374 = (inp[15]) ? node11376 : 4'b1011;
																assign node11376 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node11380 = (inp[15]) ? 4'b1111 : node11381;
															assign node11381 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node11385 = (inp[15]) ? 4'b1101 : node11386;
														assign node11386 = (inp[3]) ? node11388 : 4'b1111;
															assign node11388 = (inp[10]) ? node11390 : 4'b1111;
																assign node11390 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node11394 = (inp[10]) ? node11406 : node11395;
												assign node11395 = (inp[9]) ? node11399 : node11396;
													assign node11396 = (inp[4]) ? 4'b1111 : 4'b1011;
													assign node11399 = (inp[4]) ? node11401 : 4'b1111;
														assign node11401 = (inp[15]) ? node11403 : 4'b1001;
															assign node11403 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node11406 = (inp[3]) ? node11424 : node11407;
													assign node11407 = (inp[9]) ? node11415 : node11408;
														assign node11408 = (inp[4]) ? 4'b1111 : node11409;
															assign node11409 = (inp[0]) ? 4'b1011 : node11410;
																assign node11410 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node11415 = (inp[4]) ? node11421 : node11416;
															assign node11416 = (inp[15]) ? 4'b1111 : node11417;
																assign node11417 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node11421 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node11424 = (inp[15]) ? node11430 : node11425;
														assign node11425 = (inp[4]) ? node11427 : 4'b1001;
															assign node11427 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node11430 = (inp[0]) ? node11436 : node11431;
															assign node11431 = (inp[9]) ? node11433 : 4'b1011;
																assign node11433 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node11436 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node11439 = (inp[8]) ? node11517 : node11440;
										assign node11440 = (inp[0]) ? node11482 : node11441;
											assign node11441 = (inp[15]) ? node11467 : node11442;
												assign node11442 = (inp[3]) ? node11454 : node11443;
													assign node11443 = (inp[4]) ? node11449 : node11444;
														assign node11444 = (inp[12]) ? 4'b1011 : node11445;
															assign node11445 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node11449 = (inp[12]) ? node11451 : 4'b1101;
															assign node11451 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node11454 = (inp[9]) ? node11462 : node11455;
														assign node11455 = (inp[4]) ? node11459 : node11456;
															assign node11456 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node11459 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node11462 = (inp[10]) ? 4'b1101 : node11463;
															assign node11463 = (inp[4]) ? 4'b1101 : 4'b1001;
												assign node11467 = (inp[9]) ? node11475 : node11468;
													assign node11468 = (inp[4]) ? node11470 : 4'b1001;
														assign node11470 = (inp[12]) ? 4'b1111 : node11471;
															assign node11471 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node11475 = (inp[4]) ? node11477 : 4'b1111;
														assign node11477 = (inp[10]) ? 4'b1011 : node11478;
															assign node11478 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node11482 = (inp[15]) ? node11498 : node11483;
												assign node11483 = (inp[3]) ? node11491 : node11484;
													assign node11484 = (inp[9]) ? 4'b1111 : node11485;
														assign node11485 = (inp[4]) ? node11487 : 4'b1001;
															assign node11487 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node11491 = (inp[12]) ? node11493 : 4'b1011;
														assign node11493 = (inp[10]) ? node11495 : 4'b1011;
															assign node11495 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node11498 = (inp[12]) ? node11510 : node11499;
													assign node11499 = (inp[10]) ? node11501 : 4'b1101;
														assign node11501 = (inp[4]) ? node11507 : node11502;
															assign node11502 = (inp[9]) ? 4'b1101 : node11503;
																assign node11503 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node11507 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node11510 = (inp[4]) ? 4'b1001 : node11511;
														assign node11511 = (inp[9]) ? 4'b1101 : node11512;
															assign node11512 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node11517 = (inp[12]) ? node11575 : node11518;
											assign node11518 = (inp[0]) ? node11548 : node11519;
												assign node11519 = (inp[15]) ? node11535 : node11520;
													assign node11520 = (inp[9]) ? 4'b1100 : node11521;
														assign node11521 = (inp[3]) ? node11527 : node11522;
															assign node11522 = (inp[4]) ? node11524 : 4'b1010;
																assign node11524 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node11527 = (inp[10]) ? node11531 : node11528;
																assign node11528 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node11531 = (inp[4]) ? 4'b1100 : 4'b1000;
													assign node11535 = (inp[3]) ? node11541 : node11536;
														assign node11536 = (inp[10]) ? node11538 : 4'b1000;
															assign node11538 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node11541 = (inp[10]) ? 4'b1010 : node11542;
															assign node11542 = (inp[9]) ? node11544 : 4'b1110;
																assign node11544 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node11548 = (inp[15]) ? node11560 : node11549;
													assign node11549 = (inp[9]) ? node11551 : 4'b1110;
														assign node11551 = (inp[10]) ? node11557 : node11552;
															assign node11552 = (inp[4]) ? 4'b1110 : node11553;
																assign node11553 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node11557 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node11560 = (inp[3]) ? node11570 : node11561;
														assign node11561 = (inp[4]) ? node11567 : node11562;
															assign node11562 = (inp[10]) ? 4'b1010 : node11563;
																assign node11563 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node11567 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node11570 = (inp[9]) ? 4'b1100 : node11571;
															assign node11571 = (inp[10]) ? 4'b1000 : 4'b1100;
											assign node11575 = (inp[0]) ? node11605 : node11576;
												assign node11576 = (inp[15]) ? node11592 : node11577;
													assign node11577 = (inp[3]) ? node11585 : node11578;
														assign node11578 = (inp[9]) ? node11582 : node11579;
															assign node11579 = (inp[4]) ? 4'b1100 : 4'b1010;
															assign node11582 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node11585 = (inp[9]) ? node11589 : node11586;
															assign node11586 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node11589 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node11592 = (inp[10]) ? node11598 : node11593;
														assign node11593 = (inp[9]) ? node11595 : 4'b1010;
															assign node11595 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node11598 = (inp[4]) ? node11602 : node11599;
															assign node11599 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node11602 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node11605 = (inp[15]) ? node11617 : node11606;
													assign node11606 = (inp[10]) ? node11612 : node11607;
														assign node11607 = (inp[4]) ? 4'b1110 : node11608;
															assign node11608 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node11612 = (inp[9]) ? node11614 : 4'b1110;
															assign node11614 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node11617 = (inp[9]) ? node11621 : node11618;
														assign node11618 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node11621 = (inp[4]) ? 4'b1000 : 4'b1100;
							assign node11624 = (inp[9]) ? node12076 : node11625;
								assign node11625 = (inp[4]) ? node11887 : node11626;
									assign node11626 = (inp[10]) ? node11752 : node11627;
										assign node11627 = (inp[12]) ? node11689 : node11628;
											assign node11628 = (inp[0]) ? node11662 : node11629;
												assign node11629 = (inp[3]) ? node11649 : node11630;
													assign node11630 = (inp[15]) ? node11644 : node11631;
														assign node11631 = (inp[2]) ? node11637 : node11632;
															assign node11632 = (inp[8]) ? node11634 : 4'b1111;
																assign node11634 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node11637 = (inp[7]) ? node11641 : node11638;
																assign node11638 = (inp[8]) ? 4'b1111 : 4'b1110;
																assign node11641 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node11644 = (inp[8]) ? node11646 : 4'b1101;
															assign node11646 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node11649 = (inp[15]) ? node11659 : node11650;
														assign node11650 = (inp[2]) ? node11652 : 4'b1101;
															assign node11652 = (inp[8]) ? node11656 : node11653;
																assign node11653 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node11656 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node11659 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node11662 = (inp[8]) ? node11678 : node11663;
													assign node11663 = (inp[2]) ? node11667 : node11664;
														assign node11664 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node11667 = (inp[7]) ? node11675 : node11668;
															assign node11668 = (inp[15]) ? node11672 : node11669;
																assign node11669 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node11672 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node11675 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node11678 = (inp[2]) ? node11682 : node11679;
														assign node11679 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node11682 = (inp[7]) ? node11684 : 4'b1111;
															assign node11684 = (inp[3]) ? 4'b1110 : node11685;
																assign node11685 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node11689 = (inp[15]) ? node11719 : node11690;
												assign node11690 = (inp[2]) ? node11702 : node11691;
													assign node11691 = (inp[8]) ? 4'b1011 : node11692;
														assign node11692 = (inp[7]) ? node11698 : node11693;
															assign node11693 = (inp[3]) ? node11695 : 4'b1011;
																assign node11695 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node11698 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node11702 = (inp[3]) ? node11708 : node11703;
														assign node11703 = (inp[0]) ? node11705 : 4'b1010;
															assign node11705 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node11708 = (inp[0]) ? node11714 : node11709;
															assign node11709 = (inp[8]) ? node11711 : 4'b1001;
																assign node11711 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node11714 = (inp[7]) ? 4'b1010 : node11715;
																assign node11715 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node11719 = (inp[2]) ? node11733 : node11720;
													assign node11720 = (inp[3]) ? node11728 : node11721;
														assign node11721 = (inp[7]) ? node11725 : node11722;
															assign node11722 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node11725 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node11728 = (inp[7]) ? 4'b1010 : node11729;
															assign node11729 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node11733 = (inp[8]) ? node11745 : node11734;
														assign node11734 = (inp[7]) ? node11740 : node11735;
															assign node11735 = (inp[3]) ? 4'b1010 : node11736;
																assign node11736 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node11740 = (inp[0]) ? 4'b1001 : node11741;
																assign node11741 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node11745 = (inp[0]) ? node11749 : node11746;
															assign node11746 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node11749 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node11752 = (inp[8]) ? node11820 : node11753;
											assign node11753 = (inp[12]) ? node11789 : node11754;
												assign node11754 = (inp[0]) ? node11774 : node11755;
													assign node11755 = (inp[2]) ? node11763 : node11756;
														assign node11756 = (inp[7]) ? 4'b1010 : node11757;
															assign node11757 = (inp[15]) ? 4'b1001 : node11758;
																assign node11758 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node11763 = (inp[7]) ? node11769 : node11764;
															assign node11764 = (inp[15]) ? node11766 : 4'b1000;
																assign node11766 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node11769 = (inp[15]) ? node11771 : 4'b1001;
																assign node11771 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node11774 = (inp[3]) ? node11778 : node11775;
														assign node11775 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node11778 = (inp[15]) ? node11786 : node11779;
															assign node11779 = (inp[2]) ? node11783 : node11780;
																assign node11780 = (inp[7]) ? 4'b1010 : 4'b1011;
																assign node11783 = (inp[7]) ? 4'b1011 : 4'b1010;
															assign node11786 = (inp[7]) ? 4'b1000 : 4'b1001;
												assign node11789 = (inp[15]) ? node11805 : node11790;
													assign node11790 = (inp[3]) ? node11802 : node11791;
														assign node11791 = (inp[0]) ? node11795 : node11792;
															assign node11792 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node11795 = (inp[2]) ? node11799 : node11796;
																assign node11796 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node11799 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node11802 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node11805 = (inp[3]) ? node11815 : node11806;
														assign node11806 = (inp[0]) ? node11812 : node11807;
															assign node11807 = (inp[7]) ? 4'b1000 : node11808;
																assign node11808 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node11812 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node11815 = (inp[7]) ? node11817 : 4'b1011;
															assign node11817 = (inp[2]) ? 4'b1001 : 4'b1000;
											assign node11820 = (inp[3]) ? node11858 : node11821;
												assign node11821 = (inp[15]) ? node11839 : node11822;
													assign node11822 = (inp[0]) ? node11830 : node11823;
														assign node11823 = (inp[12]) ? 4'b1010 : node11824;
															assign node11824 = (inp[7]) ? 4'b1011 : node11825;
																assign node11825 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node11830 = (inp[12]) ? 4'b1000 : node11831;
															assign node11831 = (inp[2]) ? node11835 : node11832;
																assign node11832 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node11835 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node11839 = (inp[0]) ? node11843 : node11840;
														assign node11840 = (inp[12]) ? 4'b1001 : 4'b1000;
														assign node11843 = (inp[12]) ? node11851 : node11844;
															assign node11844 = (inp[7]) ? node11848 : node11845;
																assign node11845 = (inp[2]) ? 4'b1011 : 4'b1010;
																assign node11848 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node11851 = (inp[2]) ? node11855 : node11852;
																assign node11852 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node11855 = (inp[7]) ? 4'b1010 : 4'b1011;
												assign node11858 = (inp[12]) ? node11880 : node11859;
													assign node11859 = (inp[7]) ? node11869 : node11860;
														assign node11860 = (inp[2]) ? node11862 : 4'b1000;
															assign node11862 = (inp[15]) ? node11866 : node11863;
																assign node11863 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node11866 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node11869 = (inp[2]) ? node11875 : node11870;
															assign node11870 = (inp[0]) ? 4'b1011 : node11871;
																assign node11871 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node11875 = (inp[0]) ? node11877 : 4'b1010;
																assign node11877 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node11880 = (inp[7]) ? node11884 : node11881;
														assign node11881 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node11884 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node11887 = (inp[12]) ? node11981 : node11888;
										assign node11888 = (inp[10]) ? node11940 : node11889;
											assign node11889 = (inp[15]) ? node11907 : node11890;
												assign node11890 = (inp[3]) ? node11900 : node11891;
													assign node11891 = (inp[0]) ? node11893 : 4'b1010;
														assign node11893 = (inp[2]) ? 4'b1000 : node11894;
															assign node11894 = (inp[7]) ? node11896 : 4'b1001;
																assign node11896 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node11900 = (inp[0]) ? node11904 : node11901;
														assign node11901 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node11904 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node11907 = (inp[0]) ? node11923 : node11908;
													assign node11908 = (inp[3]) ? node11918 : node11909;
														assign node11909 = (inp[7]) ? 4'b1001 : node11910;
															assign node11910 = (inp[2]) ? node11914 : node11911;
																assign node11911 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node11914 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node11918 = (inp[2]) ? node11920 : 4'b1010;
															assign node11920 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node11923 = (inp[3]) ? node11937 : node11924;
														assign node11924 = (inp[7]) ? node11932 : node11925;
															assign node11925 = (inp[8]) ? node11929 : node11926;
																assign node11926 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node11929 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node11932 = (inp[2]) ? node11934 : 4'b1011;
																assign node11934 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node11937 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node11940 = (inp[0]) ? node11960 : node11941;
												assign node11941 = (inp[15]) ? node11951 : node11942;
													assign node11942 = (inp[7]) ? node11948 : node11943;
														assign node11943 = (inp[2]) ? node11945 : 4'b1101;
															assign node11945 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node11948 = (inp[3]) ? 4'b1100 : 4'b1101;
													assign node11951 = (inp[2]) ? 4'b1111 : node11952;
														assign node11952 = (inp[7]) ? node11956 : node11953;
															assign node11953 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node11956 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node11960 = (inp[15]) ? node11968 : node11961;
													assign node11961 = (inp[7]) ? 4'b1110 : node11962;
														assign node11962 = (inp[2]) ? node11964 : 4'b1111;
															assign node11964 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node11968 = (inp[8]) ? node11974 : node11969;
														assign node11969 = (inp[2]) ? node11971 : 4'b1100;
															assign node11971 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node11974 = (inp[7]) ? node11978 : node11975;
															assign node11975 = (inp[3]) ? 4'b1101 : 4'b1100;
															assign node11978 = (inp[3]) ? 4'b1100 : 4'b1101;
										assign node11981 = (inp[10]) ? node12035 : node11982;
											assign node11982 = (inp[8]) ? node12008 : node11983;
												assign node11983 = (inp[7]) ? node11995 : node11984;
													assign node11984 = (inp[2]) ? node11988 : node11985;
														assign node11985 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node11988 = (inp[3]) ? 4'b1100 : node11989;
															assign node11989 = (inp[15]) ? 4'b1110 : node11990;
																assign node11990 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node11995 = (inp[2]) ? node12001 : node11996;
														assign node11996 = (inp[0]) ? node11998 : 4'b1100;
															assign node11998 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node12001 = (inp[3]) ? 4'b1101 : node12002;
															assign node12002 = (inp[0]) ? node12004 : 4'b1111;
																assign node12004 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node12008 = (inp[3]) ? node12018 : node12009;
													assign node12009 = (inp[0]) ? node12015 : node12010;
														assign node12010 = (inp[2]) ? 4'b1101 : node12011;
															assign node12011 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node12015 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node12018 = (inp[0]) ? node12026 : node12019;
														assign node12019 = (inp[15]) ? 4'b1111 : node12020;
															assign node12020 = (inp[2]) ? node12022 : 4'b1100;
																assign node12022 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node12026 = (inp[15]) ? node12028 : 4'b1111;
															assign node12028 = (inp[2]) ? node12032 : node12029;
																assign node12029 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node12032 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node12035 = (inp[2]) ? node12053 : node12036;
												assign node12036 = (inp[7]) ? node12044 : node12037;
													assign node12037 = (inp[8]) ? node12039 : 4'b1101;
														assign node12039 = (inp[15]) ? 4'b1100 : node12040;
															assign node12040 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node12044 = (inp[8]) ? 4'b1111 : node12045;
														assign node12045 = (inp[15]) ? node12049 : node12046;
															assign node12046 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node12049 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node12053 = (inp[15]) ? node12067 : node12054;
													assign node12054 = (inp[0]) ? node12060 : node12055;
														assign node12055 = (inp[7]) ? node12057 : 4'b1101;
															assign node12057 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node12060 = (inp[7]) ? node12064 : node12061;
															assign node12061 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node12064 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node12067 = (inp[0]) ? node12069 : 4'b1110;
														assign node12069 = (inp[3]) ? node12073 : node12070;
															assign node12070 = (inp[7]) ? 4'b1101 : 4'b1100;
															assign node12073 = (inp[7]) ? 4'b1100 : 4'b1101;
								assign node12076 = (inp[4]) ? node12278 : node12077;
									assign node12077 = (inp[10]) ? node12175 : node12078;
										assign node12078 = (inp[12]) ? node12132 : node12079;
											assign node12079 = (inp[3]) ? node12107 : node12080;
												assign node12080 = (inp[0]) ? node12100 : node12081;
													assign node12081 = (inp[15]) ? node12087 : node12082;
														assign node12082 = (inp[2]) ? node12084 : 4'b1011;
															assign node12084 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node12087 = (inp[7]) ? node12095 : node12088;
															assign node12088 = (inp[2]) ? node12092 : node12089;
																assign node12089 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node12092 = (inp[8]) ? 4'b1001 : 4'b1000;
															assign node12095 = (inp[8]) ? node12097 : 4'b1000;
																assign node12097 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node12100 = (inp[15]) ? 4'b1011 : node12101;
														assign node12101 = (inp[8]) ? 4'b1001 : node12102;
															assign node12102 = (inp[7]) ? 4'b1001 : 4'b1000;
												assign node12107 = (inp[8]) ? node12125 : node12108;
													assign node12108 = (inp[0]) ? node12116 : node12109;
														assign node12109 = (inp[15]) ? node12111 : 4'b1000;
															assign node12111 = (inp[7]) ? node12113 : 4'b1011;
																assign node12113 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node12116 = (inp[15]) ? 4'b1000 : node12117;
															assign node12117 = (inp[7]) ? node12121 : node12118;
																assign node12118 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node12121 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node12125 = (inp[7]) ? node12129 : node12126;
														assign node12126 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node12129 = (inp[2]) ? 4'b1000 : 4'b1001;
											assign node12132 = (inp[7]) ? node12146 : node12133;
												assign node12133 = (inp[8]) ? node12137 : node12134;
													assign node12134 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node12137 = (inp[2]) ? node12141 : node12138;
														assign node12138 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node12141 = (inp[15]) ? 4'b1111 : node12142;
															assign node12142 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node12146 = (inp[8]) ? node12162 : node12147;
													assign node12147 = (inp[2]) ? node12155 : node12148;
														assign node12148 = (inp[15]) ? node12152 : node12149;
															assign node12149 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node12152 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node12155 = (inp[3]) ? node12157 : 4'b1101;
															assign node12157 = (inp[0]) ? node12159 : 4'b1111;
																assign node12159 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node12162 = (inp[2]) ? node12172 : node12163;
														assign node12163 = (inp[3]) ? node12167 : node12164;
															assign node12164 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node12167 = (inp[0]) ? 4'b1101 : node12168;
																assign node12168 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node12172 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node12175 = (inp[3]) ? node12235 : node12176;
											assign node12176 = (inp[7]) ? node12204 : node12177;
												assign node12177 = (inp[0]) ? node12193 : node12178;
													assign node12178 = (inp[15]) ? node12188 : node12179;
														assign node12179 = (inp[12]) ? 4'b1100 : node12180;
															assign node12180 = (inp[2]) ? node12184 : node12181;
																assign node12181 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node12184 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node12188 = (inp[8]) ? 4'b1111 : node12189;
															assign node12189 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node12193 = (inp[15]) ? 4'b1100 : node12194;
														assign node12194 = (inp[12]) ? 4'b1111 : node12195;
															assign node12195 = (inp[2]) ? node12199 : node12196;
																assign node12196 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node12199 = (inp[8]) ? 4'b1111 : 4'b1110;
												assign node12204 = (inp[12]) ? node12212 : node12205;
													assign node12205 = (inp[0]) ? node12209 : node12206;
														assign node12206 = (inp[2]) ? 4'b1100 : 4'b1111;
														assign node12209 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node12212 = (inp[15]) ? node12222 : node12213;
														assign node12213 = (inp[0]) ? 4'b1111 : node12214;
															assign node12214 = (inp[2]) ? node12218 : node12215;
																assign node12215 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node12218 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node12222 = (inp[0]) ? node12228 : node12223;
															assign node12223 = (inp[8]) ? 4'b1111 : node12224;
																assign node12224 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node12228 = (inp[8]) ? node12232 : node12229;
																assign node12229 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node12232 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node12235 = (inp[7]) ? node12259 : node12236;
												assign node12236 = (inp[12]) ? node12248 : node12237;
													assign node12237 = (inp[15]) ? node12241 : node12238;
														assign node12238 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node12241 = (inp[0]) ? node12243 : 4'b1111;
															assign node12243 = (inp[2]) ? 4'b1101 : node12244;
																assign node12244 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node12248 = (inp[0]) ? node12252 : node12249;
														assign node12249 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node12252 = (inp[8]) ? node12256 : node12253;
															assign node12253 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node12256 = (inp[2]) ? 4'b1111 : 4'b1110;
												assign node12259 = (inp[8]) ? node12267 : node12260;
													assign node12260 = (inp[2]) ? 4'b1111 : node12261;
														assign node12261 = (inp[0]) ? node12263 : 4'b1110;
															assign node12263 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node12267 = (inp[2]) ? node12271 : node12268;
														assign node12268 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node12271 = (inp[0]) ? node12275 : node12272;
															assign node12272 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node12275 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node12278 = (inp[12]) ? node12376 : node12279;
										assign node12279 = (inp[10]) ? node12329 : node12280;
											assign node12280 = (inp[15]) ? node12304 : node12281;
												assign node12281 = (inp[0]) ? node12287 : node12282;
													assign node12282 = (inp[3]) ? 4'b1101 : node12283;
														assign node12283 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node12287 = (inp[3]) ? node12299 : node12288;
														assign node12288 = (inp[8]) ? node12294 : node12289;
															assign node12289 = (inp[7]) ? node12291 : 4'b1110;
																assign node12291 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node12294 = (inp[2]) ? node12296 : 4'b1111;
																assign node12296 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node12299 = (inp[7]) ? 4'b1111 : node12300;
															assign node12300 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node12304 = (inp[0]) ? node12314 : node12305;
													assign node12305 = (inp[7]) ? node12307 : 4'b1110;
														assign node12307 = (inp[8]) ? node12311 : node12308;
															assign node12308 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node12311 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node12314 = (inp[8]) ? node12324 : node12315;
														assign node12315 = (inp[3]) ? 4'b1100 : node12316;
															assign node12316 = (inp[2]) ? node12320 : node12317;
																assign node12317 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node12320 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node12324 = (inp[3]) ? 4'b1101 : node12325;
															assign node12325 = (inp[7]) ? 4'b1101 : 4'b1100;
											assign node12329 = (inp[0]) ? node12345 : node12330;
												assign node12330 = (inp[15]) ? node12336 : node12331;
													assign node12331 = (inp[2]) ? node12333 : 4'b1001;
														assign node12333 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node12336 = (inp[2]) ? node12338 : 4'b1011;
														assign node12338 = (inp[7]) ? node12342 : node12339;
															assign node12339 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node12342 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node12345 = (inp[15]) ? node12363 : node12346;
													assign node12346 = (inp[3]) ? node12356 : node12347;
														assign node12347 = (inp[7]) ? node12349 : 4'b1010;
															assign node12349 = (inp[2]) ? node12353 : node12350;
																assign node12350 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node12353 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node12356 = (inp[2]) ? 4'b1011 : node12357;
															assign node12357 = (inp[8]) ? node12359 : 4'b1011;
																assign node12359 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node12363 = (inp[8]) ? node12369 : node12364;
														assign node12364 = (inp[2]) ? 4'b1001 : node12365;
															assign node12365 = (inp[3]) ? 4'b1000 : 4'b1001;
														assign node12369 = (inp[7]) ? node12373 : node12370;
															assign node12370 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node12373 = (inp[2]) ? 4'b1000 : 4'b1001;
										assign node12376 = (inp[2]) ? node12440 : node12377;
											assign node12377 = (inp[3]) ? node12411 : node12378;
												assign node12378 = (inp[10]) ? node12394 : node12379;
													assign node12379 = (inp[7]) ? node12385 : node12380;
														assign node12380 = (inp[15]) ? 4'b1001 : node12381;
															assign node12381 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node12385 = (inp[8]) ? node12391 : node12386;
															assign node12386 = (inp[15]) ? node12388 : 4'b1000;
																assign node12388 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node12391 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node12394 = (inp[15]) ? node12402 : node12395;
														assign node12395 = (inp[0]) ? node12397 : 4'b1001;
															assign node12397 = (inp[8]) ? node12399 : 4'b1010;
																assign node12399 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node12402 = (inp[0]) ? 4'b1001 : node12403;
															assign node12403 = (inp[7]) ? node12407 : node12404;
																assign node12404 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node12407 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node12411 = (inp[15]) ? node12423 : node12412;
													assign node12412 = (inp[0]) ? node12418 : node12413;
														assign node12413 = (inp[8]) ? node12415 : 4'b1000;
															assign node12415 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node12418 = (inp[7]) ? 4'b1010 : node12419;
															assign node12419 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node12423 = (inp[0]) ? node12435 : node12424;
														assign node12424 = (inp[10]) ? node12430 : node12425;
															assign node12425 = (inp[8]) ? 4'b1011 : node12426;
																assign node12426 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node12430 = (inp[8]) ? 4'b1010 : node12431;
																assign node12431 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node12435 = (inp[8]) ? 4'b1000 : node12436;
															assign node12436 = (inp[7]) ? 4'b1000 : 4'b1001;
											assign node12440 = (inp[10]) ? node12472 : node12441;
												assign node12441 = (inp[8]) ? node12459 : node12442;
													assign node12442 = (inp[7]) ? node12454 : node12443;
														assign node12443 = (inp[3]) ? node12449 : node12444;
															assign node12444 = (inp[0]) ? 4'b1000 : node12445;
																assign node12445 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node12449 = (inp[15]) ? node12451 : 4'b1010;
																assign node12451 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node12454 = (inp[15]) ? 4'b1001 : node12455;
															assign node12455 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node12459 = (inp[7]) ? node12467 : node12460;
														assign node12460 = (inp[15]) ? node12464 : node12461;
															assign node12461 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node12464 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node12467 = (inp[15]) ? node12469 : 4'b1010;
															assign node12469 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node12472 = (inp[0]) ? node12486 : node12473;
													assign node12473 = (inp[15]) ? node12479 : node12474;
														assign node12474 = (inp[8]) ? node12476 : 4'b1001;
															assign node12476 = (inp[7]) ? 4'b1000 : 4'b1001;
														assign node12479 = (inp[3]) ? node12481 : 4'b1011;
															assign node12481 = (inp[7]) ? node12483 : 4'b1010;
																assign node12483 = (inp[8]) ? 4'b1010 : 4'b1011;
													assign node12486 = (inp[15]) ? node12488 : 4'b1010;
														assign node12488 = (inp[3]) ? node12490 : 4'b1000;
															assign node12490 = (inp[7]) ? 4'b1001 : 4'b1000;
			assign node12493 = (inp[6]) ? node18743 : node12494;
				assign node12494 = (inp[13]) ? node15692 : node12495;
					assign node12495 = (inp[1]) ? node14201 : node12496;
						assign node12496 = (inp[7]) ? node13370 : node12497;
							assign node12497 = (inp[5]) ? node12917 : node12498;
								assign node12498 = (inp[15]) ? node12704 : node12499;
									assign node12499 = (inp[0]) ? node12605 : node12500;
										assign node12500 = (inp[3]) ? node12554 : node12501;
											assign node12501 = (inp[4]) ? node12521 : node12502;
												assign node12502 = (inp[2]) ? node12512 : node12503;
													assign node12503 = (inp[8]) ? node12509 : node12504;
														assign node12504 = (inp[12]) ? node12506 : 4'b0011;
															assign node12506 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node12509 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node12512 = (inp[8]) ? 4'b0011 : node12513;
														assign node12513 = (inp[9]) ? node12517 : node12514;
															assign node12514 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node12517 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node12521 = (inp[9]) ? node12537 : node12522;
													assign node12522 = (inp[10]) ? node12530 : node12523;
														assign node12523 = (inp[2]) ? node12527 : node12524;
															assign node12524 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node12527 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node12530 = (inp[12]) ? node12532 : 4'b0011;
															assign node12532 = (inp[2]) ? node12534 : 4'b0111;
																assign node12534 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node12537 = (inp[12]) ? node12551 : node12538;
														assign node12538 = (inp[10]) ? node12544 : node12539;
															assign node12539 = (inp[2]) ? node12541 : 4'b0111;
																assign node12541 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node12544 = (inp[8]) ? node12548 : node12545;
																assign node12545 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node12548 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node12551 = (inp[10]) ? 4'b0011 : 4'b0110;
											assign node12554 = (inp[9]) ? node12582 : node12555;
												assign node12555 = (inp[4]) ? node12569 : node12556;
													assign node12556 = (inp[10]) ? node12566 : node12557;
														assign node12557 = (inp[12]) ? node12559 : 4'b0111;
															assign node12559 = (inp[8]) ? node12563 : node12560;
																assign node12560 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node12563 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node12566 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node12569 = (inp[10]) ? node12579 : node12570;
														assign node12570 = (inp[12]) ? 4'b0010 : node12571;
															assign node12571 = (inp[2]) ? node12575 : node12572;
																assign node12572 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node12575 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node12579 = (inp[12]) ? 4'b0101 : 4'b0011;
												assign node12582 = (inp[4]) ? node12596 : node12583;
													assign node12583 = (inp[10]) ? node12587 : node12584;
														assign node12584 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node12587 = (inp[12]) ? node12591 : node12588;
															assign node12588 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node12591 = (inp[2]) ? 4'b0100 : node12592;
																assign node12592 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node12596 = (inp[10]) ? node12602 : node12597;
														assign node12597 = (inp[2]) ? 4'b0101 : node12598;
															assign node12598 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node12602 = (inp[2]) ? 4'b0000 : 4'b0001;
										assign node12605 = (inp[3]) ? node12651 : node12606;
											assign node12606 = (inp[10]) ? node12634 : node12607;
												assign node12607 = (inp[8]) ? node12625 : node12608;
													assign node12608 = (inp[2]) ? node12618 : node12609;
														assign node12609 = (inp[12]) ? 4'b0001 : node12610;
															assign node12610 = (inp[9]) ? node12614 : node12611;
																assign node12611 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node12614 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node12618 = (inp[4]) ? node12622 : node12619;
															assign node12619 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node12622 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node12625 = (inp[2]) ? node12627 : 4'b0000;
														assign node12627 = (inp[4]) ? node12631 : node12628;
															assign node12628 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node12631 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node12634 = (inp[12]) ? 4'b0101 : node12635;
													assign node12635 = (inp[2]) ? node12643 : node12636;
														assign node12636 = (inp[8]) ? node12638 : 4'b0001;
															assign node12638 = (inp[4]) ? 4'b0000 : node12639;
																assign node12639 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node12643 = (inp[8]) ? node12645 : 4'b0100;
															assign node12645 = (inp[9]) ? node12647 : 4'b0001;
																assign node12647 = (inp[4]) ? 4'b0101 : 4'b0001;
											assign node12651 = (inp[4]) ? node12685 : node12652;
												assign node12652 = (inp[12]) ? node12664 : node12653;
													assign node12653 = (inp[9]) ? node12655 : 4'b0101;
														assign node12655 = (inp[10]) ? node12661 : node12656;
															assign node12656 = (inp[8]) ? 4'b0001 : node12657;
																assign node12657 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node12661 = (inp[2]) ? 4'b0001 : 4'b0000;
													assign node12664 = (inp[10]) ? node12676 : node12665;
														assign node12665 = (inp[9]) ? node12671 : node12666;
															assign node12666 = (inp[2]) ? node12668 : 4'b0100;
																assign node12668 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node12671 = (inp[2]) ? 4'b0001 : node12672;
																assign node12672 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node12676 = (inp[9]) ? node12680 : node12677;
															assign node12677 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node12680 = (inp[8]) ? 4'b0110 : node12681;
																assign node12681 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node12685 = (inp[9]) ? node12691 : node12686;
													assign node12686 = (inp[2]) ? 4'b0111 : node12687;
														assign node12687 = (inp[8]) ? 4'b0000 : 4'b0001;
													assign node12691 = (inp[12]) ? node12697 : node12692;
														assign node12692 = (inp[2]) ? node12694 : 4'b0111;
															assign node12694 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node12697 = (inp[10]) ? node12701 : node12698;
															assign node12698 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node12701 = (inp[2]) ? 4'b0010 : 4'b0011;
									assign node12704 = (inp[0]) ? node12816 : node12705;
										assign node12705 = (inp[3]) ? node12755 : node12706;
											assign node12706 = (inp[10]) ? node12728 : node12707;
												assign node12707 = (inp[12]) ? node12717 : node12708;
													assign node12708 = (inp[9]) ? node12714 : node12709;
														assign node12709 = (inp[4]) ? node12711 : 4'b0100;
															assign node12711 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node12714 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node12717 = (inp[8]) ? node12725 : node12718;
														assign node12718 = (inp[2]) ? node12720 : 4'b0101;
															assign node12720 = (inp[9]) ? node12722 : 4'b0100;
																assign node12722 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node12725 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node12728 = (inp[4]) ? node12742 : node12729;
													assign node12729 = (inp[2]) ? node12735 : node12730;
														assign node12730 = (inp[8]) ? 4'b0000 : node12731;
															assign node12731 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node12735 = (inp[8]) ? 4'b0101 : node12736;
															assign node12736 = (inp[9]) ? node12738 : 4'b0000;
																assign node12738 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node12742 = (inp[9]) ? node12750 : node12743;
														assign node12743 = (inp[12]) ? node12745 : 4'b0001;
															assign node12745 = (inp[2]) ? 4'b0101 : node12746;
																assign node12746 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node12750 = (inp[12]) ? 4'b0001 : node12751;
															assign node12751 = (inp[2]) ? 4'b0100 : 4'b0101;
											assign node12755 = (inp[4]) ? node12785 : node12756;
												assign node12756 = (inp[9]) ? node12772 : node12757;
													assign node12757 = (inp[12]) ? node12767 : node12758;
														assign node12758 = (inp[10]) ? node12760 : 4'b0100;
															assign node12760 = (inp[2]) ? node12764 : node12761;
																assign node12761 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node12764 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node12767 = (inp[10]) ? 4'b0000 : node12768;
															assign node12768 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node12772 = (inp[8]) ? node12782 : node12773;
														assign node12773 = (inp[2]) ? node12777 : node12774;
															assign node12774 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node12777 = (inp[10]) ? node12779 : 4'b0000;
																assign node12779 = (inp[12]) ? 4'b0110 : 4'b0000;
														assign node12782 = (inp[2]) ? 4'b0001 : 4'b0000;
												assign node12785 = (inp[9]) ? node12801 : node12786;
													assign node12786 = (inp[10]) ? node12794 : node12787;
														assign node12787 = (inp[8]) ? node12791 : node12788;
															assign node12788 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node12791 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node12794 = (inp[12]) ? node12796 : 4'b0000;
															assign node12796 = (inp[8]) ? node12798 : 4'b0110;
																assign node12798 = (inp[2]) ? 4'b0111 : 4'b0110;
													assign node12801 = (inp[12]) ? node12807 : node12802;
														assign node12802 = (inp[8]) ? 4'b0110 : node12803;
															assign node12803 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node12807 = (inp[10]) ? node12813 : node12808;
															assign node12808 = (inp[8]) ? node12810 : 4'b0110;
																assign node12810 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node12813 = (inp[2]) ? 4'b0010 : 4'b0011;
										assign node12816 = (inp[3]) ? node12862 : node12817;
											assign node12817 = (inp[2]) ? node12843 : node12818;
												assign node12818 = (inp[8]) ? node12830 : node12819;
													assign node12819 = (inp[12]) ? node12827 : node12820;
														assign node12820 = (inp[10]) ? 4'b0111 : node12821;
															assign node12821 = (inp[9]) ? node12823 : 4'b0011;
																assign node12823 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node12827 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node12830 = (inp[12]) ? node12838 : node12831;
														assign node12831 = (inp[4]) ? node12835 : node12832;
															assign node12832 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node12835 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node12838 = (inp[9]) ? 4'b0110 : node12839;
															assign node12839 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node12843 = (inp[8]) ? node12851 : node12844;
													assign node12844 = (inp[4]) ? 4'b0110 : node12845;
														assign node12845 = (inp[9]) ? 4'b0010 : node12846;
															assign node12846 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node12851 = (inp[4]) ? node12857 : node12852;
														assign node12852 = (inp[9]) ? 4'b0011 : node12853;
															assign node12853 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node12857 = (inp[9]) ? node12859 : 4'b0011;
															assign node12859 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node12862 = (inp[4]) ? node12892 : node12863;
												assign node12863 = (inp[9]) ? node12877 : node12864;
													assign node12864 = (inp[10]) ? node12870 : node12865;
														assign node12865 = (inp[8]) ? 4'b0110 : node12866;
															assign node12866 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node12870 = (inp[12]) ? node12872 : 4'b0110;
															assign node12872 = (inp[2]) ? node12874 : 4'b0011;
																assign node12874 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node12877 = (inp[12]) ? node12883 : node12878;
														assign node12878 = (inp[10]) ? 4'b0010 : node12879;
															assign node12879 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node12883 = (inp[10]) ? node12887 : node12884;
															assign node12884 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node12887 = (inp[8]) ? node12889 : 4'b0101;
																assign node12889 = (inp[2]) ? 4'b0101 : 4'b0100;
												assign node12892 = (inp[9]) ? node12904 : node12893;
													assign node12893 = (inp[12]) ? node12895 : 4'b0011;
														assign node12895 = (inp[10]) ? node12897 : 4'b0011;
															assign node12897 = (inp[2]) ? node12901 : node12898;
																assign node12898 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node12901 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node12904 = (inp[12]) ? node12910 : node12905;
														assign node12905 = (inp[8]) ? node12907 : 4'b0100;
															assign node12907 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node12910 = (inp[8]) ? node12914 : node12911;
															assign node12911 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node12914 = (inp[2]) ? 4'b0101 : 4'b0100;
								assign node12917 = (inp[3]) ? node13137 : node12918;
									assign node12918 = (inp[10]) ? node13012 : node12919;
										assign node12919 = (inp[12]) ? node12963 : node12920;
											assign node12920 = (inp[4]) ? node12944 : node12921;
												assign node12921 = (inp[9]) ? node12937 : node12922;
													assign node12922 = (inp[15]) ? node12934 : node12923;
														assign node12923 = (inp[0]) ? node12929 : node12924;
															assign node12924 = (inp[8]) ? node12926 : 4'b0111;
																assign node12926 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node12929 = (inp[8]) ? 4'b0100 : node12930;
																assign node12930 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node12934 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node12937 = (inp[2]) ? 4'b0001 : node12938;
														assign node12938 = (inp[0]) ? node12940 : 4'b0011;
															assign node12940 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node12944 = (inp[9]) ? node12950 : node12945;
													assign node12945 = (inp[8]) ? 4'b0001 : node12946;
														assign node12946 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node12950 = (inp[2]) ? node12958 : node12951;
														assign node12951 = (inp[8]) ? node12953 : 4'b0101;
															assign node12953 = (inp[15]) ? node12955 : 4'b0100;
																assign node12955 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node12958 = (inp[15]) ? node12960 : 4'b0101;
															assign node12960 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node12963 = (inp[15]) ? node12989 : node12964;
												assign node12964 = (inp[0]) ? node12976 : node12965;
													assign node12965 = (inp[4]) ? node12973 : node12966;
														assign node12966 = (inp[9]) ? node12968 : 4'b0110;
															assign node12968 = (inp[8]) ? 4'b0011 : node12969;
																assign node12969 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node12973 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node12976 = (inp[2]) ? node12980 : node12977;
														assign node12977 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node12980 = (inp[8]) ? node12982 : 4'b0110;
															assign node12982 = (inp[4]) ? node12986 : node12983;
																assign node12983 = (inp[9]) ? 4'b0001 : 4'b0101;
																assign node12986 = (inp[9]) ? 4'b0111 : 4'b0001;
												assign node12989 = (inp[8]) ? node12997 : node12990;
													assign node12990 = (inp[2]) ? 4'b0000 : node12991;
														assign node12991 = (inp[9]) ? 4'b0101 : node12992;
															assign node12992 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node12997 = (inp[2]) ? node13005 : node12998;
														assign node12998 = (inp[9]) ? node13002 : node12999;
															assign node12999 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node13002 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node13005 = (inp[0]) ? node13007 : 4'b0101;
															assign node13007 = (inp[4]) ? node13009 : 4'b0011;
																assign node13009 = (inp[9]) ? 4'b0101 : 4'b0011;
										assign node13012 = (inp[9]) ? node13076 : node13013;
											assign node13013 = (inp[15]) ? node13041 : node13014;
												assign node13014 = (inp[0]) ? node13026 : node13015;
													assign node13015 = (inp[4]) ? node13017 : 4'b0011;
														assign node13017 = (inp[12]) ? node13019 : 4'b0011;
															assign node13019 = (inp[2]) ? node13023 : node13020;
																assign node13020 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node13023 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node13026 = (inp[4]) ? node13036 : node13027;
														assign node13027 = (inp[12]) ? node13033 : node13028;
															assign node13028 = (inp[2]) ? node13030 : 4'b0101;
																assign node13030 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node13033 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node13036 = (inp[12]) ? 4'b0111 : node13037;
															assign node13037 = (inp[2]) ? 4'b0000 : 4'b0001;
												assign node13041 = (inp[0]) ? node13059 : node13042;
													assign node13042 = (inp[8]) ? node13050 : node13043;
														assign node13043 = (inp[2]) ? 4'b0000 : node13044;
															assign node13044 = (inp[4]) ? 4'b0001 : node13045;
																assign node13045 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node13050 = (inp[2]) ? 4'b0001 : node13051;
															assign node13051 = (inp[4]) ? node13055 : node13052;
																assign node13052 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node13055 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node13059 = (inp[4]) ? node13067 : node13060;
														assign node13060 = (inp[12]) ? node13062 : 4'b0111;
															assign node13062 = (inp[2]) ? 4'b0010 : node13063;
																assign node13063 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node13067 = (inp[12]) ? node13071 : node13068;
															assign node13068 = (inp[8]) ? 4'b0011 : 4'b0010;
															assign node13071 = (inp[2]) ? node13073 : 4'b0101;
																assign node13073 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node13076 = (inp[8]) ? node13106 : node13077;
												assign node13077 = (inp[2]) ? node13085 : node13078;
													assign node13078 = (inp[12]) ? node13082 : node13079;
														assign node13079 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node13082 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node13085 = (inp[12]) ? node13099 : node13086;
														assign node13086 = (inp[4]) ? node13092 : node13087;
															assign node13087 = (inp[0]) ? node13089 : 4'b0010;
																assign node13089 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node13092 = (inp[0]) ? node13096 : node13093;
																assign node13093 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node13096 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node13099 = (inp[4]) ? 4'b0000 : node13100;
															assign node13100 = (inp[15]) ? 4'b0100 : node13101;
																assign node13101 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node13106 = (inp[2]) ? node13124 : node13107;
													assign node13107 = (inp[0]) ? node13113 : node13108;
														assign node13108 = (inp[12]) ? node13110 : 4'b0110;
															assign node13110 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node13113 = (inp[12]) ? node13117 : node13114;
															assign node13114 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node13117 = (inp[15]) ? node13121 : node13118;
																assign node13118 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node13121 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node13124 = (inp[12]) ? node13132 : node13125;
														assign node13125 = (inp[4]) ? 4'b0111 : node13126;
															assign node13126 = (inp[0]) ? 4'b0001 : node13127;
																assign node13127 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node13132 = (inp[15]) ? 4'b0001 : node13133;
															assign node13133 = (inp[0]) ? 4'b0111 : 4'b0101;
									assign node13137 = (inp[4]) ? node13243 : node13138;
										assign node13138 = (inp[9]) ? node13196 : node13139;
											assign node13139 = (inp[12]) ? node13171 : node13140;
												assign node13140 = (inp[10]) ? node13158 : node13141;
													assign node13141 = (inp[8]) ? node13155 : node13142;
														assign node13142 = (inp[2]) ? node13150 : node13143;
															assign node13143 = (inp[15]) ? node13147 : node13144;
																assign node13144 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node13147 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node13150 = (inp[0]) ? 4'b0100 : node13151;
																assign node13151 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node13155 = (inp[2]) ? 4'b0101 : 4'b0100;
													assign node13158 = (inp[0]) ? node13168 : node13159;
														assign node13159 = (inp[15]) ? node13163 : node13160;
															assign node13160 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node13163 = (inp[8]) ? node13165 : 4'b0111;
																assign node13165 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node13168 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node13171 = (inp[10]) ? node13183 : node13172;
													assign node13172 = (inp[15]) ? node13176 : node13173;
														assign node13173 = (inp[0]) ? 4'b0110 : 4'b0101;
														assign node13176 = (inp[0]) ? 4'b0101 : node13177;
															assign node13177 = (inp[8]) ? 4'b0111 : node13178;
																assign node13178 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node13183 = (inp[15]) ? node13187 : node13184;
														assign node13184 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node13187 = (inp[0]) ? node13189 : 4'b0010;
															assign node13189 = (inp[2]) ? node13193 : node13190;
																assign node13190 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node13193 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node13196 = (inp[10]) ? node13216 : node13197;
												assign node13197 = (inp[15]) ? node13209 : node13198;
													assign node13198 = (inp[0]) ? node13204 : node13199;
														assign node13199 = (inp[12]) ? node13201 : 4'b0000;
															assign node13201 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node13204 = (inp[8]) ? 4'b0011 : node13205;
															assign node13205 = (inp[12]) ? 4'b0011 : 4'b0010;
													assign node13209 = (inp[0]) ? 4'b0001 : node13210;
														assign node13210 = (inp[12]) ? node13212 : 4'b0011;
															assign node13212 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node13216 = (inp[12]) ? node13226 : node13217;
													assign node13217 = (inp[15]) ? node13221 : node13218;
														assign node13218 = (inp[0]) ? 4'b0010 : 4'b0001;
														assign node13221 = (inp[0]) ? 4'b0001 : node13222;
															assign node13222 = (inp[2]) ? 4'b0011 : 4'b0010;
													assign node13226 = (inp[15]) ? node13236 : node13227;
														assign node13227 = (inp[0]) ? node13233 : node13228;
															assign node13228 = (inp[8]) ? 4'b0101 : node13229;
																assign node13229 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node13233 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node13236 = (inp[8]) ? node13240 : node13237;
															assign node13237 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node13240 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node13243 = (inp[9]) ? node13297 : node13244;
											assign node13244 = (inp[10]) ? node13276 : node13245;
												assign node13245 = (inp[12]) ? node13261 : node13246;
													assign node13246 = (inp[0]) ? node13254 : node13247;
														assign node13247 = (inp[2]) ? node13251 : node13248;
															assign node13248 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node13251 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node13254 = (inp[15]) ? 4'b0000 : node13255;
															assign node13255 = (inp[2]) ? 4'b0010 : node13256;
																assign node13256 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node13261 = (inp[15]) ? node13271 : node13262;
														assign node13262 = (inp[0]) ? node13266 : node13263;
															assign node13263 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node13266 = (inp[2]) ? 4'b0010 : node13267;
																assign node13267 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node13271 = (inp[8]) ? node13273 : 4'b0001;
															assign node13273 = (inp[2]) ? 4'b0011 : 4'b0010;
												assign node13276 = (inp[12]) ? node13286 : node13277;
													assign node13277 = (inp[15]) ? node13279 : 4'b0011;
														assign node13279 = (inp[0]) ? 4'b0000 : node13280;
															assign node13280 = (inp[2]) ? node13282 : 4'b0010;
																assign node13282 = (inp[8]) ? 4'b0011 : 4'b0010;
													assign node13286 = (inp[2]) ? node13288 : 4'b0110;
														assign node13288 = (inp[8]) ? node13294 : node13289;
															assign node13289 = (inp[15]) ? node13291 : 4'b0110;
																assign node13291 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node13294 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node13297 = (inp[12]) ? node13333 : node13298;
												assign node13298 = (inp[10]) ? node13320 : node13299;
													assign node13299 = (inp[15]) ? node13309 : node13300;
														assign node13300 = (inp[0]) ? node13302 : 4'b0100;
															assign node13302 = (inp[8]) ? node13306 : node13303;
																assign node13303 = (inp[2]) ? 4'b0110 : 4'b0111;
																assign node13306 = (inp[2]) ? 4'b0111 : 4'b0110;
														assign node13309 = (inp[0]) ? node13315 : node13310;
															assign node13310 = (inp[2]) ? 4'b0111 : node13311;
																assign node13311 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node13315 = (inp[2]) ? 4'b0100 : node13316;
																assign node13316 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node13320 = (inp[0]) ? node13328 : node13321;
														assign node13321 = (inp[15]) ? node13323 : 4'b0101;
															assign node13323 = (inp[2]) ? 4'b0111 : node13324;
																assign node13324 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node13328 = (inp[15]) ? 4'b0101 : node13329;
															assign node13329 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node13333 = (inp[10]) ? node13347 : node13334;
													assign node13334 = (inp[2]) ? node13338 : node13335;
														assign node13335 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node13338 = (inp[8]) ? node13342 : node13339;
															assign node13339 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node13342 = (inp[0]) ? node13344 : 4'b0111;
																assign node13344 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node13347 = (inp[15]) ? node13361 : node13348;
														assign node13348 = (inp[0]) ? node13354 : node13349;
															assign node13349 = (inp[2]) ? node13351 : 4'b0001;
																assign node13351 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node13354 = (inp[2]) ? node13358 : node13355;
																assign node13355 = (inp[8]) ? 4'b0010 : 4'b0011;
																assign node13358 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node13361 = (inp[0]) ? node13363 : 4'b0011;
															assign node13363 = (inp[2]) ? node13367 : node13364;
																assign node13364 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node13367 = (inp[8]) ? 4'b0001 : 4'b0000;
							assign node13370 = (inp[15]) ? node13772 : node13371;
								assign node13371 = (inp[0]) ? node13563 : node13372;
									assign node13372 = (inp[3]) ? node13470 : node13373;
										assign node13373 = (inp[5]) ? node13421 : node13374;
											assign node13374 = (inp[8]) ? node13400 : node13375;
												assign node13375 = (inp[2]) ? node13387 : node13376;
													assign node13376 = (inp[9]) ? 4'b0010 : node13377;
														assign node13377 = (inp[10]) ? node13381 : node13378;
															assign node13378 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node13381 = (inp[12]) ? node13383 : 4'b0110;
																assign node13383 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node13387 = (inp[10]) ? node13393 : node13388;
														assign node13388 = (inp[12]) ? node13390 : 4'b0011;
															assign node13390 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node13393 = (inp[4]) ? node13395 : 4'b0111;
															assign node13395 = (inp[12]) ? 4'b0111 : node13396;
																assign node13396 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node13400 = (inp[2]) ? node13408 : node13401;
													assign node13401 = (inp[12]) ? node13403 : 4'b0111;
														assign node13403 = (inp[9]) ? 4'b0011 : node13404;
															assign node13404 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node13408 = (inp[12]) ? 4'b0110 : node13409;
														assign node13409 = (inp[10]) ? node13415 : node13410;
															assign node13410 = (inp[9]) ? node13412 : 4'b0110;
																assign node13412 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node13415 = (inp[9]) ? node13417 : 4'b0010;
																assign node13417 = (inp[4]) ? 4'b0110 : 4'b0010;
											assign node13421 = (inp[10]) ? node13445 : node13422;
												assign node13422 = (inp[4]) ? node13436 : node13423;
													assign node13423 = (inp[9]) ? node13429 : node13424;
														assign node13424 = (inp[8]) ? node13426 : 4'b0110;
															assign node13426 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node13429 = (inp[12]) ? 4'b0010 : node13430;
															assign node13430 = (inp[2]) ? node13432 : 4'b0011;
																assign node13432 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node13436 = (inp[9]) ? 4'b0101 : node13437;
														assign node13437 = (inp[12]) ? node13439 : 4'b0010;
															assign node13439 = (inp[2]) ? node13441 : 4'b0011;
																assign node13441 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node13445 = (inp[12]) ? node13457 : node13446;
													assign node13446 = (inp[9]) ? node13454 : node13447;
														assign node13447 = (inp[4]) ? node13451 : node13448;
															assign node13448 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node13451 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node13454 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node13457 = (inp[2]) ? node13465 : node13458;
														assign node13458 = (inp[8]) ? node13460 : 4'b0100;
															assign node13460 = (inp[9]) ? node13462 : 4'b0101;
																assign node13462 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node13465 = (inp[8]) ? node13467 : 4'b0011;
															assign node13467 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node13470 = (inp[5]) ? node13520 : node13471;
											assign node13471 = (inp[4]) ? node13491 : node13472;
												assign node13472 = (inp[9]) ? node13482 : node13473;
													assign node13473 = (inp[10]) ? node13477 : node13474;
														assign node13474 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node13477 = (inp[12]) ? 4'b0010 : node13478;
															assign node13478 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node13482 = (inp[12]) ? 4'b0101 : node13483;
														assign node13483 = (inp[10]) ? 4'b0010 : node13484;
															assign node13484 = (inp[2]) ? node13486 : 4'b0010;
																assign node13486 = (inp[8]) ? 4'b0010 : 4'b0011;
												assign node13491 = (inp[9]) ? node13507 : node13492;
													assign node13492 = (inp[10]) ? node13498 : node13493;
														assign node13493 = (inp[8]) ? 4'b0010 : node13494;
															assign node13494 = (inp[2]) ? 4'b0011 : 4'b0010;
														assign node13498 = (inp[12]) ? node13502 : node13499;
															assign node13499 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node13502 = (inp[2]) ? 4'b0100 : node13503;
																assign node13503 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node13507 = (inp[12]) ? node13515 : node13508;
														assign node13508 = (inp[2]) ? node13512 : node13509;
															assign node13509 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node13512 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node13515 = (inp[10]) ? node13517 : 4'b0100;
															assign node13517 = (inp[2]) ? 4'b0001 : 4'b0000;
											assign node13520 = (inp[9]) ? node13538 : node13521;
												assign node13521 = (inp[4]) ? node13529 : node13522;
													assign node13522 = (inp[8]) ? node13526 : node13523;
														assign node13523 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node13526 = (inp[2]) ? 4'b0100 : 4'b0101;
													assign node13529 = (inp[10]) ? node13531 : 4'b0001;
														assign node13531 = (inp[2]) ? node13535 : node13532;
															assign node13532 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node13535 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node13538 = (inp[4]) ? node13550 : node13539;
													assign node13539 = (inp[12]) ? node13547 : node13540;
														assign node13540 = (inp[10]) ? node13542 : 4'b0001;
															assign node13542 = (inp[8]) ? 4'b0000 : node13543;
																assign node13543 = (inp[2]) ? 4'b0001 : 4'b0000;
														assign node13547 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node13550 = (inp[12]) ? node13556 : node13551;
														assign node13551 = (inp[2]) ? node13553 : 4'b0100;
															assign node13553 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node13556 = (inp[10]) ? 4'b0000 : node13557;
															assign node13557 = (inp[2]) ? 4'b0100 : node13558;
																assign node13558 = (inp[8]) ? 4'b0101 : 4'b0100;
									assign node13563 = (inp[3]) ? node13675 : node13564;
										assign node13564 = (inp[5]) ? node13616 : node13565;
											assign node13565 = (inp[8]) ? node13595 : node13566;
												assign node13566 = (inp[2]) ? node13582 : node13567;
													assign node13567 = (inp[9]) ? node13573 : node13568;
														assign node13568 = (inp[10]) ? node13570 : 4'b0100;
															assign node13570 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node13573 = (inp[4]) ? node13579 : node13574;
															assign node13574 = (inp[12]) ? node13576 : 4'b0000;
																assign node13576 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node13579 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node13582 = (inp[4]) ? node13588 : node13583;
														assign node13583 = (inp[9]) ? node13585 : 4'b0101;
															assign node13585 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node13588 = (inp[12]) ? node13590 : 4'b0001;
															assign node13590 = (inp[10]) ? node13592 : 4'b0101;
																assign node13592 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node13595 = (inp[2]) ? node13599 : node13596;
													assign node13596 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node13599 = (inp[4]) ? node13611 : node13600;
														assign node13600 = (inp[9]) ? node13606 : node13601;
															assign node13601 = (inp[10]) ? node13603 : 4'b0100;
																assign node13603 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node13606 = (inp[10]) ? node13608 : 4'b0000;
																assign node13608 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node13611 = (inp[9]) ? node13613 : 4'b0000;
															assign node13613 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node13616 = (inp[9]) ? node13650 : node13617;
												assign node13617 = (inp[4]) ? node13639 : node13618;
													assign node13618 = (inp[10]) ? node13632 : node13619;
														assign node13619 = (inp[12]) ? node13627 : node13620;
															assign node13620 = (inp[8]) ? node13624 : node13621;
																assign node13621 = (inp[2]) ? 4'b0101 : 4'b0100;
																assign node13624 = (inp[2]) ? 4'b0100 : 4'b0101;
															assign node13627 = (inp[8]) ? node13629 : 4'b0100;
																assign node13629 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node13632 = (inp[12]) ? node13634 : 4'b0100;
															assign node13634 = (inp[8]) ? node13636 : 4'b0000;
																assign node13636 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node13639 = (inp[10]) ? node13645 : node13640;
														assign node13640 = (inp[8]) ? node13642 : 4'b0001;
															assign node13642 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node13645 = (inp[12]) ? node13647 : 4'b0000;
															assign node13647 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node13650 = (inp[4]) ? node13660 : node13651;
													assign node13651 = (inp[2]) ? node13655 : node13652;
														assign node13652 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node13655 = (inp[10]) ? node13657 : 4'b0001;
															assign node13657 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node13660 = (inp[12]) ? node13668 : node13661;
														assign node13661 = (inp[8]) ? node13665 : node13662;
															assign node13662 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node13665 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node13668 = (inp[10]) ? 4'b0011 : node13669;
															assign node13669 = (inp[2]) ? 4'b0111 : node13670;
																assign node13670 = (inp[8]) ? 4'b0111 : 4'b0110;
										assign node13675 = (inp[5]) ? node13735 : node13676;
											assign node13676 = (inp[4]) ? node13700 : node13677;
												assign node13677 = (inp[9]) ? node13687 : node13678;
													assign node13678 = (inp[2]) ? node13684 : node13679;
														assign node13679 = (inp[8]) ? 4'b0101 : node13680;
															assign node13680 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node13684 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node13687 = (inp[12]) ? node13695 : node13688;
														assign node13688 = (inp[8]) ? node13692 : node13689;
															assign node13689 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node13692 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node13695 = (inp[10]) ? node13697 : 4'b0000;
															assign node13697 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node13700 = (inp[9]) ? node13718 : node13701;
													assign node13701 = (inp[12]) ? node13709 : node13702;
														assign node13702 = (inp[8]) ? node13706 : node13703;
															assign node13703 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node13706 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node13709 = (inp[10]) ? node13713 : node13710;
															assign node13710 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node13713 = (inp[2]) ? node13715 : 4'b0110;
																assign node13715 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node13718 = (inp[12]) ? node13724 : node13719;
														assign node13719 = (inp[8]) ? 4'b0111 : node13720;
															assign node13720 = (inp[10]) ? 4'b0111 : 4'b0110;
														assign node13724 = (inp[10]) ? node13730 : node13725;
															assign node13725 = (inp[8]) ? 4'b0110 : node13726;
																assign node13726 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node13730 = (inp[2]) ? node13732 : 4'b0010;
																assign node13732 = (inp[8]) ? 4'b0010 : 4'b0011;
											assign node13735 = (inp[8]) ? node13751 : node13736;
												assign node13736 = (inp[2]) ? node13746 : node13737;
													assign node13737 = (inp[9]) ? node13739 : 4'b0010;
														assign node13739 = (inp[4]) ? 4'b0110 : node13740;
															assign node13740 = (inp[10]) ? node13742 : 4'b0010;
																assign node13742 = (inp[12]) ? 4'b0110 : 4'b0010;
													assign node13746 = (inp[4]) ? 4'b0111 : node13747;
														assign node13747 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node13751 = (inp[2]) ? node13761 : node13752;
													assign node13752 = (inp[9]) ? node13758 : node13753;
														assign node13753 = (inp[4]) ? node13755 : 4'b0111;
															assign node13755 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node13758 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node13761 = (inp[10]) ? node13763 : 4'b0010;
														assign node13763 = (inp[4]) ? 4'b0010 : node13764;
															assign node13764 = (inp[12]) ? node13768 : node13765;
																assign node13765 = (inp[9]) ? 4'b0010 : 4'b0110;
																assign node13768 = (inp[9]) ? 4'b0110 : 4'b0010;
								assign node13772 = (inp[0]) ? node13994 : node13773;
									assign node13773 = (inp[5]) ? node13875 : node13774;
										assign node13774 = (inp[3]) ? node13818 : node13775;
											assign node13775 = (inp[10]) ? node13793 : node13776;
												assign node13776 = (inp[8]) ? node13780 : node13777;
													assign node13777 = (inp[2]) ? 4'b0101 : 4'b0000;
													assign node13780 = (inp[2]) ? node13786 : node13781;
														assign node13781 = (inp[4]) ? 4'b0101 : node13782;
															assign node13782 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node13786 = (inp[12]) ? 4'b0100 : node13787;
															assign node13787 = (inp[9]) ? 4'b0100 : node13788;
																assign node13788 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node13793 = (inp[12]) ? node13805 : node13794;
													assign node13794 = (inp[8]) ? node13802 : node13795;
														assign node13795 = (inp[2]) ? node13797 : 4'b0100;
															assign node13797 = (inp[4]) ? node13799 : 4'b0101;
																assign node13799 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node13802 = (inp[2]) ? 4'b0100 : 4'b0001;
													assign node13805 = (inp[4]) ? node13811 : node13806;
														assign node13806 = (inp[9]) ? node13808 : 4'b0001;
															assign node13808 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node13811 = (inp[9]) ? 4'b0001 : node13812;
															assign node13812 = (inp[2]) ? node13814 : 4'b0101;
																assign node13814 = (inp[8]) ? 4'b0100 : 4'b0101;
											assign node13818 = (inp[4]) ? node13856 : node13819;
												assign node13819 = (inp[9]) ? node13835 : node13820;
													assign node13820 = (inp[10]) ? node13826 : node13821;
														assign node13821 = (inp[8]) ? 4'b0101 : node13822;
															assign node13822 = (inp[2]) ? 4'b0101 : 4'b0100;
														assign node13826 = (inp[12]) ? node13830 : node13827;
															assign node13827 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node13830 = (inp[2]) ? 4'b0000 : node13831;
																assign node13831 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node13835 = (inp[10]) ? node13845 : node13836;
														assign node13836 = (inp[12]) ? node13838 : 4'b0001;
															assign node13838 = (inp[8]) ? node13842 : node13839;
																assign node13839 = (inp[2]) ? 4'b0001 : 4'b0000;
																assign node13842 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node13845 = (inp[12]) ? node13851 : node13846;
															assign node13846 = (inp[8]) ? 4'b0001 : node13847;
																assign node13847 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node13851 = (inp[8]) ? node13853 : 4'b0110;
																assign node13853 = (inp[2]) ? 4'b0110 : 4'b0111;
												assign node13856 = (inp[9]) ? node13870 : node13857;
													assign node13857 = (inp[12]) ? node13865 : node13858;
														assign node13858 = (inp[8]) ? node13862 : node13859;
															assign node13859 = (inp[2]) ? 4'b0001 : 4'b0000;
															assign node13862 = (inp[10]) ? 4'b0000 : 4'b0001;
														assign node13865 = (inp[10]) ? 4'b0111 : node13866;
															assign node13866 = (inp[2]) ? 4'b0000 : 4'b0001;
													assign node13870 = (inp[8]) ? 4'b0110 : node13871;
														assign node13871 = (inp[2]) ? 4'b0111 : 4'b0110;
										assign node13875 = (inp[3]) ? node13935 : node13876;
											assign node13876 = (inp[4]) ? node13904 : node13877;
												assign node13877 = (inp[9]) ? node13889 : node13878;
													assign node13878 = (inp[10]) ? node13886 : node13879;
														assign node13879 = (inp[8]) ? node13883 : node13880;
															assign node13880 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node13883 = (inp[2]) ? 4'b0100 : 4'b0101;
														assign node13886 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node13889 = (inp[12]) ? node13897 : node13890;
														assign node13890 = (inp[2]) ? node13894 : node13891;
															assign node13891 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node13894 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node13897 = (inp[10]) ? node13901 : node13898;
															assign node13898 = (inp[2]) ? 4'b0000 : 4'b0001;
															assign node13901 = (inp[8]) ? 4'b0110 : 4'b0111;
												assign node13904 = (inp[9]) ? node13918 : node13905;
													assign node13905 = (inp[12]) ? node13911 : node13906;
														assign node13906 = (inp[8]) ? node13908 : 4'b0000;
															assign node13908 = (inp[2]) ? 4'b0000 : 4'b0001;
														assign node13911 = (inp[10]) ? node13913 : 4'b0001;
															assign node13913 = (inp[2]) ? node13915 : 4'b0110;
																assign node13915 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node13918 = (inp[10]) ? node13932 : node13919;
														assign node13919 = (inp[12]) ? node13927 : node13920;
															assign node13920 = (inp[8]) ? node13924 : node13921;
																assign node13921 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node13924 = (inp[2]) ? 4'b0110 : 4'b0111;
															assign node13927 = (inp[2]) ? node13929 : 4'b0110;
																assign node13929 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node13932 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node13935 = (inp[12]) ? node13963 : node13936;
												assign node13936 = (inp[10]) ? node13946 : node13937;
													assign node13937 = (inp[9]) ? node13943 : node13938;
														assign node13938 = (inp[4]) ? 4'b0010 : node13939;
															assign node13939 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node13943 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node13946 = (inp[8]) ? node13952 : node13947;
														assign node13947 = (inp[2]) ? node13949 : 4'b0110;
															assign node13949 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node13952 = (inp[2]) ? node13960 : node13953;
															assign node13953 = (inp[9]) ? node13957 : node13954;
																assign node13954 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node13957 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node13960 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node13963 = (inp[9]) ? node13983 : node13964;
													assign node13964 = (inp[8]) ? node13976 : node13965;
														assign node13965 = (inp[2]) ? node13973 : node13966;
															assign node13966 = (inp[10]) ? node13970 : node13967;
																assign node13967 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node13970 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node13973 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node13976 = (inp[2]) ? node13978 : 4'b0011;
															assign node13978 = (inp[4]) ? node13980 : 4'b0010;
																assign node13980 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node13983 = (inp[2]) ? node13987 : node13984;
														assign node13984 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node13987 = (inp[8]) ? 4'b0010 : node13988;
															assign node13988 = (inp[4]) ? node13990 : 4'b0111;
																assign node13990 = (inp[10]) ? 4'b0011 : 4'b0111;
									assign node13994 = (inp[3]) ? node14122 : node13995;
										assign node13995 = (inp[5]) ? node14063 : node13996;
											assign node13996 = (inp[4]) ? node14028 : node13997;
												assign node13997 = (inp[9]) ? node14009 : node13998;
													assign node13998 = (inp[10]) ? node14000 : 4'b0110;
														assign node14000 = (inp[12]) ? 4'b0011 : node14001;
															assign node14001 = (inp[8]) ? node14005 : node14002;
																assign node14002 = (inp[2]) ? 4'b0111 : 4'b0110;
																assign node14005 = (inp[2]) ? 4'b0110 : 4'b0111;
													assign node14009 = (inp[10]) ? node14021 : node14010;
														assign node14010 = (inp[12]) ? node14016 : node14011;
															assign node14011 = (inp[2]) ? node14013 : 4'b0011;
																assign node14013 = (inp[8]) ? 4'b0010 : 4'b0011;
															assign node14016 = (inp[2]) ? node14018 : 4'b0010;
																assign node14018 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node14021 = (inp[12]) ? node14023 : 4'b0010;
															assign node14023 = (inp[8]) ? 4'b0110 : node14024;
																assign node14024 = (inp[2]) ? 4'b0111 : 4'b0110;
												assign node14028 = (inp[9]) ? node14046 : node14029;
													assign node14029 = (inp[10]) ? node14035 : node14030;
														assign node14030 = (inp[8]) ? node14032 : 4'b0011;
															assign node14032 = (inp[2]) ? 4'b0010 : 4'b0011;
														assign node14035 = (inp[12]) ? node14041 : node14036;
															assign node14036 = (inp[8]) ? node14038 : 4'b0011;
																assign node14038 = (inp[2]) ? 4'b0010 : 4'b0011;
															assign node14041 = (inp[2]) ? 4'b0111 : node14042;
																assign node14042 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node14046 = (inp[12]) ? node14054 : node14047;
														assign node14047 = (inp[10]) ? node14049 : 4'b0111;
															assign node14049 = (inp[8]) ? node14051 : 4'b0110;
																assign node14051 = (inp[2]) ? 4'b0110 : 4'b0111;
														assign node14054 = (inp[10]) ? node14060 : node14055;
															assign node14055 = (inp[8]) ? 4'b0110 : node14056;
																assign node14056 = (inp[2]) ? 4'b0111 : 4'b0110;
															assign node14060 = (inp[2]) ? 4'b0010 : 4'b0011;
											assign node14063 = (inp[9]) ? node14095 : node14064;
												assign node14064 = (inp[4]) ? node14076 : node14065;
													assign node14065 = (inp[10]) ? node14073 : node14066;
														assign node14066 = (inp[2]) ? node14070 : node14067;
															assign node14067 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node14070 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node14073 = (inp[8]) ? 4'b0110 : 4'b0010;
													assign node14076 = (inp[12]) ? node14086 : node14077;
														assign node14077 = (inp[10]) ? node14079 : 4'b0010;
															assign node14079 = (inp[2]) ? node14083 : node14080;
																assign node14080 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node14083 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node14086 = (inp[10]) ? node14092 : node14087;
															assign node14087 = (inp[8]) ? 4'b0011 : node14088;
																assign node14088 = (inp[2]) ? 4'b0011 : 4'b0010;
															assign node14092 = (inp[8]) ? 4'b0100 : 4'b0101;
												assign node14095 = (inp[4]) ? node14105 : node14096;
													assign node14096 = (inp[12]) ? node14102 : node14097;
														assign node14097 = (inp[2]) ? 4'b0011 : node14098;
															assign node14098 = (inp[8]) ? 4'b0011 : 4'b0010;
														assign node14102 = (inp[10]) ? 4'b0100 : 4'b0010;
													assign node14105 = (inp[10]) ? node14113 : node14106;
														assign node14106 = (inp[2]) ? node14110 : node14107;
															assign node14107 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node14110 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node14113 = (inp[12]) ? node14117 : node14114;
															assign node14114 = (inp[2]) ? 4'b0101 : 4'b0100;
															assign node14117 = (inp[2]) ? node14119 : 4'b0001;
																assign node14119 = (inp[8]) ? 4'b0000 : 4'b0001;
										assign node14122 = (inp[5]) ? node14162 : node14123;
											assign node14123 = (inp[9]) ? node14147 : node14124;
												assign node14124 = (inp[10]) ? node14132 : node14125;
													assign node14125 = (inp[4]) ? node14127 : 4'b0111;
														assign node14127 = (inp[8]) ? node14129 : 4'b0011;
															assign node14129 = (inp[2]) ? 4'b0010 : 4'b0011;
													assign node14132 = (inp[2]) ? node14140 : node14133;
														assign node14133 = (inp[12]) ? node14137 : node14134;
															assign node14134 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node14137 = (inp[4]) ? 4'b0100 : 4'b0010;
														assign node14140 = (inp[8]) ? 4'b0010 : node14141;
															assign node14141 = (inp[4]) ? node14143 : 4'b0011;
																assign node14143 = (inp[12]) ? 4'b0101 : 4'b0011;
												assign node14147 = (inp[4]) ? node14153 : node14148;
													assign node14148 = (inp[10]) ? 4'b0100 : node14149;
														assign node14149 = (inp[12]) ? 4'b0010 : 4'b0011;
													assign node14153 = (inp[8]) ? node14155 : 4'b0100;
														assign node14155 = (inp[2]) ? 4'b0100 : node14156;
															assign node14156 = (inp[12]) ? node14158 : 4'b0101;
																assign node14158 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node14162 = (inp[10]) ? node14178 : node14163;
												assign node14163 = (inp[2]) ? node14171 : node14164;
													assign node14164 = (inp[8]) ? node14166 : 4'b0000;
														assign node14166 = (inp[9]) ? 4'b0001 : node14167;
															assign node14167 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node14171 = (inp[8]) ? 4'b0100 : node14172;
														assign node14172 = (inp[4]) ? node14174 : 4'b0001;
															assign node14174 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node14178 = (inp[8]) ? node14194 : node14179;
													assign node14179 = (inp[2]) ? node14181 : 4'b0100;
														assign node14181 = (inp[4]) ? node14189 : node14182;
															assign node14182 = (inp[9]) ? node14186 : node14183;
																assign node14183 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node14186 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node14189 = (inp[9]) ? node14191 : 4'b0101;
																assign node14191 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node14194 = (inp[2]) ? node14198 : node14195;
														assign node14195 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node14198 = (inp[4]) ? 4'b0000 : 4'b0100;
						assign node14201 = (inp[2]) ? node14947 : node14202;
							assign node14202 = (inp[8]) ? node14572 : node14203;
								assign node14203 = (inp[7]) ? node14387 : node14204;
									assign node14204 = (inp[5]) ? node14322 : node14205;
										assign node14205 = (inp[10]) ? node14249 : node14206;
											assign node14206 = (inp[15]) ? node14232 : node14207;
												assign node14207 = (inp[0]) ? node14215 : node14208;
													assign node14208 = (inp[3]) ? node14212 : node14209;
														assign node14209 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node14212 = (inp[4]) ? 4'b0101 : 4'b0111;
													assign node14215 = (inp[3]) ? node14227 : node14216;
														assign node14216 = (inp[12]) ? node14222 : node14217;
															assign node14217 = (inp[4]) ? node14219 : 4'b0101;
																assign node14219 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node14222 = (inp[9]) ? node14224 : 4'b0001;
																assign node14224 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node14227 = (inp[4]) ? 4'b0111 : node14228;
															assign node14228 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node14232 = (inp[0]) ? node14240 : node14233;
													assign node14233 = (inp[3]) ? node14235 : 4'b0101;
														assign node14235 = (inp[9]) ? 4'b0001 : node14236;
															assign node14236 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node14240 = (inp[9]) ? node14244 : node14241;
														assign node14241 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node14244 = (inp[4]) ? node14246 : 4'b0011;
															assign node14246 = (inp[12]) ? 4'b0101 : 4'b0111;
											assign node14249 = (inp[3]) ? node14287 : node14250;
												assign node14250 = (inp[12]) ? node14272 : node14251;
													assign node14251 = (inp[0]) ? node14265 : node14252;
														assign node14252 = (inp[15]) ? node14260 : node14253;
															assign node14253 = (inp[9]) ? node14257 : node14254;
																assign node14254 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node14257 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node14260 = (inp[4]) ? 4'b0001 : node14261;
																assign node14261 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node14265 = (inp[15]) ? node14267 : 4'b0101;
															assign node14267 = (inp[4]) ? node14269 : 4'b0111;
																assign node14269 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node14272 = (inp[4]) ? node14280 : node14273;
														assign node14273 = (inp[15]) ? node14277 : node14274;
															assign node14274 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node14277 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node14280 = (inp[9]) ? 4'b0001 : node14281;
															assign node14281 = (inp[15]) ? node14283 : 4'b0101;
																assign node14283 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node14287 = (inp[0]) ? node14303 : node14288;
													assign node14288 = (inp[9]) ? node14300 : node14289;
														assign node14289 = (inp[4]) ? node14297 : node14290;
															assign node14290 = (inp[15]) ? node14294 : node14291;
																assign node14291 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node14294 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node14297 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node14300 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node14303 = (inp[12]) ? node14315 : node14304;
														assign node14304 = (inp[15]) ? node14310 : node14305;
															assign node14305 = (inp[4]) ? 4'b0001 : node14306;
																assign node14306 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node14310 = (inp[4]) ? node14312 : 4'b0011;
																assign node14312 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node14315 = (inp[15]) ? 4'b0101 : node14316;
															assign node14316 = (inp[4]) ? node14318 : 4'b0111;
																assign node14318 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node14322 = (inp[4]) ? node14358 : node14323;
											assign node14323 = (inp[3]) ? node14339 : node14324;
												assign node14324 = (inp[12]) ? node14330 : node14325;
													assign node14325 = (inp[10]) ? node14327 : 4'b0011;
														assign node14327 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node14330 = (inp[9]) ? node14336 : node14331;
														assign node14331 = (inp[0]) ? 4'b0111 : node14332;
															assign node14332 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node14336 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node14339 = (inp[9]) ? node14351 : node14340;
													assign node14340 = (inp[10]) ? node14346 : node14341;
														assign node14341 = (inp[0]) ? 4'b0111 : node14342;
															assign node14342 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node14346 = (inp[12]) ? node14348 : 4'b0101;
															assign node14348 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node14351 = (inp[0]) ? node14353 : 4'b0111;
														assign node14353 = (inp[12]) ? node14355 : 4'b0001;
															assign node14355 = (inp[10]) ? 4'b0101 : 4'b0001;
											assign node14358 = (inp[9]) ? node14368 : node14359;
												assign node14359 = (inp[12]) ? node14365 : node14360;
													assign node14360 = (inp[15]) ? 4'b0011 : node14361;
														assign node14361 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node14365 = (inp[10]) ? 4'b0111 : 4'b0011;
												assign node14368 = (inp[10]) ? node14376 : node14369;
													assign node14369 = (inp[0]) ? node14373 : node14370;
														assign node14370 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node14373 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node14376 = (inp[12]) ? node14382 : node14377;
														assign node14377 = (inp[0]) ? 4'b0111 : node14378;
															assign node14378 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node14382 = (inp[3]) ? 4'b0011 : node14383;
															assign node14383 = (inp[0]) ? 4'b0011 : 4'b0001;
									assign node14387 = (inp[9]) ? node14479 : node14388;
										assign node14388 = (inp[4]) ? node14424 : node14389;
											assign node14389 = (inp[12]) ? node14409 : node14390;
												assign node14390 = (inp[10]) ? node14396 : node14391;
													assign node14391 = (inp[5]) ? node14393 : 4'b0100;
														assign node14393 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node14396 = (inp[0]) ? node14402 : node14397;
														assign node14397 = (inp[3]) ? 4'b0110 : node14398;
															assign node14398 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node14402 = (inp[15]) ? node14404 : 4'b0100;
															assign node14404 = (inp[3]) ? node14406 : 4'b0110;
																assign node14406 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node14409 = (inp[10]) ? node14417 : node14410;
													assign node14410 = (inp[5]) ? node14412 : 4'b0110;
														assign node14412 = (inp[3]) ? node14414 : 4'b0100;
															assign node14414 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node14417 = (inp[0]) ? 4'b0010 : node14418;
														assign node14418 = (inp[15]) ? 4'b0000 : node14419;
															assign node14419 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node14424 = (inp[10]) ? node14452 : node14425;
												assign node14425 = (inp[12]) ? node14437 : node14426;
													assign node14426 = (inp[5]) ? node14428 : 4'b0010;
														assign node14428 = (inp[3]) ? node14430 : 4'b0000;
															assign node14430 = (inp[0]) ? node14434 : node14431;
																assign node14431 = (inp[15]) ? 4'b0010 : 4'b0000;
																assign node14434 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node14437 = (inp[5]) ? node14443 : node14438;
														assign node14438 = (inp[0]) ? 4'b0000 : node14439;
															assign node14439 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node14443 = (inp[0]) ? node14445 : 4'b0010;
															assign node14445 = (inp[15]) ? node14449 : node14446;
																assign node14446 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node14449 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node14452 = (inp[12]) ? node14466 : node14453;
													assign node14453 = (inp[0]) ? node14459 : node14454;
														assign node14454 = (inp[15]) ? node14456 : 4'b0010;
															assign node14456 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node14459 = (inp[5]) ? node14461 : 4'b0000;
															assign node14461 = (inp[15]) ? 4'b0010 : node14462;
																assign node14462 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node14466 = (inp[15]) ? node14472 : node14467;
														assign node14467 = (inp[0]) ? 4'b0100 : node14468;
															assign node14468 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node14472 = (inp[5]) ? 4'b0110 : node14473;
															assign node14473 = (inp[3]) ? 4'b0110 : node14474;
																assign node14474 = (inp[0]) ? 4'b0110 : 4'b0100;
										assign node14479 = (inp[4]) ? node14527 : node14480;
											assign node14480 = (inp[10]) ? node14502 : node14481;
												assign node14481 = (inp[15]) ? node14491 : node14482;
													assign node14482 = (inp[0]) ? node14488 : node14483;
														assign node14483 = (inp[3]) ? node14485 : 4'b0010;
															assign node14485 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node14488 = (inp[12]) ? 4'b0010 : 4'b0000;
													assign node14491 = (inp[0]) ? node14497 : node14492;
														assign node14492 = (inp[5]) ? node14494 : 4'b0000;
															assign node14494 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node14497 = (inp[3]) ? node14499 : 4'b0010;
															assign node14499 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node14502 = (inp[12]) ? node14512 : node14503;
													assign node14503 = (inp[0]) ? node14509 : node14504;
														assign node14504 = (inp[15]) ? 4'b0000 : node14505;
															assign node14505 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node14509 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node14512 = (inp[0]) ? node14520 : node14513;
														assign node14513 = (inp[15]) ? 4'b0110 : node14514;
															assign node14514 = (inp[5]) ? 4'b0100 : node14515;
																assign node14515 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node14520 = (inp[15]) ? 4'b0100 : node14521;
															assign node14521 = (inp[3]) ? 4'b0110 : node14522;
																assign node14522 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node14527 = (inp[10]) ? node14541 : node14528;
												assign node14528 = (inp[0]) ? node14534 : node14529;
													assign node14529 = (inp[15]) ? 4'b0110 : node14530;
														assign node14530 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node14534 = (inp[15]) ? 4'b0100 : node14535;
														assign node14535 = (inp[3]) ? 4'b0110 : node14536;
															assign node14536 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node14541 = (inp[12]) ? node14559 : node14542;
													assign node14542 = (inp[0]) ? node14554 : node14543;
														assign node14543 = (inp[15]) ? node14549 : node14544;
															assign node14544 = (inp[5]) ? 4'b0100 : node14545;
																assign node14545 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node14549 = (inp[5]) ? 4'b0110 : node14550;
																assign node14550 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node14554 = (inp[15]) ? 4'b0100 : node14555;
															assign node14555 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node14559 = (inp[15]) ? node14567 : node14560;
														assign node14560 = (inp[5]) ? 4'b0000 : node14561;
															assign node14561 = (inp[0]) ? 4'b0000 : node14562;
																assign node14562 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node14567 = (inp[0]) ? node14569 : 4'b0010;
															assign node14569 = (inp[5]) ? 4'b0000 : 4'b0010;
								assign node14572 = (inp[7]) ? node14770 : node14573;
									assign node14573 = (inp[15]) ? node14661 : node14574;
										assign node14574 = (inp[0]) ? node14610 : node14575;
											assign node14575 = (inp[3]) ? node14591 : node14576;
												assign node14576 = (inp[9]) ? node14584 : node14577;
													assign node14577 = (inp[4]) ? node14579 : 4'b0110;
														assign node14579 = (inp[5]) ? 4'b0010 : node14580;
															assign node14580 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node14584 = (inp[10]) ? node14586 : 4'b0010;
														assign node14586 = (inp[5]) ? node14588 : 4'b0010;
															assign node14588 = (inp[12]) ? 4'b0000 : 4'b0100;
												assign node14591 = (inp[5]) ? node14599 : node14592;
													assign node14592 = (inp[10]) ? node14594 : 4'b0010;
														assign node14594 = (inp[12]) ? 4'b0100 : node14595;
															assign node14595 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node14599 = (inp[4]) ? 4'b0100 : node14600;
														assign node14600 = (inp[9]) ? node14604 : node14601;
															assign node14601 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node14604 = (inp[10]) ? node14606 : 4'b0000;
																assign node14606 = (inp[12]) ? 4'b0100 : 4'b0000;
											assign node14610 = (inp[3]) ? node14636 : node14611;
												assign node14611 = (inp[12]) ? node14617 : node14612;
													assign node14612 = (inp[4]) ? 4'b0000 : node14613;
														assign node14613 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node14617 = (inp[5]) ? node14627 : node14618;
														assign node14618 = (inp[10]) ? node14620 : 4'b0100;
															assign node14620 = (inp[9]) ? node14624 : node14621;
																assign node14621 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node14624 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node14627 = (inp[10]) ? node14633 : node14628;
															assign node14628 = (inp[9]) ? 4'b0000 : node14629;
																assign node14629 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node14633 = (inp[4]) ? 4'b0110 : 4'b0000;
												assign node14636 = (inp[5]) ? node14650 : node14637;
													assign node14637 = (inp[4]) ? node14645 : node14638;
														assign node14638 = (inp[9]) ? 4'b0000 : node14639;
															assign node14639 = (inp[12]) ? node14641 : 4'b0100;
																assign node14641 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node14645 = (inp[12]) ? 4'b0110 : node14646;
															assign node14646 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node14650 = (inp[12]) ? node14656 : node14651;
														assign node14651 = (inp[9]) ? node14653 : 4'b0110;
															assign node14653 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node14656 = (inp[4]) ? node14658 : 4'b0010;
															assign node14658 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node14661 = (inp[0]) ? node14717 : node14662;
											assign node14662 = (inp[5]) ? node14690 : node14663;
												assign node14663 = (inp[3]) ? node14681 : node14664;
													assign node14664 = (inp[12]) ? node14670 : node14665;
														assign node14665 = (inp[4]) ? node14667 : 4'b0000;
															assign node14667 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node14670 = (inp[10]) ? node14676 : node14671;
															assign node14671 = (inp[4]) ? 4'b0000 : node14672;
																assign node14672 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node14676 = (inp[9]) ? 4'b0100 : node14677;
																assign node14677 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node14681 = (inp[12]) ? node14687 : node14682;
														assign node14682 = (inp[10]) ? node14684 : 4'b0110;
															assign node14684 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node14687 = (inp[10]) ? 4'b0010 : 4'b0000;
												assign node14690 = (inp[3]) ? node14708 : node14691;
													assign node14691 = (inp[9]) ? node14701 : node14692;
														assign node14692 = (inp[12]) ? node14696 : node14693;
															assign node14693 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node14696 = (inp[4]) ? node14698 : 4'b0000;
																assign node14698 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node14701 = (inp[4]) ? node14703 : 4'b0000;
															assign node14703 = (inp[10]) ? node14705 : 4'b0110;
																assign node14705 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node14708 = (inp[12]) ? node14710 : 4'b0110;
														assign node14710 = (inp[9]) ? node14712 : 4'b0010;
															assign node14712 = (inp[4]) ? node14714 : 4'b0110;
																assign node14714 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node14717 = (inp[5]) ? node14743 : node14718;
												assign node14718 = (inp[3]) ? node14730 : node14719;
													assign node14719 = (inp[9]) ? node14727 : node14720;
														assign node14720 = (inp[4]) ? 4'b0010 : node14721;
															assign node14721 = (inp[10]) ? node14723 : 4'b0110;
																assign node14723 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node14727 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node14730 = (inp[4]) ? node14738 : node14731;
														assign node14731 = (inp[9]) ? 4'b0010 : node14732;
															assign node14732 = (inp[12]) ? node14734 : 4'b0110;
																assign node14734 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node14738 = (inp[12]) ? 4'b0100 : node14739;
															assign node14739 = (inp[9]) ? 4'b0100 : 4'b0010;
												assign node14743 = (inp[3]) ? node14755 : node14744;
													assign node14744 = (inp[4]) ? node14748 : node14745;
														assign node14745 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node14748 = (inp[9]) ? 4'b0100 : node14749;
															assign node14749 = (inp[10]) ? node14751 : 4'b0010;
																assign node14751 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node14755 = (inp[4]) ? node14759 : node14756;
														assign node14756 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node14759 = (inp[9]) ? node14765 : node14760;
															assign node14760 = (inp[12]) ? node14762 : 4'b0000;
																assign node14762 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node14765 = (inp[12]) ? node14767 : 4'b0100;
																assign node14767 = (inp[10]) ? 4'b0000 : 4'b0100;
									assign node14770 = (inp[5]) ? node14858 : node14771;
										assign node14771 = (inp[9]) ? node14825 : node14772;
											assign node14772 = (inp[4]) ? node14796 : node14773;
												assign node14773 = (inp[10]) ? node14787 : node14774;
													assign node14774 = (inp[12]) ? node14782 : node14775;
														assign node14775 = (inp[15]) ? node14779 : node14776;
															assign node14776 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node14779 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node14782 = (inp[0]) ? 4'b1001 : node14783;
															assign node14783 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node14787 = (inp[12]) ? 4'b1011 : node14788;
														assign node14788 = (inp[0]) ? node14792 : node14789;
															assign node14789 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node14792 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node14796 = (inp[12]) ? node14810 : node14797;
													assign node14797 = (inp[10]) ? node14805 : node14798;
														assign node14798 = (inp[15]) ? node14802 : node14799;
															assign node14799 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node14802 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node14805 = (inp[3]) ? node14807 : 4'b1101;
															assign node14807 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node14810 = (inp[10]) ? node14818 : node14811;
														assign node14811 = (inp[0]) ? 4'b1101 : node14812;
															assign node14812 = (inp[15]) ? node14814 : 4'b1101;
																assign node14814 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node14818 = (inp[15]) ? node14820 : 4'b1111;
															assign node14820 = (inp[3]) ? node14822 : 4'b1111;
																assign node14822 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node14825 = (inp[4]) ? node14841 : node14826;
												assign node14826 = (inp[12]) ? node14832 : node14827;
													assign node14827 = (inp[10]) ? 4'b1111 : node14828;
														assign node14828 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node14832 = (inp[0]) ? node14834 : 4'b1111;
														assign node14834 = (inp[3]) ? node14838 : node14835;
															assign node14835 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node14838 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node14841 = (inp[3]) ? node14849 : node14842;
													assign node14842 = (inp[0]) ? node14846 : node14843;
														assign node14843 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node14846 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node14849 = (inp[10]) ? node14853 : node14850;
														assign node14850 = (inp[15]) ? 4'b1011 : 4'b1111;
														assign node14853 = (inp[15]) ? node14855 : 4'b1011;
															assign node14855 = (inp[12]) ? 4'b1011 : 4'b1001;
										assign node14858 = (inp[10]) ? node14908 : node14859;
											assign node14859 = (inp[15]) ? node14871 : node14860;
												assign node14860 = (inp[9]) ? 4'b1101 : node14861;
													assign node14861 = (inp[4]) ? node14867 : node14862;
														assign node14862 = (inp[0]) ? 4'b1111 : node14863;
															assign node14863 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node14867 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node14871 = (inp[0]) ? node14891 : node14872;
													assign node14872 = (inp[3]) ? node14886 : node14873;
														assign node14873 = (inp[12]) ? node14881 : node14874;
															assign node14874 = (inp[4]) ? node14878 : node14875;
																assign node14875 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node14878 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node14881 = (inp[9]) ? node14883 : 4'b1111;
																assign node14883 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node14886 = (inp[4]) ? 4'b1011 : node14887;
															assign node14887 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node14891 = (inp[3]) ? node14899 : node14892;
														assign node14892 = (inp[4]) ? 4'b1101 : node14893;
															assign node14893 = (inp[9]) ? 4'b1101 : node14894;
																assign node14894 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node14899 = (inp[9]) ? 4'b1001 : node14900;
															assign node14900 = (inp[4]) ? node14904 : node14901;
																assign node14901 = (inp[12]) ? 4'b1001 : 4'b1101;
																assign node14904 = (inp[12]) ? 4'b1101 : 4'b1001;
											assign node14908 = (inp[15]) ? node14926 : node14909;
												assign node14909 = (inp[0]) ? node14919 : node14910;
													assign node14910 = (inp[9]) ? node14916 : node14911;
														assign node14911 = (inp[4]) ? 4'b1101 : node14912;
															assign node14912 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node14916 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node14919 = (inp[9]) ? node14923 : node14920;
														assign node14920 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node14923 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node14926 = (inp[0]) ? node14938 : node14927;
													assign node14927 = (inp[3]) ? node14931 : node14928;
														assign node14928 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node14931 = (inp[12]) ? 4'b1011 : node14932;
															assign node14932 = (inp[4]) ? node14934 : 4'b1111;
																assign node14934 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node14938 = (inp[9]) ? node14944 : node14939;
														assign node14939 = (inp[4]) ? 4'b1101 : node14940;
															assign node14940 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node14944 = (inp[4]) ? 4'b1001 : 4'b1101;
							assign node14947 = (inp[8]) ? node15307 : node14948;
								assign node14948 = (inp[7]) ? node15134 : node14949;
									assign node14949 = (inp[4]) ? node15049 : node14950;
										assign node14950 = (inp[9]) ? node15000 : node14951;
											assign node14951 = (inp[12]) ? node14977 : node14952;
												assign node14952 = (inp[5]) ? node14966 : node14953;
													assign node14953 = (inp[3]) ? node14959 : node14954;
														assign node14954 = (inp[0]) ? 4'b0110 : node14955;
															assign node14955 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node14959 = (inp[0]) ? node14963 : node14960;
															assign node14960 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node14963 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node14966 = (inp[3]) ? 4'b0100 : node14967;
														assign node14967 = (inp[10]) ? node14973 : node14968;
															assign node14968 = (inp[0]) ? 4'b0100 : node14969;
																assign node14969 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node14973 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node14977 = (inp[10]) ? node14989 : node14978;
													assign node14978 = (inp[3]) ? node14984 : node14979;
														assign node14979 = (inp[5]) ? node14981 : 4'b0100;
															assign node14981 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node14984 = (inp[0]) ? node14986 : 4'b0110;
															assign node14986 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node14989 = (inp[0]) ? node14997 : node14990;
														assign node14990 = (inp[15]) ? node14994 : node14991;
															assign node14991 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node14994 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node14997 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node15000 = (inp[12]) ? node15030 : node15001;
												assign node15001 = (inp[3]) ? node15015 : node15002;
													assign node15002 = (inp[5]) ? node15010 : node15003;
														assign node15003 = (inp[0]) ? node15007 : node15004;
															assign node15004 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node15007 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node15010 = (inp[15]) ? 4'b0000 : node15011;
															assign node15011 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node15015 = (inp[15]) ? node15025 : node15016;
														assign node15016 = (inp[10]) ? node15020 : node15017;
															assign node15017 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node15020 = (inp[5]) ? node15022 : 4'b0010;
																assign node15022 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node15025 = (inp[5]) ? 4'b0010 : node15026;
															assign node15026 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node15030 = (inp[10]) ? node15040 : node15031;
													assign node15031 = (inp[15]) ? 4'b0000 : node15032;
														assign node15032 = (inp[0]) ? 4'b0000 : node15033;
															assign node15033 = (inp[5]) ? node15035 : 4'b0010;
																assign node15035 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node15040 = (inp[3]) ? node15042 : 4'b0110;
														assign node15042 = (inp[15]) ? node15046 : node15043;
															assign node15043 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node15046 = (inp[0]) ? 4'b0100 : 4'b0110;
										assign node15049 = (inp[9]) ? node15105 : node15050;
											assign node15050 = (inp[12]) ? node15076 : node15051;
												assign node15051 = (inp[5]) ? node15059 : node15052;
													assign node15052 = (inp[10]) ? 4'b0000 : node15053;
														assign node15053 = (inp[15]) ? 4'b0010 : node15054;
															assign node15054 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node15059 = (inp[10]) ? node15061 : 4'b0010;
														assign node15061 = (inp[15]) ? node15069 : node15062;
															assign node15062 = (inp[0]) ? node15066 : node15063;
																assign node15063 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node15066 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node15069 = (inp[0]) ? node15073 : node15070;
																assign node15070 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node15073 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node15076 = (inp[10]) ? node15090 : node15077;
													assign node15077 = (inp[3]) ? node15085 : node15078;
														assign node15078 = (inp[15]) ? node15082 : node15079;
															assign node15079 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node15082 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node15085 = (inp[5]) ? node15087 : 4'b0000;
															assign node15087 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node15090 = (inp[0]) ? node15096 : node15091;
														assign node15091 = (inp[5]) ? node15093 : 4'b0100;
															assign node15093 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node15096 = (inp[15]) ? node15102 : node15097;
															assign node15097 = (inp[5]) ? 4'b0110 : node15098;
																assign node15098 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node15102 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node15105 = (inp[12]) ? node15123 : node15106;
												assign node15106 = (inp[15]) ? node15116 : node15107;
													assign node15107 = (inp[0]) ? node15113 : node15108;
														assign node15108 = (inp[3]) ? 4'b0100 : node15109;
															assign node15109 = (inp[10]) ? 4'b0110 : 4'b0100;
														assign node15113 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node15116 = (inp[0]) ? node15118 : 4'b0110;
														assign node15118 = (inp[3]) ? 4'b0100 : node15119;
															assign node15119 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node15123 = (inp[10]) ? node15131 : node15124;
													assign node15124 = (inp[15]) ? 4'b0100 : node15125;
														assign node15125 = (inp[5]) ? 4'b0110 : node15126;
															assign node15126 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node15131 = (inp[15]) ? 4'b0010 : 4'b0000;
									assign node15134 = (inp[9]) ? node15222 : node15135;
										assign node15135 = (inp[4]) ? node15177 : node15136;
											assign node15136 = (inp[12]) ? node15160 : node15137;
												assign node15137 = (inp[10]) ? node15155 : node15138;
													assign node15138 = (inp[5]) ? node15146 : node15139;
														assign node15139 = (inp[3]) ? 4'b1101 : node15140;
															assign node15140 = (inp[15]) ? node15142 : 4'b1101;
																assign node15142 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node15146 = (inp[15]) ? 4'b1111 : node15147;
															assign node15147 = (inp[0]) ? node15151 : node15148;
																assign node15148 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node15151 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node15155 = (inp[5]) ? 4'b1011 : node15156;
														assign node15156 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node15160 = (inp[0]) ? node15172 : node15161;
													assign node15161 = (inp[10]) ? node15167 : node15162;
														assign node15162 = (inp[15]) ? node15164 : 4'b1011;
															assign node15164 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node15167 = (inp[5]) ? node15169 : 4'b1001;
															assign node15169 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node15172 = (inp[3]) ? node15174 : 4'b1011;
														assign node15174 = (inp[10]) ? 4'b1011 : 4'b1001;
											assign node15177 = (inp[10]) ? node15201 : node15178;
												assign node15178 = (inp[12]) ? node15190 : node15179;
													assign node15179 = (inp[5]) ? node15181 : 4'b1011;
														assign node15181 = (inp[3]) ? node15183 : 4'b1011;
															assign node15183 = (inp[0]) ? node15187 : node15184;
																assign node15184 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node15187 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node15190 = (inp[15]) ? node15196 : node15191;
														assign node15191 = (inp[0]) ? node15193 : 4'b1101;
															assign node15193 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node15196 = (inp[0]) ? node15198 : 4'b1111;
															assign node15198 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node15201 = (inp[15]) ? node15207 : node15202;
													assign node15202 = (inp[0]) ? 4'b1111 : node15203;
														assign node15203 = (inp[12]) ? 4'b1111 : 4'b1101;
													assign node15207 = (inp[3]) ? 4'b1101 : node15208;
														assign node15208 = (inp[12]) ? node15214 : node15209;
															assign node15209 = (inp[5]) ? node15211 : 4'b1101;
																assign node15211 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node15214 = (inp[0]) ? node15218 : node15215;
																assign node15215 = (inp[5]) ? 4'b1111 : 4'b1101;
																assign node15218 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node15222 = (inp[4]) ? node15268 : node15223;
											assign node15223 = (inp[10]) ? node15251 : node15224;
												assign node15224 = (inp[12]) ? node15242 : node15225;
													assign node15225 = (inp[5]) ? node15233 : node15226;
														assign node15226 = (inp[0]) ? node15230 : node15227;
															assign node15227 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node15230 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node15233 = (inp[0]) ? 4'b1011 : node15234;
															assign node15234 = (inp[15]) ? node15238 : node15235;
																assign node15235 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node15238 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node15242 = (inp[0]) ? node15248 : node15243;
														assign node15243 = (inp[15]) ? node15245 : 4'b1101;
															assign node15245 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node15248 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node15251 = (inp[15]) ? node15263 : node15252;
													assign node15252 = (inp[0]) ? node15258 : node15253;
														assign node15253 = (inp[3]) ? 4'b1101 : node15254;
															assign node15254 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node15258 = (inp[12]) ? node15260 : 4'b1111;
															assign node15260 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node15263 = (inp[0]) ? 4'b1101 : node15264;
														assign node15264 = (inp[3]) ? 4'b1111 : 4'b1101;
											assign node15268 = (inp[10]) ? node15288 : node15269;
												assign node15269 = (inp[12]) ? node15281 : node15270;
													assign node15270 = (inp[3]) ? 4'b1101 : node15271;
														assign node15271 = (inp[15]) ? node15273 : 4'b1111;
															assign node15273 = (inp[5]) ? node15277 : node15274;
																assign node15274 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node15277 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node15281 = (inp[3]) ? node15283 : 4'b1011;
														assign node15283 = (inp[0]) ? 4'b1001 : node15284;
															assign node15284 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node15288 = (inp[3]) ? node15296 : node15289;
													assign node15289 = (inp[12]) ? node15291 : 4'b1001;
														assign node15291 = (inp[15]) ? node15293 : 4'b1001;
															assign node15293 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node15296 = (inp[12]) ? node15302 : node15297;
														assign node15297 = (inp[5]) ? node15299 : 4'b1011;
															assign node15299 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node15302 = (inp[15]) ? 4'b1001 : node15303;
															assign node15303 = (inp[0]) ? 4'b1011 : 4'b1001;
								assign node15307 = (inp[7]) ? node15479 : node15308;
									assign node15308 = (inp[4]) ? node15396 : node15309;
										assign node15309 = (inp[9]) ? node15343 : node15310;
											assign node15310 = (inp[12]) ? node15324 : node15311;
												assign node15311 = (inp[10]) ? node15317 : node15312;
													assign node15312 = (inp[0]) ? node15314 : 4'b1111;
														assign node15314 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node15317 = (inp[5]) ? node15319 : 4'b1001;
														assign node15319 = (inp[0]) ? node15321 : 4'b1011;
															assign node15321 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node15324 = (inp[15]) ? node15332 : node15325;
													assign node15325 = (inp[0]) ? node15327 : 4'b1011;
														assign node15327 = (inp[5]) ? node15329 : 4'b1001;
															assign node15329 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node15332 = (inp[0]) ? node15338 : node15333;
														assign node15333 = (inp[5]) ? node15335 : 4'b1001;
															assign node15335 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node15338 = (inp[3]) ? node15340 : 4'b1011;
															assign node15340 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node15343 = (inp[12]) ? node15373 : node15344;
												assign node15344 = (inp[10]) ? node15358 : node15345;
													assign node15345 = (inp[15]) ? node15353 : node15346;
														assign node15346 = (inp[0]) ? node15350 : node15347;
															assign node15347 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node15350 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node15353 = (inp[0]) ? node15355 : 4'b1001;
															assign node15355 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node15358 = (inp[5]) ? node15368 : node15359;
														assign node15359 = (inp[0]) ? 4'b1101 : node15360;
															assign node15360 = (inp[15]) ? node15364 : node15361;
																assign node15361 = (inp[3]) ? 4'b1101 : 4'b1111;
																assign node15364 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node15368 = (inp[3]) ? node15370 : 4'b1111;
															assign node15370 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node15373 = (inp[5]) ? node15387 : node15374;
													assign node15374 = (inp[3]) ? node15380 : node15375;
														assign node15375 = (inp[15]) ? node15377 : 4'b1111;
															assign node15377 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node15380 = (inp[10]) ? 4'b1101 : node15381;
															assign node15381 = (inp[0]) ? 4'b1111 : node15382;
																assign node15382 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node15387 = (inp[10]) ? node15389 : 4'b1101;
														assign node15389 = (inp[0]) ? node15393 : node15390;
															assign node15390 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node15393 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node15396 = (inp[9]) ? node15436 : node15397;
											assign node15397 = (inp[12]) ? node15415 : node15398;
												assign node15398 = (inp[10]) ? node15406 : node15399;
													assign node15399 = (inp[5]) ? 4'b1011 : node15400;
														assign node15400 = (inp[0]) ? 4'b1001 : node15401;
															assign node15401 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node15406 = (inp[3]) ? 4'b1101 : node15407;
														assign node15407 = (inp[5]) ? 4'b1111 : node15408;
															assign node15408 = (inp[0]) ? node15410 : 4'b1111;
																assign node15410 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node15415 = (inp[10]) ? node15427 : node15416;
													assign node15416 = (inp[15]) ? node15422 : node15417;
														assign node15417 = (inp[0]) ? node15419 : 4'b1101;
															assign node15419 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node15422 = (inp[3]) ? node15424 : 4'b1111;
															assign node15424 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node15427 = (inp[3]) ? node15429 : 4'b1111;
														assign node15429 = (inp[0]) ? node15433 : node15430;
															assign node15430 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node15433 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node15436 = (inp[12]) ? node15466 : node15437;
												assign node15437 = (inp[10]) ? node15459 : node15438;
													assign node15438 = (inp[3]) ? node15452 : node15439;
														assign node15439 = (inp[0]) ? node15447 : node15440;
															assign node15440 = (inp[5]) ? node15444 : node15441;
																assign node15441 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node15444 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node15447 = (inp[15]) ? node15449 : 4'b1101;
																assign node15449 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node15452 = (inp[5]) ? node15454 : 4'b1111;
															assign node15454 = (inp[15]) ? node15456 : 4'b1111;
																assign node15456 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node15459 = (inp[3]) ? node15461 : 4'b1001;
														assign node15461 = (inp[0]) ? 4'b1011 : node15462;
															assign node15462 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node15466 = (inp[3]) ? node15468 : 4'b1011;
													assign node15468 = (inp[10]) ? node15474 : node15469;
														assign node15469 = (inp[15]) ? 4'b1011 : node15470;
															assign node15470 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node15474 = (inp[15]) ? 4'b1001 : node15475;
															assign node15475 = (inp[0]) ? 4'b1011 : 4'b1001;
									assign node15479 = (inp[10]) ? node15597 : node15480;
										assign node15480 = (inp[3]) ? node15546 : node15481;
											assign node15481 = (inp[4]) ? node15513 : node15482;
												assign node15482 = (inp[15]) ? node15502 : node15483;
													assign node15483 = (inp[0]) ? node15489 : node15484;
														assign node15484 = (inp[12]) ? 4'b1100 : node15485;
															assign node15485 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node15489 = (inp[5]) ? node15497 : node15490;
															assign node15490 = (inp[9]) ? node15494 : node15491;
																assign node15491 = (inp[12]) ? 4'b1000 : 4'b1100;
																assign node15494 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node15497 = (inp[12]) ? node15499 : 4'b1000;
																assign node15499 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node15502 = (inp[0]) ? node15504 : 4'b1100;
														assign node15504 = (inp[5]) ? 4'b1110 : node15505;
															assign node15505 = (inp[9]) ? node15509 : node15506;
																assign node15506 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node15509 = (inp[12]) ? 4'b1110 : 4'b1010;
												assign node15513 = (inp[9]) ? node15529 : node15514;
													assign node15514 = (inp[12]) ? node15516 : 4'b1000;
														assign node15516 = (inp[0]) ? node15524 : node15517;
															assign node15517 = (inp[15]) ? node15521 : node15518;
																assign node15518 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node15521 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node15524 = (inp[5]) ? node15526 : 4'b1100;
																assign node15526 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node15529 = (inp[12]) ? node15539 : node15530;
														assign node15530 = (inp[0]) ? node15532 : 4'b1100;
															assign node15532 = (inp[15]) ? node15536 : node15533;
																assign node15533 = (inp[5]) ? 4'b1110 : 4'b1100;
																assign node15536 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node15539 = (inp[0]) ? node15541 : 4'b1000;
															assign node15541 = (inp[15]) ? 4'b1000 : node15542;
																assign node15542 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node15546 = (inp[12]) ? node15572 : node15547;
												assign node15547 = (inp[9]) ? node15561 : node15548;
													assign node15548 = (inp[4]) ? node15556 : node15549;
														assign node15549 = (inp[15]) ? node15551 : 4'b1110;
															assign node15551 = (inp[0]) ? 4'b1100 : node15552;
																assign node15552 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node15556 = (inp[0]) ? node15558 : 4'b1000;
															assign node15558 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node15561 = (inp[4]) ? node15567 : node15562;
														assign node15562 = (inp[5]) ? 4'b1010 : node15563;
															assign node15563 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node15567 = (inp[5]) ? 4'b1110 : node15568;
															assign node15568 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node15572 = (inp[9]) ? node15584 : node15573;
													assign node15573 = (inp[4]) ? 4'b1100 : node15574;
														assign node15574 = (inp[0]) ? node15576 : 4'b1000;
															assign node15576 = (inp[5]) ? node15580 : node15577;
																assign node15577 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node15580 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node15584 = (inp[4]) ? node15590 : node15585;
														assign node15585 = (inp[0]) ? 4'b1100 : node15586;
															assign node15586 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node15590 = (inp[0]) ? node15594 : node15591;
															assign node15591 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node15594 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node15597 = (inp[0]) ? node15649 : node15598;
											assign node15598 = (inp[12]) ? node15628 : node15599;
												assign node15599 = (inp[15]) ? node15609 : node15600;
													assign node15600 = (inp[3]) ? 4'b1100 : node15601;
														assign node15601 = (inp[5]) ? node15605 : node15602;
															assign node15602 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node15605 = (inp[9]) ? 4'b1000 : 4'b1010;
													assign node15609 = (inp[5]) ? node15619 : node15610;
														assign node15610 = (inp[4]) ? node15616 : node15611;
															assign node15611 = (inp[9]) ? node15613 : 4'b1000;
																assign node15613 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node15616 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node15619 = (inp[3]) ? node15621 : 4'b1110;
															assign node15621 = (inp[4]) ? node15625 : node15622;
																assign node15622 = (inp[9]) ? 4'b1110 : 4'b1010;
																assign node15625 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node15628 = (inp[9]) ? node15638 : node15629;
													assign node15629 = (inp[4]) ? 4'b1110 : node15630;
														assign node15630 = (inp[15]) ? node15632 : 4'b1010;
															assign node15632 = (inp[5]) ? node15634 : 4'b1000;
																assign node15634 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node15638 = (inp[4]) ? node15640 : 4'b1110;
														assign node15640 = (inp[15]) ? node15644 : node15641;
															assign node15641 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node15644 = (inp[3]) ? 4'b1010 : node15645;
																assign node15645 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node15649 = (inp[12]) ? node15671 : node15650;
												assign node15650 = (inp[9]) ? node15658 : node15651;
													assign node15651 = (inp[4]) ? 4'b1110 : node15652;
														assign node15652 = (inp[5]) ? node15654 : 4'b1010;
															assign node15654 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node15658 = (inp[4]) ? node15668 : node15659;
														assign node15659 = (inp[5]) ? node15665 : node15660;
															assign node15660 = (inp[3]) ? 4'b1110 : node15661;
																assign node15661 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node15665 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node15668 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node15671 = (inp[3]) ? node15683 : node15672;
													assign node15672 = (inp[15]) ? node15676 : node15673;
														assign node15673 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node15676 = (inp[5]) ? 4'b1010 : node15677;
															assign node15677 = (inp[4]) ? node15679 : 4'b1110;
																assign node15679 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node15683 = (inp[15]) ? node15687 : node15684;
														assign node15684 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node15687 = (inp[9]) ? node15689 : 4'b1100;
															assign node15689 = (inp[4]) ? 4'b1000 : 4'b1100;
					assign node15692 = (inp[1]) ? node17174 : node15693;
						assign node15693 = (inp[2]) ? node16439 : node15694;
							assign node15694 = (inp[8]) ? node16058 : node15695;
								assign node15695 = (inp[7]) ? node15867 : node15696;
									assign node15696 = (inp[9]) ? node15778 : node15697;
										assign node15697 = (inp[4]) ? node15735 : node15698;
											assign node15698 = (inp[10]) ? node15716 : node15699;
												assign node15699 = (inp[15]) ? node15707 : node15700;
													assign node15700 = (inp[0]) ? 4'b0101 : node15701;
														assign node15701 = (inp[5]) ? node15703 : 4'b0111;
															assign node15703 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node15707 = (inp[0]) ? node15711 : node15708;
														assign node15708 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node15711 = (inp[5]) ? node15713 : 4'b0111;
															assign node15713 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node15716 = (inp[12]) ? node15728 : node15717;
													assign node15717 = (inp[5]) ? node15719 : 4'b0111;
														assign node15719 = (inp[0]) ? node15721 : 4'b0111;
															assign node15721 = (inp[15]) ? node15725 : node15722;
																assign node15722 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node15725 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node15728 = (inp[5]) ? node15730 : 4'b0001;
														assign node15730 = (inp[15]) ? 4'b0011 : node15731;
															assign node15731 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node15735 = (inp[10]) ? node15757 : node15736;
												assign node15736 = (inp[5]) ? node15742 : node15737;
													assign node15737 = (inp[15]) ? node15739 : 4'b0011;
														assign node15739 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node15742 = (inp[15]) ? node15748 : node15743;
														assign node15743 = (inp[0]) ? node15745 : 4'b0001;
															assign node15745 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node15748 = (inp[12]) ? node15752 : node15749;
															assign node15749 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node15752 = (inp[3]) ? node15754 : 4'b0011;
																assign node15754 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node15757 = (inp[12]) ? node15767 : node15758;
													assign node15758 = (inp[0]) ? 4'b0011 : node15759;
														assign node15759 = (inp[15]) ? node15763 : node15760;
															assign node15760 = (inp[5]) ? 4'b0001 : 4'b0011;
															assign node15763 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node15767 = (inp[15]) ? node15769 : 4'b0101;
														assign node15769 = (inp[0]) ? node15773 : node15770;
															assign node15770 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node15773 = (inp[3]) ? 4'b0101 : node15774;
																assign node15774 = (inp[5]) ? 4'b0101 : 4'b0111;
										assign node15778 = (inp[4]) ? node15824 : node15779;
											assign node15779 = (inp[12]) ? node15803 : node15780;
												assign node15780 = (inp[10]) ? node15788 : node15781;
													assign node15781 = (inp[3]) ? node15783 : 4'b0011;
														assign node15783 = (inp[0]) ? 4'b0011 : node15784;
															assign node15784 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node15788 = (inp[0]) ? node15794 : node15789;
														assign node15789 = (inp[15]) ? 4'b0001 : node15790;
															assign node15790 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node15794 = (inp[3]) ? node15796 : 4'b0011;
															assign node15796 = (inp[5]) ? node15800 : node15797;
																assign node15797 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node15800 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node15803 = (inp[10]) ? node15817 : node15804;
													assign node15804 = (inp[0]) ? node15812 : node15805;
														assign node15805 = (inp[3]) ? node15809 : node15806;
															assign node15806 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node15809 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node15812 = (inp[15]) ? node15814 : 4'b0001;
															assign node15814 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node15817 = (inp[5]) ? 4'b0101 : node15818;
														assign node15818 = (inp[15]) ? 4'b0111 : node15819;
															assign node15819 = (inp[0]) ? 4'b0111 : 4'b0101;
											assign node15824 = (inp[12]) ? node15850 : node15825;
												assign node15825 = (inp[5]) ? node15843 : node15826;
													assign node15826 = (inp[0]) ? node15832 : node15827;
														assign node15827 = (inp[3]) ? 4'b0101 : node15828;
															assign node15828 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node15832 = (inp[10]) ? node15838 : node15833;
															assign node15833 = (inp[15]) ? node15835 : 4'b0111;
																assign node15835 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node15838 = (inp[15]) ? 4'b0111 : node15839;
																assign node15839 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node15843 = (inp[10]) ? 4'b0101 : node15844;
														assign node15844 = (inp[15]) ? node15846 : 4'b0101;
															assign node15846 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node15850 = (inp[10]) ? node15856 : node15851;
													assign node15851 = (inp[0]) ? 4'b0101 : node15852;
														assign node15852 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node15856 = (inp[0]) ? node15862 : node15857;
														assign node15857 = (inp[5]) ? node15859 : 4'b0011;
															assign node15859 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node15862 = (inp[15]) ? 4'b0001 : node15863;
															assign node15863 = (inp[5]) ? 4'b0011 : 4'b0001;
									assign node15867 = (inp[5]) ? node15951 : node15868;
										assign node15868 = (inp[3]) ? node15902 : node15869;
											assign node15869 = (inp[15]) ? node15883 : node15870;
												assign node15870 = (inp[0]) ? node15878 : node15871;
													assign node15871 = (inp[9]) ? 4'b0110 : node15872;
														assign node15872 = (inp[10]) ? 4'b0010 : node15873;
															assign node15873 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node15878 = (inp[10]) ? node15880 : 4'b0100;
														assign node15880 = (inp[12]) ? 4'b0100 : 4'b0000;
												assign node15883 = (inp[0]) ? node15891 : node15884;
													assign node15884 = (inp[9]) ? 4'b0000 : node15885;
														assign node15885 = (inp[4]) ? node15887 : 4'b0100;
															assign node15887 = (inp[12]) ? 4'b0100 : 4'b0000;
													assign node15891 = (inp[12]) ? node15897 : node15892;
														assign node15892 = (inp[9]) ? 4'b0110 : node15893;
															assign node15893 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node15897 = (inp[4]) ? node15899 : 4'b0010;
															assign node15899 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node15902 = (inp[4]) ? node15924 : node15903;
												assign node15903 = (inp[9]) ? node15913 : node15904;
													assign node15904 = (inp[12]) ? node15910 : node15905;
														assign node15905 = (inp[10]) ? 4'b0110 : node15906;
															assign node15906 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node15910 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node15913 = (inp[10]) ? node15917 : node15914;
														assign node15914 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node15917 = (inp[12]) ? node15921 : node15918;
															assign node15918 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node15921 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node15924 = (inp[9]) ? node15942 : node15925;
													assign node15925 = (inp[12]) ? node15933 : node15926;
														assign node15926 = (inp[10]) ? node15928 : 4'b0010;
															assign node15928 = (inp[15]) ? node15930 : 4'b0000;
																assign node15930 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node15933 = (inp[10]) ? node15935 : 4'b0010;
															assign node15935 = (inp[0]) ? node15939 : node15936;
																assign node15936 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node15939 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node15942 = (inp[12]) ? node15948 : node15943;
														assign node15943 = (inp[0]) ? node15945 : 4'b0110;
															assign node15945 = (inp[10]) ? 4'b0110 : 4'b0100;
														assign node15948 = (inp[10]) ? 4'b0010 : 4'b0110;
										assign node15951 = (inp[4]) ? node16005 : node15952;
											assign node15952 = (inp[9]) ? node15982 : node15953;
												assign node15953 = (inp[10]) ? node15965 : node15954;
													assign node15954 = (inp[3]) ? node15960 : node15955;
														assign node15955 = (inp[12]) ? 4'b0110 : node15956;
															assign node15956 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node15960 = (inp[0]) ? 4'b0100 : node15961;
															assign node15961 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node15965 = (inp[12]) ? node15973 : node15966;
														assign node15966 = (inp[3]) ? node15968 : 4'b0100;
															assign node15968 = (inp[0]) ? 4'b0110 : node15969;
																assign node15969 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node15973 = (inp[0]) ? 4'b0000 : node15974;
															assign node15974 = (inp[15]) ? node15978 : node15975;
																assign node15975 = (inp[3]) ? 4'b0000 : 4'b0010;
																assign node15978 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node15982 = (inp[10]) ? node15996 : node15983;
													assign node15983 = (inp[15]) ? node15989 : node15984;
														assign node15984 = (inp[0]) ? 4'b0010 : node15985;
															assign node15985 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node15989 = (inp[0]) ? node15993 : node15990;
															assign node15990 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node15993 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node15996 = (inp[12]) ? node16002 : node15997;
														assign node15997 = (inp[3]) ? 4'b0000 : node15998;
															assign node15998 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node16002 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node16005 = (inp[9]) ? node16029 : node16006;
												assign node16006 = (inp[10]) ? node16016 : node16007;
													assign node16007 = (inp[0]) ? node16009 : 4'b0000;
														assign node16009 = (inp[3]) ? node16013 : node16010;
															assign node16010 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node16013 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node16016 = (inp[12]) ? node16024 : node16017;
														assign node16017 = (inp[0]) ? node16019 : 4'b0010;
															assign node16019 = (inp[15]) ? node16021 : 4'b0010;
																assign node16021 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node16024 = (inp[15]) ? 4'b0110 : node16025;
															assign node16025 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node16029 = (inp[12]) ? node16045 : node16030;
													assign node16030 = (inp[3]) ? node16040 : node16031;
														assign node16031 = (inp[10]) ? node16033 : 4'b0100;
															assign node16033 = (inp[15]) ? node16037 : node16034;
																assign node16034 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node16037 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node16040 = (inp[15]) ? 4'b0110 : node16041;
															assign node16041 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node16045 = (inp[10]) ? node16053 : node16046;
														assign node16046 = (inp[15]) ? node16050 : node16047;
															assign node16047 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node16050 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node16053 = (inp[15]) ? node16055 : 4'b0000;
															assign node16055 = (inp[0]) ? 4'b0000 : 4'b0010;
								assign node16058 = (inp[7]) ? node16254 : node16059;
									assign node16059 = (inp[15]) ? node16163 : node16060;
										assign node16060 = (inp[12]) ? node16114 : node16061;
											assign node16061 = (inp[10]) ? node16081 : node16062;
												assign node16062 = (inp[3]) ? node16072 : node16063;
													assign node16063 = (inp[0]) ? node16069 : node16064;
														assign node16064 = (inp[9]) ? 4'b0110 : node16065;
															assign node16065 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node16069 = (inp[4]) ? 4'b0110 : 4'b0000;
													assign node16072 = (inp[5]) ? 4'b0110 : node16073;
														assign node16073 = (inp[9]) ? node16077 : node16074;
															assign node16074 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node16077 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node16081 = (inp[0]) ? node16103 : node16082;
													assign node16082 = (inp[3]) ? node16092 : node16083;
														assign node16083 = (inp[4]) ? node16087 : node16084;
															assign node16084 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node16087 = (inp[5]) ? 4'b0100 : node16088;
																assign node16088 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node16092 = (inp[5]) ? node16098 : node16093;
															assign node16093 = (inp[9]) ? node16095 : 4'b0010;
																assign node16095 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node16098 = (inp[4]) ? node16100 : 4'b0000;
																assign node16100 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node16103 = (inp[5]) ? node16109 : node16104;
														assign node16104 = (inp[3]) ? node16106 : 4'b0000;
															assign node16106 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node16109 = (inp[4]) ? 4'b0110 : node16110;
															assign node16110 = (inp[9]) ? 4'b0000 : 4'b0100;
											assign node16114 = (inp[5]) ? node16140 : node16115;
												assign node16115 = (inp[0]) ? node16127 : node16116;
													assign node16116 = (inp[3]) ? node16122 : node16117;
														assign node16117 = (inp[4]) ? node16119 : 4'b0010;
															assign node16119 = (inp[10]) ? 4'b0110 : 4'b0010;
														assign node16122 = (inp[9]) ? node16124 : 4'b0100;
															assign node16124 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node16127 = (inp[9]) ? node16133 : node16128;
														assign node16128 = (inp[4]) ? 4'b0000 : node16129;
															assign node16129 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node16133 = (inp[10]) ? node16137 : node16134;
															assign node16134 = (inp[3]) ? 4'b0000 : 4'b0100;
															assign node16137 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node16140 = (inp[0]) ? node16146 : node16141;
													assign node16141 = (inp[10]) ? node16143 : 4'b0100;
														assign node16143 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node16146 = (inp[3]) ? node16154 : node16147;
														assign node16147 = (inp[10]) ? 4'b0010 : node16148;
															assign node16148 = (inp[9]) ? 4'b0000 : node16149;
																assign node16149 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node16154 = (inp[10]) ? 4'b0110 : node16155;
															assign node16155 = (inp[9]) ? node16159 : node16156;
																assign node16156 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node16159 = (inp[4]) ? 4'b0110 : 4'b0010;
										assign node16163 = (inp[0]) ? node16217 : node16164;
											assign node16164 = (inp[3]) ? node16190 : node16165;
												assign node16165 = (inp[5]) ? node16179 : node16166;
													assign node16166 = (inp[10]) ? node16172 : node16167;
														assign node16167 = (inp[12]) ? node16169 : 4'b0000;
															assign node16169 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node16172 = (inp[4]) ? node16174 : 4'b0100;
															assign node16174 = (inp[9]) ? node16176 : 4'b0100;
																assign node16176 = (inp[12]) ? 4'b0000 : 4'b0100;
													assign node16179 = (inp[9]) ? node16185 : node16180;
														assign node16180 = (inp[10]) ? 4'b0000 : node16181;
															assign node16181 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node16185 = (inp[4]) ? 4'b0110 : node16186;
															assign node16186 = (inp[10]) ? 4'b0110 : 4'b0000;
												assign node16190 = (inp[4]) ? node16206 : node16191;
													assign node16191 = (inp[5]) ? node16199 : node16192;
														assign node16192 = (inp[12]) ? node16194 : 4'b0000;
															assign node16194 = (inp[10]) ? node16196 : 4'b0000;
																assign node16196 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node16199 = (inp[9]) ? node16203 : node16200;
															assign node16200 = (inp[10]) ? 4'b0010 : 4'b0110;
															assign node16203 = (inp[10]) ? 4'b0110 : 4'b0010;
													assign node16206 = (inp[9]) ? node16212 : node16207;
														assign node16207 = (inp[10]) ? 4'b0110 : node16208;
															assign node16208 = (inp[12]) ? 4'b0000 : 4'b0010;
														assign node16212 = (inp[12]) ? node16214 : 4'b0110;
															assign node16214 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node16217 = (inp[5]) ? node16233 : node16218;
												assign node16218 = (inp[4]) ? node16228 : node16219;
													assign node16219 = (inp[9]) ? node16223 : node16220;
														assign node16220 = (inp[3]) ? 4'b0110 : 4'b0010;
														assign node16223 = (inp[12]) ? node16225 : 4'b0010;
															assign node16225 = (inp[3]) ? 4'b0010 : 4'b0110;
													assign node16228 = (inp[9]) ? node16230 : 4'b0010;
														assign node16230 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node16233 = (inp[3]) ? node16247 : node16234;
													assign node16234 = (inp[9]) ? node16242 : node16235;
														assign node16235 = (inp[4]) ? 4'b0010 : node16236;
															assign node16236 = (inp[12]) ? node16238 : 4'b0110;
																assign node16238 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node16242 = (inp[12]) ? 4'b0100 : node16243;
															assign node16243 = (inp[4]) ? 4'b0100 : 4'b0010;
													assign node16247 = (inp[10]) ? node16249 : 4'b0000;
														assign node16249 = (inp[9]) ? node16251 : 4'b0000;
															assign node16251 = (inp[12]) ? 4'b0100 : 4'b0000;
									assign node16254 = (inp[3]) ? node16368 : node16255;
										assign node16255 = (inp[4]) ? node16319 : node16256;
											assign node16256 = (inp[9]) ? node16282 : node16257;
												assign node16257 = (inp[12]) ? node16267 : node16258;
													assign node16258 = (inp[10]) ? 4'b1011 : node16259;
														assign node16259 = (inp[15]) ? node16263 : node16260;
															assign node16260 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node16263 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node16267 = (inp[5]) ? node16277 : node16268;
														assign node16268 = (inp[10]) ? node16270 : 4'b1011;
															assign node16270 = (inp[0]) ? node16274 : node16271;
																assign node16271 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node16274 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node16277 = (inp[15]) ? node16279 : 4'b1001;
															assign node16279 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node16282 = (inp[10]) ? node16298 : node16283;
													assign node16283 = (inp[12]) ? node16289 : node16284;
														assign node16284 = (inp[15]) ? node16286 : 4'b1001;
															assign node16286 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node16289 = (inp[15]) ? node16291 : 4'b1111;
															assign node16291 = (inp[5]) ? node16295 : node16292;
																assign node16292 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node16295 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node16298 = (inp[12]) ? node16312 : node16299;
														assign node16299 = (inp[5]) ? node16305 : node16300;
															assign node16300 = (inp[15]) ? 4'b1111 : node16301;
																assign node16301 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node16305 = (inp[0]) ? node16309 : node16306;
																assign node16306 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node16309 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node16312 = (inp[5]) ? node16314 : 4'b1101;
															assign node16314 = (inp[15]) ? node16316 : 4'b1111;
																assign node16316 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node16319 = (inp[9]) ? node16341 : node16320;
												assign node16320 = (inp[12]) ? node16330 : node16321;
													assign node16321 = (inp[10]) ? node16323 : 4'b1001;
														assign node16323 = (inp[0]) ? node16325 : 4'b1101;
															assign node16325 = (inp[15]) ? 4'b1111 : node16326;
																assign node16326 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node16330 = (inp[5]) ? node16336 : node16331;
														assign node16331 = (inp[10]) ? 4'b1101 : node16332;
															assign node16332 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node16336 = (inp[0]) ? 4'b1111 : node16337;
															assign node16337 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node16341 = (inp[10]) ? node16357 : node16342;
													assign node16342 = (inp[12]) ? node16350 : node16343;
														assign node16343 = (inp[5]) ? 4'b1101 : node16344;
															assign node16344 = (inp[15]) ? 4'b1101 : node16345;
																assign node16345 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node16350 = (inp[15]) ? node16354 : node16351;
															assign node16351 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node16354 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node16357 = (inp[0]) ? node16365 : node16358;
														assign node16358 = (inp[15]) ? node16362 : node16359;
															assign node16359 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node16362 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node16365 = (inp[15]) ? 4'b1011 : 4'b1001;
										assign node16368 = (inp[4]) ? node16398 : node16369;
											assign node16369 = (inp[9]) ? node16387 : node16370;
												assign node16370 = (inp[10]) ? node16378 : node16371;
													assign node16371 = (inp[12]) ? 4'b1001 : node16372;
														assign node16372 = (inp[15]) ? node16374 : 4'b1101;
															assign node16374 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node16378 = (inp[15]) ? node16382 : node16379;
														assign node16379 = (inp[12]) ? 4'b1001 : 4'b1011;
														assign node16382 = (inp[5]) ? node16384 : 4'b1001;
															assign node16384 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node16387 = (inp[12]) ? node16393 : node16388;
													assign node16388 = (inp[10]) ? 4'b1101 : node16389;
														assign node16389 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node16393 = (inp[5]) ? 4'b1101 : node16394;
														assign node16394 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node16398 = (inp[9]) ? node16422 : node16399;
												assign node16399 = (inp[10]) ? node16411 : node16400;
													assign node16400 = (inp[12]) ? node16406 : node16401;
														assign node16401 = (inp[0]) ? node16403 : 4'b1001;
															assign node16403 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node16406 = (inp[0]) ? 4'b1101 : node16407;
															assign node16407 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node16411 = (inp[5]) ? node16413 : 4'b1101;
														assign node16413 = (inp[12]) ? 4'b1111 : node16414;
															assign node16414 = (inp[0]) ? node16418 : node16415;
																assign node16415 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node16418 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node16422 = (inp[10]) ? node16434 : node16423;
													assign node16423 = (inp[12]) ? node16431 : node16424;
														assign node16424 = (inp[5]) ? node16426 : 4'b1111;
															assign node16426 = (inp[0]) ? 4'b1101 : node16427;
																assign node16427 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node16431 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node16434 = (inp[5]) ? 4'b1001 : node16435;
														assign node16435 = (inp[15]) ? 4'b1011 : 4'b1001;
							assign node16439 = (inp[8]) ? node16785 : node16440;
								assign node16440 = (inp[7]) ? node16596 : node16441;
									assign node16441 = (inp[12]) ? node16491 : node16442;
										assign node16442 = (inp[0]) ? node16468 : node16443;
											assign node16443 = (inp[4]) ? node16459 : node16444;
												assign node16444 = (inp[9]) ? node16454 : node16445;
													assign node16445 = (inp[15]) ? node16451 : node16446;
														assign node16446 = (inp[5]) ? node16448 : 4'b0110;
															assign node16448 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node16451 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node16454 = (inp[10]) ? 4'b0000 : node16455;
														assign node16455 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node16459 = (inp[9]) ? node16465 : node16460;
													assign node16460 = (inp[15]) ? node16462 : 4'b0010;
														assign node16462 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node16465 = (inp[15]) ? 4'b0110 : 4'b0100;
											assign node16468 = (inp[15]) ? node16482 : node16469;
												assign node16469 = (inp[3]) ? node16475 : node16470;
													assign node16470 = (inp[4]) ? node16472 : 4'b0000;
														assign node16472 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node16475 = (inp[10]) ? node16477 : 4'b0000;
														assign node16477 = (inp[4]) ? 4'b0110 : node16478;
															assign node16478 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node16482 = (inp[3]) ? 4'b0010 : node16483;
													assign node16483 = (inp[4]) ? node16487 : node16484;
														assign node16484 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node16487 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node16491 = (inp[5]) ? node16545 : node16492;
											assign node16492 = (inp[0]) ? node16512 : node16493;
												assign node16493 = (inp[15]) ? node16505 : node16494;
													assign node16494 = (inp[9]) ? node16500 : node16495;
														assign node16495 = (inp[3]) ? node16497 : 4'b0010;
															assign node16497 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node16500 = (inp[10]) ? 4'b0110 : node16501;
															assign node16501 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node16505 = (inp[10]) ? node16507 : 4'b0000;
														assign node16507 = (inp[3]) ? node16509 : 4'b0000;
															assign node16509 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node16512 = (inp[15]) ? node16530 : node16513;
													assign node16513 = (inp[9]) ? node16523 : node16514;
														assign node16514 = (inp[3]) ? 4'b0100 : node16515;
															assign node16515 = (inp[10]) ? node16519 : node16516;
																assign node16516 = (inp[4]) ? 4'b0000 : 4'b0100;
																assign node16519 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node16523 = (inp[4]) ? 4'b0010 : node16524;
															assign node16524 = (inp[10]) ? node16526 : 4'b0000;
																assign node16526 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node16530 = (inp[9]) ? node16542 : node16531;
														assign node16531 = (inp[3]) ? node16537 : node16532;
															assign node16532 = (inp[4]) ? node16534 : 4'b0110;
																assign node16534 = (inp[10]) ? 4'b0110 : 4'b0010;
															assign node16537 = (inp[10]) ? 4'b0010 : node16538;
																assign node16538 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node16542 = (inp[3]) ? 4'b0100 : 4'b0010;
											assign node16545 = (inp[9]) ? node16575 : node16546;
												assign node16546 = (inp[3]) ? node16566 : node16547;
													assign node16547 = (inp[15]) ? node16555 : node16548;
														assign node16548 = (inp[10]) ? node16552 : node16549;
															assign node16549 = (inp[4]) ? 4'b0000 : 4'b0110;
															assign node16552 = (inp[0]) ? 4'b0110 : 4'b0010;
														assign node16555 = (inp[4]) ? node16559 : node16556;
															assign node16556 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node16559 = (inp[10]) ? node16563 : node16560;
																assign node16560 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node16563 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node16566 = (inp[4]) ? node16572 : node16567;
														assign node16567 = (inp[15]) ? 4'b0000 : node16568;
															assign node16568 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node16572 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node16575 = (inp[3]) ? node16591 : node16576;
													assign node16576 = (inp[10]) ? node16584 : node16577;
														assign node16577 = (inp[4]) ? 4'b0100 : node16578;
															assign node16578 = (inp[0]) ? 4'b0000 : node16579;
																assign node16579 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node16584 = (inp[15]) ? node16588 : node16585;
															assign node16585 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node16588 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node16591 = (inp[10]) ? node16593 : 4'b0010;
														assign node16593 = (inp[15]) ? 4'b0100 : 4'b0000;
									assign node16596 = (inp[3]) ? node16694 : node16597;
										assign node16597 = (inp[4]) ? node16653 : node16598;
											assign node16598 = (inp[9]) ? node16622 : node16599;
												assign node16599 = (inp[10]) ? node16611 : node16600;
													assign node16600 = (inp[12]) ? node16606 : node16601;
														assign node16601 = (inp[0]) ? node16603 : 4'b1101;
															assign node16603 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node16606 = (inp[5]) ? 4'b1011 : node16607;
															assign node16607 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node16611 = (inp[12]) ? 4'b1001 : node16612;
														assign node16612 = (inp[5]) ? 4'b1011 : node16613;
															assign node16613 = (inp[0]) ? node16617 : node16614;
																assign node16614 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node16617 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node16622 = (inp[12]) ? node16634 : node16623;
													assign node16623 = (inp[10]) ? node16629 : node16624;
														assign node16624 = (inp[15]) ? 4'b1011 : node16625;
															assign node16625 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node16629 = (inp[15]) ? node16631 : 4'b1101;
															assign node16631 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node16634 = (inp[15]) ? node16644 : node16635;
														assign node16635 = (inp[10]) ? node16641 : node16636;
															assign node16636 = (inp[0]) ? node16638 : 4'b1111;
																assign node16638 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node16641 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node16644 = (inp[10]) ? node16646 : 4'b1101;
															assign node16646 = (inp[5]) ? node16650 : node16647;
																assign node16647 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node16650 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node16653 = (inp[9]) ? node16671 : node16654;
												assign node16654 = (inp[10]) ? node16664 : node16655;
													assign node16655 = (inp[12]) ? node16661 : node16656;
														assign node16656 = (inp[15]) ? node16658 : 4'b1011;
															assign node16658 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node16661 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node16664 = (inp[0]) ? 4'b1111 : node16665;
														assign node16665 = (inp[15]) ? node16667 : 4'b1111;
															assign node16667 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node16671 = (inp[10]) ? node16689 : node16672;
													assign node16672 = (inp[12]) ? node16680 : node16673;
														assign node16673 = (inp[0]) ? 4'b1101 : node16674;
															assign node16674 = (inp[15]) ? node16676 : 4'b1111;
																assign node16676 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node16680 = (inp[5]) ? 4'b1011 : node16681;
															assign node16681 = (inp[0]) ? node16685 : node16682;
																assign node16682 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node16685 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node16689 = (inp[5]) ? 4'b1011 : node16690;
														assign node16690 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node16694 = (inp[10]) ? node16758 : node16695;
											assign node16695 = (inp[12]) ? node16727 : node16696;
												assign node16696 = (inp[15]) ? node16714 : node16697;
													assign node16697 = (inp[0]) ? node16707 : node16698;
														assign node16698 = (inp[5]) ? node16704 : node16699;
															assign node16699 = (inp[9]) ? 4'b1011 : node16700;
																assign node16700 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node16704 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node16707 = (inp[5]) ? node16709 : 4'b1001;
															assign node16709 = (inp[4]) ? node16711 : 4'b1011;
																assign node16711 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node16714 = (inp[4]) ? node16724 : node16715;
														assign node16715 = (inp[9]) ? node16719 : node16716;
															assign node16716 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node16719 = (inp[5]) ? 4'b1001 : node16720;
																assign node16720 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node16724 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node16727 = (inp[5]) ? node16747 : node16728;
													assign node16728 = (inp[9]) ? node16740 : node16729;
														assign node16729 = (inp[4]) ? node16735 : node16730;
															assign node16730 = (inp[15]) ? node16732 : 4'b1001;
																assign node16732 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node16735 = (inp[0]) ? node16737 : 4'b1111;
																assign node16737 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node16740 = (inp[4]) ? 4'b1001 : node16741;
															assign node16741 = (inp[15]) ? 4'b1101 : node16742;
																assign node16742 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node16747 = (inp[15]) ? node16755 : node16748;
														assign node16748 = (inp[9]) ? node16752 : node16749;
															assign node16749 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node16752 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node16755 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node16758 = (inp[0]) ? node16776 : node16759;
												assign node16759 = (inp[15]) ? node16769 : node16760;
													assign node16760 = (inp[5]) ? node16764 : node16761;
														assign node16761 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node16764 = (inp[9]) ? 4'b1001 : node16765;
															assign node16765 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node16769 = (inp[9]) ? node16773 : node16770;
														assign node16770 = (inp[5]) ? 4'b1111 : 4'b1001;
														assign node16773 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node16776 = (inp[15]) ? node16778 : 4'b1011;
													assign node16778 = (inp[9]) ? node16782 : node16779;
														assign node16779 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node16782 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node16785 = (inp[7]) ? node16961 : node16786;
									assign node16786 = (inp[0]) ? node16868 : node16787;
										assign node16787 = (inp[10]) ? node16841 : node16788;
											assign node16788 = (inp[4]) ? node16814 : node16789;
												assign node16789 = (inp[15]) ? node16799 : node16790;
													assign node16790 = (inp[5]) ? node16796 : node16791;
														assign node16791 = (inp[9]) ? node16793 : 4'b1111;
															assign node16793 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node16796 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node16799 = (inp[3]) ? node16805 : node16800;
														assign node16800 = (inp[12]) ? node16802 : 4'b1101;
															assign node16802 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node16805 = (inp[5]) ? node16809 : node16806;
															assign node16806 = (inp[12]) ? 4'b1111 : 4'b1001;
															assign node16809 = (inp[12]) ? node16811 : 4'b1111;
																assign node16811 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node16814 = (inp[5]) ? node16830 : node16815;
													assign node16815 = (inp[12]) ? node16819 : node16816;
														assign node16816 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node16819 = (inp[9]) ? node16823 : node16820;
															assign node16820 = (inp[3]) ? 4'b1111 : 4'b1101;
															assign node16823 = (inp[15]) ? node16827 : node16824;
																assign node16824 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node16827 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node16830 = (inp[15]) ? node16836 : node16831;
														assign node16831 = (inp[12]) ? 4'b1101 : node16832;
															assign node16832 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node16836 = (inp[12]) ? 4'b1011 : node16837;
															assign node16837 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node16841 = (inp[9]) ? node16855 : node16842;
												assign node16842 = (inp[4]) ? node16846 : node16843;
													assign node16843 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node16846 = (inp[15]) ? node16850 : node16847;
														assign node16847 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node16850 = (inp[5]) ? 4'b1111 : node16851;
															assign node16851 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node16855 = (inp[4]) ? node16865 : node16856;
													assign node16856 = (inp[15]) ? node16860 : node16857;
														assign node16857 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node16860 = (inp[3]) ? 4'b1111 : node16861;
															assign node16861 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node16865 = (inp[5]) ? 4'b1001 : 4'b1011;
										assign node16868 = (inp[10]) ? node16932 : node16869;
											assign node16869 = (inp[3]) ? node16907 : node16870;
												assign node16870 = (inp[15]) ? node16888 : node16871;
													assign node16871 = (inp[12]) ? node16877 : node16872;
														assign node16872 = (inp[9]) ? node16874 : 4'b1001;
															assign node16874 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node16877 = (inp[5]) ? node16883 : node16878;
															assign node16878 = (inp[4]) ? node16880 : 4'b1101;
																assign node16880 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node16883 = (inp[9]) ? 4'b1111 : node16884;
																assign node16884 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node16888 = (inp[5]) ? node16894 : node16889;
														assign node16889 = (inp[4]) ? 4'b1011 : node16890;
															assign node16890 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node16894 = (inp[9]) ? node16900 : node16895;
															assign node16895 = (inp[12]) ? node16897 : 4'b1011;
																assign node16897 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node16900 = (inp[4]) ? node16904 : node16901;
																assign node16901 = (inp[12]) ? 4'b1101 : 4'b1011;
																assign node16904 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node16907 = (inp[5]) ? node16929 : node16908;
													assign node16908 = (inp[12]) ? node16916 : node16909;
														assign node16909 = (inp[9]) ? node16913 : node16910;
															assign node16910 = (inp[15]) ? 4'b1011 : 4'b1101;
															assign node16913 = (inp[15]) ? 4'b1101 : 4'b1001;
														assign node16916 = (inp[15]) ? node16922 : node16917;
															assign node16917 = (inp[9]) ? node16919 : 4'b1111;
																assign node16919 = (inp[4]) ? 4'b1011 : 4'b1111;
															assign node16922 = (inp[9]) ? node16926 : node16923;
																assign node16923 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node16926 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node16929 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node16932 = (inp[9]) ? node16948 : node16933;
												assign node16933 = (inp[4]) ? node16941 : node16934;
													assign node16934 = (inp[12]) ? 4'b1001 : node16935;
														assign node16935 = (inp[15]) ? 4'b1011 : node16936;
															assign node16936 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node16941 = (inp[12]) ? 4'b1101 : node16942;
														assign node16942 = (inp[15]) ? 4'b1101 : node16943;
															assign node16943 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node16948 = (inp[4]) ? node16954 : node16949;
													assign node16949 = (inp[5]) ? node16951 : 4'b1101;
														assign node16951 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node16954 = (inp[15]) ? node16956 : 4'b1011;
														assign node16956 = (inp[3]) ? 4'b1001 : node16957;
															assign node16957 = (inp[5]) ? 4'b1001 : 4'b1011;
									assign node16961 = (inp[12]) ? node17071 : node16962;
										assign node16962 = (inp[0]) ? node17010 : node16963;
											assign node16963 = (inp[9]) ? node16987 : node16964;
												assign node16964 = (inp[5]) ? node16974 : node16965;
													assign node16965 = (inp[4]) ? node16967 : 4'b1110;
														assign node16967 = (inp[10]) ? node16969 : 4'b1000;
															assign node16969 = (inp[15]) ? node16971 : 4'b1100;
																assign node16971 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node16974 = (inp[15]) ? node16980 : node16975;
														assign node16975 = (inp[10]) ? 4'b1100 : node16976;
															assign node16976 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node16980 = (inp[3]) ? 4'b1010 : node16981;
															assign node16981 = (inp[4]) ? 4'b1000 : node16982;
																assign node16982 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node16987 = (inp[3]) ? node17003 : node16988;
													assign node16988 = (inp[10]) ? node16994 : node16989;
														assign node16989 = (inp[4]) ? node16991 : 4'b1010;
															assign node16991 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node16994 = (inp[4]) ? node16996 : 4'b1110;
															assign node16996 = (inp[15]) ? node17000 : node16997;
																assign node16997 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node17000 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node17003 = (inp[15]) ? node17005 : 4'b1100;
														assign node17005 = (inp[4]) ? node17007 : 4'b1110;
															assign node17007 = (inp[10]) ? 4'b1010 : 4'b1110;
											assign node17010 = (inp[15]) ? node17046 : node17011;
												assign node17011 = (inp[3]) ? node17027 : node17012;
													assign node17012 = (inp[5]) ? node17020 : node17013;
														assign node17013 = (inp[4]) ? node17017 : node17014;
															assign node17014 = (inp[10]) ? 4'b1000 : 4'b1100;
															assign node17017 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node17020 = (inp[4]) ? node17022 : 4'b1100;
															assign node17022 = (inp[9]) ? node17024 : 4'b1110;
																assign node17024 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node17027 = (inp[5]) ? node17035 : node17028;
														assign node17028 = (inp[9]) ? node17030 : 4'b1110;
															assign node17030 = (inp[10]) ? node17032 : 4'b1110;
																assign node17032 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node17035 = (inp[10]) ? node17041 : node17036;
															assign node17036 = (inp[9]) ? node17038 : 4'b1110;
																assign node17038 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node17041 = (inp[9]) ? 4'b1010 : node17042;
																assign node17042 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node17046 = (inp[5]) ? node17062 : node17047;
													assign node17047 = (inp[9]) ? node17057 : node17048;
														assign node17048 = (inp[3]) ? 4'b1010 : node17049;
															assign node17049 = (inp[10]) ? node17053 : node17050;
																assign node17050 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node17053 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node17057 = (inp[3]) ? node17059 : 4'b1010;
															assign node17059 = (inp[4]) ? 4'b1000 : 4'b1010;
													assign node17062 = (inp[4]) ? node17066 : node17063;
														assign node17063 = (inp[9]) ? 4'b1100 : 4'b1110;
														assign node17066 = (inp[10]) ? 4'b1000 : node17067;
															assign node17067 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node17071 = (inp[10]) ? node17125 : node17072;
											assign node17072 = (inp[4]) ? node17096 : node17073;
												assign node17073 = (inp[9]) ? node17087 : node17074;
													assign node17074 = (inp[0]) ? node17080 : node17075;
														assign node17075 = (inp[15]) ? node17077 : 4'b1010;
															assign node17077 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node17080 = (inp[15]) ? 4'b1000 : node17081;
															assign node17081 = (inp[5]) ? node17083 : 4'b1000;
																assign node17083 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node17087 = (inp[5]) ? node17089 : 4'b1100;
														assign node17089 = (inp[15]) ? node17093 : node17090;
															assign node17090 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node17093 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node17096 = (inp[9]) ? node17112 : node17097;
													assign node17097 = (inp[0]) ? node17107 : node17098;
														assign node17098 = (inp[15]) ? node17102 : node17099;
															assign node17099 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node17102 = (inp[3]) ? 4'b1110 : node17103;
																assign node17103 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node17107 = (inp[5]) ? node17109 : 4'b1100;
															assign node17109 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node17112 = (inp[3]) ? 4'b1010 : node17113;
														assign node17113 = (inp[5]) ? node17119 : node17114;
															assign node17114 = (inp[0]) ? 4'b1000 : node17115;
																assign node17115 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node17119 = (inp[0]) ? 4'b1010 : node17120;
																assign node17120 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node17125 = (inp[9]) ? node17147 : node17126;
												assign node17126 = (inp[4]) ? node17144 : node17127;
													assign node17127 = (inp[0]) ? node17137 : node17128;
														assign node17128 = (inp[3]) ? node17132 : node17129;
															assign node17129 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node17132 = (inp[15]) ? node17134 : 4'b1000;
																assign node17134 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node17137 = (inp[15]) ? node17141 : node17138;
															assign node17138 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node17141 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node17144 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node17147 = (inp[4]) ? node17161 : node17148;
													assign node17148 = (inp[15]) ? node17156 : node17149;
														assign node17149 = (inp[0]) ? 4'b1110 : node17150;
															assign node17150 = (inp[3]) ? 4'b1100 : node17151;
																assign node17151 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node17156 = (inp[0]) ? 4'b1100 : node17157;
															assign node17157 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node17161 = (inp[5]) ? node17167 : node17162;
														assign node17162 = (inp[0]) ? node17164 : 4'b1010;
															assign node17164 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node17167 = (inp[0]) ? node17171 : node17168;
															assign node17168 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node17171 = (inp[3]) ? 4'b1000 : 4'b1010;
						assign node17174 = (inp[7]) ? node17962 : node17175;
							assign node17175 = (inp[3]) ? node17605 : node17176;
								assign node17176 = (inp[8]) ? node17382 : node17177;
									assign node17177 = (inp[2]) ? node17283 : node17178;
										assign node17178 = (inp[5]) ? node17228 : node17179;
											assign node17179 = (inp[0]) ? node17195 : node17180;
												assign node17180 = (inp[15]) ? node17188 : node17181;
													assign node17181 = (inp[4]) ? 4'b1111 : node17182;
														assign node17182 = (inp[9]) ? 4'b1111 : node17183;
															assign node17183 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node17188 = (inp[4]) ? node17190 : 4'b1101;
														assign node17190 = (inp[12]) ? node17192 : 4'b1001;
															assign node17192 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node17195 = (inp[15]) ? node17211 : node17196;
													assign node17196 = (inp[10]) ? node17204 : node17197;
														assign node17197 = (inp[9]) ? node17199 : 4'b1001;
															assign node17199 = (inp[12]) ? node17201 : 4'b1001;
																assign node17201 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node17204 = (inp[4]) ? node17208 : node17205;
															assign node17205 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node17208 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node17211 = (inp[9]) ? node17223 : node17212;
														assign node17212 = (inp[4]) ? node17218 : node17213;
															assign node17213 = (inp[10]) ? 4'b1011 : node17214;
																assign node17214 = (inp[12]) ? 4'b1011 : 4'b1111;
															assign node17218 = (inp[10]) ? 4'b1111 : node17219;
																assign node17219 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node17223 = (inp[12]) ? node17225 : 4'b1011;
															assign node17225 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node17228 = (inp[15]) ? node17256 : node17229;
												assign node17229 = (inp[4]) ? node17243 : node17230;
													assign node17230 = (inp[0]) ? node17236 : node17231;
														assign node17231 = (inp[9]) ? node17233 : 4'b1011;
															assign node17233 = (inp[12]) ? 4'b1101 : 4'b1011;
														assign node17236 = (inp[12]) ? 4'b1001 : node17237;
															assign node17237 = (inp[9]) ? 4'b1001 : node17238;
																assign node17238 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node17243 = (inp[0]) ? node17247 : node17244;
														assign node17244 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node17247 = (inp[12]) ? node17253 : node17248;
															assign node17248 = (inp[9]) ? node17250 : 4'b1001;
																assign node17250 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node17253 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node17256 = (inp[0]) ? node17272 : node17257;
													assign node17257 = (inp[9]) ? node17267 : node17258;
														assign node17258 = (inp[4]) ? node17264 : node17259;
															assign node17259 = (inp[12]) ? 4'b1001 : node17260;
																assign node17260 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node17264 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node17267 = (inp[12]) ? 4'b1111 : node17268;
															assign node17268 = (inp[10]) ? 4'b1011 : 4'b1001;
													assign node17272 = (inp[4]) ? node17274 : 4'b1101;
														assign node17274 = (inp[10]) ? node17280 : node17275;
															assign node17275 = (inp[12]) ? 4'b1101 : node17276;
																assign node17276 = (inp[9]) ? 4'b1101 : 4'b1011;
															assign node17280 = (inp[9]) ? 4'b1001 : 4'b1101;
										assign node17283 = (inp[12]) ? node17329 : node17284;
											assign node17284 = (inp[5]) ? node17298 : node17285;
												assign node17285 = (inp[15]) ? node17289 : node17286;
													assign node17286 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node17289 = (inp[0]) ? 4'b1010 : node17290;
														assign node17290 = (inp[9]) ? node17292 : 4'b1000;
															assign node17292 = (inp[10]) ? node17294 : 4'b1100;
																assign node17294 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node17298 = (inp[9]) ? node17318 : node17299;
													assign node17299 = (inp[4]) ? node17307 : node17300;
														assign node17300 = (inp[10]) ? 4'b1010 : node17301;
															assign node17301 = (inp[15]) ? node17303 : 4'b1110;
																assign node17303 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node17307 = (inp[10]) ? node17315 : node17308;
															assign node17308 = (inp[0]) ? node17312 : node17309;
																assign node17309 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node17312 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node17315 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node17318 = (inp[0]) ? node17326 : node17319;
														assign node17319 = (inp[10]) ? node17323 : node17320;
															assign node17320 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node17323 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node17326 = (inp[4]) ? 4'b1110 : 4'b1000;
											assign node17329 = (inp[5]) ? node17351 : node17330;
												assign node17330 = (inp[4]) ? node17342 : node17331;
													assign node17331 = (inp[9]) ? node17333 : 4'b1010;
														assign node17333 = (inp[10]) ? 4'b1110 : node17334;
															assign node17334 = (inp[0]) ? node17338 : node17335;
																assign node17335 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node17338 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node17342 = (inp[10]) ? node17346 : node17343;
														assign node17343 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node17346 = (inp[0]) ? node17348 : 4'b1100;
															assign node17348 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node17351 = (inp[10]) ? node17363 : node17352;
													assign node17352 = (inp[0]) ? node17354 : 4'b1010;
														assign node17354 = (inp[9]) ? node17358 : node17355;
															assign node17355 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node17358 = (inp[15]) ? 4'b1000 : node17359;
																assign node17359 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node17363 = (inp[0]) ? node17375 : node17364;
														assign node17364 = (inp[15]) ? node17368 : node17365;
															assign node17365 = (inp[9]) ? 4'b1000 : 4'b1010;
															assign node17368 = (inp[4]) ? node17372 : node17369;
																assign node17369 = (inp[9]) ? 4'b1110 : 4'b1000;
																assign node17372 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node17375 = (inp[4]) ? 4'b1100 : node17376;
															assign node17376 = (inp[9]) ? node17378 : 4'b1010;
																assign node17378 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node17382 = (inp[2]) ? node17498 : node17383;
										assign node17383 = (inp[4]) ? node17441 : node17384;
											assign node17384 = (inp[9]) ? node17412 : node17385;
												assign node17385 = (inp[10]) ? node17405 : node17386;
													assign node17386 = (inp[12]) ? node17400 : node17387;
														assign node17387 = (inp[5]) ? node17395 : node17388;
															assign node17388 = (inp[15]) ? node17392 : node17389;
																assign node17389 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node17392 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node17395 = (inp[15]) ? node17397 : 4'b1100;
																assign node17397 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node17400 = (inp[15]) ? 4'b1000 : node17401;
															assign node17401 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node17405 = (inp[15]) ? node17409 : node17406;
														assign node17406 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node17409 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node17412 = (inp[10]) ? node17424 : node17413;
													assign node17413 = (inp[12]) ? node17417 : node17414;
														assign node17414 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node17417 = (inp[15]) ? node17419 : 4'b1100;
															assign node17419 = (inp[5]) ? node17421 : 4'b1110;
																assign node17421 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node17424 = (inp[5]) ? node17434 : node17425;
														assign node17425 = (inp[12]) ? node17427 : 4'b1110;
															assign node17427 = (inp[0]) ? node17431 : node17428;
																assign node17428 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node17431 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node17434 = (inp[0]) ? node17438 : node17435;
															assign node17435 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node17438 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node17441 = (inp[9]) ? node17469 : node17442;
												assign node17442 = (inp[10]) ? node17450 : node17443;
													assign node17443 = (inp[12]) ? node17447 : node17444;
														assign node17444 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node17447 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node17450 = (inp[0]) ? node17456 : node17451;
														assign node17451 = (inp[5]) ? node17453 : 4'b1100;
															assign node17453 = (inp[12]) ? 4'b1100 : 4'b1110;
														assign node17456 = (inp[12]) ? node17464 : node17457;
															assign node17457 = (inp[15]) ? node17461 : node17458;
																assign node17458 = (inp[5]) ? 4'b1110 : 4'b1100;
																assign node17461 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node17464 = (inp[5]) ? node17466 : 4'b1110;
																assign node17466 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node17469 = (inp[12]) ? node17481 : node17470;
													assign node17470 = (inp[10]) ? node17474 : node17471;
														assign node17471 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node17474 = (inp[15]) ? 4'b1000 : node17475;
															assign node17475 = (inp[0]) ? node17477 : 4'b1000;
																assign node17477 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node17481 = (inp[10]) ? node17491 : node17482;
														assign node17482 = (inp[0]) ? node17484 : 4'b1010;
															assign node17484 = (inp[15]) ? node17488 : node17485;
																assign node17485 = (inp[5]) ? 4'b1010 : 4'b1000;
																assign node17488 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node17491 = (inp[0]) ? 4'b1010 : node17492;
															assign node17492 = (inp[15]) ? 4'b1000 : node17493;
																assign node17493 = (inp[5]) ? 4'b1000 : 4'b1010;
										assign node17498 = (inp[10]) ? node17570 : node17499;
											assign node17499 = (inp[15]) ? node17525 : node17500;
												assign node17500 = (inp[0]) ? node17516 : node17501;
													assign node17501 = (inp[12]) ? 4'b1111 : node17502;
														assign node17502 = (inp[5]) ? node17510 : node17503;
															assign node17503 = (inp[9]) ? node17507 : node17504;
																assign node17504 = (inp[4]) ? 4'b1011 : 4'b1111;
																assign node17507 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node17510 = (inp[4]) ? node17512 : 4'b1011;
																assign node17512 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node17516 = (inp[12]) ? node17518 : 4'b1001;
														assign node17518 = (inp[5]) ? node17522 : node17519;
															assign node17519 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node17522 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node17525 = (inp[0]) ? node17551 : node17526;
													assign node17526 = (inp[5]) ? node17540 : node17527;
														assign node17527 = (inp[12]) ? node17533 : node17528;
															assign node17528 = (inp[9]) ? 4'b1001 : node17529;
																assign node17529 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node17533 = (inp[4]) ? node17537 : node17534;
																assign node17534 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node17537 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node17540 = (inp[4]) ? node17546 : node17541;
															assign node17541 = (inp[9]) ? 4'b1001 : node17542;
																assign node17542 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node17546 = (inp[12]) ? 4'b1111 : node17547;
																assign node17547 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node17551 = (inp[5]) ? node17561 : node17552;
														assign node17552 = (inp[4]) ? 4'b1011 : node17553;
															assign node17553 = (inp[9]) ? node17557 : node17554;
																assign node17554 = (inp[12]) ? 4'b1011 : 4'b1111;
																assign node17557 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node17561 = (inp[12]) ? node17563 : 4'b1111;
															assign node17563 = (inp[9]) ? node17567 : node17564;
																assign node17564 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node17567 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node17570 = (inp[0]) ? node17596 : node17571;
												assign node17571 = (inp[4]) ? node17581 : node17572;
													assign node17572 = (inp[9]) ? node17576 : node17573;
														assign node17573 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node17576 = (inp[15]) ? node17578 : 4'b1101;
															assign node17578 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node17581 = (inp[9]) ? node17593 : node17582;
														assign node17582 = (inp[12]) ? node17588 : node17583;
															assign node17583 = (inp[15]) ? 4'b1101 : node17584;
																assign node17584 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node17588 = (inp[15]) ? node17590 : 4'b1101;
																assign node17590 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node17593 = (inp[12]) ? 4'b1011 : 4'b1001;
												assign node17596 = (inp[9]) ? node17602 : node17597;
													assign node17597 = (inp[12]) ? node17599 : 4'b1111;
														assign node17599 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node17602 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node17605 = (inp[2]) ? node17787 : node17606;
									assign node17606 = (inp[8]) ? node17706 : node17607;
										assign node17607 = (inp[12]) ? node17661 : node17608;
											assign node17608 = (inp[10]) ? node17632 : node17609;
												assign node17609 = (inp[9]) ? node17621 : node17610;
													assign node17610 = (inp[4]) ? node17614 : node17611;
														assign node17611 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node17614 = (inp[0]) ? 4'b1001 : node17615;
															assign node17615 = (inp[15]) ? 4'b1001 : node17616;
																assign node17616 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node17621 = (inp[4]) ? node17627 : node17622;
														assign node17622 = (inp[15]) ? node17624 : 4'b1001;
															assign node17624 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node17627 = (inp[0]) ? 4'b1111 : node17628;
															assign node17628 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node17632 = (inp[5]) ? node17648 : node17633;
													assign node17633 = (inp[15]) ? 4'b1011 : node17634;
														assign node17634 = (inp[0]) ? node17642 : node17635;
															assign node17635 = (inp[9]) ? node17639 : node17636;
																assign node17636 = (inp[4]) ? 4'b1101 : 4'b1011;
																assign node17639 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node17642 = (inp[9]) ? 4'b1111 : node17643;
																assign node17643 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node17648 = (inp[0]) ? node17658 : node17649;
														assign node17649 = (inp[15]) ? node17651 : 4'b1001;
															assign node17651 = (inp[4]) ? node17655 : node17652;
																assign node17652 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node17655 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node17658 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node17661 = (inp[0]) ? node17683 : node17662;
												assign node17662 = (inp[15]) ? node17672 : node17663;
													assign node17663 = (inp[10]) ? node17665 : 4'b1101;
														assign node17665 = (inp[4]) ? node17669 : node17666;
															assign node17666 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node17669 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node17672 = (inp[10]) ? node17674 : 4'b1011;
														assign node17674 = (inp[5]) ? node17680 : node17675;
															assign node17675 = (inp[4]) ? node17677 : 4'b1001;
																assign node17677 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node17680 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node17683 = (inp[15]) ? node17691 : node17684;
													assign node17684 = (inp[9]) ? node17688 : node17685;
														assign node17685 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node17688 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node17691 = (inp[10]) ? node17697 : node17692;
														assign node17692 = (inp[5]) ? node17694 : 4'b1101;
															assign node17694 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node17697 = (inp[9]) ? node17703 : node17698;
															assign node17698 = (inp[4]) ? 4'b1101 : node17699;
																assign node17699 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node17703 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node17706 = (inp[4]) ? node17748 : node17707;
											assign node17707 = (inp[9]) ? node17727 : node17708;
												assign node17708 = (inp[12]) ? node17720 : node17709;
													assign node17709 = (inp[10]) ? node17715 : node17710;
														assign node17710 = (inp[0]) ? 4'b1110 : node17711;
															assign node17711 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node17715 = (inp[0]) ? node17717 : 4'b1010;
															assign node17717 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node17720 = (inp[15]) ? node17722 : 4'b1010;
														assign node17722 = (inp[10]) ? 4'b1000 : node17723;
															assign node17723 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node17727 = (inp[12]) ? node17741 : node17728;
													assign node17728 = (inp[10]) ? node17736 : node17729;
														assign node17729 = (inp[0]) ? 4'b1010 : node17730;
															assign node17730 = (inp[5]) ? node17732 : 4'b1010;
																assign node17732 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node17736 = (inp[0]) ? 4'b1110 : node17737;
															assign node17737 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node17741 = (inp[0]) ? node17745 : node17742;
														assign node17742 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node17745 = (inp[10]) ? 4'b1110 : 4'b1100;
											assign node17748 = (inp[9]) ? node17770 : node17749;
												assign node17749 = (inp[12]) ? node17761 : node17750;
													assign node17750 = (inp[10]) ? node17756 : node17751;
														assign node17751 = (inp[5]) ? node17753 : 4'b1000;
															assign node17753 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node17756 = (inp[15]) ? node17758 : 4'b1100;
															assign node17758 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node17761 = (inp[5]) ? 4'b1110 : node17762;
														assign node17762 = (inp[15]) ? node17766 : node17763;
															assign node17763 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node17766 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node17770 = (inp[10]) ? node17780 : node17771;
													assign node17771 = (inp[12]) ? node17775 : node17772;
														assign node17772 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node17775 = (inp[5]) ? node17777 : 4'b1000;
															assign node17777 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node17780 = (inp[15]) ? node17784 : node17781;
														assign node17781 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node17784 = (inp[0]) ? 4'b1000 : 4'b1010;
									assign node17787 = (inp[8]) ? node17889 : node17788;
										assign node17788 = (inp[9]) ? node17836 : node17789;
											assign node17789 = (inp[4]) ? node17817 : node17790;
												assign node17790 = (inp[12]) ? node17804 : node17791;
													assign node17791 = (inp[10]) ? node17799 : node17792;
														assign node17792 = (inp[15]) ? node17794 : 4'b1100;
															assign node17794 = (inp[0]) ? node17796 : 4'b1110;
																assign node17796 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node17799 = (inp[5]) ? 4'b1000 : node17800;
															assign node17800 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node17804 = (inp[5]) ? node17810 : node17805;
														assign node17805 = (inp[0]) ? 4'b1000 : node17806;
															assign node17806 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node17810 = (inp[10]) ? 4'b1000 : node17811;
															assign node17811 = (inp[15]) ? node17813 : 4'b1010;
																assign node17813 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node17817 = (inp[12]) ? node17829 : node17818;
													assign node17818 = (inp[10]) ? node17824 : node17819;
														assign node17819 = (inp[5]) ? 4'b1000 : node17820;
															assign node17820 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node17824 = (inp[5]) ? node17826 : 4'b1100;
															assign node17826 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node17829 = (inp[0]) ? node17833 : node17830;
														assign node17830 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node17833 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node17836 = (inp[4]) ? node17868 : node17837;
												assign node17837 = (inp[12]) ? node17857 : node17838;
													assign node17838 = (inp[10]) ? node17846 : node17839;
														assign node17839 = (inp[5]) ? 4'b1000 : node17840;
															assign node17840 = (inp[0]) ? node17842 : 4'b1000;
																assign node17842 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node17846 = (inp[5]) ? node17852 : node17847;
															assign node17847 = (inp[15]) ? 4'b1110 : node17848;
																assign node17848 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node17852 = (inp[15]) ? node17854 : 4'b1110;
																assign node17854 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node17857 = (inp[10]) ? node17863 : node17858;
														assign node17858 = (inp[0]) ? node17860 : 4'b1110;
															assign node17860 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node17863 = (inp[0]) ? node17865 : 4'b1100;
															assign node17865 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node17868 = (inp[12]) ? node17878 : node17869;
													assign node17869 = (inp[10]) ? 4'b1010 : node17870;
														assign node17870 = (inp[5]) ? node17872 : 4'b1100;
															assign node17872 = (inp[15]) ? 4'b1110 : node17873;
																assign node17873 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node17878 = (inp[10]) ? node17884 : node17879;
														assign node17879 = (inp[0]) ? node17881 : 4'b1010;
															assign node17881 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node17884 = (inp[0]) ? node17886 : 4'b1000;
															assign node17886 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node17889 = (inp[15]) ? node17923 : node17890;
											assign node17890 = (inp[0]) ? node17906 : node17891;
												assign node17891 = (inp[12]) ? node17903 : node17892;
													assign node17892 = (inp[5]) ? node17894 : 4'b1101;
														assign node17894 = (inp[9]) ? 4'b1101 : node17895;
															assign node17895 = (inp[4]) ? node17899 : node17896;
																assign node17896 = (inp[10]) ? 4'b1001 : 4'b1101;
																assign node17899 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node17903 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node17906 = (inp[4]) ? node17918 : node17907;
													assign node17907 = (inp[5]) ? 4'b1111 : node17908;
														assign node17908 = (inp[9]) ? node17914 : node17909;
															assign node17909 = (inp[10]) ? 4'b1001 : node17910;
																assign node17910 = (inp[12]) ? 4'b1001 : 4'b1101;
															assign node17914 = (inp[12]) ? 4'b1111 : 4'b1001;
													assign node17918 = (inp[10]) ? node17920 : 4'b1111;
														assign node17920 = (inp[9]) ? 4'b1011 : 4'b1111;
											assign node17923 = (inp[0]) ? node17941 : node17924;
												assign node17924 = (inp[5]) ? node17934 : node17925;
													assign node17925 = (inp[9]) ? node17931 : node17926;
														assign node17926 = (inp[10]) ? node17928 : 4'b1001;
															assign node17928 = (inp[4]) ? 4'b1111 : 4'b1001;
														assign node17931 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node17934 = (inp[9]) ? 4'b1011 : node17935;
														assign node17935 = (inp[10]) ? node17937 : 4'b1011;
															assign node17937 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node17941 = (inp[5]) ? node17951 : node17942;
													assign node17942 = (inp[9]) ? node17948 : node17943;
														assign node17943 = (inp[10]) ? node17945 : 4'b1011;
															assign node17945 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node17948 = (inp[4]) ? 4'b1001 : 4'b1101;
													assign node17951 = (inp[12]) ? 4'b1001 : node17952;
														assign node17952 = (inp[10]) ? 4'b1001 : node17953;
															assign node17953 = (inp[4]) ? node17957 : node17954;
																assign node17954 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node17957 = (inp[9]) ? 4'b1101 : 4'b1001;
							assign node17962 = (inp[4]) ? node18338 : node17963;
								assign node17963 = (inp[9]) ? node18141 : node17964;
									assign node17964 = (inp[10]) ? node18056 : node17965;
										assign node17965 = (inp[12]) ? node18011 : node17966;
											assign node17966 = (inp[2]) ? node17992 : node17967;
												assign node17967 = (inp[8]) ? node17973 : node17968;
													assign node17968 = (inp[3]) ? node17970 : 4'b1110;
														assign node17970 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node17973 = (inp[3]) ? node17979 : node17974;
														assign node17974 = (inp[0]) ? node17976 : 4'b1111;
															assign node17976 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node17979 = (inp[0]) ? node17987 : node17980;
															assign node17980 = (inp[5]) ? node17984 : node17981;
																assign node17981 = (inp[15]) ? 4'b1101 : 4'b1111;
																assign node17984 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node17987 = (inp[15]) ? 4'b1101 : node17988;
																assign node17988 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node17992 = (inp[8]) ? node18002 : node17993;
													assign node17993 = (inp[0]) ? node17999 : node17994;
														assign node17994 = (inp[3]) ? 4'b1101 : node17995;
															assign node17995 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node17999 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node18002 = (inp[0]) ? node18004 : 4'b1110;
														assign node18004 = (inp[5]) ? node18006 : 4'b1100;
															assign node18006 = (inp[3]) ? node18008 : 4'b1100;
																assign node18008 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node18011 = (inp[5]) ? node18031 : node18012;
												assign node18012 = (inp[15]) ? node18022 : node18013;
													assign node18013 = (inp[0]) ? node18019 : node18014;
														assign node18014 = (inp[8]) ? 4'b1010 : node18015;
															assign node18015 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node18019 = (inp[3]) ? 4'b1000 : 4'b1001;
													assign node18022 = (inp[0]) ? 4'b1010 : node18023;
														assign node18023 = (inp[3]) ? 4'b1001 : node18024;
															assign node18024 = (inp[2]) ? node18026 : 4'b1000;
																assign node18026 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node18031 = (inp[2]) ? node18045 : node18032;
													assign node18032 = (inp[8]) ? node18038 : node18033;
														assign node18033 = (inp[3]) ? 4'b1010 : node18034;
															assign node18034 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node18038 = (inp[3]) ? node18042 : node18039;
															assign node18039 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node18042 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node18045 = (inp[8]) ? node18047 : 4'b1001;
														assign node18047 = (inp[0]) ? node18049 : 4'b1010;
															assign node18049 = (inp[15]) ? node18053 : node18050;
																assign node18050 = (inp[3]) ? 4'b1010 : 4'b1000;
																assign node18053 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node18056 = (inp[3]) ? node18090 : node18057;
											assign node18057 = (inp[8]) ? node18075 : node18058;
												assign node18058 = (inp[2]) ? node18066 : node18059;
													assign node18059 = (inp[5]) ? node18061 : 4'b1010;
														assign node18061 = (inp[0]) ? node18063 : 4'b1000;
															assign node18063 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node18066 = (inp[5]) ? node18072 : node18067;
														assign node18067 = (inp[0]) ? 4'b1011 : node18068;
															assign node18068 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node18072 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node18075 = (inp[2]) ? node18083 : node18076;
													assign node18076 = (inp[5]) ? 4'b1001 : node18077;
														assign node18077 = (inp[12]) ? node18079 : 4'b1001;
															assign node18079 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node18083 = (inp[15]) ? node18087 : node18084;
														assign node18084 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node18087 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node18090 = (inp[12]) ? node18116 : node18091;
												assign node18091 = (inp[0]) ? node18099 : node18092;
													assign node18092 = (inp[8]) ? node18096 : node18093;
														assign node18093 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node18096 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node18099 = (inp[2]) ? node18107 : node18100;
														assign node18100 = (inp[8]) ? node18102 : 4'b1010;
															assign node18102 = (inp[5]) ? 4'b1011 : node18103;
																assign node18103 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node18107 = (inp[8]) ? 4'b1010 : node18108;
															assign node18108 = (inp[5]) ? node18112 : node18109;
																assign node18109 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node18112 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node18116 = (inp[0]) ? node18130 : node18117;
													assign node18117 = (inp[8]) ? node18127 : node18118;
														assign node18118 = (inp[2]) ? node18122 : node18119;
															assign node18119 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node18122 = (inp[5]) ? node18124 : 4'b1001;
																assign node18124 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node18127 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node18130 = (inp[15]) ? node18134 : node18131;
														assign node18131 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node18134 = (inp[5]) ? 4'b1001 : node18135;
															assign node18135 = (inp[8]) ? node18137 : 4'b1011;
																assign node18137 = (inp[2]) ? 4'b1010 : 4'b1011;
									assign node18141 = (inp[10]) ? node18247 : node18142;
										assign node18142 = (inp[12]) ? node18188 : node18143;
											assign node18143 = (inp[3]) ? node18167 : node18144;
												assign node18144 = (inp[0]) ? node18156 : node18145;
													assign node18145 = (inp[15]) ? node18153 : node18146;
														assign node18146 = (inp[2]) ? node18150 : node18147;
															assign node18147 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node18150 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node18153 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node18156 = (inp[15]) ? node18162 : node18157;
														assign node18157 = (inp[2]) ? 4'b1001 : node18158;
															assign node18158 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node18162 = (inp[2]) ? node18164 : 4'b1010;
															assign node18164 = (inp[5]) ? 4'b1011 : 4'b1010;
												assign node18167 = (inp[2]) ? node18173 : node18168;
													assign node18168 = (inp[8]) ? 4'b1001 : node18169;
														assign node18169 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node18173 = (inp[8]) ? node18175 : 4'b1001;
														assign node18175 = (inp[15]) ? node18183 : node18176;
															assign node18176 = (inp[0]) ? node18180 : node18177;
																assign node18177 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node18180 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node18183 = (inp[5]) ? 4'b1010 : node18184;
																assign node18184 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node18188 = (inp[3]) ? node18222 : node18189;
												assign node18189 = (inp[5]) ? node18201 : node18190;
													assign node18190 = (inp[15]) ? node18196 : node18191;
														assign node18191 = (inp[2]) ? node18193 : 4'b1110;
															assign node18193 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node18196 = (inp[0]) ? node18198 : 4'b1101;
															assign node18198 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node18201 = (inp[0]) ? node18211 : node18202;
														assign node18202 = (inp[15]) ? 4'b1111 : node18203;
															assign node18203 = (inp[2]) ? node18207 : node18204;
																assign node18204 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node18207 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node18211 = (inp[15]) ? node18217 : node18212;
															assign node18212 = (inp[8]) ? node18214 : 4'b1111;
																assign node18214 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node18217 = (inp[2]) ? node18219 : 4'b1100;
																assign node18219 = (inp[8]) ? 4'b1100 : 4'b1101;
												assign node18222 = (inp[15]) ? node18232 : node18223;
													assign node18223 = (inp[0]) ? 4'b1111 : node18224;
														assign node18224 = (inp[2]) ? node18228 : node18225;
															assign node18225 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node18228 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node18232 = (inp[0]) ? node18242 : node18233;
														assign node18233 = (inp[5]) ? node18237 : node18234;
															assign node18234 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node18237 = (inp[8]) ? node18239 : 4'b1110;
																assign node18239 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node18242 = (inp[8]) ? node18244 : 4'b1100;
															assign node18244 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node18247 = (inp[3]) ? node18307 : node18248;
											assign node18248 = (inp[5]) ? node18276 : node18249;
												assign node18249 = (inp[0]) ? node18261 : node18250;
													assign node18250 = (inp[15]) ? node18256 : node18251;
														assign node18251 = (inp[2]) ? node18253 : 4'b1110;
															assign node18253 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node18256 = (inp[2]) ? node18258 : 4'b1100;
															assign node18258 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node18261 = (inp[15]) ? node18263 : 4'b1100;
														assign node18263 = (inp[12]) ? node18271 : node18264;
															assign node18264 = (inp[8]) ? node18268 : node18265;
																assign node18265 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node18268 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node18271 = (inp[8]) ? node18273 : 4'b1110;
																assign node18273 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node18276 = (inp[15]) ? node18288 : node18277;
													assign node18277 = (inp[0]) ? node18285 : node18278;
														assign node18278 = (inp[8]) ? node18282 : node18279;
															assign node18279 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node18282 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node18285 = (inp[12]) ? 4'b1110 : 4'b1111;
													assign node18288 = (inp[0]) ? node18300 : node18289;
														assign node18289 = (inp[12]) ? node18295 : node18290;
															assign node18290 = (inp[2]) ? node18292 : 4'b1111;
																assign node18292 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node18295 = (inp[8]) ? node18297 : 4'b1110;
																assign node18297 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node18300 = (inp[2]) ? node18304 : node18301;
															assign node18301 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node18304 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node18307 = (inp[2]) ? node18323 : node18308;
												assign node18308 = (inp[8]) ? node18316 : node18309;
													assign node18309 = (inp[15]) ? node18313 : node18310;
														assign node18310 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node18313 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node18316 = (inp[0]) ? node18320 : node18317;
														assign node18317 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node18320 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node18323 = (inp[8]) ? node18331 : node18324;
													assign node18324 = (inp[15]) ? node18328 : node18325;
														assign node18325 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node18328 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node18331 = (inp[15]) ? node18335 : node18332;
														assign node18332 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node18335 = (inp[0]) ? 4'b1100 : 4'b1110;
								assign node18338 = (inp[9]) ? node18542 : node18339;
									assign node18339 = (inp[12]) ? node18435 : node18340;
										assign node18340 = (inp[10]) ? node18384 : node18341;
											assign node18341 = (inp[8]) ? node18367 : node18342;
												assign node18342 = (inp[2]) ? node18364 : node18343;
													assign node18343 = (inp[5]) ? node18355 : node18344;
														assign node18344 = (inp[3]) ? node18350 : node18345;
															assign node18345 = (inp[0]) ? node18347 : 4'b1000;
																assign node18347 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node18350 = (inp[15]) ? 4'b1010 : node18351;
																assign node18351 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node18355 = (inp[15]) ? node18357 : 4'b1010;
															assign node18357 = (inp[0]) ? node18361 : node18358;
																assign node18358 = (inp[3]) ? 4'b1010 : 4'b1000;
																assign node18361 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node18364 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node18367 = (inp[2]) ? node18375 : node18368;
													assign node18368 = (inp[3]) ? 4'b1001 : node18369;
														assign node18369 = (inp[5]) ? node18371 : 4'b1001;
															assign node18371 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node18375 = (inp[5]) ? node18381 : node18376;
														assign node18376 = (inp[0]) ? node18378 : 4'b1000;
															assign node18378 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node18381 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node18384 = (inp[8]) ? node18408 : node18385;
												assign node18385 = (inp[2]) ? node18401 : node18386;
													assign node18386 = (inp[5]) ? node18388 : 4'b1110;
														assign node18388 = (inp[3]) ? node18396 : node18389;
															assign node18389 = (inp[15]) ? node18393 : node18390;
																assign node18390 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node18393 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node18396 = (inp[0]) ? 4'b1100 : node18397;
																assign node18397 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node18401 = (inp[15]) ? node18403 : 4'b1101;
														assign node18403 = (inp[3]) ? 4'b1101 : node18404;
															assign node18404 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node18408 = (inp[2]) ? node18422 : node18409;
													assign node18409 = (inp[3]) ? 4'b1111 : node18410;
														assign node18410 = (inp[0]) ? node18416 : node18411;
															assign node18411 = (inp[5]) ? node18413 : 4'b1101;
																assign node18413 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node18416 = (inp[15]) ? 4'b1111 : node18417;
																assign node18417 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node18422 = (inp[15]) ? 4'b1110 : node18423;
														assign node18423 = (inp[0]) ? node18429 : node18424;
															assign node18424 = (inp[5]) ? 4'b1100 : node18425;
																assign node18425 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node18429 = (inp[3]) ? 4'b1110 : node18430;
																assign node18430 = (inp[5]) ? 4'b1110 : 4'b1100;
										assign node18435 = (inp[5]) ? node18479 : node18436;
											assign node18436 = (inp[0]) ? node18458 : node18437;
												assign node18437 = (inp[15]) ? node18445 : node18438;
													assign node18438 = (inp[3]) ? 4'b1100 : node18439;
														assign node18439 = (inp[2]) ? 4'b1110 : node18440;
															assign node18440 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node18445 = (inp[3]) ? node18451 : node18446;
														assign node18446 = (inp[2]) ? 4'b1100 : node18447;
															assign node18447 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node18451 = (inp[2]) ? node18455 : node18452;
															assign node18452 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node18455 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node18458 = (inp[15]) ? node18470 : node18459;
													assign node18459 = (inp[3]) ? node18467 : node18460;
														assign node18460 = (inp[8]) ? node18464 : node18461;
															assign node18461 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node18464 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node18467 = (inp[10]) ? 4'b1110 : 4'b1111;
													assign node18470 = (inp[3]) ? node18476 : node18471;
														assign node18471 = (inp[2]) ? node18473 : 4'b1110;
															assign node18473 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node18476 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node18479 = (inp[10]) ? node18519 : node18480;
												assign node18480 = (inp[3]) ? node18498 : node18481;
													assign node18481 = (inp[0]) ? node18489 : node18482;
														assign node18482 = (inp[15]) ? node18484 : 4'b1100;
															assign node18484 = (inp[2]) ? 4'b1110 : node18485;
																assign node18485 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node18489 = (inp[15]) ? node18495 : node18490;
															assign node18490 = (inp[8]) ? node18492 : 4'b1111;
																assign node18492 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node18495 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node18498 = (inp[15]) ? node18510 : node18499;
														assign node18499 = (inp[0]) ? node18505 : node18500;
															assign node18500 = (inp[8]) ? 4'b1101 : node18501;
																assign node18501 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node18505 = (inp[8]) ? node18507 : 4'b1111;
																assign node18507 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node18510 = (inp[0]) ? node18514 : node18511;
															assign node18511 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node18514 = (inp[8]) ? node18516 : 4'b1101;
																assign node18516 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node18519 = (inp[2]) ? node18533 : node18520;
													assign node18520 = (inp[8]) ? node18528 : node18521;
														assign node18521 = (inp[0]) ? node18525 : node18522;
															assign node18522 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node18525 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node18528 = (inp[15]) ? node18530 : 4'b1101;
															assign node18530 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node18533 = (inp[8]) ? node18535 : 4'b1111;
														assign node18535 = (inp[15]) ? node18539 : node18536;
															assign node18536 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node18539 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node18542 = (inp[12]) ? node18646 : node18543;
										assign node18543 = (inp[10]) ? node18605 : node18544;
											assign node18544 = (inp[15]) ? node18574 : node18545;
												assign node18545 = (inp[0]) ? node18563 : node18546;
													assign node18546 = (inp[3]) ? node18556 : node18547;
														assign node18547 = (inp[5]) ? node18553 : node18548;
															assign node18548 = (inp[2]) ? node18550 : 4'b1110;
																assign node18550 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node18553 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node18556 = (inp[8]) ? node18560 : node18557;
															assign node18557 = (inp[2]) ? 4'b1101 : 4'b1100;
															assign node18560 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node18563 = (inp[3]) ? node18567 : node18564;
														assign node18564 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node18567 = (inp[2]) ? node18571 : node18568;
															assign node18568 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node18571 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node18574 = (inp[0]) ? node18586 : node18575;
													assign node18575 = (inp[3]) ? 4'b1110 : node18576;
														assign node18576 = (inp[5]) ? 4'b1110 : node18577;
															assign node18577 = (inp[2]) ? node18581 : node18578;
																assign node18578 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node18581 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node18586 = (inp[5]) ? node18594 : node18587;
														assign node18587 = (inp[3]) ? node18591 : node18588;
															assign node18588 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node18591 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node18594 = (inp[3]) ? node18600 : node18595;
															assign node18595 = (inp[2]) ? node18597 : 4'b1101;
																assign node18597 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node18600 = (inp[8]) ? 4'b1101 : node18601;
																assign node18601 = (inp[2]) ? 4'b1101 : 4'b1100;
											assign node18605 = (inp[8]) ? node18621 : node18606;
												assign node18606 = (inp[2]) ? node18616 : node18607;
													assign node18607 = (inp[0]) ? node18613 : node18608;
														assign node18608 = (inp[3]) ? node18610 : 4'b1010;
															assign node18610 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node18613 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node18616 = (inp[3]) ? node18618 : 4'b1001;
														assign node18618 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node18621 = (inp[2]) ? node18637 : node18622;
													assign node18622 = (inp[15]) ? node18628 : node18623;
														assign node18623 = (inp[0]) ? 4'b1011 : node18624;
															assign node18624 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node18628 = (inp[5]) ? 4'b1001 : node18629;
															assign node18629 = (inp[3]) ? node18633 : node18630;
																assign node18630 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node18633 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node18637 = (inp[15]) ? node18639 : 4'b1000;
														assign node18639 = (inp[3]) ? 4'b1010 : node18640;
															assign node18640 = (inp[5]) ? 4'b1010 : node18641;
																assign node18641 = (inp[0]) ? 4'b1010 : 4'b1000;
										assign node18646 = (inp[0]) ? node18704 : node18647;
											assign node18647 = (inp[15]) ? node18675 : node18648;
												assign node18648 = (inp[5]) ? node18660 : node18649;
													assign node18649 = (inp[3]) ? node18655 : node18650;
														assign node18650 = (inp[8]) ? 4'b1010 : node18651;
															assign node18651 = (inp[10]) ? 4'b1010 : 4'b1011;
														assign node18655 = (inp[8]) ? 4'b1000 : node18656;
															assign node18656 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node18660 = (inp[3]) ? node18670 : node18661;
														assign node18661 = (inp[10]) ? node18667 : node18662;
															assign node18662 = (inp[8]) ? node18664 : 4'b1000;
																assign node18664 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node18667 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node18670 = (inp[8]) ? 4'b1001 : node18671;
															assign node18671 = (inp[10]) ? 4'b1000 : 4'b1001;
												assign node18675 = (inp[5]) ? node18685 : node18676;
													assign node18676 = (inp[3]) ? 4'b1011 : node18677;
														assign node18677 = (inp[8]) ? node18681 : node18678;
															assign node18678 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node18681 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node18685 = (inp[10]) ? node18697 : node18686;
														assign node18686 = (inp[3]) ? node18692 : node18687;
															assign node18687 = (inp[2]) ? 4'b1011 : node18688;
																assign node18688 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node18692 = (inp[8]) ? node18694 : 4'b1011;
																assign node18694 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node18697 = (inp[2]) ? node18701 : node18698;
															assign node18698 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node18701 = (inp[8]) ? 4'b1010 : 4'b1011;
											assign node18704 = (inp[15]) ? node18720 : node18705;
												assign node18705 = (inp[3]) ? node18713 : node18706;
													assign node18706 = (inp[8]) ? node18710 : node18707;
														assign node18707 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node18710 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node18713 = (inp[8]) ? node18717 : node18714;
														assign node18714 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node18717 = (inp[2]) ? 4'b1010 : 4'b1011;
												assign node18720 = (inp[3]) ? node18732 : node18721;
													assign node18721 = (inp[5]) ? node18727 : node18722;
														assign node18722 = (inp[2]) ? node18724 : 4'b1010;
															assign node18724 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node18727 = (inp[8]) ? 4'b1000 : node18728;
															assign node18728 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node18732 = (inp[5]) ? node18738 : node18733;
														assign node18733 = (inp[8]) ? 4'b1001 : node18734;
															assign node18734 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node18738 = (inp[2]) ? node18740 : 4'b1000;
															assign node18740 = (inp[8]) ? 4'b1000 : 4'b1001;
				assign node18743 = (inp[13]) ? node21813 : node18744;
					assign node18744 = (inp[1]) ? node20392 : node18745;
						assign node18745 = (inp[15]) ? node19547 : node18746;
							assign node18746 = (inp[0]) ? node19166 : node18747;
								assign node18747 = (inp[5]) ? node18977 : node18748;
									assign node18748 = (inp[3]) ? node18854 : node18749;
										assign node18749 = (inp[12]) ? node18811 : node18750;
											assign node18750 = (inp[10]) ? node18782 : node18751;
												assign node18751 = (inp[9]) ? node18763 : node18752;
													assign node18752 = (inp[4]) ? node18758 : node18753;
														assign node18753 = (inp[8]) ? 4'b1111 : node18754;
															assign node18754 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node18758 = (inp[2]) ? 4'b1011 : node18759;
															assign node18759 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node18763 = (inp[4]) ? node18775 : node18764;
														assign node18764 = (inp[8]) ? node18770 : node18765;
															assign node18765 = (inp[7]) ? node18767 : 4'b1011;
																assign node18767 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node18770 = (inp[7]) ? node18772 : 4'b1010;
																assign node18772 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node18775 = (inp[2]) ? node18777 : 4'b1111;
															assign node18777 = (inp[8]) ? 4'b1110 : node18778;
																assign node18778 = (inp[7]) ? 4'b1111 : 4'b1110;
												assign node18782 = (inp[2]) ? node18796 : node18783;
													assign node18783 = (inp[7]) ? node18789 : node18784;
														assign node18784 = (inp[8]) ? node18786 : 4'b1111;
															assign node18786 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node18789 = (inp[8]) ? node18791 : 4'b1010;
															assign node18791 = (inp[9]) ? node18793 : 4'b1111;
																assign node18793 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node18796 = (inp[9]) ? node18804 : node18797;
														assign node18797 = (inp[4]) ? node18799 : 4'b1010;
															assign node18799 = (inp[8]) ? node18801 : 4'b1110;
																assign node18801 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node18804 = (inp[4]) ? 4'b1010 : node18805;
															assign node18805 = (inp[7]) ? node18807 : 4'b1111;
																assign node18807 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node18811 = (inp[8]) ? node18829 : node18812;
												assign node18812 = (inp[7]) ? node18824 : node18813;
													assign node18813 = (inp[2]) ? node18817 : node18814;
														assign node18814 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node18817 = (inp[4]) ? node18821 : node18818;
															assign node18818 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node18821 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node18824 = (inp[2]) ? node18826 : 4'b1110;
														assign node18826 = (inp[4]) ? 4'b1111 : 4'b1011;
												assign node18829 = (inp[7]) ? node18845 : node18830;
													assign node18830 = (inp[2]) ? node18834 : node18831;
														assign node18831 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node18834 = (inp[10]) ? node18840 : node18835;
															assign node18835 = (inp[9]) ? 4'b1111 : node18836;
																assign node18836 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node18840 = (inp[9]) ? node18842 : 4'b1111;
																assign node18842 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node18845 = (inp[2]) ? node18847 : 4'b1011;
														assign node18847 = (inp[4]) ? node18851 : node18848;
															assign node18848 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node18851 = (inp[9]) ? 4'b1010 : 4'b1110;
										assign node18854 = (inp[4]) ? node18916 : node18855;
											assign node18855 = (inp[9]) ? node18887 : node18856;
												assign node18856 = (inp[10]) ? node18874 : node18857;
													assign node18857 = (inp[12]) ? node18869 : node18858;
														assign node18858 = (inp[8]) ? node18864 : node18859;
															assign node18859 = (inp[2]) ? node18861 : 4'b1111;
																assign node18861 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node18864 = (inp[2]) ? node18866 : 4'b1110;
																assign node18866 = (inp[7]) ? 4'b1110 : 4'b1111;
														assign node18869 = (inp[2]) ? 4'b1010 : node18870;
															assign node18870 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node18874 = (inp[12]) ? node18880 : node18875;
														assign node18875 = (inp[8]) ? node18877 : 4'b1010;
															assign node18877 = (inp[2]) ? 4'b1011 : 4'b1010;
														assign node18880 = (inp[2]) ? node18882 : 4'b1011;
															assign node18882 = (inp[7]) ? node18884 : 4'b1010;
																assign node18884 = (inp[8]) ? 4'b1010 : 4'b1011;
												assign node18887 = (inp[10]) ? node18903 : node18888;
													assign node18888 = (inp[12]) ? node18900 : node18889;
														assign node18889 = (inp[7]) ? node18895 : node18890;
															assign node18890 = (inp[8]) ? 4'b1011 : node18891;
																assign node18891 = (inp[2]) ? 4'b1010 : 4'b1011;
															assign node18895 = (inp[2]) ? node18897 : 4'b1010;
																assign node18897 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node18900 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node18903 = (inp[7]) ? node18909 : node18904;
														assign node18904 = (inp[12]) ? node18906 : 4'b1100;
															assign node18906 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node18909 = (inp[12]) ? node18911 : 4'b1101;
															assign node18911 = (inp[2]) ? node18913 : 4'b1100;
																assign node18913 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node18916 = (inp[9]) ? node18956 : node18917;
												assign node18917 = (inp[10]) ? node18937 : node18918;
													assign node18918 = (inp[12]) ? node18932 : node18919;
														assign node18919 = (inp[2]) ? node18927 : node18920;
															assign node18920 = (inp[7]) ? node18924 : node18921;
																assign node18921 = (inp[8]) ? 4'b1010 : 4'b1011;
																assign node18924 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node18927 = (inp[7]) ? node18929 : 4'b1011;
																assign node18929 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node18932 = (inp[8]) ? 4'b1101 : node18933;
															assign node18933 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node18937 = (inp[7]) ? node18943 : node18938;
														assign node18938 = (inp[12]) ? 4'b1101 : node18939;
															assign node18939 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node18943 = (inp[12]) ? node18951 : node18944;
															assign node18944 = (inp[2]) ? node18948 : node18945;
																assign node18945 = (inp[8]) ? 4'b1101 : 4'b1100;
																assign node18948 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node18951 = (inp[2]) ? 4'b1100 : node18952;
																assign node18952 = (inp[8]) ? 4'b1101 : 4'b1100;
												assign node18956 = (inp[10]) ? node18968 : node18957;
													assign node18957 = (inp[12]) ? node18959 : 4'b1100;
														assign node18959 = (inp[8]) ? 4'b1000 : node18960;
															assign node18960 = (inp[7]) ? node18964 : node18961;
																assign node18961 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node18964 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node18968 = (inp[12]) ? node18970 : 4'b1001;
														assign node18970 = (inp[7]) ? node18974 : node18971;
															assign node18971 = (inp[2]) ? 4'b1001 : 4'b1000;
															assign node18974 = (inp[2]) ? 4'b1000 : 4'b1001;
									assign node18977 = (inp[3]) ? node19067 : node18978;
										assign node18978 = (inp[9]) ? node19024 : node18979;
											assign node18979 = (inp[4]) ? node18995 : node18980;
												assign node18980 = (inp[12]) ? node18988 : node18981;
													assign node18981 = (inp[10]) ? node18983 : 4'b1111;
														assign node18983 = (inp[2]) ? 4'b1011 : node18984;
															assign node18984 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node18988 = (inp[8]) ? 4'b1010 : node18989;
														assign node18989 = (inp[7]) ? 4'b1011 : node18990;
															assign node18990 = (inp[10]) ? 4'b1011 : 4'b1010;
												assign node18995 = (inp[10]) ? node19011 : node18996;
													assign node18996 = (inp[12]) ? node19004 : node18997;
														assign node18997 = (inp[2]) ? 4'b1010 : node18998;
															assign node18998 = (inp[7]) ? 4'b1010 : node18999;
																assign node18999 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node19004 = (inp[2]) ? 4'b1100 : node19005;
															assign node19005 = (inp[7]) ? 4'b1101 : node19006;
																assign node19006 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node19011 = (inp[2]) ? node19019 : node19012;
														assign node19012 = (inp[7]) ? node19016 : node19013;
															assign node19013 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node19016 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node19019 = (inp[7]) ? node19021 : 4'b1100;
															assign node19021 = (inp[8]) ? 4'b1100 : 4'b1101;
											assign node19024 = (inp[4]) ? node19046 : node19025;
												assign node19025 = (inp[10]) ? node19035 : node19026;
													assign node19026 = (inp[12]) ? node19030 : node19027;
														assign node19027 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node19030 = (inp[2]) ? node19032 : 4'b1101;
															assign node19032 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node19035 = (inp[8]) ? node19037 : 4'b1100;
														assign node19037 = (inp[12]) ? 4'b1100 : node19038;
															assign node19038 = (inp[7]) ? node19042 : node19039;
																assign node19039 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node19042 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node19046 = (inp[10]) ? node19060 : node19047;
													assign node19047 = (inp[12]) ? node19053 : node19048;
														assign node19048 = (inp[7]) ? node19050 : 4'b1101;
															assign node19050 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node19053 = (inp[7]) ? 4'b1000 : node19054;
															assign node19054 = (inp[2]) ? 4'b1000 : node19055;
																assign node19055 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node19060 = (inp[2]) ? node19062 : 4'b1001;
														assign node19062 = (inp[8]) ? 4'b1000 : node19063;
															assign node19063 = (inp[7]) ? 4'b1001 : 4'b1000;
										assign node19067 = (inp[8]) ? node19119 : node19068;
											assign node19068 = (inp[4]) ? node19104 : node19069;
												assign node19069 = (inp[9]) ? node19085 : node19070;
													assign node19070 = (inp[10]) ? node19080 : node19071;
														assign node19071 = (inp[12]) ? 4'b1001 : node19072;
															assign node19072 = (inp[2]) ? node19076 : node19073;
																assign node19073 = (inp[7]) ? 4'b1100 : 4'b1101;
																assign node19076 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node19080 = (inp[2]) ? 4'b1000 : node19081;
															assign node19081 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node19085 = (inp[10]) ? node19097 : node19086;
														assign node19086 = (inp[12]) ? node19092 : node19087;
															assign node19087 = (inp[7]) ? 4'b1000 : node19088;
																assign node19088 = (inp[2]) ? 4'b1000 : 4'b1001;
															assign node19092 = (inp[7]) ? 4'b1100 : node19093;
																assign node19093 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node19097 = (inp[2]) ? node19101 : node19098;
															assign node19098 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node19101 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node19104 = (inp[9]) ? node19110 : node19105;
													assign node19105 = (inp[10]) ? 4'b1101 : node19106;
														assign node19106 = (inp[12]) ? 4'b1100 : 4'b1000;
													assign node19110 = (inp[2]) ? node19116 : node19111;
														assign node19111 = (inp[12]) ? 4'b1001 : node19112;
															assign node19112 = (inp[7]) ? 4'b1100 : 4'b1101;
														assign node19116 = (inp[7]) ? 4'b1001 : 4'b1000;
											assign node19119 = (inp[7]) ? node19147 : node19120;
												assign node19120 = (inp[2]) ? node19136 : node19121;
													assign node19121 = (inp[12]) ? node19129 : node19122;
														assign node19122 = (inp[9]) ? 4'b1000 : node19123;
															assign node19123 = (inp[10]) ? node19125 : 4'b1000;
																assign node19125 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node19129 = (inp[4]) ? node19133 : node19130;
															assign node19130 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node19133 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node19136 = (inp[4]) ? node19142 : node19137;
														assign node19137 = (inp[9]) ? 4'b1101 : node19138;
															assign node19138 = (inp[12]) ? 4'b1001 : 4'b1101;
														assign node19142 = (inp[10]) ? 4'b1001 : node19143;
															assign node19143 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node19147 = (inp[2]) ? node19161 : node19148;
													assign node19148 = (inp[12]) ? node19154 : node19149;
														assign node19149 = (inp[9]) ? node19151 : 4'b1001;
															assign node19151 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node19154 = (inp[4]) ? node19158 : node19155;
															assign node19155 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node19158 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node19161 = (inp[4]) ? 4'b1000 : node19162;
														assign node19162 = (inp[9]) ? 4'b1100 : 4'b1000;
								assign node19166 = (inp[5]) ? node19354 : node19167;
									assign node19167 = (inp[3]) ? node19261 : node19168;
										assign node19168 = (inp[10]) ? node19212 : node19169;
											assign node19169 = (inp[4]) ? node19181 : node19170;
												assign node19170 = (inp[12]) ? node19174 : node19171;
													assign node19171 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node19174 = (inp[8]) ? 4'b1100 : node19175;
														assign node19175 = (inp[7]) ? node19177 : 4'b1101;
															assign node19177 = (inp[2]) ? 4'b1101 : 4'b1100;
												assign node19181 = (inp[7]) ? node19201 : node19182;
													assign node19182 = (inp[12]) ? node19192 : node19183;
														assign node19183 = (inp[9]) ? node19185 : 4'b1001;
															assign node19185 = (inp[8]) ? node19189 : node19186;
																assign node19186 = (inp[2]) ? 4'b1100 : 4'b1101;
																assign node19189 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node19192 = (inp[9]) ? node19196 : node19193;
															assign node19193 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node19196 = (inp[2]) ? node19198 : 4'b1001;
																assign node19198 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node19201 = (inp[9]) ? node19205 : node19202;
														assign node19202 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node19205 = (inp[12]) ? node19209 : node19206;
															assign node19206 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node19209 = (inp[8]) ? 4'b1000 : 4'b1001;
											assign node19212 = (inp[7]) ? node19232 : node19213;
												assign node19213 = (inp[4]) ? node19219 : node19214;
													assign node19214 = (inp[9]) ? 4'b1100 : node19215;
														assign node19215 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node19219 = (inp[9]) ? node19225 : node19220;
														assign node19220 = (inp[2]) ? 4'b1101 : node19221;
															assign node19221 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node19225 = (inp[2]) ? node19229 : node19226;
															assign node19226 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node19229 = (inp[8]) ? 4'b1001 : 4'b1000;
												assign node19232 = (inp[4]) ? node19250 : node19233;
													assign node19233 = (inp[9]) ? node19241 : node19234;
														assign node19234 = (inp[12]) ? 4'b1000 : node19235;
															assign node19235 = (inp[2]) ? 4'b1000 : node19236;
																assign node19236 = (inp[8]) ? 4'b1001 : 4'b1000;
														assign node19241 = (inp[12]) ? node19245 : node19242;
															assign node19242 = (inp[8]) ? 4'b1100 : 4'b1101;
															assign node19245 = (inp[8]) ? node19247 : 4'b1100;
																assign node19247 = (inp[2]) ? 4'b1100 : 4'b1101;
													assign node19250 = (inp[9]) ? node19258 : node19251;
														assign node19251 = (inp[2]) ? node19255 : node19252;
															assign node19252 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node19255 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node19258 = (inp[12]) ? 4'b1000 : 4'b1001;
										assign node19261 = (inp[4]) ? node19305 : node19262;
											assign node19262 = (inp[9]) ? node19278 : node19263;
												assign node19263 = (inp[12]) ? node19267 : node19264;
													assign node19264 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node19267 = (inp[8]) ? node19273 : node19268;
														assign node19268 = (inp[2]) ? node19270 : 4'b1000;
															assign node19270 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node19273 = (inp[7]) ? node19275 : 4'b1001;
															assign node19275 = (inp[2]) ? 4'b1000 : 4'b1001;
												assign node19278 = (inp[12]) ? node19296 : node19279;
													assign node19279 = (inp[10]) ? node19289 : node19280;
														assign node19280 = (inp[7]) ? 4'b1001 : node19281;
															assign node19281 = (inp[8]) ? node19285 : node19282;
																assign node19282 = (inp[2]) ? 4'b1000 : 4'b1001;
																assign node19285 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node19289 = (inp[8]) ? 4'b1111 : node19290;
															assign node19290 = (inp[7]) ? 4'b1110 : node19291;
																assign node19291 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node19296 = (inp[8]) ? node19298 : 4'b1111;
														assign node19298 = (inp[2]) ? node19302 : node19299;
															assign node19299 = (inp[7]) ? 4'b1111 : 4'b1110;
															assign node19302 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node19305 = (inp[9]) ? node19339 : node19306;
												assign node19306 = (inp[10]) ? node19324 : node19307;
													assign node19307 = (inp[12]) ? node19317 : node19308;
														assign node19308 = (inp[8]) ? 4'b1000 : node19309;
															assign node19309 = (inp[2]) ? node19313 : node19310;
																assign node19310 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node19313 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node19317 = (inp[2]) ? 4'b1111 : node19318;
															assign node19318 = (inp[7]) ? node19320 : 4'b1110;
																assign node19320 = (inp[8]) ? 4'b1111 : 4'b1110;
													assign node19324 = (inp[2]) ? node19332 : node19325;
														assign node19325 = (inp[12]) ? 4'b1110 : node19326;
															assign node19326 = (inp[7]) ? node19328 : 4'b1111;
																assign node19328 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node19332 = (inp[12]) ? 4'b1111 : node19333;
															assign node19333 = (inp[8]) ? node19335 : 4'b1110;
																assign node19335 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node19339 = (inp[10]) ? node19345 : node19340;
													assign node19340 = (inp[12]) ? 4'b1011 : node19341;
														assign node19341 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node19345 = (inp[7]) ? node19349 : node19346;
														assign node19346 = (inp[12]) ? 4'b1010 : 4'b1011;
														assign node19349 = (inp[2]) ? node19351 : 4'b1011;
															assign node19351 = (inp[8]) ? 4'b1010 : 4'b1011;
									assign node19354 = (inp[3]) ? node19458 : node19355;
										assign node19355 = (inp[9]) ? node19397 : node19356;
											assign node19356 = (inp[4]) ? node19376 : node19357;
												assign node19357 = (inp[12]) ? node19367 : node19358;
													assign node19358 = (inp[10]) ? 4'b1000 : node19359;
														assign node19359 = (inp[7]) ? node19361 : 4'b1100;
															assign node19361 = (inp[2]) ? node19363 : 4'b1100;
																assign node19363 = (inp[8]) ? 4'b1100 : 4'b1101;
													assign node19367 = (inp[2]) ? 4'b1000 : node19368;
														assign node19368 = (inp[10]) ? 4'b1001 : node19369;
															assign node19369 = (inp[7]) ? 4'b1000 : node19370;
																assign node19370 = (inp[8]) ? 4'b1000 : 4'b1001;
												assign node19376 = (inp[10]) ? node19388 : node19377;
													assign node19377 = (inp[12]) ? 4'b1110 : node19378;
														assign node19378 = (inp[2]) ? node19380 : 4'b1000;
															assign node19380 = (inp[8]) ? node19384 : node19381;
																assign node19381 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node19384 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node19388 = (inp[7]) ? node19390 : 4'b1110;
														assign node19390 = (inp[2]) ? node19394 : node19391;
															assign node19391 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node19394 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node19397 = (inp[4]) ? node19433 : node19398;
												assign node19398 = (inp[12]) ? node19412 : node19399;
													assign node19399 = (inp[10]) ? node19407 : node19400;
														assign node19400 = (inp[7]) ? 4'b1001 : node19401;
															assign node19401 = (inp[8]) ? node19403 : 4'b1000;
																assign node19403 = (inp[2]) ? 4'b1001 : 4'b1000;
														assign node19407 = (inp[8]) ? 4'b1111 : node19408;
															assign node19408 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node19412 = (inp[8]) ? node19424 : node19413;
														assign node19413 = (inp[10]) ? node19419 : node19414;
															assign node19414 = (inp[7]) ? 4'b1111 : node19415;
																assign node19415 = (inp[2]) ? 4'b1110 : 4'b1111;
															assign node19419 = (inp[7]) ? node19421 : 4'b1111;
																assign node19421 = (inp[2]) ? 4'b1111 : 4'b1110;
														assign node19424 = (inp[10]) ? 4'b1110 : node19425;
															assign node19425 = (inp[7]) ? node19429 : node19426;
																assign node19426 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node19429 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node19433 = (inp[10]) ? node19445 : node19434;
													assign node19434 = (inp[12]) ? node19438 : node19435;
														assign node19435 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node19438 = (inp[7]) ? 4'b1010 : node19439;
															assign node19439 = (inp[8]) ? 4'b1011 : node19440;
																assign node19440 = (inp[2]) ? 4'b1010 : 4'b1011;
													assign node19445 = (inp[8]) ? node19453 : node19446;
														assign node19446 = (inp[2]) ? node19450 : node19447;
															assign node19447 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node19450 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node19453 = (inp[2]) ? node19455 : 4'b1010;
															assign node19455 = (inp[7]) ? 4'b1010 : 4'b1011;
										assign node19458 = (inp[9]) ? node19498 : node19459;
											assign node19459 = (inp[4]) ? node19469 : node19460;
												assign node19460 = (inp[10]) ? node19466 : node19461;
													assign node19461 = (inp[12]) ? 4'b1010 : node19462;
														assign node19462 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node19466 = (inp[7]) ? 4'b1011 : 4'b1010;
												assign node19469 = (inp[10]) ? node19483 : node19470;
													assign node19470 = (inp[12]) ? node19478 : node19471;
														assign node19471 = (inp[8]) ? node19473 : 4'b1011;
															assign node19473 = (inp[2]) ? node19475 : 4'b1010;
																assign node19475 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node19478 = (inp[2]) ? 4'b1111 : node19479;
															assign node19479 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node19483 = (inp[7]) ? node19487 : node19484;
														assign node19484 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node19487 = (inp[12]) ? node19493 : node19488;
															assign node19488 = (inp[8]) ? 4'b1110 : node19489;
																assign node19489 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node19493 = (inp[2]) ? 4'b1111 : node19494;
																assign node19494 = (inp[8]) ? 4'b1111 : 4'b1110;
											assign node19498 = (inp[4]) ? node19516 : node19499;
												assign node19499 = (inp[12]) ? node19509 : node19500;
													assign node19500 = (inp[10]) ? 4'b1110 : node19501;
														assign node19501 = (inp[8]) ? 4'b1011 : node19502;
															assign node19502 = (inp[2]) ? node19504 : 4'b1010;
																assign node19504 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node19509 = (inp[8]) ? node19511 : 4'b1111;
														assign node19511 = (inp[2]) ? node19513 : 4'b1111;
															assign node19513 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node19516 = (inp[10]) ? node19530 : node19517;
													assign node19517 = (inp[12]) ? node19525 : node19518;
														assign node19518 = (inp[8]) ? node19522 : node19519;
															assign node19519 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node19522 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node19525 = (inp[8]) ? 4'b1011 : node19526;
															assign node19526 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node19530 = (inp[12]) ? node19538 : node19531;
														assign node19531 = (inp[7]) ? 4'b1011 : node19532;
															assign node19532 = (inp[8]) ? 4'b1011 : node19533;
																assign node19533 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node19538 = (inp[8]) ? 4'b1010 : node19539;
															assign node19539 = (inp[7]) ? node19543 : node19540;
																assign node19540 = (inp[2]) ? 4'b1010 : 4'b1011;
																assign node19543 = (inp[2]) ? 4'b1011 : 4'b1010;
							assign node19547 = (inp[10]) ? node19991 : node19548;
								assign node19548 = (inp[12]) ? node19774 : node19549;
									assign node19549 = (inp[0]) ? node19671 : node19550;
										assign node19550 = (inp[5]) ? node19614 : node19551;
											assign node19551 = (inp[4]) ? node19581 : node19552;
												assign node19552 = (inp[9]) ? node19568 : node19553;
													assign node19553 = (inp[3]) ? node19563 : node19554;
														assign node19554 = (inp[7]) ? 4'b1100 : node19555;
															assign node19555 = (inp[2]) ? node19559 : node19556;
																assign node19556 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node19559 = (inp[8]) ? 4'b1101 : 4'b1100;
														assign node19563 = (inp[2]) ? node19565 : 4'b1101;
															assign node19565 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node19568 = (inp[8]) ? node19574 : node19569;
														assign node19569 = (inp[3]) ? node19571 : 4'b1000;
															assign node19571 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node19574 = (inp[3]) ? node19576 : 4'b1001;
															assign node19576 = (inp[7]) ? 4'b1000 : node19577;
																assign node19577 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node19581 = (inp[9]) ? node19605 : node19582;
													assign node19582 = (inp[2]) ? node19598 : node19583;
														assign node19583 = (inp[3]) ? node19591 : node19584;
															assign node19584 = (inp[8]) ? node19588 : node19585;
																assign node19585 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node19588 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node19591 = (inp[8]) ? node19595 : node19592;
																assign node19592 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node19595 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node19598 = (inp[8]) ? node19602 : node19599;
															assign node19599 = (inp[7]) ? 4'b1001 : 4'b1000;
															assign node19602 = (inp[7]) ? 4'b1000 : 4'b1001;
													assign node19605 = (inp[3]) ? node19611 : node19606;
														assign node19606 = (inp[2]) ? node19608 : 4'b1101;
															assign node19608 = (inp[8]) ? 4'b1100 : 4'b1101;
														assign node19611 = (inp[8]) ? 4'b1110 : 4'b1111;
											assign node19614 = (inp[3]) ? node19642 : node19615;
												assign node19615 = (inp[9]) ? node19631 : node19616;
													assign node19616 = (inp[4]) ? node19624 : node19617;
														assign node19617 = (inp[8]) ? 4'b1100 : node19618;
															assign node19618 = (inp[7]) ? 4'b1101 : node19619;
																assign node19619 = (inp[2]) ? 4'b1100 : 4'b1101;
														assign node19624 = (inp[8]) ? 4'b1000 : node19625;
															assign node19625 = (inp[7]) ? 4'b1000 : node19626;
																assign node19626 = (inp[2]) ? 4'b1000 : 4'b1001;
													assign node19631 = (inp[4]) ? node19633 : 4'b1001;
														assign node19633 = (inp[2]) ? node19635 : 4'b1111;
															assign node19635 = (inp[8]) ? node19639 : node19636;
																assign node19636 = (inp[7]) ? 4'b1111 : 4'b1110;
																assign node19639 = (inp[7]) ? 4'b1110 : 4'b1111;
												assign node19642 = (inp[4]) ? node19652 : node19643;
													assign node19643 = (inp[9]) ? node19645 : 4'b1111;
														assign node19645 = (inp[2]) ? 4'b1010 : node19646;
															assign node19646 = (inp[7]) ? node19648 : 4'b1011;
																assign node19648 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node19652 = (inp[9]) ? node19662 : node19653;
														assign node19653 = (inp[2]) ? node19655 : 4'b1010;
															assign node19655 = (inp[7]) ? node19659 : node19656;
																assign node19656 = (inp[8]) ? 4'b1011 : 4'b1010;
																assign node19659 = (inp[8]) ? 4'b1010 : 4'b1011;
														assign node19662 = (inp[2]) ? 4'b1111 : node19663;
															assign node19663 = (inp[8]) ? node19667 : node19664;
																assign node19664 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node19667 = (inp[7]) ? 4'b1111 : 4'b1110;
										assign node19671 = (inp[5]) ? node19721 : node19672;
											assign node19672 = (inp[3]) ? node19690 : node19673;
												assign node19673 = (inp[2]) ? node19683 : node19674;
													assign node19674 = (inp[7]) ? 4'b1011 : node19675;
														assign node19675 = (inp[8]) ? node19677 : 4'b1011;
															assign node19677 = (inp[9]) ? node19679 : 4'b1010;
																assign node19679 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node19683 = (inp[4]) ? 4'b1111 : node19684;
														assign node19684 = (inp[9]) ? 4'b1010 : node19685;
															assign node19685 = (inp[8]) ? 4'b1110 : 4'b1111;
												assign node19690 = (inp[9]) ? node19710 : node19691;
													assign node19691 = (inp[4]) ? node19705 : node19692;
														assign node19692 = (inp[2]) ? node19700 : node19693;
															assign node19693 = (inp[7]) ? node19697 : node19694;
																assign node19694 = (inp[8]) ? 4'b1110 : 4'b1111;
																assign node19697 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node19700 = (inp[8]) ? 4'b1111 : node19701;
																assign node19701 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node19705 = (inp[8]) ? 4'b1011 : node19706;
															assign node19706 = (inp[7]) ? 4'b1011 : 4'b1010;
													assign node19710 = (inp[4]) ? node19712 : 4'b1011;
														assign node19712 = (inp[2]) ? node19714 : 4'b1101;
															assign node19714 = (inp[8]) ? node19718 : node19715;
																assign node19715 = (inp[7]) ? 4'b1101 : 4'b1100;
																assign node19718 = (inp[7]) ? 4'b1100 : 4'b1101;
											assign node19721 = (inp[3]) ? node19751 : node19722;
												assign node19722 = (inp[4]) ? node19740 : node19723;
													assign node19723 = (inp[9]) ? node19733 : node19724;
														assign node19724 = (inp[8]) ? 4'b1111 : node19725;
															assign node19725 = (inp[2]) ? node19729 : node19726;
																assign node19726 = (inp[7]) ? 4'b1110 : 4'b1111;
																assign node19729 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node19733 = (inp[2]) ? 4'b1010 : node19734;
															assign node19734 = (inp[8]) ? 4'b1011 : node19735;
																assign node19735 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node19740 = (inp[9]) ? node19744 : node19741;
														assign node19741 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node19744 = (inp[8]) ? 4'b1100 : node19745;
															assign node19745 = (inp[2]) ? 4'b1100 : node19746;
																assign node19746 = (inp[7]) ? 4'b1100 : 4'b1101;
												assign node19751 = (inp[9]) ? node19763 : node19752;
													assign node19752 = (inp[4]) ? node19754 : 4'b1100;
														assign node19754 = (inp[2]) ? 4'b1000 : node19755;
															assign node19755 = (inp[8]) ? node19759 : node19756;
																assign node19756 = (inp[7]) ? 4'b1000 : 4'b1001;
																assign node19759 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node19763 = (inp[4]) ? node19771 : node19764;
														assign node19764 = (inp[2]) ? 4'b1001 : node19765;
															assign node19765 = (inp[8]) ? node19767 : 4'b1001;
																assign node19767 = (inp[7]) ? 4'b1001 : 4'b1000;
														assign node19771 = (inp[7]) ? 4'b1101 : 4'b1100;
									assign node19774 = (inp[7]) ? node19876 : node19775;
										assign node19775 = (inp[5]) ? node19845 : node19776;
											assign node19776 = (inp[0]) ? node19814 : node19777;
												assign node19777 = (inp[3]) ? node19799 : node19778;
													assign node19778 = (inp[4]) ? node19786 : node19779;
														assign node19779 = (inp[9]) ? 4'b1100 : node19780;
															assign node19780 = (inp[2]) ? 4'b1001 : node19781;
																assign node19781 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node19786 = (inp[9]) ? node19794 : node19787;
															assign node19787 = (inp[2]) ? node19791 : node19788;
																assign node19788 = (inp[8]) ? 4'b1100 : 4'b1101;
																assign node19791 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node19794 = (inp[2]) ? node19796 : 4'b1001;
																assign node19796 = (inp[8]) ? 4'b1001 : 4'b1000;
													assign node19799 = (inp[9]) ? node19807 : node19800;
														assign node19800 = (inp[4]) ? 4'b1111 : node19801;
															assign node19801 = (inp[8]) ? 4'b1000 : node19802;
																assign node19802 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node19807 = (inp[4]) ? node19811 : node19808;
															assign node19808 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node19811 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node19814 = (inp[3]) ? node19826 : node19815;
													assign node19815 = (inp[8]) ? node19823 : node19816;
														assign node19816 = (inp[2]) ? 4'b1010 : node19817;
															assign node19817 = (inp[9]) ? 4'b1111 : node19818;
																assign node19818 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node19823 = (inp[2]) ? 4'b1011 : 4'b1010;
													assign node19826 = (inp[9]) ? node19834 : node19827;
														assign node19827 = (inp[4]) ? node19829 : 4'b1011;
															assign node19829 = (inp[8]) ? node19831 : 4'b1101;
																assign node19831 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node19834 = (inp[4]) ? node19838 : node19835;
															assign node19835 = (inp[8]) ? 4'b1101 : 4'b1100;
															assign node19838 = (inp[2]) ? node19842 : node19839;
																assign node19839 = (inp[8]) ? 4'b1000 : 4'b1001;
																assign node19842 = (inp[8]) ? 4'b1001 : 4'b1000;
											assign node19845 = (inp[0]) ? node19859 : node19846;
												assign node19846 = (inp[8]) ? node19854 : node19847;
													assign node19847 = (inp[2]) ? node19849 : 4'b1111;
														assign node19849 = (inp[9]) ? 4'b1110 : node19850;
															assign node19850 = (inp[4]) ? 4'b1110 : 4'b1000;
													assign node19854 = (inp[9]) ? 4'b1111 : node19855;
														assign node19855 = (inp[4]) ? 4'b1111 : 4'b1001;
												assign node19859 = (inp[9]) ? node19871 : node19860;
													assign node19860 = (inp[4]) ? node19868 : node19861;
														assign node19861 = (inp[2]) ? node19865 : node19862;
															assign node19862 = (inp[8]) ? 4'b1000 : 4'b1001;
															assign node19865 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node19868 = (inp[2]) ? 4'b1101 : 4'b1100;
													assign node19871 = (inp[8]) ? 4'b1101 : node19872;
														assign node19872 = (inp[2]) ? 4'b1100 : 4'b1101;
										assign node19876 = (inp[8]) ? node19934 : node19877;
											assign node19877 = (inp[2]) ? node19897 : node19878;
												assign node19878 = (inp[9]) ? node19886 : node19879;
													assign node19879 = (inp[4]) ? node19881 : 4'b1010;
														assign node19881 = (inp[5]) ? node19883 : 4'b1110;
															assign node19883 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node19886 = (inp[4]) ? node19892 : node19887;
														assign node19887 = (inp[0]) ? 4'b1100 : node19888;
															assign node19888 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node19892 = (inp[5]) ? 4'b1010 : node19893;
															assign node19893 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node19897 = (inp[3]) ? node19919 : node19898;
													assign node19898 = (inp[0]) ? node19912 : node19899;
														assign node19899 = (inp[5]) ? node19905 : node19900;
															assign node19900 = (inp[4]) ? node19902 : 4'b1101;
																assign node19902 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node19905 = (inp[9]) ? node19909 : node19906;
																assign node19906 = (inp[4]) ? 4'b1111 : 4'b1001;
																assign node19909 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node19912 = (inp[5]) ? node19916 : node19913;
															assign node19913 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node19916 = (inp[9]) ? 4'b1001 : 4'b1011;
													assign node19919 = (inp[5]) ? node19927 : node19920;
														assign node19920 = (inp[9]) ? node19924 : node19921;
															assign node19921 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node19924 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node19927 = (inp[0]) ? node19929 : 4'b1011;
															assign node19929 = (inp[9]) ? 4'b1001 : node19930;
																assign node19930 = (inp[4]) ? 4'b1101 : 4'b1001;
											assign node19934 = (inp[2]) ? node19968 : node19935;
												assign node19935 = (inp[0]) ? node19951 : node19936;
													assign node19936 = (inp[3]) ? node19944 : node19937;
														assign node19937 = (inp[9]) ? node19941 : node19938;
															assign node19938 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node19941 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node19944 = (inp[9]) ? node19948 : node19945;
															assign node19945 = (inp[4]) ? 4'b1111 : 4'b1001;
															assign node19948 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node19951 = (inp[3]) ? node19959 : node19952;
														assign node19952 = (inp[5]) ? 4'b1101 : node19953;
															assign node19953 = (inp[9]) ? 4'b1011 : node19954;
																assign node19954 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node19959 = (inp[9]) ? node19965 : node19960;
															assign node19960 = (inp[4]) ? 4'b1101 : node19961;
																assign node19961 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node19965 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node19968 = (inp[5]) ? node19986 : node19969;
													assign node19969 = (inp[0]) ? node19977 : node19970;
														assign node19970 = (inp[3]) ? 4'b1110 : node19971;
															assign node19971 = (inp[9]) ? 4'b1100 : node19972;
																assign node19972 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node19977 = (inp[3]) ? node19983 : node19978;
															assign node19978 = (inp[9]) ? node19980 : 4'b1110;
																assign node19980 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node19983 = (inp[9]) ? 4'b1100 : 4'b1010;
													assign node19986 = (inp[4]) ? node19988 : 4'b1010;
														assign node19988 = (inp[0]) ? 4'b1100 : 4'b1010;
								assign node19991 = (inp[0]) ? node20213 : node19992;
									assign node19992 = (inp[5]) ? node20112 : node19993;
										assign node19993 = (inp[3]) ? node20049 : node19994;
											assign node19994 = (inp[12]) ? node20018 : node19995;
												assign node19995 = (inp[8]) ? node20013 : node19996;
													assign node19996 = (inp[2]) ? node20010 : node19997;
														assign node19997 = (inp[7]) ? node20005 : node19998;
															assign node19998 = (inp[9]) ? node20002 : node19999;
																assign node19999 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node20002 = (inp[4]) ? 4'b1001 : 4'b1101;
															assign node20005 = (inp[9]) ? node20007 : 4'b1000;
																assign node20007 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node20010 = (inp[7]) ? 4'b1101 : 4'b1100;
													assign node20013 = (inp[2]) ? 4'b1001 : node20014;
														assign node20014 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node20018 = (inp[8]) ? node20036 : node20019;
													assign node20019 = (inp[4]) ? node20027 : node20020;
														assign node20020 = (inp[2]) ? node20024 : node20021;
															assign node20021 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node20024 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node20027 = (inp[9]) ? node20033 : node20028;
															assign node20028 = (inp[2]) ? 4'b1100 : node20029;
																assign node20029 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node20033 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node20036 = (inp[7]) ? node20044 : node20037;
														assign node20037 = (inp[2]) ? 4'b1101 : node20038;
															assign node20038 = (inp[4]) ? 4'b1100 : node20039;
																assign node20039 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node20044 = (inp[9]) ? node20046 : 4'b1000;
															assign node20046 = (inp[4]) ? 4'b1000 : 4'b1100;
											assign node20049 = (inp[4]) ? node20083 : node20050;
												assign node20050 = (inp[9]) ? node20068 : node20051;
													assign node20051 = (inp[12]) ? node20061 : node20052;
														assign node20052 = (inp[2]) ? node20054 : 4'b1001;
															assign node20054 = (inp[7]) ? node20058 : node20055;
																assign node20055 = (inp[8]) ? 4'b1001 : 4'b1000;
																assign node20058 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node20061 = (inp[7]) ? 4'b1000 : node20062;
															assign node20062 = (inp[8]) ? node20064 : 4'b1001;
																assign node20064 = (inp[2]) ? 4'b1001 : 4'b1000;
													assign node20068 = (inp[12]) ? node20074 : node20069;
														assign node20069 = (inp[2]) ? 4'b1110 : node20070;
															assign node20070 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node20074 = (inp[7]) ? node20076 : 4'b1111;
															assign node20076 = (inp[8]) ? node20080 : node20077;
																assign node20077 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node20080 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node20083 = (inp[9]) ? node20099 : node20084;
													assign node20084 = (inp[7]) ? node20092 : node20085;
														assign node20085 = (inp[2]) ? node20089 : node20086;
															assign node20086 = (inp[8]) ? 4'b1110 : 4'b1111;
															assign node20089 = (inp[8]) ? 4'b1111 : 4'b1110;
														assign node20092 = (inp[2]) ? node20096 : node20093;
															assign node20093 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node20096 = (inp[8]) ? 4'b1110 : 4'b1111;
													assign node20099 = (inp[2]) ? node20105 : node20100;
														assign node20100 = (inp[7]) ? node20102 : 4'b1010;
															assign node20102 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node20105 = (inp[8]) ? node20109 : node20106;
															assign node20106 = (inp[12]) ? 4'b1010 : 4'b1011;
															assign node20109 = (inp[12]) ? 4'b1011 : 4'b1010;
										assign node20112 = (inp[4]) ? node20164 : node20113;
											assign node20113 = (inp[9]) ? node20143 : node20114;
												assign node20114 = (inp[3]) ? node20128 : node20115;
													assign node20115 = (inp[8]) ? node20121 : node20116;
														assign node20116 = (inp[7]) ? 4'b1001 : node20117;
															assign node20117 = (inp[2]) ? 4'b1000 : 4'b1001;
														assign node20121 = (inp[12]) ? node20125 : node20122;
															assign node20122 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node20125 = (inp[7]) ? 4'b1001 : 4'b1000;
													assign node20128 = (inp[12]) ? node20138 : node20129;
														assign node20129 = (inp[2]) ? node20131 : 4'b1011;
															assign node20131 = (inp[8]) ? node20135 : node20132;
																assign node20132 = (inp[7]) ? 4'b1011 : 4'b1010;
																assign node20135 = (inp[7]) ? 4'b1010 : 4'b1011;
														assign node20138 = (inp[2]) ? 4'b1010 : node20139;
															assign node20139 = (inp[8]) ? 4'b1011 : 4'b1010;
												assign node20143 = (inp[3]) ? node20155 : node20144;
													assign node20144 = (inp[12]) ? node20146 : 4'b1111;
														assign node20146 = (inp[8]) ? node20148 : 4'b1111;
															assign node20148 = (inp[7]) ? node20152 : node20149;
																assign node20149 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node20152 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node20155 = (inp[8]) ? 4'b1111 : node20156;
														assign node20156 = (inp[12]) ? 4'b1111 : node20157;
															assign node20157 = (inp[2]) ? 4'b1110 : node20158;
																assign node20158 = (inp[7]) ? 4'b1110 : 4'b1111;
											assign node20164 = (inp[9]) ? node20198 : node20165;
												assign node20165 = (inp[3]) ? node20185 : node20166;
													assign node20166 = (inp[7]) ? node20172 : node20167;
														assign node20167 = (inp[12]) ? node20169 : 4'b1110;
															assign node20169 = (inp[8]) ? 4'b1110 : 4'b1111;
														assign node20172 = (inp[12]) ? node20178 : node20173;
															assign node20173 = (inp[2]) ? 4'b1111 : node20174;
																assign node20174 = (inp[8]) ? 4'b1111 : 4'b1110;
															assign node20178 = (inp[8]) ? node20182 : node20179;
																assign node20179 = (inp[2]) ? 4'b1111 : 4'b1110;
																assign node20182 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node20185 = (inp[8]) ? node20191 : node20186;
														assign node20186 = (inp[2]) ? node20188 : 4'b1111;
															assign node20188 = (inp[7]) ? 4'b1111 : 4'b1110;
														assign node20191 = (inp[7]) ? node20195 : node20192;
															assign node20192 = (inp[2]) ? 4'b1111 : 4'b1110;
															assign node20195 = (inp[2]) ? 4'b1110 : 4'b1111;
												assign node20198 = (inp[7]) ? node20204 : node20199;
													assign node20199 = (inp[8]) ? node20201 : 4'b1011;
														assign node20201 = (inp[3]) ? 4'b1010 : 4'b1011;
													assign node20204 = (inp[3]) ? 4'b1010 : node20205;
														assign node20205 = (inp[2]) ? node20209 : node20206;
															assign node20206 = (inp[8]) ? 4'b1011 : 4'b1010;
															assign node20209 = (inp[8]) ? 4'b1010 : 4'b1011;
									assign node20213 = (inp[3]) ? node20311 : node20214;
										assign node20214 = (inp[5]) ? node20258 : node20215;
											assign node20215 = (inp[8]) ? node20235 : node20216;
												assign node20216 = (inp[4]) ? node20230 : node20217;
													assign node20217 = (inp[9]) ? node20225 : node20218;
														assign node20218 = (inp[2]) ? node20222 : node20219;
															assign node20219 = (inp[7]) ? 4'b1010 : 4'b1011;
															assign node20222 = (inp[7]) ? 4'b1011 : 4'b1010;
														assign node20225 = (inp[7]) ? 4'b1110 : node20226;
															assign node20226 = (inp[2]) ? 4'b1110 : 4'b1111;
													assign node20230 = (inp[9]) ? node20232 : 4'b1110;
														assign node20232 = (inp[2]) ? 4'b1011 : 4'b1010;
												assign node20235 = (inp[4]) ? node20247 : node20236;
													assign node20236 = (inp[9]) ? node20242 : node20237;
														assign node20237 = (inp[7]) ? node20239 : 4'b1010;
															assign node20239 = (inp[2]) ? 4'b1010 : 4'b1011;
														assign node20242 = (inp[2]) ? 4'b1111 : node20243;
															assign node20243 = (inp[7]) ? 4'b1111 : 4'b1110;
													assign node20247 = (inp[9]) ? node20253 : node20248;
														assign node20248 = (inp[12]) ? node20250 : 4'b1111;
															assign node20250 = (inp[2]) ? 4'b1110 : 4'b1111;
														assign node20253 = (inp[7]) ? node20255 : 4'b1011;
															assign node20255 = (inp[2]) ? 4'b1010 : 4'b1011;
											assign node20258 = (inp[9]) ? node20286 : node20259;
												assign node20259 = (inp[4]) ? node20277 : node20260;
													assign node20260 = (inp[12]) ? node20266 : node20261;
														assign node20261 = (inp[7]) ? 4'b1011 : node20262;
															assign node20262 = (inp[8]) ? 4'b1011 : 4'b1010;
														assign node20266 = (inp[8]) ? node20272 : node20267;
															assign node20267 = (inp[7]) ? node20269 : 4'b1011;
																assign node20269 = (inp[2]) ? 4'b1011 : 4'b1010;
															assign node20272 = (inp[2]) ? node20274 : 4'b1010;
																assign node20274 = (inp[7]) ? 4'b1010 : 4'b1011;
													assign node20277 = (inp[2]) ? 4'b1101 : node20278;
														assign node20278 = (inp[12]) ? node20280 : 4'b1100;
															assign node20280 = (inp[8]) ? node20282 : 4'b1101;
																assign node20282 = (inp[7]) ? 4'b1101 : 4'b1100;
												assign node20286 = (inp[4]) ? node20296 : node20287;
													assign node20287 = (inp[2]) ? node20289 : 4'b1100;
														assign node20289 = (inp[12]) ? node20291 : 4'b1101;
															assign node20291 = (inp[7]) ? 4'b1100 : node20292;
																assign node20292 = (inp[8]) ? 4'b1101 : 4'b1100;
													assign node20296 = (inp[12]) ? node20298 : 4'b1000;
														assign node20298 = (inp[2]) ? node20304 : node20299;
															assign node20299 = (inp[8]) ? 4'b1000 : node20300;
																assign node20300 = (inp[7]) ? 4'b1000 : 4'b1001;
															assign node20304 = (inp[8]) ? node20308 : node20305;
																assign node20305 = (inp[7]) ? 4'b1001 : 4'b1000;
																assign node20308 = (inp[7]) ? 4'b1000 : 4'b1001;
										assign node20311 = (inp[9]) ? node20347 : node20312;
											assign node20312 = (inp[4]) ? node20330 : node20313;
												assign node20313 = (inp[5]) ? node20327 : node20314;
													assign node20314 = (inp[2]) ? node20320 : node20315;
														assign node20315 = (inp[7]) ? node20317 : 4'b1010;
															assign node20317 = (inp[12]) ? 4'b1010 : 4'b1011;
														assign node20320 = (inp[12]) ? 4'b1011 : node20321;
															assign node20321 = (inp[7]) ? 4'b1011 : node20322;
																assign node20322 = (inp[8]) ? 4'b1011 : 4'b1010;
													assign node20327 = (inp[2]) ? 4'b1001 : 4'b1000;
												assign node20330 = (inp[12]) ? node20336 : node20331;
													assign node20331 = (inp[5]) ? 4'b1101 : node20332;
														assign node20332 = (inp[7]) ? 4'b1100 : 4'b1101;
													assign node20336 = (inp[8]) ? node20342 : node20337;
														assign node20337 = (inp[7]) ? node20339 : 4'b1101;
															assign node20339 = (inp[2]) ? 4'b1101 : 4'b1100;
														assign node20342 = (inp[7]) ? node20344 : 4'b1100;
															assign node20344 = (inp[2]) ? 4'b1100 : 4'b1101;
											assign node20347 = (inp[4]) ? node20377 : node20348;
												assign node20348 = (inp[8]) ? node20362 : node20349;
													assign node20349 = (inp[12]) ? node20357 : node20350;
														assign node20350 = (inp[2]) ? node20354 : node20351;
															assign node20351 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node20354 = (inp[7]) ? 4'b1101 : 4'b1100;
														assign node20357 = (inp[7]) ? 4'b1101 : node20358;
															assign node20358 = (inp[5]) ? 4'b1101 : 4'b1100;
													assign node20362 = (inp[12]) ? 4'b1100 : node20363;
														assign node20363 = (inp[5]) ? node20369 : node20364;
															assign node20364 = (inp[2]) ? node20366 : 4'b1100;
																assign node20366 = (inp[7]) ? 4'b1100 : 4'b1101;
															assign node20369 = (inp[7]) ? node20373 : node20370;
																assign node20370 = (inp[2]) ? 4'b1101 : 4'b1100;
																assign node20373 = (inp[2]) ? 4'b1100 : 4'b1101;
												assign node20377 = (inp[2]) ? node20383 : node20378;
													assign node20378 = (inp[7]) ? 4'b1001 : node20379;
														assign node20379 = (inp[8]) ? 4'b1000 : 4'b1001;
													assign node20383 = (inp[5]) ? node20387 : node20384;
														assign node20384 = (inp[8]) ? 4'b1000 : 4'b1001;
														assign node20387 = (inp[7]) ? 4'b1000 : node20388;
															assign node20388 = (inp[8]) ? 4'b1001 : 4'b1000;
						assign node20392 = (inp[7]) ? node21070 : node20393;
							assign node20393 = (inp[8]) ? node20763 : node20394;
								assign node20394 = (inp[2]) ? node20592 : node20395;
									assign node20395 = (inp[3]) ? node20491 : node20396;
										assign node20396 = (inp[5]) ? node20434 : node20397;
											assign node20397 = (inp[12]) ? node20423 : node20398;
												assign node20398 = (inp[15]) ? node20408 : node20399;
													assign node20399 = (inp[0]) ? node20403 : node20400;
														assign node20400 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node20403 = (inp[9]) ? 4'b1101 : node20404;
															assign node20404 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node20408 = (inp[0]) ? node20414 : node20409;
														assign node20409 = (inp[10]) ? 4'b1101 : node20410;
															assign node20410 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node20414 = (inp[9]) ? node20416 : 4'b1011;
															assign node20416 = (inp[4]) ? node20420 : node20417;
																assign node20417 = (inp[10]) ? 4'b1111 : 4'b1011;
																assign node20420 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node20423 = (inp[4]) ? node20427 : node20424;
													assign node20424 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node20427 = (inp[9]) ? 4'b1011 : node20428;
														assign node20428 = (inp[0]) ? node20430 : 4'b1111;
															assign node20430 = (inp[15]) ? 4'b1111 : 4'b1101;
											assign node20434 = (inp[12]) ? node20466 : node20435;
												assign node20435 = (inp[15]) ? node20453 : node20436;
													assign node20436 = (inp[4]) ? node20446 : node20437;
														assign node20437 = (inp[9]) ? node20441 : node20438;
															assign node20438 = (inp[10]) ? 4'b1011 : 4'b1111;
															assign node20441 = (inp[10]) ? node20443 : 4'b1001;
																assign node20443 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node20446 = (inp[0]) ? node20448 : 4'b1011;
															assign node20448 = (inp[10]) ? node20450 : 4'b1111;
																assign node20450 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node20453 = (inp[10]) ? node20455 : 4'b1101;
														assign node20455 = (inp[4]) ? node20461 : node20456;
															assign node20456 = (inp[9]) ? 4'b1111 : node20457;
																assign node20457 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node20461 = (inp[9]) ? node20463 : 4'b1101;
																assign node20463 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node20466 = (inp[10]) ? node20472 : node20467;
													assign node20467 = (inp[4]) ? 4'b1001 : node20468;
														assign node20468 = (inp[0]) ? 4'b1111 : 4'b1011;
													assign node20472 = (inp[9]) ? node20480 : node20473;
														assign node20473 = (inp[4]) ? 4'b1101 : node20474;
															assign node20474 = (inp[15]) ? node20476 : 4'b1001;
																assign node20476 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node20480 = (inp[4]) ? node20486 : node20481;
															assign node20481 = (inp[0]) ? 4'b1101 : node20482;
																assign node20482 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node20486 = (inp[15]) ? 4'b1011 : node20487;
																assign node20487 = (inp[0]) ? 4'b1011 : 4'b1001;
										assign node20491 = (inp[12]) ? node20545 : node20492;
											assign node20492 = (inp[0]) ? node20520 : node20493;
												assign node20493 = (inp[15]) ? node20505 : node20494;
													assign node20494 = (inp[9]) ? 4'b1101 : node20495;
														assign node20495 = (inp[5]) ? node20499 : node20496;
															assign node20496 = (inp[4]) ? 4'b1101 : 4'b1011;
															assign node20499 = (inp[4]) ? node20501 : 4'b1101;
																assign node20501 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node20505 = (inp[5]) ? node20513 : node20506;
														assign node20506 = (inp[10]) ? 4'b1001 : node20507;
															assign node20507 = (inp[9]) ? 4'b1001 : node20508;
																assign node20508 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node20513 = (inp[4]) ? 4'b1011 : node20514;
															assign node20514 = (inp[10]) ? 4'b1111 : node20515;
																assign node20515 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node20520 = (inp[15]) ? node20536 : node20521;
													assign node20521 = (inp[5]) ? node20531 : node20522;
														assign node20522 = (inp[4]) ? node20526 : node20523;
															assign node20523 = (inp[9]) ? 4'b1111 : 4'b1001;
															assign node20526 = (inp[10]) ? node20528 : 4'b1111;
																assign node20528 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node20531 = (inp[10]) ? 4'b1011 : node20532;
															assign node20532 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node20536 = (inp[9]) ? node20538 : 4'b1101;
														assign node20538 = (inp[10]) ? node20542 : node20539;
															assign node20539 = (inp[5]) ? 4'b1001 : 4'b1011;
															assign node20542 = (inp[4]) ? 4'b1001 : 4'b1101;
											assign node20545 = (inp[10]) ? node20573 : node20546;
												assign node20546 = (inp[5]) ? node20554 : node20547;
													assign node20547 = (inp[9]) ? node20551 : node20548;
														assign node20548 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node20551 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node20554 = (inp[15]) ? node20562 : node20555;
														assign node20555 = (inp[0]) ? node20557 : 4'b1101;
															assign node20557 = (inp[4]) ? 4'b1011 : node20558;
																assign node20558 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node20562 = (inp[0]) ? node20566 : node20563;
															assign node20563 = (inp[4]) ? 4'b1111 : 4'b1011;
															assign node20566 = (inp[9]) ? node20570 : node20567;
																assign node20567 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node20570 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node20573 = (inp[5]) ? node20583 : node20574;
													assign node20574 = (inp[4]) ? node20580 : node20575;
														assign node20575 = (inp[15]) ? 4'b1011 : node20576;
															assign node20576 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node20580 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node20583 = (inp[0]) ? node20587 : node20584;
														assign node20584 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node20587 = (inp[4]) ? 4'b1001 : node20588;
															assign node20588 = (inp[15]) ? 4'b1101 : 4'b1111;
									assign node20592 = (inp[15]) ? node20682 : node20593;
										assign node20593 = (inp[3]) ? node20631 : node20594;
											assign node20594 = (inp[0]) ? node20608 : node20595;
												assign node20595 = (inp[5]) ? node20599 : node20596;
													assign node20596 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node20599 = (inp[9]) ? node20605 : node20600;
														assign node20600 = (inp[12]) ? node20602 : 4'b1010;
															assign node20602 = (inp[4]) ? 4'b1100 : 4'b1010;
														assign node20605 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node20608 = (inp[5]) ? node20620 : node20609;
													assign node20609 = (inp[12]) ? node20611 : 4'b1100;
														assign node20611 = (inp[10]) ? node20617 : node20612;
															assign node20612 = (inp[9]) ? node20614 : 4'b1100;
																assign node20614 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node20617 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node20620 = (inp[4]) ? node20628 : node20621;
														assign node20621 = (inp[10]) ? node20625 : node20622;
															assign node20622 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node20625 = (inp[9]) ? 4'b1110 : 4'b1000;
														assign node20628 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node20631 = (inp[0]) ? node20651 : node20632;
												assign node20632 = (inp[4]) ? node20644 : node20633;
													assign node20633 = (inp[9]) ? node20639 : node20634;
														assign node20634 = (inp[5]) ? 4'b1000 : node20635;
															assign node20635 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node20639 = (inp[10]) ? 4'b1100 : node20640;
															assign node20640 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node20644 = (inp[9]) ? node20648 : node20645;
														assign node20645 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node20648 = (inp[10]) ? 4'b1000 : 4'b1100;
												assign node20651 = (inp[5]) ? node20667 : node20652;
													assign node20652 = (inp[9]) ? node20664 : node20653;
														assign node20653 = (inp[4]) ? node20659 : node20654;
															assign node20654 = (inp[10]) ? 4'b1000 : node20655;
																assign node20655 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node20659 = (inp[12]) ? 4'b1110 : node20660;
																assign node20660 = (inp[10]) ? 4'b1110 : 4'b1000;
														assign node20664 = (inp[10]) ? 4'b1110 : 4'b1010;
													assign node20667 = (inp[9]) ? node20673 : node20668;
														assign node20668 = (inp[4]) ? node20670 : 4'b1010;
															assign node20670 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node20673 = (inp[4]) ? node20677 : node20674;
															assign node20674 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node20677 = (inp[10]) ? 4'b1010 : node20678;
																assign node20678 = (inp[12]) ? 4'b1010 : 4'b1110;
										assign node20682 = (inp[9]) ? node20714 : node20683;
											assign node20683 = (inp[4]) ? node20699 : node20684;
												assign node20684 = (inp[0]) ? node20692 : node20685;
													assign node20685 = (inp[5]) ? 4'b1010 : node20686;
														assign node20686 = (inp[12]) ? 4'b1000 : node20687;
															assign node20687 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node20692 = (inp[5]) ? node20696 : node20693;
														assign node20693 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node20696 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node20699 = (inp[12]) ? node20707 : node20700;
													assign node20700 = (inp[10]) ? node20704 : node20701;
														assign node20701 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node20704 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node20707 = (inp[0]) ? node20709 : 4'b1110;
														assign node20709 = (inp[3]) ? 4'b1100 : node20710;
															assign node20710 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node20714 = (inp[4]) ? node20738 : node20715;
												assign node20715 = (inp[10]) ? node20727 : node20716;
													assign node20716 = (inp[12]) ? node20722 : node20717;
														assign node20717 = (inp[5]) ? node20719 : 4'b1010;
															assign node20719 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node20722 = (inp[3]) ? 4'b1100 : node20723;
															assign node20723 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node20727 = (inp[12]) ? node20735 : node20728;
														assign node20728 = (inp[3]) ? 4'b1100 : node20729;
															assign node20729 = (inp[0]) ? node20731 : 4'b1100;
																assign node20731 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node20735 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node20738 = (inp[12]) ? node20752 : node20739;
													assign node20739 = (inp[10]) ? node20749 : node20740;
														assign node20740 = (inp[5]) ? node20746 : node20741;
															assign node20741 = (inp[3]) ? 4'b1100 : node20742;
																assign node20742 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node20746 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node20749 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node20752 = (inp[0]) ? node20758 : node20753;
														assign node20753 = (inp[3]) ? 4'b1010 : node20754;
															assign node20754 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node20758 = (inp[3]) ? 4'b1000 : node20759;
															assign node20759 = (inp[5]) ? 4'b1000 : 4'b1010;
								assign node20763 = (inp[2]) ? node20921 : node20764;
									assign node20764 = (inp[9]) ? node20834 : node20765;
										assign node20765 = (inp[4]) ? node20799 : node20766;
											assign node20766 = (inp[12]) ? node20786 : node20767;
												assign node20767 = (inp[10]) ? node20781 : node20768;
													assign node20768 = (inp[3]) ? node20776 : node20769;
														assign node20769 = (inp[0]) ? node20773 : node20770;
															assign node20770 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node20773 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node20776 = (inp[15]) ? node20778 : 4'b1100;
															assign node20778 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node20781 = (inp[15]) ? 4'b1000 : node20782;
														assign node20782 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node20786 = (inp[0]) ? node20794 : node20787;
													assign node20787 = (inp[15]) ? 4'b1000 : node20788;
														assign node20788 = (inp[3]) ? node20790 : 4'b1010;
															assign node20790 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node20794 = (inp[15]) ? 4'b1010 : node20795;
														assign node20795 = (inp[5]) ? 4'b1010 : 4'b1000;
											assign node20799 = (inp[10]) ? node20817 : node20800;
												assign node20800 = (inp[12]) ? node20808 : node20801;
													assign node20801 = (inp[0]) ? node20803 : 4'b1000;
														assign node20803 = (inp[3]) ? 4'b1010 : node20804;
															assign node20804 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node20808 = (inp[15]) ? node20812 : node20809;
														assign node20809 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node20812 = (inp[0]) ? 4'b1100 : node20813;
															assign node20813 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node20817 = (inp[15]) ? node20825 : node20818;
													assign node20818 = (inp[0]) ? 4'b1110 : node20819;
														assign node20819 = (inp[5]) ? 4'b1100 : node20820;
															assign node20820 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node20825 = (inp[5]) ? node20831 : node20826;
														assign node20826 = (inp[0]) ? node20828 : 4'b1100;
															assign node20828 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node20831 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node20834 = (inp[4]) ? node20874 : node20835;
											assign node20835 = (inp[10]) ? node20857 : node20836;
												assign node20836 = (inp[12]) ? node20852 : node20837;
													assign node20837 = (inp[0]) ? node20847 : node20838;
														assign node20838 = (inp[3]) ? node20842 : node20839;
															assign node20839 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node20842 = (inp[15]) ? node20844 : 4'b1000;
																assign node20844 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node20847 = (inp[5]) ? 4'b1000 : node20848;
															assign node20848 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node20852 = (inp[5]) ? node20854 : 4'b1100;
														assign node20854 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node20857 = (inp[5]) ? node20869 : node20858;
													assign node20858 = (inp[0]) ? node20866 : node20859;
														assign node20859 = (inp[3]) ? node20863 : node20860;
															assign node20860 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node20863 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node20866 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node20869 = (inp[3]) ? node20871 : 4'b1100;
														assign node20871 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node20874 = (inp[10]) ? node20896 : node20875;
												assign node20875 = (inp[12]) ? node20885 : node20876;
													assign node20876 = (inp[15]) ? node20882 : node20877;
														assign node20877 = (inp[3]) ? node20879 : 4'b1100;
															assign node20879 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node20882 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node20885 = (inp[15]) ? node20891 : node20886;
														assign node20886 = (inp[0]) ? node20888 : 4'b1000;
															assign node20888 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node20891 = (inp[0]) ? node20893 : 4'b1010;
															assign node20893 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node20896 = (inp[3]) ? node20908 : node20897;
													assign node20897 = (inp[0]) ? node20903 : node20898;
														assign node20898 = (inp[5]) ? node20900 : 4'b1010;
															assign node20900 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node20903 = (inp[5]) ? node20905 : 4'b1000;
															assign node20905 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node20908 = (inp[5]) ? node20914 : node20909;
														assign node20909 = (inp[0]) ? node20911 : 4'b1000;
															assign node20911 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node20914 = (inp[0]) ? node20918 : node20915;
															assign node20915 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node20918 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node20921 = (inp[0]) ? node20991 : node20922;
										assign node20922 = (inp[9]) ? node20956 : node20923;
											assign node20923 = (inp[4]) ? node20935 : node20924;
												assign node20924 = (inp[12]) ? 4'b0001 : node20925;
													assign node20925 = (inp[10]) ? node20929 : node20926;
														assign node20926 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node20929 = (inp[15]) ? 4'b0001 : node20930;
															assign node20930 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node20935 = (inp[10]) ? node20947 : node20936;
													assign node20936 = (inp[12]) ? node20942 : node20937;
														assign node20937 = (inp[15]) ? 4'b0001 : node20938;
															assign node20938 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node20942 = (inp[15]) ? node20944 : 4'b0101;
															assign node20944 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node20947 = (inp[15]) ? node20953 : node20948;
														assign node20948 = (inp[3]) ? 4'b0101 : node20949;
															assign node20949 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node20953 = (inp[5]) ? 4'b0111 : 4'b0101;
											assign node20956 = (inp[4]) ? node20980 : node20957;
												assign node20957 = (inp[12]) ? node20969 : node20958;
													assign node20958 = (inp[10]) ? node20964 : node20959;
														assign node20959 = (inp[5]) ? node20961 : 4'b0011;
															assign node20961 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node20964 = (inp[15]) ? node20966 : 4'b0101;
															assign node20966 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node20969 = (inp[15]) ? node20975 : node20970;
														assign node20970 = (inp[5]) ? 4'b0101 : node20971;
															assign node20971 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node20975 = (inp[3]) ? 4'b0111 : node20976;
															assign node20976 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node20980 = (inp[15]) ? node20986 : node20981;
													assign node20981 = (inp[10]) ? 4'b0001 : node20982;
														assign node20982 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node20986 = (inp[5]) ? 4'b0011 : node20987;
														assign node20987 = (inp[3]) ? 4'b0011 : 4'b0001;
										assign node20991 = (inp[5]) ? node21029 : node20992;
											assign node20992 = (inp[15]) ? node21008 : node20993;
												assign node20993 = (inp[9]) ? node20997 : node20994;
													assign node20994 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node20997 = (inp[3]) ? node20999 : 4'b0101;
														assign node20999 = (inp[4]) ? node21005 : node21000;
															assign node21000 = (inp[12]) ? 4'b0111 : node21001;
																assign node21001 = (inp[10]) ? 4'b0111 : 4'b0001;
															assign node21005 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node21008 = (inp[3]) ? node21020 : node21009;
													assign node21009 = (inp[4]) ? node21011 : 4'b0111;
														assign node21011 = (inp[10]) ? node21017 : node21012;
															assign node21012 = (inp[12]) ? 4'b0011 : node21013;
																assign node21013 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node21017 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node21020 = (inp[9]) ? node21022 : 4'b0011;
														assign node21022 = (inp[4]) ? node21024 : 4'b0101;
															assign node21024 = (inp[10]) ? 4'b0001 : node21025;
																assign node21025 = (inp[12]) ? 4'b0001 : 4'b0101;
											assign node21029 = (inp[15]) ? node21047 : node21030;
												assign node21030 = (inp[4]) ? node21038 : node21031;
													assign node21031 = (inp[3]) ? 4'b0011 : node21032;
														assign node21032 = (inp[9]) ? node21034 : 4'b0001;
															assign node21034 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node21038 = (inp[9]) ? node21044 : node21039;
														assign node21039 = (inp[10]) ? 4'b0111 : node21040;
															assign node21040 = (inp[3]) ? 4'b0011 : 4'b0111;
														assign node21044 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node21047 = (inp[3]) ? node21059 : node21048;
													assign node21048 = (inp[4]) ? node21050 : 4'b0011;
														assign node21050 = (inp[9]) ? node21054 : node21051;
															assign node21051 = (inp[10]) ? 4'b0101 : 4'b0011;
															assign node21054 = (inp[10]) ? 4'b0001 : node21055;
																assign node21055 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node21059 = (inp[10]) ? node21065 : node21060;
														assign node21060 = (inp[4]) ? node21062 : 4'b0001;
															assign node21062 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node21065 = (inp[4]) ? node21067 : 4'b0101;
															assign node21067 = (inp[9]) ? 4'b0001 : 4'b0101;
							assign node21070 = (inp[2]) ? node21434 : node21071;
								assign node21071 = (inp[8]) ? node21241 : node21072;
									assign node21072 = (inp[4]) ? node21160 : node21073;
										assign node21073 = (inp[9]) ? node21113 : node21074;
											assign node21074 = (inp[12]) ? node21096 : node21075;
												assign node21075 = (inp[10]) ? node21089 : node21076;
													assign node21076 = (inp[3]) ? node21082 : node21077;
														assign node21077 = (inp[15]) ? node21079 : 4'b1100;
															assign node21079 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node21082 = (inp[15]) ? node21084 : 4'b1110;
															assign node21084 = (inp[0]) ? node21086 : 4'b1100;
																assign node21086 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node21089 = (inp[5]) ? 4'b1010 : node21090;
														assign node21090 = (inp[0]) ? 4'b1000 : node21091;
															assign node21091 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node21096 = (inp[0]) ? node21102 : node21097;
													assign node21097 = (inp[15]) ? 4'b1000 : node21098;
														assign node21098 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node21102 = (inp[10]) ? 4'b1010 : node21103;
														assign node21103 = (inp[3]) ? node21105 : 4'b1010;
															assign node21105 = (inp[5]) ? node21109 : node21106;
																assign node21106 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node21109 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node21113 = (inp[12]) ? node21135 : node21114;
												assign node21114 = (inp[10]) ? node21124 : node21115;
													assign node21115 = (inp[15]) ? 4'b1000 : node21116;
														assign node21116 = (inp[5]) ? node21118 : 4'b1010;
															assign node21118 = (inp[0]) ? node21120 : 4'b1000;
																assign node21120 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node21124 = (inp[5]) ? node21130 : node21125;
														assign node21125 = (inp[3]) ? node21127 : 4'b1100;
															assign node21127 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node21130 = (inp[3]) ? node21132 : 4'b1110;
															assign node21132 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node21135 = (inp[15]) ? node21151 : node21136;
													assign node21136 = (inp[10]) ? node21144 : node21137;
														assign node21137 = (inp[3]) ? 4'b1100 : node21138;
															assign node21138 = (inp[0]) ? node21140 : 4'b1110;
																assign node21140 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node21144 = (inp[3]) ? 4'b1110 : node21145;
															assign node21145 = (inp[0]) ? node21147 : 4'b1110;
																assign node21147 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node21151 = (inp[5]) ? node21157 : node21152;
														assign node21152 = (inp[0]) ? node21154 : 4'b1100;
															assign node21154 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node21157 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node21160 = (inp[9]) ? node21204 : node21161;
											assign node21161 = (inp[10]) ? node21187 : node21162;
												assign node21162 = (inp[12]) ? node21180 : node21163;
													assign node21163 = (inp[3]) ? node21173 : node21164;
														assign node21164 = (inp[5]) ? node21166 : 4'b1000;
															assign node21166 = (inp[0]) ? node21170 : node21167;
																assign node21167 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node21170 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node21173 = (inp[5]) ? 4'b1010 : node21174;
															assign node21174 = (inp[15]) ? node21176 : 4'b1010;
																assign node21176 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node21180 = (inp[15]) ? node21182 : 4'b1110;
														assign node21182 = (inp[0]) ? 4'b1100 : node21183;
															assign node21183 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node21187 = (inp[3]) ? node21191 : node21188;
													assign node21188 = (inp[12]) ? 4'b1110 : 4'b1100;
													assign node21191 = (inp[12]) ? node21199 : node21192;
														assign node21192 = (inp[5]) ? 4'b1110 : node21193;
															assign node21193 = (inp[15]) ? 4'b1110 : node21194;
																assign node21194 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node21199 = (inp[0]) ? 4'b1100 : node21200;
															assign node21200 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node21204 = (inp[12]) ? node21222 : node21205;
												assign node21205 = (inp[10]) ? node21211 : node21206;
													assign node21206 = (inp[5]) ? 4'b1100 : node21207;
														assign node21207 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node21211 = (inp[15]) ? node21219 : node21212;
														assign node21212 = (inp[5]) ? 4'b1000 : node21213;
															assign node21213 = (inp[0]) ? 4'b1010 : node21214;
																assign node21214 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node21219 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node21222 = (inp[0]) ? node21230 : node21223;
													assign node21223 = (inp[15]) ? 4'b1010 : node21224;
														assign node21224 = (inp[3]) ? 4'b1000 : node21225;
															assign node21225 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node21230 = (inp[15]) ? node21236 : node21231;
														assign node21231 = (inp[10]) ? 4'b1010 : node21232;
															assign node21232 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node21236 = (inp[5]) ? 4'b1000 : node21237;
															assign node21237 = (inp[10]) ? 4'b1000 : 4'b1010;
									assign node21241 = (inp[5]) ? node21341 : node21242;
										assign node21242 = (inp[10]) ? node21294 : node21243;
											assign node21243 = (inp[12]) ? node21273 : node21244;
												assign node21244 = (inp[3]) ? node21256 : node21245;
													assign node21245 = (inp[0]) ? node21249 : node21246;
														assign node21246 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node21249 = (inp[15]) ? node21251 : 4'b0001;
															assign node21251 = (inp[4]) ? 4'b0111 : node21252;
																assign node21252 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node21256 = (inp[4]) ? node21264 : node21257;
														assign node21257 = (inp[9]) ? 4'b0001 : node21258;
															assign node21258 = (inp[15]) ? node21260 : 4'b0101;
																assign node21260 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node21264 = (inp[9]) ? node21268 : node21265;
															assign node21265 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node21268 = (inp[0]) ? node21270 : 4'b0111;
																assign node21270 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node21273 = (inp[15]) ? node21283 : node21274;
													assign node21274 = (inp[4]) ? node21278 : node21275;
														assign node21275 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node21278 = (inp[3]) ? 4'b0011 : node21279;
															assign node21279 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node21283 = (inp[0]) ? node21291 : node21284;
														assign node21284 = (inp[3]) ? 4'b0011 : node21285;
															assign node21285 = (inp[4]) ? node21287 : 4'b0001;
																assign node21287 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node21291 = (inp[3]) ? 4'b0101 : 4'b0011;
											assign node21294 = (inp[9]) ? node21318 : node21295;
												assign node21295 = (inp[4]) ? node21307 : node21296;
													assign node21296 = (inp[3]) ? node21304 : node21297;
														assign node21297 = (inp[12]) ? 4'b0001 : node21298;
															assign node21298 = (inp[15]) ? 4'b0011 : node21299;
																assign node21299 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node21304 = (inp[12]) ? 4'b0011 : 4'b0001;
													assign node21307 = (inp[12]) ? node21313 : node21308;
														assign node21308 = (inp[0]) ? node21310 : 4'b0111;
															assign node21310 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node21313 = (inp[3]) ? 4'b0101 : node21314;
															assign node21314 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node21318 = (inp[4]) ? node21336 : node21319;
													assign node21319 = (inp[12]) ? node21327 : node21320;
														assign node21320 = (inp[15]) ? 4'b0101 : node21321;
															assign node21321 = (inp[0]) ? node21323 : 4'b0101;
																assign node21323 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node21327 = (inp[15]) ? 4'b0111 : node21328;
															assign node21328 = (inp[3]) ? node21332 : node21329;
																assign node21329 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node21332 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node21336 = (inp[0]) ? node21338 : 4'b0001;
														assign node21338 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node21341 = (inp[15]) ? node21393 : node21342;
											assign node21342 = (inp[0]) ? node21370 : node21343;
												assign node21343 = (inp[12]) ? node21361 : node21344;
													assign node21344 = (inp[3]) ? node21354 : node21345;
														assign node21345 = (inp[9]) ? 4'b0101 : node21346;
															assign node21346 = (inp[4]) ? node21350 : node21347;
																assign node21347 = (inp[10]) ? 4'b0011 : 4'b0111;
																assign node21350 = (inp[10]) ? 4'b0101 : 4'b0011;
														assign node21354 = (inp[10]) ? node21356 : 4'b0101;
															assign node21356 = (inp[4]) ? node21358 : 4'b0101;
																assign node21358 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node21361 = (inp[3]) ? 4'b0001 : node21362;
														assign node21362 = (inp[4]) ? node21366 : node21363;
															assign node21363 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node21366 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node21370 = (inp[4]) ? node21386 : node21371;
													assign node21371 = (inp[3]) ? node21381 : node21372;
														assign node21372 = (inp[10]) ? node21378 : node21373;
															assign node21373 = (inp[9]) ? 4'b0001 : node21374;
																assign node21374 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node21378 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node21381 = (inp[10]) ? 4'b0011 : node21382;
															assign node21382 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node21386 = (inp[12]) ? node21390 : node21387;
														assign node21387 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node21390 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node21393 = (inp[0]) ? node21415 : node21394;
												assign node21394 = (inp[4]) ? node21408 : node21395;
													assign node21395 = (inp[3]) ? node21405 : node21396;
														assign node21396 = (inp[9]) ? node21402 : node21397;
															assign node21397 = (inp[12]) ? 4'b0001 : node21398;
																assign node21398 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node21402 = (inp[10]) ? 4'b0111 : 4'b0001;
														assign node21405 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node21408 = (inp[9]) ? node21410 : 4'b0111;
														assign node21410 = (inp[10]) ? 4'b0011 : node21411;
															assign node21411 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node21415 = (inp[9]) ? node21429 : node21416;
													assign node21416 = (inp[4]) ? node21424 : node21417;
														assign node21417 = (inp[3]) ? node21419 : 4'b0011;
															assign node21419 = (inp[10]) ? 4'b0001 : node21420;
																assign node21420 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node21424 = (inp[10]) ? 4'b0101 : node21425;
															assign node21425 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node21429 = (inp[4]) ? 4'b0001 : node21430;
														assign node21430 = (inp[10]) ? 4'b0101 : 4'b0001;
								assign node21434 = (inp[8]) ? node21632 : node21435;
									assign node21435 = (inp[3]) ? node21531 : node21436;
										assign node21436 = (inp[0]) ? node21484 : node21437;
											assign node21437 = (inp[15]) ? node21463 : node21438;
												assign node21438 = (inp[5]) ? node21454 : node21439;
													assign node21439 = (inp[12]) ? node21445 : node21440;
														assign node21440 = (inp[4]) ? node21442 : 4'b0111;
															assign node21442 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node21445 = (inp[10]) ? node21449 : node21446;
															assign node21446 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node21449 = (inp[9]) ? node21451 : 4'b0111;
																assign node21451 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node21454 = (inp[10]) ? 4'b0101 : node21455;
														assign node21455 = (inp[12]) ? node21459 : node21456;
															assign node21456 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node21459 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node21463 = (inp[5]) ? node21473 : node21464;
													assign node21464 = (inp[10]) ? node21466 : 4'b0101;
														assign node21466 = (inp[4]) ? node21470 : node21467;
															assign node21467 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node21470 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node21473 = (inp[4]) ? node21479 : node21474;
														assign node21474 = (inp[9]) ? node21476 : 4'b0001;
															assign node21476 = (inp[10]) ? 4'b0111 : 4'b0001;
														assign node21479 = (inp[10]) ? 4'b0011 : node21480;
															assign node21480 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node21484 = (inp[15]) ? node21500 : node21485;
												assign node21485 = (inp[5]) ? node21491 : node21486;
													assign node21486 = (inp[9]) ? 4'b0001 : node21487;
														assign node21487 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node21491 = (inp[9]) ? node21497 : node21492;
														assign node21492 = (inp[4]) ? 4'b0111 : node21493;
															assign node21493 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node21497 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node21500 = (inp[5]) ? node21518 : node21501;
													assign node21501 = (inp[4]) ? node21513 : node21502;
														assign node21502 = (inp[9]) ? node21508 : node21503;
															assign node21503 = (inp[10]) ? 4'b0011 : node21504;
																assign node21504 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node21508 = (inp[12]) ? 4'b0111 : node21509;
																assign node21509 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node21513 = (inp[10]) ? node21515 : 4'b0111;
															assign node21515 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node21518 = (inp[9]) ? node21528 : node21519;
														assign node21519 = (inp[12]) ? 4'b0011 : node21520;
															assign node21520 = (inp[10]) ? node21524 : node21521;
																assign node21521 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node21524 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node21528 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node21531 = (inp[10]) ? node21597 : node21532;
											assign node21532 = (inp[9]) ? node21568 : node21533;
												assign node21533 = (inp[0]) ? node21547 : node21534;
													assign node21534 = (inp[15]) ? node21540 : node21535;
														assign node21535 = (inp[5]) ? 4'b0101 : node21536;
															assign node21536 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node21540 = (inp[5]) ? node21542 : 4'b0101;
															assign node21542 = (inp[4]) ? node21544 : 4'b0011;
																assign node21544 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node21547 = (inp[15]) ? node21557 : node21548;
														assign node21548 = (inp[5]) ? node21550 : 4'b0001;
															assign node21550 = (inp[12]) ? node21554 : node21551;
																assign node21551 = (inp[4]) ? 4'b0011 : 4'b0111;
																assign node21554 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node21557 = (inp[5]) ? node21563 : node21558;
															assign node21558 = (inp[12]) ? node21560 : 4'b0011;
																assign node21560 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node21563 = (inp[12]) ? 4'b0001 : node21564;
																assign node21564 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node21568 = (inp[4]) ? node21586 : node21569;
													assign node21569 = (inp[12]) ? node21583 : node21570;
														assign node21570 = (inp[5]) ? node21578 : node21571;
															assign node21571 = (inp[15]) ? node21575 : node21572;
																assign node21572 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node21575 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node21578 = (inp[15]) ? node21580 : 4'b0011;
																assign node21580 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node21583 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node21586 = (inp[12]) ? node21590 : node21587;
														assign node21587 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node21590 = (inp[0]) ? node21594 : node21591;
															assign node21591 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node21594 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node21597 = (inp[4]) ? node21613 : node21598;
												assign node21598 = (inp[9]) ? node21606 : node21599;
													assign node21599 = (inp[15]) ? node21603 : node21600;
														assign node21600 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node21603 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node21606 = (inp[0]) ? node21610 : node21607;
														assign node21607 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node21610 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node21613 = (inp[9]) ? node21623 : node21614;
													assign node21614 = (inp[12]) ? node21618 : node21615;
														assign node21615 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node21618 = (inp[0]) ? 4'b0101 : node21619;
															assign node21619 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node21623 = (inp[5]) ? node21625 : 4'b0011;
														assign node21625 = (inp[15]) ? node21629 : node21626;
															assign node21626 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node21629 = (inp[0]) ? 4'b0001 : 4'b0011;
									assign node21632 = (inp[4]) ? node21726 : node21633;
										assign node21633 = (inp[9]) ? node21685 : node21634;
											assign node21634 = (inp[12]) ? node21654 : node21635;
												assign node21635 = (inp[10]) ? node21645 : node21636;
													assign node21636 = (inp[5]) ? node21638 : 4'b0110;
														assign node21638 = (inp[15]) ? 4'b0100 : node21639;
															assign node21639 = (inp[3]) ? node21641 : 4'b0110;
																assign node21641 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node21645 = (inp[3]) ? node21647 : 4'b0010;
														assign node21647 = (inp[0]) ? 4'b0000 : node21648;
															assign node21648 = (inp[5]) ? 4'b0010 : node21649;
																assign node21649 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node21654 = (inp[10]) ? node21674 : node21655;
													assign node21655 = (inp[5]) ? node21663 : node21656;
														assign node21656 = (inp[15]) ? node21660 : node21657;
															assign node21657 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node21660 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node21663 = (inp[3]) ? node21669 : node21664;
															assign node21664 = (inp[15]) ? 4'b0010 : node21665;
																assign node21665 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node21669 = (inp[15]) ? node21671 : 4'b0000;
																assign node21671 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node21674 = (inp[0]) ? node21680 : node21675;
														assign node21675 = (inp[15]) ? 4'b0000 : node21676;
															assign node21676 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node21680 = (inp[15]) ? node21682 : 4'b0000;
															assign node21682 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node21685 = (inp[12]) ? node21713 : node21686;
												assign node21686 = (inp[10]) ? node21704 : node21687;
													assign node21687 = (inp[5]) ? node21695 : node21688;
														assign node21688 = (inp[0]) ? node21692 : node21689;
															assign node21689 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node21692 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node21695 = (inp[15]) ? node21697 : 4'b0000;
															assign node21697 = (inp[0]) ? node21701 : node21698;
																assign node21698 = (inp[3]) ? 4'b0010 : 4'b0000;
																assign node21701 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node21704 = (inp[15]) ? node21706 : 4'b0100;
														assign node21706 = (inp[3]) ? 4'b0100 : node21707;
															assign node21707 = (inp[5]) ? node21709 : 4'b0110;
																assign node21709 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node21713 = (inp[15]) ? node21717 : node21714;
													assign node21714 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node21717 = (inp[5]) ? 4'b0110 : node21718;
														assign node21718 = (inp[0]) ? node21722 : node21719;
															assign node21719 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node21722 = (inp[3]) ? 4'b0100 : 4'b0110;
										assign node21726 = (inp[9]) ? node21772 : node21727;
											assign node21727 = (inp[12]) ? node21751 : node21728;
												assign node21728 = (inp[10]) ? node21740 : node21729;
													assign node21729 = (inp[5]) ? node21735 : node21730;
														assign node21730 = (inp[3]) ? node21732 : 4'b0000;
															assign node21732 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node21735 = (inp[15]) ? node21737 : 4'b0010;
															assign node21737 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node21740 = (inp[3]) ? node21746 : node21741;
														assign node21741 = (inp[15]) ? 4'b0100 : node21742;
															assign node21742 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node21746 = (inp[15]) ? 4'b0110 : node21747;
															assign node21747 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node21751 = (inp[0]) ? node21759 : node21752;
													assign node21752 = (inp[15]) ? node21756 : node21753;
														assign node21753 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node21756 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node21759 = (inp[15]) ? node21765 : node21760;
														assign node21760 = (inp[3]) ? 4'b0110 : node21761;
															assign node21761 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node21765 = (inp[10]) ? node21767 : 4'b0100;
															assign node21767 = (inp[3]) ? 4'b0100 : node21768;
																assign node21768 = (inp[5]) ? 4'b0100 : 4'b0110;
											assign node21772 = (inp[10]) ? node21796 : node21773;
												assign node21773 = (inp[12]) ? node21785 : node21774;
													assign node21774 = (inp[0]) ? node21776 : 4'b0110;
														assign node21776 = (inp[5]) ? 4'b0100 : node21777;
															assign node21777 = (inp[3]) ? node21781 : node21778;
																assign node21778 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node21781 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node21785 = (inp[0]) ? node21791 : node21786;
														assign node21786 = (inp[15]) ? 4'b0010 : node21787;
															assign node21787 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node21791 = (inp[15]) ? 4'b0000 : node21792;
															assign node21792 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node21796 = (inp[12]) ? node21808 : node21797;
													assign node21797 = (inp[0]) ? node21801 : node21798;
														assign node21798 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node21801 = (inp[15]) ? node21803 : 4'b0010;
															assign node21803 = (inp[5]) ? 4'b0000 : node21804;
																assign node21804 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node21808 = (inp[3]) ? 4'b0010 : node21809;
														assign node21809 = (inp[0]) ? 4'b0010 : 4'b0000;
					assign node21813 = (inp[1]) ? node23267 : node21814;
						assign node21814 = (inp[7]) ? node22528 : node21815;
							assign node21815 = (inp[8]) ? node22147 : node21816;
								assign node21816 = (inp[2]) ? node21962 : node21817;
									assign node21817 = (inp[9]) ? node21891 : node21818;
										assign node21818 = (inp[4]) ? node21856 : node21819;
											assign node21819 = (inp[12]) ? node21841 : node21820;
												assign node21820 = (inp[10]) ? node21830 : node21821;
													assign node21821 = (inp[15]) ? node21827 : node21822;
														assign node21822 = (inp[3]) ? node21824 : 4'b1111;
															assign node21824 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node21827 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node21830 = (inp[3]) ? node21836 : node21831;
														assign node21831 = (inp[15]) ? 4'b1011 : node21832;
															assign node21832 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node21836 = (inp[15]) ? node21838 : 4'b1001;
															assign node21838 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node21841 = (inp[3]) ? node21851 : node21842;
													assign node21842 = (inp[5]) ? node21848 : node21843;
														assign node21843 = (inp[10]) ? 4'b1011 : node21844;
															assign node21844 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node21848 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node21851 = (inp[0]) ? node21853 : 4'b1001;
														assign node21853 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node21856 = (inp[12]) ? node21874 : node21857;
												assign node21857 = (inp[10]) ? node21865 : node21858;
													assign node21858 = (inp[0]) ? node21860 : 4'b1011;
														assign node21860 = (inp[5]) ? 4'b1001 : node21861;
															assign node21861 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node21865 = (inp[0]) ? 4'b1101 : node21866;
														assign node21866 = (inp[15]) ? node21868 : 4'b1101;
															assign node21868 = (inp[3]) ? 4'b1111 : node21869;
																assign node21869 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node21874 = (inp[15]) ? node21884 : node21875;
													assign node21875 = (inp[0]) ? node21879 : node21876;
														assign node21876 = (inp[10]) ? 4'b1111 : 4'b1101;
														assign node21879 = (inp[5]) ? 4'b1111 : node21880;
															assign node21880 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node21884 = (inp[0]) ? node21888 : node21885;
														assign node21885 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node21888 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node21891 = (inp[4]) ? node21917 : node21892;
											assign node21892 = (inp[12]) ? node21906 : node21893;
												assign node21893 = (inp[10]) ? node21901 : node21894;
													assign node21894 = (inp[15]) ? 4'b1001 : node21895;
														assign node21895 = (inp[5]) ? node21897 : 4'b1011;
															assign node21897 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node21901 = (inp[5]) ? 4'b1111 : node21902;
														assign node21902 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node21906 = (inp[15]) ? node21912 : node21907;
													assign node21907 = (inp[0]) ? node21909 : 4'b1101;
														assign node21909 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node21912 = (inp[5]) ? node21914 : 4'b1111;
														assign node21914 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node21917 = (inp[12]) ? node21935 : node21918;
												assign node21918 = (inp[10]) ? node21924 : node21919;
													assign node21919 = (inp[0]) ? 4'b1101 : node21920;
														assign node21920 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node21924 = (inp[5]) ? 4'b1001 : node21925;
														assign node21925 = (inp[0]) ? 4'b1011 : node21926;
															assign node21926 = (inp[3]) ? node21930 : node21927;
																assign node21927 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node21930 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node21935 = (inp[3]) ? node21949 : node21936;
													assign node21936 = (inp[0]) ? node21942 : node21937;
														assign node21937 = (inp[5]) ? node21939 : 4'b1011;
															assign node21939 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node21942 = (inp[15]) ? node21946 : node21943;
															assign node21943 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node21946 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node21949 = (inp[10]) ? node21957 : node21950;
														assign node21950 = (inp[5]) ? node21952 : 4'b1001;
															assign node21952 = (inp[0]) ? 4'b1011 : node21953;
																assign node21953 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node21957 = (inp[0]) ? node21959 : 4'b1001;
															assign node21959 = (inp[15]) ? 4'b1001 : 4'b1011;
									assign node21962 = (inp[3]) ? node22050 : node21963;
										assign node21963 = (inp[0]) ? node22007 : node21964;
											assign node21964 = (inp[15]) ? node21984 : node21965;
												assign node21965 = (inp[4]) ? node21975 : node21966;
													assign node21966 = (inp[5]) ? 4'b1010 : node21967;
														assign node21967 = (inp[10]) ? node21971 : node21968;
															assign node21968 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node21971 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node21975 = (inp[5]) ? node21981 : node21976;
														assign node21976 = (inp[12]) ? node21978 : 4'b1110;
															assign node21978 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node21981 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node21984 = (inp[5]) ? node21996 : node21985;
													assign node21985 = (inp[4]) ? node21991 : node21986;
														assign node21986 = (inp[9]) ? node21988 : 4'b1000;
															assign node21988 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node21991 = (inp[9]) ? node21993 : 4'b1100;
															assign node21993 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node21996 = (inp[4]) ? 4'b1010 : node21997;
														assign node21997 = (inp[9]) ? node22003 : node21998;
															assign node21998 = (inp[10]) ? 4'b1000 : node21999;
																assign node21999 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node22003 = (inp[12]) ? 4'b1110 : 4'b1000;
											assign node22007 = (inp[15]) ? node22027 : node22008;
												assign node22008 = (inp[5]) ? node22018 : node22009;
													assign node22009 = (inp[10]) ? node22011 : 4'b1100;
														assign node22011 = (inp[9]) ? node22015 : node22012;
															assign node22012 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node22015 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node22018 = (inp[10]) ? 4'b1110 : node22019;
														assign node22019 = (inp[9]) ? 4'b1010 : node22020;
															assign node22020 = (inp[12]) ? 4'b1000 : node22021;
																assign node22021 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node22027 = (inp[5]) ? node22039 : node22028;
													assign node22028 = (inp[4]) ? node22036 : node22029;
														assign node22029 = (inp[9]) ? 4'b1110 : node22030;
															assign node22030 = (inp[10]) ? 4'b1010 : node22031;
																assign node22031 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node22036 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node22039 = (inp[4]) ? node22043 : node22040;
														assign node22040 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node22043 = (inp[9]) ? node22045 : 4'b1100;
															assign node22045 = (inp[12]) ? 4'b1000 : node22046;
																assign node22046 = (inp[10]) ? 4'b1000 : 4'b1100;
										assign node22050 = (inp[15]) ? node22084 : node22051;
											assign node22051 = (inp[0]) ? node22063 : node22052;
												assign node22052 = (inp[9]) ? 4'b1100 : node22053;
													assign node22053 = (inp[4]) ? 4'b1100 : node22054;
														assign node22054 = (inp[5]) ? node22058 : node22055;
															assign node22055 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node22058 = (inp[12]) ? 4'b1000 : 4'b1100;
												assign node22063 = (inp[5]) ? node22071 : node22064;
													assign node22064 = (inp[9]) ? node22066 : 4'b1110;
														assign node22066 = (inp[12]) ? 4'b1010 : node22067;
															assign node22067 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node22071 = (inp[10]) ? node22079 : node22072;
														assign node22072 = (inp[9]) ? node22074 : 4'b1010;
															assign node22074 = (inp[12]) ? 4'b1110 : node22075;
																assign node22075 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node22079 = (inp[4]) ? node22081 : 4'b1110;
															assign node22081 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node22084 = (inp[0]) ? node22106 : node22085;
												assign node22085 = (inp[4]) ? node22095 : node22086;
													assign node22086 = (inp[9]) ? 4'b1110 : node22087;
														assign node22087 = (inp[5]) ? node22091 : node22088;
															assign node22088 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node22091 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node22095 = (inp[9]) ? node22101 : node22096;
														assign node22096 = (inp[10]) ? 4'b1110 : node22097;
															assign node22097 = (inp[12]) ? 4'b1110 : 4'b1010;
														assign node22101 = (inp[12]) ? 4'b1010 : node22102;
															assign node22102 = (inp[5]) ? 4'b1110 : 4'b1010;
												assign node22106 = (inp[5]) ? node22124 : node22107;
													assign node22107 = (inp[9]) ? node22115 : node22108;
														assign node22108 = (inp[12]) ? 4'b1010 : node22109;
															assign node22109 = (inp[10]) ? 4'b1100 : node22110;
																assign node22110 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node22115 = (inp[4]) ? node22119 : node22116;
															assign node22116 = (inp[10]) ? 4'b1100 : 4'b1010;
															assign node22119 = (inp[12]) ? 4'b1000 : node22120;
																assign node22120 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node22124 = (inp[12]) ? node22134 : node22125;
														assign node22125 = (inp[10]) ? node22127 : 4'b1100;
															assign node22127 = (inp[9]) ? node22131 : node22128;
																assign node22128 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node22131 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node22134 = (inp[10]) ? node22140 : node22135;
															assign node22135 = (inp[9]) ? node22137 : 4'b1000;
																assign node22137 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node22140 = (inp[9]) ? node22144 : node22141;
																assign node22141 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node22144 = (inp[4]) ? 4'b1000 : 4'b1100;
								assign node22147 = (inp[2]) ? node22323 : node22148;
									assign node22148 = (inp[12]) ? node22248 : node22149;
										assign node22149 = (inp[5]) ? node22197 : node22150;
											assign node22150 = (inp[9]) ? node22174 : node22151;
												assign node22151 = (inp[0]) ? node22163 : node22152;
													assign node22152 = (inp[15]) ? node22158 : node22153;
														assign node22153 = (inp[4]) ? 4'b1100 : node22154;
															assign node22154 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node22158 = (inp[10]) ? 4'b1000 : node22159;
															assign node22159 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node22163 = (inp[15]) ? node22167 : node22164;
														assign node22164 = (inp[10]) ? 4'b1100 : 4'b1000;
														assign node22167 = (inp[3]) ? 4'b1010 : node22168;
															assign node22168 = (inp[4]) ? node22170 : 4'b1110;
																assign node22170 = (inp[10]) ? 4'b1110 : 4'b1010;
												assign node22174 = (inp[4]) ? node22186 : node22175;
													assign node22175 = (inp[10]) ? node22183 : node22176;
														assign node22176 = (inp[3]) ? 4'b1000 : node22177;
															assign node22177 = (inp[0]) ? 4'b1010 : node22178;
																assign node22178 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node22183 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node22186 = (inp[10]) ? node22188 : 4'b1110;
														assign node22188 = (inp[15]) ? 4'b1010 : node22189;
															assign node22189 = (inp[0]) ? node22193 : node22190;
																assign node22190 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node22193 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node22197 = (inp[15]) ? node22225 : node22198;
												assign node22198 = (inp[0]) ? node22216 : node22199;
													assign node22199 = (inp[9]) ? node22211 : node22200;
														assign node22200 = (inp[3]) ? node22206 : node22201;
															assign node22201 = (inp[4]) ? 4'b1100 : node22202;
																assign node22202 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node22206 = (inp[4]) ? 4'b1000 : node22207;
																assign node22207 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node22211 = (inp[4]) ? node22213 : 4'b1100;
															assign node22213 = (inp[10]) ? 4'b1000 : 4'b1100;
													assign node22216 = (inp[3]) ? node22220 : node22217;
														assign node22217 = (inp[4]) ? 4'b1010 : 4'b1000;
														assign node22220 = (inp[10]) ? node22222 : 4'b1010;
															assign node22222 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node22225 = (inp[0]) ? node22239 : node22226;
													assign node22226 = (inp[4]) ? node22232 : node22227;
														assign node22227 = (inp[3]) ? 4'b1110 : node22228;
															assign node22228 = (inp[10]) ? 4'b1110 : 4'b1100;
														assign node22232 = (inp[3]) ? 4'b1010 : node22233;
															assign node22233 = (inp[10]) ? node22235 : 4'b1110;
																assign node22235 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node22239 = (inp[9]) ? 4'b1100 : node22240;
														assign node22240 = (inp[4]) ? node22242 : 4'b1010;
															assign node22242 = (inp[10]) ? 4'b1100 : node22243;
																assign node22243 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node22248 = (inp[0]) ? node22292 : node22249;
											assign node22249 = (inp[15]) ? node22267 : node22250;
												assign node22250 = (inp[5]) ? node22260 : node22251;
													assign node22251 = (inp[4]) ? node22255 : node22252;
														assign node22252 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node22255 = (inp[9]) ? node22257 : 4'b1100;
															assign node22257 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node22260 = (inp[9]) ? 4'b1100 : node22261;
														assign node22261 = (inp[4]) ? 4'b1100 : node22262;
															assign node22262 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node22267 = (inp[5]) ? node22285 : node22268;
													assign node22268 = (inp[3]) ? node22280 : node22269;
														assign node22269 = (inp[10]) ? node22275 : node22270;
															assign node22270 = (inp[4]) ? 4'b1100 : node22271;
																assign node22271 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node22275 = (inp[4]) ? node22277 : 4'b1100;
																assign node22277 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node22280 = (inp[9]) ? node22282 : 4'b1000;
															assign node22282 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node22285 = (inp[4]) ? node22289 : node22286;
														assign node22286 = (inp[10]) ? 4'b1010 : 4'b1000;
														assign node22289 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node22292 = (inp[15]) ? node22312 : node22293;
												assign node22293 = (inp[5]) ? node22305 : node22294;
													assign node22294 = (inp[3]) ? node22300 : node22295;
														assign node22295 = (inp[4]) ? node22297 : 4'b1100;
															assign node22297 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node22300 = (inp[4]) ? node22302 : 4'b1000;
															assign node22302 = (inp[10]) ? 4'b1110 : 4'b1010;
													assign node22305 = (inp[9]) ? node22309 : node22306;
														assign node22306 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node22309 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node22312 = (inp[4]) ? node22320 : node22313;
													assign node22313 = (inp[9]) ? node22315 : 4'b1010;
														assign node22315 = (inp[3]) ? 4'b1100 : node22316;
															assign node22316 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node22320 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node22323 = (inp[9]) ? node22415 : node22324;
										assign node22324 = (inp[4]) ? node22362 : node22325;
											assign node22325 = (inp[10]) ? node22343 : node22326;
												assign node22326 = (inp[12]) ? node22336 : node22327;
													assign node22327 = (inp[15]) ? node22329 : 4'b0101;
														assign node22329 = (inp[3]) ? node22331 : 4'b0101;
															assign node22331 = (inp[0]) ? 4'b0111 : node22332;
																assign node22332 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node22336 = (inp[3]) ? 4'b0001 : node22337;
														assign node22337 = (inp[0]) ? node22339 : 4'b0011;
															assign node22339 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node22343 = (inp[5]) ? node22351 : node22344;
													assign node22344 = (inp[15]) ? node22348 : node22345;
														assign node22345 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node22348 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node22351 = (inp[15]) ? node22357 : node22352;
														assign node22352 = (inp[0]) ? 4'b0011 : node22353;
															assign node22353 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node22357 = (inp[0]) ? 4'b0001 : node22358;
															assign node22358 = (inp[3]) ? 4'b0011 : 4'b0001;
											assign node22362 = (inp[10]) ? node22390 : node22363;
												assign node22363 = (inp[12]) ? node22375 : node22364;
													assign node22364 = (inp[5]) ? 4'b0001 : node22365;
														assign node22365 = (inp[3]) ? node22367 : 4'b0011;
															assign node22367 = (inp[0]) ? node22371 : node22368;
																assign node22368 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node22371 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node22375 = (inp[5]) ? 4'b0101 : node22376;
														assign node22376 = (inp[15]) ? node22382 : node22377;
															assign node22377 = (inp[0]) ? 4'b0111 : node22378;
																assign node22378 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node22382 = (inp[0]) ? node22386 : node22383;
																assign node22383 = (inp[3]) ? 4'b0111 : 4'b0101;
																assign node22386 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node22390 = (inp[3]) ? node22400 : node22391;
													assign node22391 = (inp[12]) ? 4'b0101 : node22392;
														assign node22392 = (inp[0]) ? 4'b0111 : node22393;
															assign node22393 = (inp[15]) ? node22395 : 4'b0101;
																assign node22395 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node22400 = (inp[5]) ? node22410 : node22401;
														assign node22401 = (inp[12]) ? 4'b0111 : node22402;
															assign node22402 = (inp[0]) ? node22406 : node22403;
																assign node22403 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node22406 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node22410 = (inp[12]) ? node22412 : 4'b0101;
															assign node22412 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node22415 = (inp[4]) ? node22475 : node22416;
											assign node22416 = (inp[10]) ? node22442 : node22417;
												assign node22417 = (inp[12]) ? node22429 : node22418;
													assign node22418 = (inp[15]) ? 4'b0011 : node22419;
														assign node22419 = (inp[0]) ? node22425 : node22420;
															assign node22420 = (inp[5]) ? node22422 : 4'b0011;
																assign node22422 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node22425 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node22429 = (inp[3]) ? node22435 : node22430;
														assign node22430 = (inp[5]) ? node22432 : 4'b0101;
															assign node22432 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node22435 = (inp[15]) ? node22439 : node22436;
															assign node22436 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node22439 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node22442 = (inp[12]) ? node22460 : node22443;
													assign node22443 = (inp[15]) ? node22449 : node22444;
														assign node22444 = (inp[3]) ? node22446 : 4'b0111;
															assign node22446 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node22449 = (inp[0]) ? node22455 : node22450;
															assign node22450 = (inp[5]) ? 4'b0111 : node22451;
																assign node22451 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node22455 = (inp[3]) ? 4'b0101 : node22456;
																assign node22456 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node22460 = (inp[15]) ? node22470 : node22461;
														assign node22461 = (inp[0]) ? node22467 : node22462;
															assign node22462 = (inp[3]) ? 4'b0101 : node22463;
																assign node22463 = (inp[5]) ? 4'b0101 : 4'b0111;
															assign node22467 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node22470 = (inp[0]) ? node22472 : 4'b0111;
															assign node22472 = (inp[5]) ? 4'b0101 : 4'b0111;
											assign node22475 = (inp[12]) ? node22499 : node22476;
												assign node22476 = (inp[10]) ? node22486 : node22477;
													assign node22477 = (inp[0]) ? 4'b0101 : node22478;
														assign node22478 = (inp[15]) ? node22482 : node22479;
															assign node22479 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node22482 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node22486 = (inp[15]) ? node22488 : 4'b0011;
														assign node22488 = (inp[0]) ? node22494 : node22489;
															assign node22489 = (inp[3]) ? 4'b0011 : node22490;
																assign node22490 = (inp[5]) ? 4'b0011 : 4'b0001;
															assign node22494 = (inp[5]) ? 4'b0001 : node22495;
																assign node22495 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node22499 = (inp[0]) ? node22513 : node22500;
													assign node22500 = (inp[3]) ? 4'b0011 : node22501;
														assign node22501 = (inp[10]) ? node22507 : node22502;
															assign node22502 = (inp[5]) ? 4'b0011 : node22503;
																assign node22503 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node22507 = (inp[5]) ? node22509 : 4'b0011;
																assign node22509 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node22513 = (inp[10]) ? node22523 : node22514;
														assign node22514 = (inp[3]) ? 4'b0011 : node22515;
															assign node22515 = (inp[5]) ? node22519 : node22516;
																assign node22516 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node22519 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node22523 = (inp[15]) ? 4'b0001 : node22524;
															assign node22524 = (inp[3]) ? 4'b0011 : 4'b0001;
							assign node22528 = (inp[2]) ? node22888 : node22529;
								assign node22529 = (inp[8]) ? node22691 : node22530;
									assign node22530 = (inp[9]) ? node22612 : node22531;
										assign node22531 = (inp[4]) ? node22571 : node22532;
											assign node22532 = (inp[10]) ? node22554 : node22533;
												assign node22533 = (inp[12]) ? node22541 : node22534;
													assign node22534 = (inp[15]) ? node22536 : 4'b1100;
														assign node22536 = (inp[5]) ? node22538 : 4'b1110;
															assign node22538 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node22541 = (inp[5]) ? node22547 : node22542;
														assign node22542 = (inp[15]) ? node22544 : 4'b1000;
															assign node22544 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node22547 = (inp[3]) ? node22549 : 4'b1010;
															assign node22549 = (inp[15]) ? 4'b1010 : node22550;
																assign node22550 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node22554 = (inp[15]) ? node22564 : node22555;
													assign node22555 = (inp[0]) ? node22559 : node22556;
														assign node22556 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node22559 = (inp[5]) ? node22561 : 4'b1000;
															assign node22561 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node22564 = (inp[12]) ? 4'b1000 : node22565;
														assign node22565 = (inp[0]) ? 4'b1010 : node22566;
															assign node22566 = (inp[3]) ? 4'b1010 : 4'b1000;
											assign node22571 = (inp[10]) ? node22595 : node22572;
												assign node22572 = (inp[12]) ? node22582 : node22573;
													assign node22573 = (inp[15]) ? node22577 : node22574;
														assign node22574 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node22577 = (inp[0]) ? node22579 : 4'b1000;
															assign node22579 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node22582 = (inp[5]) ? node22590 : node22583;
														assign node22583 = (inp[15]) ? node22587 : node22584;
															assign node22584 = (inp[3]) ? 4'b1100 : 4'b1110;
															assign node22587 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node22590 = (inp[15]) ? node22592 : 4'b1110;
															assign node22592 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node22595 = (inp[3]) ? node22605 : node22596;
													assign node22596 = (inp[0]) ? node22598 : 4'b1110;
														assign node22598 = (inp[15]) ? node22602 : node22599;
															assign node22599 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node22602 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node22605 = (inp[15]) ? node22609 : node22606;
														assign node22606 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node22609 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node22612 = (inp[4]) ? node22648 : node22613;
											assign node22613 = (inp[10]) ? node22631 : node22614;
												assign node22614 = (inp[12]) ? node22626 : node22615;
													assign node22615 = (inp[15]) ? node22617 : 4'b1000;
														assign node22617 = (inp[5]) ? node22621 : node22618;
															assign node22618 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node22621 = (inp[3]) ? node22623 : 4'b1000;
																assign node22623 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node22626 = (inp[15]) ? 4'b1100 : node22627;
														assign node22627 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node22631 = (inp[3]) ? node22643 : node22632;
													assign node22632 = (inp[15]) ? node22638 : node22633;
														assign node22633 = (inp[12]) ? node22635 : 4'b1110;
															assign node22635 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node22638 = (inp[0]) ? 4'b1100 : node22639;
															assign node22639 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node22643 = (inp[15]) ? 4'b1110 : node22644;
														assign node22644 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node22648 = (inp[12]) ? node22668 : node22649;
												assign node22649 = (inp[10]) ? node22659 : node22650;
													assign node22650 = (inp[5]) ? node22652 : 4'b1100;
														assign node22652 = (inp[15]) ? node22656 : node22653;
															assign node22653 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node22656 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node22659 = (inp[15]) ? node22663 : node22660;
														assign node22660 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node22663 = (inp[5]) ? node22665 : 4'b1000;
															assign node22665 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node22668 = (inp[5]) ? node22684 : node22669;
													assign node22669 = (inp[10]) ? node22677 : node22670;
														assign node22670 = (inp[0]) ? node22672 : 4'b1000;
															assign node22672 = (inp[15]) ? node22674 : 4'b1000;
																assign node22674 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node22677 = (inp[15]) ? 4'b1000 : node22678;
															assign node22678 = (inp[0]) ? node22680 : 4'b1010;
																assign node22680 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node22684 = (inp[0]) ? node22688 : node22685;
														assign node22685 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node22688 = (inp[15]) ? 4'b1000 : 4'b1010;
									assign node22691 = (inp[12]) ? node22795 : node22692;
										assign node22692 = (inp[10]) ? node22736 : node22693;
											assign node22693 = (inp[9]) ? node22723 : node22694;
												assign node22694 = (inp[4]) ? node22710 : node22695;
													assign node22695 = (inp[0]) ? node22705 : node22696;
														assign node22696 = (inp[15]) ? node22702 : node22697;
															assign node22697 = (inp[5]) ? node22699 : 4'b0111;
																assign node22699 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node22702 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node22705 = (inp[15]) ? 4'b0111 : node22706;
															assign node22706 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node22710 = (inp[5]) ? node22712 : 4'b0011;
														assign node22712 = (inp[15]) ? node22718 : node22713;
															assign node22713 = (inp[3]) ? 4'b0001 : node22714;
																assign node22714 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node22718 = (inp[0]) ? 4'b0011 : node22719;
																assign node22719 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node22723 = (inp[4]) ? node22729 : node22724;
													assign node22724 = (inp[15]) ? 4'b0001 : node22725;
														assign node22725 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node22729 = (inp[3]) ? node22731 : 4'b0101;
														assign node22731 = (inp[0]) ? 4'b0111 : node22732;
															assign node22732 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node22736 = (inp[4]) ? node22766 : node22737;
												assign node22737 = (inp[9]) ? node22753 : node22738;
													assign node22738 = (inp[0]) ? node22744 : node22739;
														assign node22739 = (inp[15]) ? 4'b0001 : node22740;
															assign node22740 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node22744 = (inp[5]) ? node22746 : 4'b0011;
															assign node22746 = (inp[15]) ? node22750 : node22747;
																assign node22747 = (inp[3]) ? 4'b0011 : 4'b0001;
																assign node22750 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node22753 = (inp[5]) ? node22761 : node22754;
														assign node22754 = (inp[3]) ? node22758 : node22755;
															assign node22755 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node22758 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node22761 = (inp[15]) ? node22763 : 4'b0111;
															assign node22763 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node22766 = (inp[9]) ? node22782 : node22767;
													assign node22767 = (inp[0]) ? node22775 : node22768;
														assign node22768 = (inp[15]) ? 4'b0111 : node22769;
															assign node22769 = (inp[3]) ? 4'b0101 : node22770;
																assign node22770 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node22775 = (inp[15]) ? 4'b0101 : node22776;
															assign node22776 = (inp[3]) ? 4'b0111 : node22777;
																assign node22777 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node22782 = (inp[15]) ? node22788 : node22783;
														assign node22783 = (inp[0]) ? node22785 : 4'b0001;
															assign node22785 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node22788 = (inp[0]) ? 4'b0001 : node22789;
															assign node22789 = (inp[3]) ? 4'b0011 : node22790;
																assign node22790 = (inp[5]) ? 4'b0011 : 4'b0001;
										assign node22795 = (inp[15]) ? node22843 : node22796;
											assign node22796 = (inp[3]) ? node22824 : node22797;
												assign node22797 = (inp[0]) ? node22809 : node22798;
													assign node22798 = (inp[5]) ? node22806 : node22799;
														assign node22799 = (inp[4]) ? node22803 : node22800;
															assign node22800 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node22803 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node22806 = (inp[9]) ? 4'b0001 : 4'b0011;
													assign node22809 = (inp[5]) ? node22817 : node22810;
														assign node22810 = (inp[10]) ? 4'b0101 : node22811;
															assign node22811 = (inp[4]) ? node22813 : 4'b0001;
																assign node22813 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node22817 = (inp[10]) ? node22819 : 4'b0111;
															assign node22819 = (inp[9]) ? node22821 : 4'b0001;
																assign node22821 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node22824 = (inp[0]) ? node22836 : node22825;
													assign node22825 = (inp[5]) ? node22831 : node22826;
														assign node22826 = (inp[4]) ? node22828 : 4'b0011;
															assign node22828 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node22831 = (inp[4]) ? 4'b0001 : node22832;
															assign node22832 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node22836 = (inp[9]) ? node22840 : node22837;
														assign node22837 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node22840 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node22843 = (inp[5]) ? node22873 : node22844;
												assign node22844 = (inp[0]) ? node22860 : node22845;
													assign node22845 = (inp[3]) ? node22853 : node22846;
														assign node22846 = (inp[9]) ? node22850 : node22847;
															assign node22847 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node22850 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node22853 = (inp[4]) ? node22857 : node22854;
															assign node22854 = (inp[9]) ? 4'b0111 : 4'b0001;
															assign node22857 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node22860 = (inp[3]) ? node22868 : node22861;
														assign node22861 = (inp[10]) ? 4'b0111 : node22862;
															assign node22862 = (inp[9]) ? node22864 : 4'b0011;
																assign node22864 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node22868 = (inp[9]) ? node22870 : 4'b0011;
															assign node22870 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node22873 = (inp[0]) ? node22883 : node22874;
													assign node22874 = (inp[4]) ? node22880 : node22875;
														assign node22875 = (inp[9]) ? 4'b0111 : node22876;
															assign node22876 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node22880 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node22883 = (inp[4]) ? 4'b0101 : node22884;
														assign node22884 = (inp[9]) ? 4'b0101 : 4'b0011;
								assign node22888 = (inp[8]) ? node23102 : node22889;
									assign node22889 = (inp[10]) ? node23013 : node22890;
										assign node22890 = (inp[15]) ? node22962 : node22891;
											assign node22891 = (inp[9]) ? node22921 : node22892;
												assign node22892 = (inp[3]) ? node22908 : node22893;
													assign node22893 = (inp[0]) ? node22903 : node22894;
														assign node22894 = (inp[5]) ? node22900 : node22895;
															assign node22895 = (inp[4]) ? node22897 : 4'b0111;
																assign node22897 = (inp[12]) ? 4'b0111 : 4'b0011;
															assign node22900 = (inp[12]) ? 4'b0101 : 4'b0111;
														assign node22903 = (inp[12]) ? node22905 : 4'b0101;
															assign node22905 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node22908 = (inp[12]) ? node22916 : node22909;
														assign node22909 = (inp[4]) ? 4'b0011 : node22910;
															assign node22910 = (inp[0]) ? 4'b0101 : node22911;
																assign node22911 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node22916 = (inp[4]) ? node22918 : 4'b0011;
															assign node22918 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node22921 = (inp[3]) ? node22949 : node22922;
													assign node22922 = (inp[0]) ? node22938 : node22923;
														assign node22923 = (inp[5]) ? node22931 : node22924;
															assign node22924 = (inp[12]) ? node22928 : node22925;
																assign node22925 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node22928 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node22931 = (inp[12]) ? node22935 : node22932;
																assign node22932 = (inp[4]) ? 4'b0101 : 4'b0011;
																assign node22935 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node22938 = (inp[5]) ? node22944 : node22939;
															assign node22939 = (inp[12]) ? node22941 : 4'b0001;
																assign node22941 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node22944 = (inp[12]) ? node22946 : 4'b0001;
																assign node22946 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node22949 = (inp[0]) ? node22955 : node22950;
														assign node22950 = (inp[4]) ? node22952 : 4'b0101;
															assign node22952 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node22955 = (inp[5]) ? node22957 : 4'b0001;
															assign node22957 = (inp[12]) ? 4'b0111 : node22958;
																assign node22958 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node22962 = (inp[4]) ? node22982 : node22963;
												assign node22963 = (inp[0]) ? node22973 : node22964;
													assign node22964 = (inp[9]) ? node22970 : node22965;
														assign node22965 = (inp[3]) ? 4'b0011 : node22966;
															assign node22966 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node22970 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node22973 = (inp[3]) ? node22979 : node22974;
														assign node22974 = (inp[9]) ? 4'b0011 : node22975;
															assign node22975 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node22979 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node22982 = (inp[0]) ? node22996 : node22983;
													assign node22983 = (inp[5]) ? node22993 : node22984;
														assign node22984 = (inp[3]) ? node22990 : node22985;
															assign node22985 = (inp[9]) ? node22987 : 4'b0001;
																assign node22987 = (inp[12]) ? 4'b0001 : 4'b0101;
															assign node22990 = (inp[12]) ? 4'b0011 : 4'b0001;
														assign node22993 = (inp[3]) ? 4'b0111 : 4'b0011;
													assign node22996 = (inp[5]) ? node23004 : node22997;
														assign node22997 = (inp[3]) ? node22999 : 4'b0111;
															assign node22999 = (inp[12]) ? 4'b0101 : node23000;
																assign node23000 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node23004 = (inp[3]) ? 4'b0101 : node23005;
															assign node23005 = (inp[9]) ? node23009 : node23006;
																assign node23006 = (inp[12]) ? 4'b0101 : 4'b0011;
																assign node23009 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node23013 = (inp[4]) ? node23061 : node23014;
											assign node23014 = (inp[9]) ? node23038 : node23015;
												assign node23015 = (inp[3]) ? node23029 : node23016;
													assign node23016 = (inp[12]) ? node23022 : node23017;
														assign node23017 = (inp[0]) ? node23019 : 4'b0001;
															assign node23019 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node23022 = (inp[15]) ? node23026 : node23023;
															assign node23023 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node23026 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node23029 = (inp[0]) ? node23031 : 4'b0011;
														assign node23031 = (inp[5]) ? node23035 : node23032;
															assign node23032 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node23035 = (inp[12]) ? 4'b0001 : 4'b0011;
												assign node23038 = (inp[0]) ? node23048 : node23039;
													assign node23039 = (inp[15]) ? node23043 : node23040;
														assign node23040 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node23043 = (inp[3]) ? 4'b0111 : node23044;
															assign node23044 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node23048 = (inp[12]) ? node23056 : node23049;
														assign node23049 = (inp[15]) ? node23053 : node23050;
															assign node23050 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node23053 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node23056 = (inp[3]) ? node23058 : 4'b0111;
															assign node23058 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node23061 = (inp[9]) ? node23081 : node23062;
												assign node23062 = (inp[15]) ? node23072 : node23063;
													assign node23063 = (inp[12]) ? node23065 : 4'b0101;
														assign node23065 = (inp[3]) ? 4'b0101 : node23066;
															assign node23066 = (inp[0]) ? node23068 : 4'b0111;
																assign node23068 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node23072 = (inp[12]) ? node23074 : 4'b0111;
														assign node23074 = (inp[3]) ? node23078 : node23075;
															assign node23075 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node23078 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node23081 = (inp[0]) ? node23093 : node23082;
													assign node23082 = (inp[15]) ? node23088 : node23083;
														assign node23083 = (inp[3]) ? 4'b0001 : node23084;
															assign node23084 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node23088 = (inp[3]) ? 4'b0011 : node23089;
															assign node23089 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node23093 = (inp[15]) ? node23097 : node23094;
														assign node23094 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node23097 = (inp[3]) ? 4'b0001 : node23098;
															assign node23098 = (inp[12]) ? 4'b0011 : 4'b0001;
									assign node23102 = (inp[5]) ? node23192 : node23103;
										assign node23103 = (inp[15]) ? node23153 : node23104;
											assign node23104 = (inp[4]) ? node23124 : node23105;
												assign node23105 = (inp[0]) ? node23115 : node23106;
													assign node23106 = (inp[10]) ? 4'b0010 : node23107;
														assign node23107 = (inp[12]) ? node23111 : node23108;
															assign node23108 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node23111 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node23115 = (inp[9]) ? node23117 : 4'b0000;
														assign node23117 = (inp[3]) ? 4'b0110 : node23118;
															assign node23118 = (inp[12]) ? 4'b0100 : node23119;
																assign node23119 = (inp[10]) ? 4'b0100 : 4'b0000;
												assign node23124 = (inp[9]) ? node23134 : node23125;
													assign node23125 = (inp[10]) ? node23129 : node23126;
														assign node23126 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node23129 = (inp[0]) ? node23131 : 4'b0100;
															assign node23131 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node23134 = (inp[12]) ? node23146 : node23135;
														assign node23135 = (inp[10]) ? node23143 : node23136;
															assign node23136 = (inp[3]) ? node23140 : node23137;
																assign node23137 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node23140 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node23143 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node23146 = (inp[0]) ? node23150 : node23147;
															assign node23147 = (inp[3]) ? 4'b0000 : 4'b0010;
															assign node23150 = (inp[3]) ? 4'b0010 : 4'b0000;
											assign node23153 = (inp[0]) ? node23175 : node23154;
												assign node23154 = (inp[3]) ? node23168 : node23155;
													assign node23155 = (inp[9]) ? node23165 : node23156;
														assign node23156 = (inp[4]) ? node23162 : node23157;
															assign node23157 = (inp[10]) ? 4'b0000 : node23158;
																assign node23158 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node23162 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node23165 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node23168 = (inp[9]) ? node23170 : 4'b0000;
														assign node23170 = (inp[12]) ? node23172 : 4'b0000;
															assign node23172 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node23175 = (inp[3]) ? node23183 : node23176;
													assign node23176 = (inp[9]) ? node23178 : 4'b0010;
														assign node23178 = (inp[4]) ? node23180 : 4'b0110;
															assign node23180 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node23183 = (inp[12]) ? node23185 : 4'b0010;
														assign node23185 = (inp[9]) ? node23189 : node23186;
															assign node23186 = (inp[4]) ? 4'b0100 : 4'b0010;
															assign node23189 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node23192 = (inp[0]) ? node23222 : node23193;
											assign node23193 = (inp[15]) ? node23205 : node23194;
												assign node23194 = (inp[4]) ? node23198 : node23195;
													assign node23195 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node23198 = (inp[9]) ? node23200 : 4'b0100;
														assign node23200 = (inp[12]) ? 4'b0000 : node23201;
															assign node23201 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node23205 = (inp[9]) ? node23215 : node23206;
													assign node23206 = (inp[4]) ? 4'b0110 : node23207;
														assign node23207 = (inp[3]) ? node23211 : node23208;
															assign node23208 = (inp[12]) ? 4'b0000 : 4'b0100;
															assign node23211 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node23215 = (inp[4]) ? node23217 : 4'b0110;
														assign node23217 = (inp[12]) ? 4'b0010 : node23218;
															assign node23218 = (inp[10]) ? 4'b0010 : 4'b0110;
											assign node23222 = (inp[15]) ? node23246 : node23223;
												assign node23223 = (inp[3]) ? node23235 : node23224;
													assign node23224 = (inp[4]) ? 4'b0110 : node23225;
														assign node23225 = (inp[9]) ? node23229 : node23226;
															assign node23226 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node23229 = (inp[10]) ? 4'b0110 : node23230;
																assign node23230 = (inp[12]) ? 4'b0110 : 4'b0000;
													assign node23235 = (inp[9]) ? node23241 : node23236;
														assign node23236 = (inp[10]) ? 4'b0110 : node23237;
															assign node23237 = (inp[12]) ? 4'b0110 : 4'b0010;
														assign node23241 = (inp[4]) ? 4'b0010 : node23242;
															assign node23242 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node23246 = (inp[9]) ? node23260 : node23247;
													assign node23247 = (inp[4]) ? node23255 : node23248;
														assign node23248 = (inp[3]) ? 4'b0000 : node23249;
															assign node23249 = (inp[12]) ? 4'b0010 : node23250;
																assign node23250 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node23255 = (inp[10]) ? 4'b0100 : node23256;
															assign node23256 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node23260 = (inp[4]) ? node23262 : 4'b0100;
														assign node23262 = (inp[10]) ? 4'b0000 : node23263;
															assign node23263 = (inp[12]) ? 4'b0000 : 4'b0100;
						assign node23267 = (inp[2]) ? node24079 : node23268;
							assign node23268 = (inp[0]) ? node23652 : node23269;
								assign node23269 = (inp[15]) ? node23473 : node23270;
									assign node23270 = (inp[3]) ? node23362 : node23271;
										assign node23271 = (inp[5]) ? node23325 : node23272;
											assign node23272 = (inp[12]) ? node23298 : node23273;
												assign node23273 = (inp[7]) ? node23287 : node23274;
													assign node23274 = (inp[8]) ? node23282 : node23275;
														assign node23275 = (inp[10]) ? 4'b0011 : node23276;
															assign node23276 = (inp[9]) ? 4'b0011 : node23277;
																assign node23277 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node23282 = (inp[4]) ? 4'b0010 : node23283;
															assign node23283 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node23287 = (inp[8]) ? node23291 : node23288;
														assign node23288 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node23291 = (inp[9]) ? 4'b0011 : node23292;
															assign node23292 = (inp[10]) ? 4'b0111 : node23293;
																assign node23293 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node23298 = (inp[7]) ? node23314 : node23299;
													assign node23299 = (inp[8]) ? node23309 : node23300;
														assign node23300 = (inp[10]) ? node23302 : 4'b0111;
															assign node23302 = (inp[4]) ? node23306 : node23303;
																assign node23303 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node23306 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node23309 = (inp[10]) ? 4'b0110 : node23310;
															assign node23310 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node23314 = (inp[8]) ? node23318 : node23315;
														assign node23315 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node23318 = (inp[10]) ? node23320 : 4'b0011;
															assign node23320 = (inp[9]) ? 4'b0111 : node23321;
																assign node23321 = (inp[4]) ? 4'b0111 : 4'b0011;
											assign node23325 = (inp[9]) ? node23347 : node23326;
												assign node23326 = (inp[4]) ? node23340 : node23327;
													assign node23327 = (inp[12]) ? node23333 : node23328;
														assign node23328 = (inp[8]) ? node23330 : 4'b0010;
															assign node23330 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node23333 = (inp[8]) ? node23337 : node23334;
															assign node23334 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node23337 = (inp[7]) ? 4'b0011 : 4'b0010;
													assign node23340 = (inp[10]) ? node23344 : node23341;
														assign node23341 = (inp[12]) ? 4'b0101 : 4'b0010;
														assign node23344 = (inp[12]) ? 4'b0100 : 4'b0101;
												assign node23347 = (inp[10]) ? node23359 : node23348;
													assign node23348 = (inp[4]) ? node23350 : 4'b0011;
														assign node23350 = (inp[12]) ? node23352 : 4'b0101;
															assign node23352 = (inp[7]) ? node23356 : node23353;
																assign node23353 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node23356 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node23359 = (inp[4]) ? 4'b0000 : 4'b0100;
										assign node23362 = (inp[5]) ? node23412 : node23363;
											assign node23363 = (inp[9]) ? node23383 : node23364;
												assign node23364 = (inp[10]) ? node23374 : node23365;
													assign node23365 = (inp[7]) ? node23371 : node23366;
														assign node23366 = (inp[8]) ? node23368 : 4'b0011;
															assign node23368 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node23371 = (inp[8]) ? 4'b0011 : 4'b0100;
													assign node23374 = (inp[12]) ? node23376 : 4'b0010;
														assign node23376 = (inp[8]) ? node23380 : node23377;
															assign node23377 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node23380 = (inp[7]) ? 4'b0011 : 4'b0010;
												assign node23383 = (inp[4]) ? node23393 : node23384;
													assign node23384 = (inp[10]) ? node23388 : node23385;
														assign node23385 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node23388 = (inp[7]) ? 4'b0100 : node23389;
															assign node23389 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node23393 = (inp[10]) ? node23401 : node23394;
														assign node23394 = (inp[12]) ? node23398 : node23395;
															assign node23395 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node23398 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node23401 = (inp[12]) ? node23407 : node23402;
															assign node23402 = (inp[7]) ? node23404 : 4'b0000;
																assign node23404 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node23407 = (inp[8]) ? 4'b0001 : node23408;
																assign node23408 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node23412 = (inp[10]) ? node23448 : node23413;
												assign node23413 = (inp[8]) ? node23433 : node23414;
													assign node23414 = (inp[7]) ? node23424 : node23415;
														assign node23415 = (inp[9]) ? 4'b0101 : node23416;
															assign node23416 = (inp[4]) ? node23420 : node23417;
																assign node23417 = (inp[12]) ? 4'b0001 : 4'b0101;
																assign node23420 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node23424 = (inp[12]) ? node23426 : 4'b0100;
															assign node23426 = (inp[9]) ? node23430 : node23427;
																assign node23427 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node23430 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node23433 = (inp[7]) ? node23445 : node23434;
														assign node23434 = (inp[12]) ? node23440 : node23435;
															assign node23435 = (inp[4]) ? 4'b0000 : node23436;
																assign node23436 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node23440 = (inp[9]) ? 4'b0100 : node23441;
																assign node23441 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node23445 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node23448 = (inp[9]) ? node23464 : node23449;
													assign node23449 = (inp[4]) ? 4'b0100 : node23450;
														assign node23450 = (inp[12]) ? node23458 : node23451;
															assign node23451 = (inp[8]) ? node23455 : node23452;
																assign node23452 = (inp[7]) ? 4'b0000 : 4'b0001;
																assign node23455 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node23458 = (inp[7]) ? node23460 : 4'b0000;
																assign node23460 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node23464 = (inp[4]) ? node23470 : node23465;
														assign node23465 = (inp[7]) ? node23467 : 4'b0100;
															assign node23467 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node23470 = (inp[7]) ? 4'b0000 : 4'b0001;
									assign node23473 = (inp[5]) ? node23555 : node23474;
										assign node23474 = (inp[3]) ? node23504 : node23475;
											assign node23475 = (inp[8]) ? node23495 : node23476;
												assign node23476 = (inp[7]) ? node23484 : node23477;
													assign node23477 = (inp[4]) ? 4'b0101 : node23478;
														assign node23478 = (inp[9]) ? node23480 : 4'b0001;
															assign node23480 = (inp[12]) ? 4'b0101 : 4'b0001;
													assign node23484 = (inp[10]) ? node23490 : node23485;
														assign node23485 = (inp[9]) ? node23487 : 4'b0000;
															assign node23487 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node23490 = (inp[9]) ? node23492 : 4'b0100;
															assign node23492 = (inp[4]) ? 4'b0000 : 4'b0100;
												assign node23495 = (inp[7]) ? 4'b0001 : node23496;
													assign node23496 = (inp[9]) ? node23498 : 4'b0000;
														assign node23498 = (inp[4]) ? node23500 : 4'b0100;
															assign node23500 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node23504 = (inp[9]) ? node23536 : node23505;
												assign node23505 = (inp[4]) ? node23517 : node23506;
													assign node23506 = (inp[7]) ? node23514 : node23507;
														assign node23507 = (inp[8]) ? node23509 : 4'b0001;
															assign node23509 = (inp[10]) ? 4'b0000 : node23510;
																assign node23510 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node23514 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node23517 = (inp[12]) ? node23527 : node23518;
														assign node23518 = (inp[10]) ? node23524 : node23519;
															assign node23519 = (inp[7]) ? node23521 : 4'b0001;
																assign node23521 = (inp[8]) ? 4'b0001 : 4'b0000;
															assign node23524 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node23527 = (inp[10]) ? 4'b0110 : node23528;
															assign node23528 = (inp[7]) ? node23532 : node23529;
																assign node23529 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node23532 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node23536 = (inp[4]) ? node23544 : node23537;
													assign node23537 = (inp[8]) ? node23541 : node23538;
														assign node23538 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node23541 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node23544 = (inp[12]) ? node23550 : node23545;
														assign node23545 = (inp[7]) ? node23547 : 4'b0111;
															assign node23547 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node23550 = (inp[8]) ? node23552 : 4'b0011;
															assign node23552 = (inp[7]) ? 4'b0011 : 4'b0010;
										assign node23555 = (inp[3]) ? node23607 : node23556;
											assign node23556 = (inp[9]) ? node23582 : node23557;
												assign node23557 = (inp[4]) ? node23569 : node23558;
													assign node23558 = (inp[12]) ? node23564 : node23559;
														assign node23559 = (inp[7]) ? node23561 : 4'b0100;
															assign node23561 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node23564 = (inp[7]) ? node23566 : 4'b0000;
															assign node23566 = (inp[10]) ? 4'b0001 : 4'b0000;
													assign node23569 = (inp[12]) ? node23577 : node23570;
														assign node23570 = (inp[10]) ? 4'b0111 : node23571;
															assign node23571 = (inp[7]) ? node23573 : 4'b0001;
																assign node23573 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node23577 = (inp[8]) ? node23579 : 4'b0111;
															assign node23579 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node23582 = (inp[4]) ? node23598 : node23583;
													assign node23583 = (inp[10]) ? node23591 : node23584;
														assign node23584 = (inp[12]) ? node23586 : 4'b0001;
															assign node23586 = (inp[7]) ? 4'b0111 : node23587;
																assign node23587 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node23591 = (inp[7]) ? node23595 : node23592;
															assign node23592 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node23595 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node23598 = (inp[12]) ? node23602 : node23599;
														assign node23599 = (inp[8]) ? 4'b0011 : 4'b0111;
														assign node23602 = (inp[8]) ? 4'b0011 : node23603;
															assign node23603 = (inp[7]) ? 4'b0010 : 4'b0011;
											assign node23607 = (inp[10]) ? node23635 : node23608;
												assign node23608 = (inp[7]) ? node23626 : node23609;
													assign node23609 = (inp[8]) ? node23619 : node23610;
														assign node23610 = (inp[9]) ? 4'b0011 : node23611;
															assign node23611 = (inp[4]) ? node23615 : node23612;
																assign node23612 = (inp[12]) ? 4'b0011 : 4'b0111;
																assign node23615 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node23619 = (inp[12]) ? 4'b0110 : node23620;
															assign node23620 = (inp[9]) ? 4'b0010 : node23621;
																assign node23621 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node23626 = (inp[8]) ? 4'b0111 : node23627;
														assign node23627 = (inp[4]) ? node23631 : node23628;
															assign node23628 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node23631 = (inp[12]) ? 4'b0110 : 4'b0010;
												assign node23635 = (inp[7]) ? node23647 : node23636;
													assign node23636 = (inp[8]) ? node23642 : node23637;
														assign node23637 = (inp[4]) ? node23639 : 4'b0111;
															assign node23639 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node23642 = (inp[9]) ? 4'b0010 : node23643;
															assign node23643 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node23647 = (inp[8]) ? node23649 : 4'b0010;
														assign node23649 = (inp[4]) ? 4'b0111 : 4'b0011;
								assign node23652 = (inp[15]) ? node23870 : node23653;
									assign node23653 = (inp[3]) ? node23759 : node23654;
										assign node23654 = (inp[5]) ? node23710 : node23655;
											assign node23655 = (inp[4]) ? node23683 : node23656;
												assign node23656 = (inp[9]) ? node23668 : node23657;
													assign node23657 = (inp[12]) ? node23663 : node23658;
														assign node23658 = (inp[8]) ? 4'b0100 : node23659;
															assign node23659 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node23663 = (inp[8]) ? 4'b0000 : node23664;
															assign node23664 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node23668 = (inp[12]) ? node23672 : node23669;
														assign node23669 = (inp[7]) ? 4'b0101 : 4'b0000;
														assign node23672 = (inp[10]) ? node23678 : node23673;
															assign node23673 = (inp[8]) ? 4'b0101 : node23674;
																assign node23674 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node23678 = (inp[8]) ? 4'b0100 : node23679;
																assign node23679 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node23683 = (inp[9]) ? node23695 : node23684;
													assign node23684 = (inp[10]) ? node23690 : node23685;
														assign node23685 = (inp[7]) ? 4'b0000 : node23686;
															assign node23686 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node23690 = (inp[7]) ? node23692 : 4'b0100;
															assign node23692 = (inp[8]) ? 4'b0101 : 4'b0100;
													assign node23695 = (inp[10]) ? node23705 : node23696;
														assign node23696 = (inp[12]) ? node23702 : node23697;
															assign node23697 = (inp[7]) ? node23699 : 4'b0101;
																assign node23699 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node23702 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node23705 = (inp[8]) ? 4'b0001 : node23706;
															assign node23706 = (inp[7]) ? 4'b0000 : 4'b0001;
											assign node23710 = (inp[4]) ? node23746 : node23711;
												assign node23711 = (inp[9]) ? node23729 : node23712;
													assign node23712 = (inp[10]) ? node23722 : node23713;
														assign node23713 = (inp[12]) ? 4'b0001 : node23714;
															assign node23714 = (inp[7]) ? node23718 : node23715;
																assign node23715 = (inp[8]) ? 4'b0100 : 4'b0101;
																assign node23718 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node23722 = (inp[7]) ? node23726 : node23723;
															assign node23723 = (inp[8]) ? 4'b0000 : 4'b0001;
															assign node23726 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node23729 = (inp[12]) ? node23737 : node23730;
														assign node23730 = (inp[10]) ? 4'b0110 : node23731;
															assign node23731 = (inp[8]) ? 4'b0001 : node23732;
																assign node23732 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node23737 = (inp[10]) ? node23741 : node23738;
															assign node23738 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node23741 = (inp[8]) ? node23743 : 4'b0110;
																assign node23743 = (inp[7]) ? 4'b0111 : 4'b0110;
												assign node23746 = (inp[9]) ? node23752 : node23747;
													assign node23747 = (inp[10]) ? 4'b0110 : node23748;
														assign node23748 = (inp[8]) ? 4'b0111 : 4'b0110;
													assign node23752 = (inp[7]) ? node23754 : 4'b0010;
														assign node23754 = (inp[8]) ? node23756 : 4'b0010;
															assign node23756 = (inp[12]) ? 4'b0011 : 4'b0111;
										assign node23759 = (inp[5]) ? node23815 : node23760;
											assign node23760 = (inp[4]) ? node23786 : node23761;
												assign node23761 = (inp[9]) ? node23771 : node23762;
													assign node23762 = (inp[10]) ? node23766 : node23763;
														assign node23763 = (inp[12]) ? 4'b0000 : 4'b0100;
														assign node23766 = (inp[8]) ? node23768 : 4'b0001;
															assign node23768 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node23771 = (inp[10]) ? node23779 : node23772;
														assign node23772 = (inp[12]) ? 4'b0110 : node23773;
															assign node23773 = (inp[7]) ? 4'b0001 : node23774;
																assign node23774 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node23779 = (inp[7]) ? node23783 : node23780;
															assign node23780 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node23783 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node23786 = (inp[9]) ? node23800 : node23787;
													assign node23787 = (inp[12]) ? node23795 : node23788;
														assign node23788 = (inp[10]) ? node23792 : node23789;
															assign node23789 = (inp[7]) ? 4'b0000 : 4'b0001;
															assign node23792 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node23795 = (inp[8]) ? node23797 : 4'b0111;
															assign node23797 = (inp[7]) ? 4'b0111 : 4'b0110;
													assign node23800 = (inp[10]) ? 4'b0010 : node23801;
														assign node23801 = (inp[12]) ? node23809 : node23802;
															assign node23802 = (inp[7]) ? node23806 : node23803;
																assign node23803 = (inp[8]) ? 4'b0110 : 4'b0111;
																assign node23806 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node23809 = (inp[7]) ? node23811 : 4'b0011;
																assign node23811 = (inp[8]) ? 4'b0011 : 4'b0010;
											assign node23815 = (inp[7]) ? node23839 : node23816;
												assign node23816 = (inp[8]) ? node23828 : node23817;
													assign node23817 = (inp[4]) ? 4'b0111 : node23818;
														assign node23818 = (inp[9]) ? node23822 : node23819;
															assign node23819 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node23822 = (inp[10]) ? 4'b0111 : node23823;
																assign node23823 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node23828 = (inp[4]) ? 4'b0010 : node23829;
														assign node23829 = (inp[12]) ? 4'b0110 : node23830;
															assign node23830 = (inp[9]) ? node23834 : node23831;
																assign node23831 = (inp[10]) ? 4'b0010 : 4'b0110;
																assign node23834 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node23839 = (inp[8]) ? node23859 : node23840;
													assign node23840 = (inp[10]) ? node23850 : node23841;
														assign node23841 = (inp[9]) ? node23843 : 4'b0010;
															assign node23843 = (inp[4]) ? node23847 : node23844;
																assign node23844 = (inp[12]) ? 4'b0110 : 4'b0010;
																assign node23847 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node23850 = (inp[12]) ? node23856 : node23851;
															assign node23851 = (inp[9]) ? node23853 : 4'b0110;
																assign node23853 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node23856 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node23859 = (inp[10]) ? node23861 : 4'b0011;
														assign node23861 = (inp[12]) ? node23865 : node23862;
															assign node23862 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node23865 = (inp[9]) ? node23867 : 4'b0011;
																assign node23867 = (inp[4]) ? 4'b0011 : 4'b0111;
									assign node23870 = (inp[3]) ? node23972 : node23871;
										assign node23871 = (inp[5]) ? node23927 : node23872;
											assign node23872 = (inp[4]) ? node23896 : node23873;
												assign node23873 = (inp[9]) ? node23883 : node23874;
													assign node23874 = (inp[12]) ? node23878 : node23875;
														assign node23875 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node23878 = (inp[7]) ? 4'b0011 : node23879;
															assign node23879 = (inp[10]) ? 4'b0010 : 4'b0011;
													assign node23883 = (inp[10]) ? node23891 : node23884;
														assign node23884 = (inp[12]) ? node23886 : 4'b0011;
															assign node23886 = (inp[7]) ? 4'b0111 : node23887;
																assign node23887 = (inp[8]) ? 4'b0110 : 4'b0111;
														assign node23891 = (inp[7]) ? node23893 : 4'b0110;
															assign node23893 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node23896 = (inp[9]) ? node23912 : node23897;
													assign node23897 = (inp[10]) ? node23905 : node23898;
														assign node23898 = (inp[12]) ? node23900 : 4'b0010;
															assign node23900 = (inp[8]) ? node23902 : 4'b0110;
																assign node23902 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node23905 = (inp[12]) ? node23909 : node23906;
															assign node23906 = (inp[8]) ? 4'b0111 : 4'b0110;
															assign node23909 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node23912 = (inp[10]) ? node23920 : node23913;
														assign node23913 = (inp[12]) ? 4'b0010 : node23914;
															assign node23914 = (inp[8]) ? 4'b0111 : node23915;
																assign node23915 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node23920 = (inp[8]) ? node23924 : node23921;
															assign node23921 = (inp[7]) ? 4'b0010 : 4'b0011;
															assign node23924 = (inp[7]) ? 4'b0011 : 4'b0010;
											assign node23927 = (inp[4]) ? node23955 : node23928;
												assign node23928 = (inp[9]) ? node23942 : node23929;
													assign node23929 = (inp[12]) ? node23937 : node23930;
														assign node23930 = (inp[10]) ? 4'b0011 : node23931;
															assign node23931 = (inp[8]) ? node23933 : 4'b0110;
																assign node23933 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node23937 = (inp[8]) ? 4'b0011 : node23938;
															assign node23938 = (inp[7]) ? 4'b0010 : 4'b0011;
													assign node23942 = (inp[12]) ? node23950 : node23943;
														assign node23943 = (inp[10]) ? 4'b0101 : node23944;
															assign node23944 = (inp[8]) ? node23946 : 4'b0010;
																assign node23946 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node23950 = (inp[10]) ? 4'b0101 : node23951;
															assign node23951 = (inp[7]) ? 4'b0100 : 4'b0101;
												assign node23955 = (inp[7]) ? node23959 : node23956;
													assign node23956 = (inp[8]) ? 4'b0100 : 4'b0101;
													assign node23959 = (inp[8]) ? node23965 : node23960;
														assign node23960 = (inp[9]) ? 4'b0000 : node23961;
															assign node23961 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node23965 = (inp[12]) ? node23969 : node23966;
															assign node23966 = (inp[9]) ? 4'b0101 : 4'b0011;
															assign node23969 = (inp[9]) ? 4'b0001 : 4'b0101;
										assign node23972 = (inp[5]) ? node24026 : node23973;
											assign node23973 = (inp[9]) ? node23999 : node23974;
												assign node23974 = (inp[4]) ? node23988 : node23975;
													assign node23975 = (inp[7]) ? node23981 : node23976;
														assign node23976 = (inp[12]) ? node23978 : 4'b0111;
															assign node23978 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node23981 = (inp[8]) ? 4'b0011 : node23982;
															assign node23982 = (inp[10]) ? 4'b0010 : node23983;
																assign node23983 = (inp[12]) ? 4'b0010 : 4'b0110;
													assign node23988 = (inp[12]) ? node23996 : node23989;
														assign node23989 = (inp[10]) ? 4'b0101 : node23990;
															assign node23990 = (inp[8]) ? node23992 : 4'b0010;
																assign node23992 = (inp[7]) ? 4'b0011 : 4'b0010;
														assign node23996 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node23999 = (inp[4]) ? node24011 : node24000;
													assign node24000 = (inp[10]) ? node24006 : node24001;
														assign node24001 = (inp[12]) ? 4'b0100 : node24002;
															assign node24002 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node24006 = (inp[8]) ? node24008 : 4'b0101;
															assign node24008 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node24011 = (inp[12]) ? node24017 : node24012;
														assign node24012 = (inp[10]) ? 4'b0001 : node24013;
															assign node24013 = (inp[8]) ? 4'b0101 : 4'b0100;
														assign node24017 = (inp[10]) ? 4'b0000 : node24018;
															assign node24018 = (inp[7]) ? node24022 : node24019;
																assign node24019 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node24022 = (inp[8]) ? 4'b0001 : 4'b0000;
											assign node24026 = (inp[9]) ? node24056 : node24027;
												assign node24027 = (inp[4]) ? node24045 : node24028;
													assign node24028 = (inp[10]) ? node24036 : node24029;
														assign node24029 = (inp[12]) ? node24031 : 4'b0100;
															assign node24031 = (inp[8]) ? 4'b0000 : node24032;
																assign node24032 = (inp[7]) ? 4'b0000 : 4'b0001;
														assign node24036 = (inp[12]) ? 4'b0001 : node24037;
															assign node24037 = (inp[7]) ? node24041 : node24038;
																assign node24038 = (inp[8]) ? 4'b0000 : 4'b0001;
																assign node24041 = (inp[8]) ? 4'b0001 : 4'b0000;
													assign node24045 = (inp[10]) ? node24051 : node24046;
														assign node24046 = (inp[7]) ? 4'b0101 : node24047;
															assign node24047 = (inp[8]) ? 4'b0000 : 4'b0001;
														assign node24051 = (inp[12]) ? node24053 : 4'b0100;
															assign node24053 = (inp[8]) ? 4'b0101 : 4'b0100;
												assign node24056 = (inp[4]) ? node24066 : node24057;
													assign node24057 = (inp[8]) ? node24063 : node24058;
														assign node24058 = (inp[10]) ? 4'b0101 : node24059;
															assign node24059 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node24063 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node24066 = (inp[10]) ? node24074 : node24067;
														assign node24067 = (inp[12]) ? 4'b0001 : node24068;
															assign node24068 = (inp[7]) ? 4'b0101 : node24069;
																assign node24069 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node24074 = (inp[8]) ? node24076 : 4'b0000;
															assign node24076 = (inp[7]) ? 4'b0001 : 4'b0000;
							assign node24079 = (inp[3]) ? node24447 : node24080;
								assign node24080 = (inp[4]) ? node24256 : node24081;
									assign node24081 = (inp[9]) ? node24163 : node24082;
										assign node24082 = (inp[12]) ? node24132 : node24083;
											assign node24083 = (inp[10]) ? node24113 : node24084;
												assign node24084 = (inp[15]) ? node24100 : node24085;
													assign node24085 = (inp[0]) ? node24095 : node24086;
														assign node24086 = (inp[5]) ? node24090 : node24087;
															assign node24087 = (inp[8]) ? 4'b0110 : 4'b0111;
															assign node24090 = (inp[8]) ? node24092 : 4'b0110;
																assign node24092 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node24095 = (inp[8]) ? node24097 : 4'b0100;
															assign node24097 = (inp[7]) ? 4'b0100 : 4'b0101;
													assign node24100 = (inp[0]) ? node24108 : node24101;
														assign node24101 = (inp[7]) ? node24105 : node24102;
															assign node24102 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node24105 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node24108 = (inp[7]) ? 4'b0111 : node24109;
															assign node24109 = (inp[8]) ? 4'b0111 : 4'b0110;
												assign node24113 = (inp[7]) ? node24121 : node24114;
													assign node24114 = (inp[8]) ? 4'b0001 : node24115;
														assign node24115 = (inp[15]) ? node24117 : 4'b0000;
															assign node24117 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node24121 = (inp[8]) ? node24127 : node24122;
														assign node24122 = (inp[5]) ? node24124 : 4'b0011;
															assign node24124 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node24127 = (inp[0]) ? node24129 : 4'b0010;
															assign node24129 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node24132 = (inp[7]) ? node24152 : node24133;
												assign node24133 = (inp[8]) ? node24143 : node24134;
													assign node24134 = (inp[10]) ? 4'b0000 : node24135;
														assign node24135 = (inp[0]) ? node24139 : node24136;
															assign node24136 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node24139 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node24143 = (inp[5]) ? node24145 : 4'b0011;
														assign node24145 = (inp[10]) ? node24149 : node24146;
															assign node24146 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node24149 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node24152 = (inp[8]) ? node24158 : node24153;
													assign node24153 = (inp[0]) ? node24155 : 4'b0001;
														assign node24155 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node24158 = (inp[15]) ? 4'b0000 : node24159;
														assign node24159 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node24163 = (inp[12]) ? node24217 : node24164;
											assign node24164 = (inp[10]) ? node24188 : node24165;
												assign node24165 = (inp[0]) ? node24179 : node24166;
													assign node24166 = (inp[15]) ? node24172 : node24167;
														assign node24167 = (inp[7]) ? node24169 : 4'b0010;
															assign node24169 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node24172 = (inp[5]) ? 4'b0001 : node24173;
															assign node24173 = (inp[8]) ? 4'b0001 : node24174;
																assign node24174 = (inp[7]) ? 4'b0001 : 4'b0000;
													assign node24179 = (inp[15]) ? node24183 : node24180;
														assign node24180 = (inp[7]) ? 4'b0001 : 4'b0000;
														assign node24183 = (inp[7]) ? 4'b0010 : node24184;
															assign node24184 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node24188 = (inp[0]) ? node24202 : node24189;
													assign node24189 = (inp[15]) ? node24199 : node24190;
														assign node24190 = (inp[5]) ? 4'b0100 : node24191;
															assign node24191 = (inp[8]) ? node24195 : node24192;
																assign node24192 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node24195 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node24199 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node24202 = (inp[15]) ? node24208 : node24203;
														assign node24203 = (inp[8]) ? 4'b0100 : node24204;
															assign node24204 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node24208 = (inp[5]) ? node24214 : node24209;
															assign node24209 = (inp[8]) ? node24211 : 4'b0111;
																assign node24211 = (inp[7]) ? 4'b0110 : 4'b0111;
															assign node24214 = (inp[8]) ? 4'b0101 : 4'b0100;
											assign node24217 = (inp[5]) ? node24233 : node24218;
												assign node24218 = (inp[7]) ? node24228 : node24219;
													assign node24219 = (inp[8]) ? node24223 : node24220;
														assign node24220 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node24223 = (inp[0]) ? node24225 : 4'b0111;
															assign node24225 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node24228 = (inp[8]) ? 4'b0100 : node24229;
														assign node24229 = (inp[10]) ? 4'b0111 : 4'b0101;
												assign node24233 = (inp[0]) ? node24247 : node24234;
													assign node24234 = (inp[15]) ? node24242 : node24235;
														assign node24235 = (inp[7]) ? node24239 : node24236;
															assign node24236 = (inp[8]) ? 4'b0101 : 4'b0100;
															assign node24239 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node24242 = (inp[7]) ? node24244 : 4'b0110;
															assign node24244 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node24247 = (inp[15]) ? 4'b0100 : node24248;
														assign node24248 = (inp[10]) ? 4'b0110 : node24249;
															assign node24249 = (inp[7]) ? node24251 : 4'b0110;
																assign node24251 = (inp[8]) ? 4'b0110 : 4'b0111;
									assign node24256 = (inp[9]) ? node24352 : node24257;
										assign node24257 = (inp[10]) ? node24303 : node24258;
											assign node24258 = (inp[12]) ? node24278 : node24259;
												assign node24259 = (inp[15]) ? node24269 : node24260;
													assign node24260 = (inp[0]) ? node24262 : 4'b0011;
														assign node24262 = (inp[8]) ? node24266 : node24263;
															assign node24263 = (inp[5]) ? 4'b0000 : 4'b0001;
															assign node24266 = (inp[7]) ? 4'b0000 : 4'b0001;
													assign node24269 = (inp[0]) ? node24275 : node24270;
														assign node24270 = (inp[7]) ? 4'b0000 : node24271;
															assign node24271 = (inp[8]) ? 4'b0001 : 4'b0000;
														assign node24275 = (inp[8]) ? 4'b0011 : 4'b0010;
												assign node24278 = (inp[7]) ? node24292 : node24279;
													assign node24279 = (inp[8]) ? node24281 : 4'b0100;
														assign node24281 = (inp[0]) ? node24287 : node24282;
															assign node24282 = (inp[5]) ? 4'b0111 : node24283;
																assign node24283 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node24287 = (inp[5]) ? 4'b0101 : node24288;
																assign node24288 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node24292 = (inp[8]) ? node24296 : node24293;
														assign node24293 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node24296 = (inp[15]) ? 4'b0110 : node24297;
															assign node24297 = (inp[5]) ? node24299 : 4'b0100;
																assign node24299 = (inp[0]) ? 4'b0110 : 4'b0100;
											assign node24303 = (inp[0]) ? node24323 : node24304;
												assign node24304 = (inp[8]) ? node24312 : node24305;
													assign node24305 = (inp[7]) ? 4'b0101 : node24306;
														assign node24306 = (inp[15]) ? node24308 : 4'b0100;
															assign node24308 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node24312 = (inp[7]) ? node24320 : node24313;
														assign node24313 = (inp[15]) ? node24317 : node24314;
															assign node24314 = (inp[12]) ? 4'b0111 : 4'b0101;
															assign node24317 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node24320 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node24323 = (inp[5]) ? node24341 : node24324;
													assign node24324 = (inp[15]) ? node24336 : node24325;
														assign node24325 = (inp[12]) ? node24331 : node24326;
															assign node24326 = (inp[8]) ? 4'b0101 : node24327;
																assign node24327 = (inp[7]) ? 4'b0101 : 4'b0100;
															assign node24331 = (inp[8]) ? node24333 : 4'b0100;
																assign node24333 = (inp[7]) ? 4'b0100 : 4'b0101;
														assign node24336 = (inp[7]) ? node24338 : 4'b0110;
															assign node24338 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node24341 = (inp[15]) ? node24349 : node24342;
														assign node24342 = (inp[12]) ? 4'b0111 : node24343;
															assign node24343 = (inp[8]) ? node24345 : 4'b0110;
																assign node24345 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node24349 = (inp[7]) ? 4'b0100 : 4'b0101;
										assign node24352 = (inp[10]) ? node24404 : node24353;
											assign node24353 = (inp[12]) ? node24379 : node24354;
												assign node24354 = (inp[0]) ? node24366 : node24355;
													assign node24355 = (inp[15]) ? node24363 : node24356;
														assign node24356 = (inp[5]) ? node24358 : 4'b0111;
															assign node24358 = (inp[7]) ? node24360 : 4'b0101;
																assign node24360 = (inp[8]) ? 4'b0100 : 4'b0101;
														assign node24363 = (inp[7]) ? 4'b0101 : 4'b0100;
													assign node24366 = (inp[8]) ? node24374 : node24367;
														assign node24367 = (inp[15]) ? node24371 : node24368;
															assign node24368 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node24371 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node24374 = (inp[5]) ? node24376 : 4'b0101;
															assign node24376 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node24379 = (inp[7]) ? node24393 : node24380;
													assign node24380 = (inp[8]) ? node24386 : node24381;
														assign node24381 = (inp[15]) ? node24383 : 4'b0010;
															assign node24383 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node24386 = (inp[0]) ? 4'b0011 : node24387;
															assign node24387 = (inp[15]) ? 4'b0001 : node24388;
																assign node24388 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node24393 = (inp[8]) ? node24395 : 4'b0011;
														assign node24395 = (inp[5]) ? 4'b0000 : node24396;
															assign node24396 = (inp[0]) ? node24400 : node24397;
																assign node24397 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node24400 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node24404 = (inp[15]) ? node24426 : node24405;
												assign node24405 = (inp[12]) ? node24415 : node24406;
													assign node24406 = (inp[7]) ? node24412 : node24407;
														assign node24407 = (inp[0]) ? node24409 : 4'b0000;
															assign node24409 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node24412 = (inp[8]) ? 4'b0010 : 4'b0011;
													assign node24415 = (inp[7]) ? node24423 : node24416;
														assign node24416 = (inp[5]) ? node24420 : node24417;
															assign node24417 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node24420 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node24423 = (inp[8]) ? 4'b0000 : 4'b0001;
												assign node24426 = (inp[7]) ? node24436 : node24427;
													assign node24427 = (inp[8]) ? 4'b0011 : node24428;
														assign node24428 = (inp[0]) ? node24432 : node24429;
															assign node24429 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node24432 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node24436 = (inp[8]) ? node24440 : node24437;
														assign node24437 = (inp[12]) ? 4'b0011 : 4'b0001;
														assign node24440 = (inp[0]) ? node24444 : node24441;
															assign node24441 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node24444 = (inp[5]) ? 4'b0000 : 4'b0010;
								assign node24447 = (inp[10]) ? node24691 : node24448;
									assign node24448 = (inp[5]) ? node24568 : node24449;
										assign node24449 = (inp[7]) ? node24505 : node24450;
											assign node24450 = (inp[8]) ? node24478 : node24451;
												assign node24451 = (inp[15]) ? node24469 : node24452;
													assign node24452 = (inp[12]) ? node24460 : node24453;
														assign node24453 = (inp[4]) ? node24457 : node24454;
															assign node24454 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node24457 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node24460 = (inp[0]) ? node24464 : node24461;
															assign node24461 = (inp[9]) ? 4'b0100 : 4'b0010;
															assign node24464 = (inp[9]) ? node24466 : 4'b0110;
																assign node24466 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node24469 = (inp[4]) ? node24471 : 4'b0010;
														assign node24471 = (inp[0]) ? node24475 : node24472;
															assign node24472 = (inp[9]) ? 4'b0010 : 4'b0000;
															assign node24475 = (inp[12]) ? 4'b0000 : 4'b0010;
												assign node24478 = (inp[12]) ? node24496 : node24479;
													assign node24479 = (inp[0]) ? node24487 : node24480;
														assign node24480 = (inp[15]) ? node24484 : node24481;
															assign node24481 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node24484 = (inp[9]) ? 4'b0111 : 4'b0101;
														assign node24487 = (inp[9]) ? node24491 : node24488;
															assign node24488 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node24491 = (inp[4]) ? node24493 : 4'b0011;
																assign node24493 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node24496 = (inp[0]) ? node24498 : 4'b0011;
														assign node24498 = (inp[4]) ? node24502 : node24499;
															assign node24499 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node24502 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node24505 = (inp[8]) ? node24541 : node24506;
												assign node24506 = (inp[12]) ? node24526 : node24507;
													assign node24507 = (inp[9]) ? node24521 : node24508;
														assign node24508 = (inp[4]) ? node24516 : node24509;
															assign node24509 = (inp[15]) ? node24513 : node24510;
																assign node24510 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node24513 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node24516 = (inp[15]) ? node24518 : 4'b0011;
																assign node24518 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node24521 = (inp[4]) ? 4'b0101 : node24522;
															assign node24522 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node24526 = (inp[0]) ? node24532 : node24527;
														assign node24527 = (inp[4]) ? node24529 : 4'b0011;
															assign node24529 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node24532 = (inp[9]) ? node24538 : node24533;
															assign node24533 = (inp[4]) ? 4'b0111 : node24534;
																assign node24534 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node24538 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node24541 = (inp[9]) ? node24555 : node24542;
													assign node24542 = (inp[15]) ? node24550 : node24543;
														assign node24543 = (inp[4]) ? node24547 : node24544;
															assign node24544 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node24547 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node24550 = (inp[12]) ? 4'b0100 : node24551;
															assign node24551 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node24555 = (inp[0]) ? node24563 : node24556;
														assign node24556 = (inp[15]) ? node24558 : 4'b0010;
															assign node24558 = (inp[4]) ? node24560 : 4'b0110;
																assign node24560 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node24563 = (inp[4]) ? 4'b0110 : node24564;
															assign node24564 = (inp[15]) ? 4'b0100 : 4'b0000;
										assign node24568 = (inp[4]) ? node24646 : node24569;
											assign node24569 = (inp[9]) ? node24609 : node24570;
												assign node24570 = (inp[12]) ? node24592 : node24571;
													assign node24571 = (inp[15]) ? node24583 : node24572;
														assign node24572 = (inp[0]) ? node24580 : node24573;
															assign node24573 = (inp[8]) ? node24577 : node24574;
																assign node24574 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node24577 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node24580 = (inp[7]) ? 4'b0111 : 4'b0110;
														assign node24583 = (inp[0]) ? 4'b0100 : node24584;
															assign node24584 = (inp[7]) ? node24588 : node24585;
																assign node24585 = (inp[8]) ? 4'b0111 : 4'b0110;
																assign node24588 = (inp[8]) ? 4'b0110 : 4'b0111;
													assign node24592 = (inp[7]) ? node24598 : node24593;
														assign node24593 = (inp[8]) ? node24595 : 4'b0010;
															assign node24595 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node24598 = (inp[8]) ? node24604 : node24599;
															assign node24599 = (inp[0]) ? node24601 : 4'b0001;
																assign node24601 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node24604 = (inp[0]) ? node24606 : 4'b0010;
																assign node24606 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node24609 = (inp[12]) ? node24625 : node24610;
													assign node24610 = (inp[15]) ? node24622 : node24611;
														assign node24611 = (inp[0]) ? node24615 : node24612;
															assign node24612 = (inp[7]) ? 4'b0001 : 4'b0000;
															assign node24615 = (inp[7]) ? node24619 : node24616;
																assign node24616 = (inp[8]) ? 4'b0011 : 4'b0010;
																assign node24619 = (inp[8]) ? 4'b0010 : 4'b0011;
														assign node24622 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node24625 = (inp[15]) ? node24637 : node24626;
														assign node24626 = (inp[0]) ? node24630 : node24627;
															assign node24627 = (inp[7]) ? 4'b0100 : 4'b0101;
															assign node24630 = (inp[8]) ? node24634 : node24631;
																assign node24631 = (inp[7]) ? 4'b0111 : 4'b0110;
																assign node24634 = (inp[7]) ? 4'b0110 : 4'b0111;
														assign node24637 = (inp[0]) ? node24639 : 4'b0111;
															assign node24639 = (inp[8]) ? node24643 : node24640;
																assign node24640 = (inp[7]) ? 4'b0101 : 4'b0100;
																assign node24643 = (inp[7]) ? 4'b0100 : 4'b0101;
											assign node24646 = (inp[9]) ? node24670 : node24647;
												assign node24647 = (inp[12]) ? node24659 : node24648;
													assign node24648 = (inp[15]) ? node24656 : node24649;
														assign node24649 = (inp[0]) ? node24651 : 4'b0001;
															assign node24651 = (inp[8]) ? node24653 : 4'b0011;
																assign node24653 = (inp[7]) ? 4'b0010 : 4'b0011;
														assign node24656 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node24659 = (inp[0]) ? node24663 : node24660;
														assign node24660 = (inp[15]) ? 4'b0111 : 4'b0100;
														assign node24663 = (inp[15]) ? node24665 : 4'b0111;
															assign node24665 = (inp[8]) ? 4'b0101 : node24666;
																assign node24666 = (inp[7]) ? 4'b0101 : 4'b0100;
												assign node24670 = (inp[12]) ? node24686 : node24671;
													assign node24671 = (inp[0]) ? node24683 : node24672;
														assign node24672 = (inp[15]) ? node24678 : node24673;
															assign node24673 = (inp[7]) ? node24675 : 4'b0101;
																assign node24675 = (inp[8]) ? 4'b0100 : 4'b0101;
															assign node24678 = (inp[7]) ? 4'b0111 : node24679;
																assign node24679 = (inp[8]) ? 4'b0111 : 4'b0110;
														assign node24683 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node24686 = (inp[15]) ? 4'b0011 : node24687;
														assign node24687 = (inp[0]) ? 4'b0011 : 4'b0001;
									assign node24691 = (inp[7]) ? node24805 : node24692;
										assign node24692 = (inp[8]) ? node24764 : node24693;
											assign node24693 = (inp[12]) ? node24739 : node24694;
												assign node24694 = (inp[5]) ? node24716 : node24695;
													assign node24695 = (inp[15]) ? node24705 : node24696;
														assign node24696 = (inp[9]) ? node24702 : node24697;
															assign node24697 = (inp[4]) ? 4'b0110 : node24698;
																assign node24698 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node24702 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node24705 = (inp[0]) ? node24711 : node24706;
															assign node24706 = (inp[9]) ? node24708 : 4'b0110;
																assign node24708 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node24711 = (inp[4]) ? 4'b0100 : node24712;
																assign node24712 = (inp[9]) ? 4'b0100 : 4'b0010;
													assign node24716 = (inp[15]) ? node24728 : node24717;
														assign node24717 = (inp[0]) ? node24725 : node24718;
															assign node24718 = (inp[9]) ? node24722 : node24719;
																assign node24719 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node24722 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node24725 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node24728 = (inp[0]) ? node24732 : node24729;
															assign node24729 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node24732 = (inp[4]) ? node24736 : node24733;
																assign node24733 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node24736 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node24739 = (inp[4]) ? node24753 : node24740;
													assign node24740 = (inp[9]) ? 4'b0100 : node24741;
														assign node24741 = (inp[5]) ? node24747 : node24742;
															assign node24742 = (inp[0]) ? node24744 : 4'b0010;
																assign node24744 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node24747 = (inp[0]) ? node24749 : 4'b0000;
																assign node24749 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node24753 = (inp[9]) ? node24759 : node24754;
														assign node24754 = (inp[15]) ? node24756 : 4'b0100;
															assign node24756 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node24759 = (inp[0]) ? node24761 : 4'b0010;
															assign node24761 = (inp[15]) ? 4'b0000 : 4'b0010;
											assign node24764 = (inp[9]) ? node24788 : node24765;
												assign node24765 = (inp[4]) ? node24781 : node24766;
													assign node24766 = (inp[5]) ? node24776 : node24767;
														assign node24767 = (inp[12]) ? 4'b0001 : node24768;
															assign node24768 = (inp[0]) ? node24772 : node24769;
																assign node24769 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node24772 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node24776 = (inp[12]) ? 4'b0011 : node24777;
															assign node24777 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node24781 = (inp[5]) ? 4'b0111 : node24782;
														assign node24782 = (inp[15]) ? 4'b0101 : node24783;
															assign node24783 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node24788 = (inp[4]) ? node24802 : node24789;
													assign node24789 = (inp[5]) ? node24795 : node24790;
														assign node24790 = (inp[15]) ? node24792 : 4'b0101;
															assign node24792 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node24795 = (inp[0]) ? node24799 : node24796;
															assign node24796 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node24799 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node24802 = (inp[5]) ? 4'b0001 : 4'b0011;
										assign node24805 = (inp[8]) ? node24839 : node24806;
											assign node24806 = (inp[0]) ? node24824 : node24807;
												assign node24807 = (inp[15]) ? node24817 : node24808;
													assign node24808 = (inp[9]) ? node24814 : node24809;
														assign node24809 = (inp[5]) ? node24811 : 4'b0011;
															assign node24811 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node24814 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node24817 = (inp[4]) ? node24821 : node24818;
														assign node24818 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node24821 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node24824 = (inp[15]) ? node24832 : node24825;
													assign node24825 = (inp[9]) ? 4'b0111 : node24826;
														assign node24826 = (inp[4]) ? 4'b0111 : node24827;
															assign node24827 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node24832 = (inp[4]) ? node24836 : node24833;
														assign node24833 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node24836 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node24839 = (inp[9]) ? node24851 : node24840;
												assign node24840 = (inp[4]) ? node24846 : node24841;
													assign node24841 = (inp[12]) ? node24843 : 4'b0000;
														assign node24843 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node24846 = (inp[0]) ? node24848 : 4'b0100;
														assign node24848 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node24851 = (inp[4]) ? node24859 : node24852;
													assign node24852 = (inp[12]) ? node24856 : node24853;
														assign node24853 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node24856 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node24859 = (inp[0]) ? node24861 : 4'b0000;
														assign node24861 = (inp[15]) ? 4'b0000 : 4'b0010;
		assign node24864 = (inp[8]) ? node33612 : node24865;
			assign node24865 = (inp[7]) ? node29327 : node24866;
				assign node24866 = (inp[6]) ? node27198 : node24867;
					assign node24867 = (inp[11]) ? node26051 : node24868;
						assign node24868 = (inp[1]) ? node25392 : node24869;
							assign node24869 = (inp[5]) ? node25041 : node24870;
								assign node24870 = (inp[4]) ? node24934 : node24871;
									assign node24871 = (inp[9]) ? node24911 : node24872;
										assign node24872 = (inp[12]) ? node24880 : node24873;
											assign node24873 = (inp[0]) ? node24877 : node24874;
												assign node24874 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node24877 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node24880 = (inp[10]) ? node24896 : node24881;
												assign node24881 = (inp[2]) ? node24887 : node24882;
													assign node24882 = (inp[15]) ? 4'b1110 : node24883;
														assign node24883 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node24887 = (inp[13]) ? node24889 : 4'b1100;
														assign node24889 = (inp[0]) ? node24893 : node24890;
															assign node24890 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node24893 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node24896 = (inp[2]) ? node24902 : node24897;
													assign node24897 = (inp[0]) ? node24899 : 4'b1000;
														assign node24899 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node24902 = (inp[13]) ? node24904 : 4'b1010;
														assign node24904 = (inp[0]) ? node24908 : node24905;
															assign node24905 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node24908 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node24911 = (inp[12]) ? node24919 : node24912;
											assign node24912 = (inp[0]) ? node24916 : node24913;
												assign node24913 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node24916 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node24919 = (inp[10]) ? node24927 : node24920;
												assign node24920 = (inp[0]) ? node24924 : node24921;
													assign node24921 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node24924 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node24927 = (inp[3]) ? node24929 : 4'b1100;
													assign node24929 = (inp[0]) ? 4'b1110 : node24930;
														assign node24930 = (inp[15]) ? 4'b1110 : 4'b1100;
									assign node24934 = (inp[9]) ? node24978 : node24935;
										assign node24935 = (inp[12]) ? node24943 : node24936;
											assign node24936 = (inp[0]) ? node24940 : node24937;
												assign node24937 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node24940 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node24943 = (inp[10]) ? node24963 : node24944;
												assign node24944 = (inp[2]) ? node24952 : node24945;
													assign node24945 = (inp[0]) ? node24949 : node24946;
														assign node24946 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node24949 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node24952 = (inp[3]) ? 4'b1010 : node24953;
														assign node24953 = (inp[13]) ? node24959 : node24954;
															assign node24954 = (inp[15]) ? node24956 : 4'b1010;
																assign node24956 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node24959 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node24963 = (inp[0]) ? node24971 : node24964;
													assign node24964 = (inp[2]) ? node24966 : 4'b1110;
														assign node24966 = (inp[3]) ? node24968 : 4'b1110;
															assign node24968 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node24971 = (inp[13]) ? node24973 : 4'b1100;
														assign node24973 = (inp[15]) ? node24975 : 4'b1110;
															assign node24975 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node24978 = (inp[12]) ? node25006 : node24979;
											assign node24979 = (inp[10]) ? node24991 : node24980;
												assign node24980 = (inp[3]) ? 4'b1100 : node24981;
													assign node24981 = (inp[2]) ? node24985 : node24982;
														assign node24982 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node24985 = (inp[0]) ? node24987 : 4'b1100;
															assign node24987 = (inp[13]) ? 4'b1100 : 4'b1110;
												assign node24991 = (inp[15]) ? node24999 : node24992;
													assign node24992 = (inp[0]) ? node24996 : node24993;
														assign node24993 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node24996 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node24999 = (inp[0]) ? node25003 : node25000;
														assign node25000 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node25003 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node25006 = (inp[10]) ? node25024 : node25007;
												assign node25007 = (inp[0]) ? node25015 : node25008;
													assign node25008 = (inp[15]) ? node25012 : node25009;
														assign node25009 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node25012 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node25015 = (inp[13]) ? node25017 : 4'b1100;
														assign node25017 = (inp[2]) ? node25019 : 4'b1110;
															assign node25019 = (inp[3]) ? node25021 : 4'b1100;
																assign node25021 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node25024 = (inp[13]) ? node25032 : node25025;
													assign node25025 = (inp[3]) ? 4'b1010 : node25026;
														assign node25026 = (inp[0]) ? 4'b1010 : node25027;
															assign node25027 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node25032 = (inp[2]) ? node25034 : 4'b1000;
														assign node25034 = (inp[3]) ? node25036 : 4'b1010;
															assign node25036 = (inp[0]) ? node25038 : 4'b1000;
																assign node25038 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node25041 = (inp[3]) ? node25231 : node25042;
									assign node25042 = (inp[10]) ? node25124 : node25043;
										assign node25043 = (inp[2]) ? node25079 : node25044;
											assign node25044 = (inp[13]) ? node25062 : node25045;
												assign node25045 = (inp[12]) ? node25053 : node25046;
													assign node25046 = (inp[15]) ? node25050 : node25047;
														assign node25047 = (inp[4]) ? 4'b1110 : 4'b1100;
														assign node25050 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node25053 = (inp[9]) ? node25059 : node25054;
														assign node25054 = (inp[0]) ? node25056 : 4'b1100;
															assign node25056 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node25059 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node25062 = (inp[12]) ? node25070 : node25063;
													assign node25063 = (inp[4]) ? node25065 : 4'b1100;
														assign node25065 = (inp[15]) ? 4'b1000 : node25066;
															assign node25066 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node25070 = (inp[9]) ? node25074 : node25071;
														assign node25071 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node25074 = (inp[4]) ? 4'b1100 : node25075;
															assign node25075 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node25079 = (inp[9]) ? node25099 : node25080;
												assign node25080 = (inp[4]) ? node25094 : node25081;
													assign node25081 = (inp[13]) ? node25089 : node25082;
														assign node25082 = (inp[0]) ? node25086 : node25083;
															assign node25083 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node25086 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node25089 = (inp[0]) ? node25091 : 4'b1110;
															assign node25091 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node25094 = (inp[12]) ? node25096 : 4'b1000;
														assign node25096 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node25099 = (inp[4]) ? node25111 : node25100;
													assign node25100 = (inp[13]) ? node25106 : node25101;
														assign node25101 = (inp[0]) ? node25103 : 4'b1010;
															assign node25103 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node25106 = (inp[15]) ? node25108 : 4'b1000;
															assign node25108 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node25111 = (inp[13]) ? node25117 : node25112;
														assign node25112 = (inp[0]) ? node25114 : 4'b1110;
															assign node25114 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node25117 = (inp[15]) ? node25121 : node25118;
															assign node25118 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node25121 = (inp[0]) ? 4'b1100 : 4'b1110;
										assign node25124 = (inp[13]) ? node25160 : node25125;
											assign node25125 = (inp[12]) ? node25147 : node25126;
												assign node25126 = (inp[2]) ? node25138 : node25127;
													assign node25127 = (inp[9]) ? node25131 : node25128;
														assign node25128 = (inp[4]) ? 4'b1010 : 4'b1100;
														assign node25131 = (inp[4]) ? node25133 : 4'b1010;
															assign node25133 = (inp[0]) ? node25135 : 4'b1100;
																assign node25135 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node25138 = (inp[15]) ? 4'b1110 : node25139;
														assign node25139 = (inp[4]) ? 4'b1110 : node25140;
															assign node25140 = (inp[9]) ? 4'b1000 : node25141;
																assign node25141 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node25147 = (inp[4]) ? node25151 : node25148;
													assign node25148 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node25151 = (inp[9]) ? node25155 : node25152;
														assign node25152 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node25155 = (inp[0]) ? node25157 : 4'b1010;
															assign node25157 = (inp[2]) ? 4'b1000 : 4'b1010;
											assign node25160 = (inp[2]) ? node25198 : node25161;
												assign node25161 = (inp[15]) ? node25181 : node25162;
													assign node25162 = (inp[9]) ? node25174 : node25163;
														assign node25163 = (inp[0]) ? node25169 : node25164;
															assign node25164 = (inp[12]) ? 4'b1100 : node25165;
																assign node25165 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node25169 = (inp[12]) ? 4'b1000 : node25170;
																assign node25170 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node25174 = (inp[12]) ? node25178 : node25175;
															assign node25175 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node25178 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node25181 = (inp[9]) ? 4'b1100 : node25182;
														assign node25182 = (inp[0]) ? node25190 : node25183;
															assign node25183 = (inp[12]) ? node25187 : node25184;
																assign node25184 = (inp[4]) ? 4'b1000 : 4'b1100;
																assign node25187 = (inp[4]) ? 4'b1110 : 4'b1000;
															assign node25190 = (inp[4]) ? node25194 : node25191;
																assign node25191 = (inp[12]) ? 4'b1010 : 4'b1110;
																assign node25194 = (inp[12]) ? 4'b1100 : 4'b1010;
												assign node25198 = (inp[0]) ? node25214 : node25199;
													assign node25199 = (inp[12]) ? node25211 : node25200;
														assign node25200 = (inp[9]) ? node25204 : node25201;
															assign node25201 = (inp[4]) ? 4'b1010 : 4'b1110;
															assign node25204 = (inp[4]) ? node25208 : node25205;
																assign node25205 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node25208 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node25211 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node25214 = (inp[12]) ? node25224 : node25215;
														assign node25215 = (inp[15]) ? node25217 : 4'b1110;
															assign node25217 = (inp[4]) ? node25221 : node25218;
																assign node25218 = (inp[9]) ? 4'b1010 : 4'b1110;
																assign node25221 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node25224 = (inp[15]) ? 4'b1000 : node25225;
															assign node25225 = (inp[4]) ? node25227 : 4'b1000;
																assign node25227 = (inp[9]) ? 4'b1010 : 4'b1110;
									assign node25231 = (inp[13]) ? node25317 : node25232;
										assign node25232 = (inp[15]) ? node25268 : node25233;
											assign node25233 = (inp[0]) ? node25245 : node25234;
												assign node25234 = (inp[9]) ? node25238 : node25235;
													assign node25235 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node25238 = (inp[4]) ? node25240 : 4'b1000;
														assign node25240 = (inp[10]) ? node25242 : 4'b1100;
															assign node25242 = (inp[2]) ? 4'b1000 : 4'b1100;
												assign node25245 = (inp[12]) ? node25253 : node25246;
													assign node25246 = (inp[2]) ? node25248 : 4'b1110;
														assign node25248 = (inp[9]) ? node25250 : 4'b1110;
															assign node25250 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node25253 = (inp[9]) ? node25263 : node25254;
														assign node25254 = (inp[2]) ? node25260 : node25255;
															assign node25255 = (inp[4]) ? node25257 : 4'b1010;
																assign node25257 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node25260 = (inp[10]) ? 4'b1010 : 4'b1110;
														assign node25263 = (inp[4]) ? node25265 : 4'b1110;
															assign node25265 = (inp[2]) ? 4'b1010 : 4'b1110;
											assign node25268 = (inp[0]) ? node25288 : node25269;
												assign node25269 = (inp[10]) ? node25275 : node25270;
													assign node25270 = (inp[4]) ? 4'b1010 : node25271;
														assign node25271 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node25275 = (inp[2]) ? node25281 : node25276;
														assign node25276 = (inp[12]) ? 4'b1110 : node25277;
															assign node25277 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node25281 = (inp[12]) ? 4'b1010 : node25282;
															assign node25282 = (inp[4]) ? 4'b1110 : node25283;
																assign node25283 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node25288 = (inp[12]) ? node25306 : node25289;
													assign node25289 = (inp[2]) ? node25295 : node25290;
														assign node25290 = (inp[4]) ? node25292 : 4'b1000;
															assign node25292 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node25295 = (inp[10]) ? node25301 : node25296;
															assign node25296 = (inp[4]) ? node25298 : 4'b1000;
																assign node25298 = (inp[9]) ? 4'b1100 : 4'b1000;
															assign node25301 = (inp[4]) ? 4'b1000 : node25302;
																assign node25302 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node25306 = (inp[4]) ? node25314 : node25307;
														assign node25307 = (inp[10]) ? node25311 : node25308;
															assign node25308 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node25311 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node25314 = (inp[2]) ? 4'b1100 : 4'b1000;
										assign node25317 = (inp[10]) ? node25343 : node25318;
											assign node25318 = (inp[4]) ? node25334 : node25319;
												assign node25319 = (inp[9]) ? node25325 : node25320;
													assign node25320 = (inp[0]) ? 4'b1110 : node25321;
														assign node25321 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node25325 = (inp[12]) ? node25327 : 4'b1010;
														assign node25327 = (inp[15]) ? node25331 : node25328;
															assign node25328 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node25331 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node25334 = (inp[9]) ? node25336 : 4'b1010;
													assign node25336 = (inp[12]) ? 4'b1110 : node25337;
														assign node25337 = (inp[0]) ? 4'b1110 : node25338;
															assign node25338 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node25343 = (inp[12]) ? node25365 : node25344;
												assign node25344 = (inp[15]) ? node25354 : node25345;
													assign node25345 = (inp[0]) ? node25351 : node25346;
														assign node25346 = (inp[4]) ? node25348 : 4'b1100;
															assign node25348 = (inp[9]) ? 4'b1100 : 4'b1000;
														assign node25351 = (inp[2]) ? 4'b1110 : 4'b1010;
													assign node25354 = (inp[0]) ? node25358 : node25355;
														assign node25355 = (inp[2]) ? 4'b1010 : 4'b1110;
														assign node25358 = (inp[4]) ? node25362 : node25359;
															assign node25359 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node25362 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node25365 = (inp[2]) ? node25381 : node25366;
													assign node25366 = (inp[15]) ? node25378 : node25367;
														assign node25367 = (inp[0]) ? node25375 : node25368;
															assign node25368 = (inp[9]) ? node25372 : node25369;
																assign node25369 = (inp[4]) ? 4'b1100 : 4'b1000;
																assign node25372 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node25375 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node25378 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node25381 = (inp[0]) ? node25385 : node25382;
														assign node25382 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node25385 = (inp[9]) ? node25389 : node25386;
															assign node25386 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node25389 = (inp[4]) ? 4'b1000 : 4'b1100;
							assign node25392 = (inp[13]) ? node25680 : node25393;
								assign node25393 = (inp[9]) ? node25541 : node25394;
									assign node25394 = (inp[4]) ? node25454 : node25395;
										assign node25395 = (inp[12]) ? node25419 : node25396;
											assign node25396 = (inp[15]) ? node25408 : node25397;
												assign node25397 = (inp[0]) ? node25403 : node25398;
													assign node25398 = (inp[3]) ? node25400 : 4'b1110;
														assign node25400 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node25403 = (inp[5]) ? node25405 : 4'b1100;
														assign node25405 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node25408 = (inp[0]) ? node25414 : node25409;
													assign node25409 = (inp[3]) ? node25411 : 4'b1100;
														assign node25411 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node25414 = (inp[3]) ? node25416 : 4'b1110;
														assign node25416 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node25419 = (inp[10]) ? node25439 : node25420;
												assign node25420 = (inp[0]) ? node25430 : node25421;
													assign node25421 = (inp[5]) ? node25423 : 4'b1110;
														assign node25423 = (inp[3]) ? node25427 : node25424;
															assign node25424 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node25427 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node25430 = (inp[3]) ? node25432 : 4'b1100;
														assign node25432 = (inp[5]) ? node25436 : node25433;
															assign node25433 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node25436 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node25439 = (inp[3]) ? node25447 : node25440;
													assign node25440 = (inp[5]) ? 4'b1010 : node25441;
														assign node25441 = (inp[15]) ? 4'b1000 : node25442;
															assign node25442 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node25447 = (inp[15]) ? 4'b1010 : node25448;
														assign node25448 = (inp[5]) ? node25450 : 4'b1010;
															assign node25450 = (inp[0]) ? 4'b1010 : 4'b1000;
										assign node25454 = (inp[12]) ? node25490 : node25455;
											assign node25455 = (inp[5]) ? node25475 : node25456;
												assign node25456 = (inp[2]) ? node25470 : node25457;
													assign node25457 = (inp[3]) ? node25465 : node25458;
														assign node25458 = (inp[10]) ? node25460 : 4'b1000;
															assign node25460 = (inp[0]) ? node25462 : 4'b1000;
																assign node25462 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node25465 = (inp[15]) ? 4'b1000 : node25466;
															assign node25466 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node25470 = (inp[0]) ? 4'b1010 : node25471;
														assign node25471 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node25475 = (inp[15]) ? node25483 : node25476;
													assign node25476 = (inp[2]) ? node25478 : 4'b1000;
														assign node25478 = (inp[3]) ? node25480 : 4'b1000;
															assign node25480 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node25483 = (inp[3]) ? node25487 : node25484;
														assign node25484 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node25487 = (inp[0]) ? 4'b1000 : 4'b1010;
											assign node25490 = (inp[10]) ? node25512 : node25491;
												assign node25491 = (inp[2]) ? node25493 : 4'b1010;
													assign node25493 = (inp[3]) ? node25503 : node25494;
														assign node25494 = (inp[5]) ? node25498 : node25495;
															assign node25495 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node25498 = (inp[15]) ? node25500 : 4'b1000;
																assign node25500 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node25503 = (inp[15]) ? 4'b1010 : node25504;
															assign node25504 = (inp[5]) ? node25508 : node25505;
																assign node25505 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node25508 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node25512 = (inp[3]) ? node25526 : node25513;
													assign node25513 = (inp[15]) ? node25519 : node25514;
														assign node25514 = (inp[5]) ? node25516 : 4'b1100;
															assign node25516 = (inp[2]) ? 4'b1110 : 4'b1100;
														assign node25519 = (inp[5]) ? node25523 : node25520;
															assign node25520 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node25523 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node25526 = (inp[5]) ? node25532 : node25527;
														assign node25527 = (inp[15]) ? node25529 : 4'b1110;
															assign node25529 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node25532 = (inp[2]) ? node25534 : 4'b1100;
															assign node25534 = (inp[0]) ? node25538 : node25535;
																assign node25535 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node25538 = (inp[15]) ? 4'b1100 : 4'b1110;
									assign node25541 = (inp[4]) ? node25605 : node25542;
										assign node25542 = (inp[12]) ? node25566 : node25543;
											assign node25543 = (inp[15]) ? node25555 : node25544;
												assign node25544 = (inp[0]) ? node25550 : node25545;
													assign node25545 = (inp[3]) ? node25547 : 4'b1010;
														assign node25547 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node25550 = (inp[3]) ? node25552 : 4'b1000;
														assign node25552 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node25555 = (inp[0]) ? node25561 : node25556;
													assign node25556 = (inp[5]) ? node25558 : 4'b1000;
														assign node25558 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node25561 = (inp[3]) ? node25563 : 4'b1010;
														assign node25563 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node25566 = (inp[10]) ? node25580 : node25567;
												assign node25567 = (inp[3]) ? node25573 : node25568;
													assign node25568 = (inp[0]) ? 4'b1010 : node25569;
														assign node25569 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node25573 = (inp[5]) ? 4'b1010 : node25574;
														assign node25574 = (inp[15]) ? node25576 : 4'b1000;
															assign node25576 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node25580 = (inp[2]) ? node25598 : node25581;
													assign node25581 = (inp[5]) ? node25591 : node25582;
														assign node25582 = (inp[3]) ? 4'b1110 : node25583;
															assign node25583 = (inp[0]) ? node25587 : node25584;
																assign node25584 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node25587 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node25591 = (inp[3]) ? 4'b1100 : node25592;
															assign node25592 = (inp[15]) ? 4'b1100 : node25593;
																assign node25593 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node25598 = (inp[0]) ? node25600 : 4'b1110;
														assign node25600 = (inp[5]) ? node25602 : 4'b1100;
															assign node25602 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node25605 = (inp[10]) ? node25645 : node25606;
											assign node25606 = (inp[3]) ? node25620 : node25607;
												assign node25607 = (inp[15]) ? node25615 : node25608;
													assign node25608 = (inp[5]) ? node25612 : node25609;
														assign node25609 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node25612 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node25615 = (inp[0]) ? 4'b1110 : node25616;
														assign node25616 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node25620 = (inp[12]) ? node25634 : node25621;
													assign node25621 = (inp[5]) ? node25627 : node25622;
														assign node25622 = (inp[15]) ? node25624 : 4'b1100;
															assign node25624 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node25627 = (inp[15]) ? node25631 : node25628;
															assign node25628 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node25631 = (inp[2]) ? 4'b1110 : 4'b1100;
													assign node25634 = (inp[2]) ? node25636 : 4'b1100;
														assign node25636 = (inp[5]) ? 4'b1100 : node25637;
															assign node25637 = (inp[0]) ? node25641 : node25638;
																assign node25638 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node25641 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node25645 = (inp[12]) ? node25663 : node25646;
												assign node25646 = (inp[3]) ? node25658 : node25647;
													assign node25647 = (inp[15]) ? node25653 : node25648;
														assign node25648 = (inp[5]) ? node25650 : 4'b1110;
															assign node25650 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node25653 = (inp[5]) ? node25655 : 4'b1100;
															assign node25655 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node25658 = (inp[2]) ? node25660 : 4'b1100;
														assign node25660 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node25663 = (inp[2]) ? node25671 : node25664;
													assign node25664 = (inp[15]) ? node25668 : node25665;
														assign node25665 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node25668 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node25671 = (inp[0]) ? node25673 : 4'b1010;
														assign node25673 = (inp[15]) ? node25677 : node25674;
															assign node25674 = (inp[3]) ? 4'b1010 : 4'b1000;
															assign node25677 = (inp[3]) ? 4'b1000 : 4'b1010;
								assign node25680 = (inp[12]) ? node25846 : node25681;
									assign node25681 = (inp[10]) ? node25775 : node25682;
										assign node25682 = (inp[9]) ? node25722 : node25683;
											assign node25683 = (inp[4]) ? node25705 : node25684;
												assign node25684 = (inp[15]) ? node25696 : node25685;
													assign node25685 = (inp[2]) ? node25687 : 4'b0110;
														assign node25687 = (inp[0]) ? node25691 : node25688;
															assign node25688 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node25691 = (inp[3]) ? node25693 : 4'b0100;
																assign node25693 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node25696 = (inp[0]) ? node25702 : node25697;
														assign node25697 = (inp[5]) ? node25699 : 4'b0100;
															assign node25699 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node25702 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node25705 = (inp[3]) ? node25709 : node25706;
													assign node25706 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node25709 = (inp[0]) ? node25717 : node25710;
														assign node25710 = (inp[5]) ? node25714 : node25711;
															assign node25711 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node25714 = (inp[2]) ? 4'b0000 : 4'b0010;
														assign node25717 = (inp[2]) ? 4'b0010 : node25718;
															assign node25718 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node25722 = (inp[4]) ? node25758 : node25723;
												assign node25723 = (inp[2]) ? node25741 : node25724;
													assign node25724 = (inp[3]) ? node25734 : node25725;
														assign node25725 = (inp[5]) ? 4'b0010 : node25726;
															assign node25726 = (inp[0]) ? node25730 : node25727;
																assign node25727 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node25730 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node25734 = (inp[5]) ? 4'b0000 : node25735;
															assign node25735 = (inp[0]) ? 4'b0000 : node25736;
																assign node25736 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node25741 = (inp[15]) ? node25753 : node25742;
														assign node25742 = (inp[0]) ? node25748 : node25743;
															assign node25743 = (inp[3]) ? node25745 : 4'b0010;
																assign node25745 = (inp[5]) ? 4'b0000 : 4'b0010;
															assign node25748 = (inp[3]) ? node25750 : 4'b0000;
																assign node25750 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node25753 = (inp[3]) ? 4'b0010 : node25754;
															assign node25754 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node25758 = (inp[5]) ? node25768 : node25759;
													assign node25759 = (inp[15]) ? node25761 : 4'b0110;
														assign node25761 = (inp[0]) ? node25765 : node25762;
															assign node25762 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node25765 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node25768 = (inp[0]) ? node25772 : node25769;
														assign node25769 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node25772 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node25775 = (inp[9]) ? node25809 : node25776;
											assign node25776 = (inp[4]) ? node25794 : node25777;
												assign node25777 = (inp[2]) ? node25785 : node25778;
													assign node25778 = (inp[15]) ? 4'b0110 : node25779;
														assign node25779 = (inp[0]) ? node25781 : 4'b0110;
															assign node25781 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node25785 = (inp[0]) ? node25789 : node25786;
														assign node25786 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node25789 = (inp[15]) ? 4'b0110 : node25790;
															assign node25790 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node25794 = (inp[15]) ? node25800 : node25795;
													assign node25795 = (inp[0]) ? node25797 : 4'b0010;
														assign node25797 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node25800 = (inp[0]) ? node25806 : node25801;
														assign node25801 = (inp[5]) ? node25803 : 4'b0000;
															assign node25803 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node25806 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node25809 = (inp[4]) ? node25823 : node25810;
												assign node25810 = (inp[15]) ? node25816 : node25811;
													assign node25811 = (inp[0]) ? 4'b0000 : node25812;
														assign node25812 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node25816 = (inp[0]) ? node25820 : node25817;
														assign node25817 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node25820 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node25823 = (inp[15]) ? node25835 : node25824;
													assign node25824 = (inp[0]) ? node25830 : node25825;
														assign node25825 = (inp[5]) ? 4'b0100 : node25826;
															assign node25826 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node25830 = (inp[5]) ? 4'b0110 : node25831;
															assign node25831 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node25835 = (inp[0]) ? node25841 : node25836;
														assign node25836 = (inp[3]) ? 4'b0110 : node25837;
															assign node25837 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node25841 = (inp[3]) ? 4'b0100 : node25842;
															assign node25842 = (inp[5]) ? 4'b0100 : 4'b0110;
									assign node25846 = (inp[3]) ? node25950 : node25847;
										assign node25847 = (inp[15]) ? node25893 : node25848;
											assign node25848 = (inp[0]) ? node25866 : node25849;
												assign node25849 = (inp[5]) ? node25859 : node25850;
													assign node25850 = (inp[2]) ? node25852 : 4'b0110;
														assign node25852 = (inp[4]) ? 4'b0010 : node25853;
															assign node25853 = (inp[10]) ? 4'b0110 : node25854;
																assign node25854 = (inp[9]) ? 4'b0010 : 4'b0110;
													assign node25859 = (inp[9]) ? 4'b0100 : node25860;
														assign node25860 = (inp[10]) ? 4'b0100 : node25861;
															assign node25861 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node25866 = (inp[5]) ? node25878 : node25867;
													assign node25867 = (inp[9]) ? node25873 : node25868;
														assign node25868 = (inp[4]) ? 4'b0000 : node25869;
															assign node25869 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node25873 = (inp[10]) ? node25875 : 4'b0100;
															assign node25875 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node25878 = (inp[10]) ? node25886 : node25879;
														assign node25879 = (inp[4]) ? node25883 : node25880;
															assign node25880 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node25883 = (inp[9]) ? 4'b0110 : 4'b0000;
														assign node25886 = (inp[4]) ? node25890 : node25887;
															assign node25887 = (inp[9]) ? 4'b0110 : 4'b0000;
															assign node25890 = (inp[9]) ? 4'b0010 : 4'b0110;
											assign node25893 = (inp[0]) ? node25923 : node25894;
												assign node25894 = (inp[5]) ? node25908 : node25895;
													assign node25895 = (inp[2]) ? node25901 : node25896;
														assign node25896 = (inp[9]) ? node25898 : 4'b0000;
															assign node25898 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node25901 = (inp[4]) ? 4'b0000 : node25902;
															assign node25902 = (inp[10]) ? 4'b0100 : node25903;
																assign node25903 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node25908 = (inp[9]) ? node25916 : node25909;
														assign node25909 = (inp[2]) ? 4'b0000 : node25910;
															assign node25910 = (inp[10]) ? 4'b0110 : node25911;
																assign node25911 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node25916 = (inp[4]) ? node25920 : node25917;
															assign node25917 = (inp[10]) ? 4'b0110 : 4'b0000;
															assign node25920 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node25923 = (inp[5]) ? node25943 : node25924;
													assign node25924 = (inp[10]) ? node25932 : node25925;
														assign node25925 = (inp[4]) ? node25929 : node25926;
															assign node25926 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node25929 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node25932 = (inp[2]) ? node25938 : node25933;
															assign node25933 = (inp[9]) ? 4'b0010 : node25934;
																assign node25934 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node25938 = (inp[9]) ? node25940 : 4'b0010;
																assign node25940 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node25943 = (inp[10]) ? node25945 : 4'b0010;
														assign node25945 = (inp[4]) ? node25947 : 4'b0010;
															assign node25947 = (inp[9]) ? 4'b0000 : 4'b0100;
										assign node25950 = (inp[0]) ? node26000 : node25951;
											assign node25951 = (inp[15]) ? node25979 : node25952;
												assign node25952 = (inp[5]) ? node25964 : node25953;
													assign node25953 = (inp[2]) ? node25959 : node25954;
														assign node25954 = (inp[10]) ? node25956 : 4'b0010;
															assign node25956 = (inp[4]) ? 4'b0000 : 4'b0010;
														assign node25959 = (inp[4]) ? 4'b0000 : node25960;
															assign node25960 = (inp[9]) ? 4'b0100 : 4'b0110;
													assign node25964 = (inp[9]) ? node25972 : node25965;
														assign node25965 = (inp[10]) ? node25969 : node25966;
															assign node25966 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node25969 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node25972 = (inp[4]) ? node25976 : node25973;
															assign node25973 = (inp[10]) ? 4'b0100 : 4'b0000;
															assign node25976 = (inp[10]) ? 4'b0000 : 4'b0100;
												assign node25979 = (inp[5]) ? node25991 : node25980;
													assign node25980 = (inp[10]) ? node25986 : node25981;
														assign node25981 = (inp[4]) ? 4'b0000 : node25982;
															assign node25982 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node25986 = (inp[4]) ? node25988 : 4'b0000;
															assign node25988 = (inp[2]) ? 4'b0110 : 4'b0010;
													assign node25991 = (inp[4]) ? 4'b0010 : node25992;
														assign node25992 = (inp[10]) ? node25996 : node25993;
															assign node25993 = (inp[9]) ? 4'b0010 : 4'b0110;
															assign node25996 = (inp[9]) ? 4'b0110 : 4'b0010;
											assign node26000 = (inp[15]) ? node26022 : node26001;
												assign node26001 = (inp[5]) ? node26011 : node26002;
													assign node26002 = (inp[9]) ? node26004 : 4'b0000;
														assign node26004 = (inp[10]) ? node26008 : node26005;
															assign node26005 = (inp[4]) ? 4'b0110 : 4'b0000;
															assign node26008 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node26011 = (inp[2]) ? node26017 : node26012;
														assign node26012 = (inp[4]) ? 4'b0110 : node26013;
															assign node26013 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node26017 = (inp[10]) ? node26019 : 4'b0010;
															assign node26019 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node26022 = (inp[5]) ? node26038 : node26023;
													assign node26023 = (inp[10]) ? node26033 : node26024;
														assign node26024 = (inp[2]) ? node26028 : node26025;
															assign node26025 = (inp[9]) ? 4'b0100 : 4'b0110;
															assign node26028 = (inp[9]) ? 4'b0010 : node26029;
																assign node26029 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node26033 = (inp[9]) ? node26035 : 4'b0100;
															assign node26035 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node26038 = (inp[4]) ? node26046 : node26039;
														assign node26039 = (inp[10]) ? node26043 : node26040;
															assign node26040 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node26043 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node26046 = (inp[2]) ? 4'b0100 : node26047;
															assign node26047 = (inp[10]) ? 4'b0000 : 4'b0100;
						assign node26051 = (inp[13]) ? node26621 : node26052;
							assign node26052 = (inp[3]) ? node26348 : node26053;
								assign node26053 = (inp[12]) ? node26177 : node26054;
									assign node26054 = (inp[5]) ? node26104 : node26055;
										assign node26055 = (inp[15]) ? node26075 : node26056;
											assign node26056 = (inp[0]) ? node26068 : node26057;
												assign node26057 = (inp[2]) ? node26063 : node26058;
													assign node26058 = (inp[9]) ? node26060 : 4'b0010;
														assign node26060 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node26063 = (inp[9]) ? node26065 : 4'b0110;
														assign node26065 = (inp[4]) ? 4'b0110 : 4'b0010;
												assign node26068 = (inp[9]) ? node26072 : node26069;
													assign node26069 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node26072 = (inp[4]) ? 4'b0100 : 4'b0000;
											assign node26075 = (inp[0]) ? node26083 : node26076;
												assign node26076 = (inp[9]) ? node26080 : node26077;
													assign node26077 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node26080 = (inp[4]) ? 4'b0100 : 4'b0000;
												assign node26083 = (inp[2]) ? node26091 : node26084;
													assign node26084 = (inp[4]) ? node26088 : node26085;
														assign node26085 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node26088 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node26091 = (inp[10]) ? node26097 : node26092;
														assign node26092 = (inp[1]) ? 4'b0010 : node26093;
															assign node26093 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node26097 = (inp[1]) ? node26099 : 4'b0010;
															assign node26099 = (inp[4]) ? node26101 : 4'b0110;
																assign node26101 = (inp[9]) ? 4'b0110 : 4'b0010;
										assign node26104 = (inp[9]) ? node26144 : node26105;
											assign node26105 = (inp[4]) ? node26119 : node26106;
												assign node26106 = (inp[2]) ? node26114 : node26107;
													assign node26107 = (inp[15]) ? node26111 : node26108;
														assign node26108 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node26111 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node26114 = (inp[0]) ? node26116 : 4'b0110;
														assign node26116 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node26119 = (inp[1]) ? node26139 : node26120;
													assign node26120 = (inp[2]) ? node26130 : node26121;
														assign node26121 = (inp[10]) ? node26123 : 4'b0010;
															assign node26123 = (inp[15]) ? node26127 : node26124;
																assign node26124 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node26127 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node26130 = (inp[10]) ? 4'b0010 : node26131;
															assign node26131 = (inp[0]) ? node26135 : node26132;
																assign node26132 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node26135 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26139 = (inp[15]) ? node26141 : 4'b0000;
														assign node26141 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node26144 = (inp[4]) ? node26170 : node26145;
												assign node26145 = (inp[1]) ? node26161 : node26146;
													assign node26146 = (inp[10]) ? node26152 : node26147;
														assign node26147 = (inp[15]) ? 4'b0000 : node26148;
															assign node26148 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node26152 = (inp[2]) ? 4'b0010 : node26153;
															assign node26153 = (inp[0]) ? node26157 : node26154;
																assign node26154 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node26157 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26161 = (inp[10]) ? node26167 : node26162;
														assign node26162 = (inp[0]) ? node26164 : 4'b0010;
															assign node26164 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node26167 = (inp[2]) ? 4'b0000 : 4'b0010;
												assign node26170 = (inp[15]) ? node26174 : node26171;
													assign node26171 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node26174 = (inp[0]) ? 4'b0100 : 4'b0110;
									assign node26177 = (inp[9]) ? node26239 : node26178;
										assign node26178 = (inp[15]) ? node26206 : node26179;
											assign node26179 = (inp[0]) ? node26189 : node26180;
												assign node26180 = (inp[4]) ? node26184 : node26181;
													assign node26181 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node26184 = (inp[10]) ? node26186 : 4'b0010;
														assign node26186 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node26189 = (inp[5]) ? node26199 : node26190;
													assign node26190 = (inp[1]) ? 4'b0100 : node26191;
														assign node26191 = (inp[4]) ? node26195 : node26192;
															assign node26192 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node26195 = (inp[10]) ? 4'b0100 : 4'b0000;
													assign node26199 = (inp[4]) ? node26203 : node26200;
														assign node26200 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node26203 = (inp[10]) ? 4'b0110 : 4'b0000;
											assign node26206 = (inp[0]) ? node26228 : node26207;
												assign node26207 = (inp[5]) ? node26221 : node26208;
													assign node26208 = (inp[2]) ? node26216 : node26209;
														assign node26209 = (inp[1]) ? node26211 : 4'b0000;
															assign node26211 = (inp[10]) ? 4'b0000 : node26212;
																assign node26212 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node26216 = (inp[10]) ? node26218 : 4'b0000;
															assign node26218 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node26221 = (inp[4]) ? node26225 : node26222;
														assign node26222 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node26225 = (inp[10]) ? 4'b0110 : 4'b0000;
												assign node26228 = (inp[5]) ? node26234 : node26229;
													assign node26229 = (inp[2]) ? 4'b0110 : node26230;
														assign node26230 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node26234 = (inp[4]) ? node26236 : 4'b0010;
														assign node26236 = (inp[10]) ? 4'b0100 : 4'b0010;
										assign node26239 = (inp[2]) ? node26299 : node26240;
											assign node26240 = (inp[1]) ? node26270 : node26241;
												assign node26241 = (inp[10]) ? node26253 : node26242;
													assign node26242 = (inp[4]) ? node26248 : node26243;
														assign node26243 = (inp[5]) ? 4'b0000 : node26244;
															assign node26244 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node26248 = (inp[15]) ? node26250 : 4'b0100;
															assign node26250 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node26253 = (inp[4]) ? node26267 : node26254;
														assign node26254 = (inp[15]) ? node26260 : node26255;
															assign node26255 = (inp[0]) ? 4'b0100 : node26256;
																assign node26256 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node26260 = (inp[0]) ? node26264 : node26261;
																assign node26261 = (inp[5]) ? 4'b0110 : 4'b0100;
																assign node26264 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node26267 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node26270 = (inp[5]) ? node26282 : node26271;
													assign node26271 = (inp[0]) ? node26275 : node26272;
														assign node26272 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node26275 = (inp[15]) ? node26279 : node26276;
															assign node26276 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node26279 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node26282 = (inp[4]) ? node26290 : node26283;
														assign node26283 = (inp[10]) ? 4'b0110 : node26284;
															assign node26284 = (inp[15]) ? node26286 : 4'b0010;
																assign node26286 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node26290 = (inp[10]) ? node26296 : node26291;
															assign node26291 = (inp[15]) ? node26293 : 4'b0110;
																assign node26293 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node26296 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node26299 = (inp[10]) ? node26321 : node26300;
												assign node26300 = (inp[4]) ? node26314 : node26301;
													assign node26301 = (inp[1]) ? node26309 : node26302;
														assign node26302 = (inp[0]) ? node26306 : node26303;
															assign node26303 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node26306 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node26309 = (inp[5]) ? node26311 : 4'b0010;
															assign node26311 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node26314 = (inp[15]) ? node26316 : 4'b0110;
														assign node26316 = (inp[5]) ? node26318 : 4'b0100;
															assign node26318 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node26321 = (inp[4]) ? node26333 : node26322;
													assign node26322 = (inp[15]) ? 4'b0110 : node26323;
														assign node26323 = (inp[1]) ? node26327 : node26324;
															assign node26324 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node26327 = (inp[5]) ? 4'b0110 : node26328;
																assign node26328 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node26333 = (inp[0]) ? node26341 : node26334;
														assign node26334 = (inp[1]) ? node26336 : 4'b0010;
															assign node26336 = (inp[15]) ? 4'b0010 : node26337;
																assign node26337 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node26341 = (inp[15]) ? node26345 : node26342;
															assign node26342 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node26345 = (inp[5]) ? 4'b0000 : 4'b0010;
								assign node26348 = (inp[9]) ? node26530 : node26349;
									assign node26349 = (inp[4]) ? node26441 : node26350;
										assign node26350 = (inp[12]) ? node26410 : node26351;
											assign node26351 = (inp[10]) ? node26377 : node26352;
												assign node26352 = (inp[0]) ? node26372 : node26353;
													assign node26353 = (inp[2]) ? node26359 : node26354;
														assign node26354 = (inp[15]) ? node26356 : 4'b0110;
															assign node26356 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node26359 = (inp[1]) ? node26365 : node26360;
															assign node26360 = (inp[15]) ? 4'b0110 : node26361;
																assign node26361 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node26365 = (inp[15]) ? node26369 : node26366;
																assign node26366 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node26369 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node26372 = (inp[2]) ? 4'b0110 : node26373;
														assign node26373 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node26377 = (inp[2]) ? node26397 : node26378;
													assign node26378 = (inp[0]) ? node26388 : node26379;
														assign node26379 = (inp[1]) ? 4'b0110 : node26380;
															assign node26380 = (inp[5]) ? node26384 : node26381;
																assign node26381 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node26384 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node26388 = (inp[1]) ? node26390 : 4'b0110;
															assign node26390 = (inp[15]) ? node26394 : node26391;
																assign node26391 = (inp[5]) ? 4'b0110 : 4'b0100;
																assign node26394 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node26397 = (inp[5]) ? node26403 : node26398;
														assign node26398 = (inp[1]) ? node26400 : 4'b0100;
															assign node26400 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node26403 = (inp[0]) ? node26407 : node26404;
															assign node26404 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node26407 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node26410 = (inp[10]) ? node26428 : node26411;
												assign node26411 = (inp[15]) ? node26423 : node26412;
													assign node26412 = (inp[1]) ? 4'b0110 : node26413;
														assign node26413 = (inp[2]) ? node26419 : node26414;
															assign node26414 = (inp[0]) ? 4'b0110 : node26415;
																assign node26415 = (inp[5]) ? 4'b0100 : 4'b0110;
															assign node26419 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node26423 = (inp[0]) ? node26425 : 4'b0100;
														assign node26425 = (inp[2]) ? 4'b0100 : 4'b0110;
												assign node26428 = (inp[15]) ? node26436 : node26429;
													assign node26429 = (inp[0]) ? node26433 : node26430;
														assign node26430 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node26433 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node26436 = (inp[0]) ? node26438 : 4'b0010;
														assign node26438 = (inp[5]) ? 4'b0000 : 4'b0010;
										assign node26441 = (inp[10]) ? node26477 : node26442;
											assign node26442 = (inp[0]) ? node26460 : node26443;
												assign node26443 = (inp[1]) ? node26451 : node26444;
													assign node26444 = (inp[5]) ? node26448 : node26445;
														assign node26445 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node26448 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26451 = (inp[12]) ? node26453 : 4'b0010;
														assign node26453 = (inp[5]) ? node26457 : node26454;
															assign node26454 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node26457 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node26460 = (inp[12]) ? node26472 : node26461;
													assign node26461 = (inp[2]) ? node26467 : node26462;
														assign node26462 = (inp[1]) ? 4'b0000 : node26463;
															assign node26463 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node26467 = (inp[1]) ? 4'b0010 : node26468;
															assign node26468 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node26472 = (inp[5]) ? 4'b0010 : node26473;
														assign node26473 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node26477 = (inp[12]) ? node26495 : node26478;
												assign node26478 = (inp[1]) ? node26488 : node26479;
													assign node26479 = (inp[15]) ? node26481 : 4'b0000;
														assign node26481 = (inp[0]) ? node26485 : node26482;
															assign node26482 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node26485 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node26488 = (inp[5]) ? node26490 : 4'b0010;
														assign node26490 = (inp[0]) ? node26492 : 4'b0010;
															assign node26492 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node26495 = (inp[2]) ? node26509 : node26496;
													assign node26496 = (inp[5]) ? node26504 : node26497;
														assign node26497 = (inp[0]) ? node26501 : node26498;
															assign node26498 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node26501 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node26504 = (inp[15]) ? 4'b0110 : node26505;
															assign node26505 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node26509 = (inp[1]) ? node26521 : node26510;
														assign node26510 = (inp[5]) ? node26516 : node26511;
															assign node26511 = (inp[15]) ? 4'b0110 : node26512;
																assign node26512 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node26516 = (inp[0]) ? 4'b0100 : node26517;
																assign node26517 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node26521 = (inp[5]) ? node26523 : 4'b0100;
															assign node26523 = (inp[15]) ? node26527 : node26524;
																assign node26524 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node26527 = (inp[0]) ? 4'b0100 : 4'b0110;
									assign node26530 = (inp[4]) ? node26590 : node26531;
										assign node26531 = (inp[10]) ? node26573 : node26532;
											assign node26532 = (inp[1]) ? node26554 : node26533;
												assign node26533 = (inp[2]) ? node26545 : node26534;
													assign node26534 = (inp[5]) ? node26540 : node26535;
														assign node26535 = (inp[15]) ? 4'b0000 : node26536;
															assign node26536 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node26540 = (inp[0]) ? 4'b0010 : node26541;
															assign node26541 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26545 = (inp[12]) ? 4'b0010 : node26546;
														assign node26546 = (inp[5]) ? 4'b0000 : node26547;
															assign node26547 = (inp[15]) ? 4'b0010 : node26548;
																assign node26548 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node26554 = (inp[5]) ? node26560 : node26555;
													assign node26555 = (inp[0]) ? 4'b0000 : node26556;
														assign node26556 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node26560 = (inp[2]) ? node26568 : node26561;
														assign node26561 = (inp[0]) ? node26565 : node26562;
															assign node26562 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node26565 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node26568 = (inp[15]) ? node26570 : 4'b0000;
															assign node26570 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node26573 = (inp[12]) ? node26585 : node26574;
												assign node26574 = (inp[5]) ? node26580 : node26575;
													assign node26575 = (inp[0]) ? node26577 : 4'b0010;
														assign node26577 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26580 = (inp[0]) ? node26582 : 4'b0000;
														assign node26582 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node26585 = (inp[0]) ? node26587 : 4'b0110;
													assign node26587 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node26590 = (inp[12]) ? node26598 : node26591;
											assign node26591 = (inp[0]) ? node26595 : node26592;
												assign node26592 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node26595 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node26598 = (inp[10]) ? node26608 : node26599;
												assign node26599 = (inp[1]) ? 4'b0100 : node26600;
													assign node26600 = (inp[15]) ? node26604 : node26601;
														assign node26601 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node26604 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node26608 = (inp[1]) ? node26610 : 4'b0000;
													assign node26610 = (inp[5]) ? node26618 : node26611;
														assign node26611 = (inp[15]) ? node26615 : node26612;
															assign node26612 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node26615 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node26618 = (inp[15]) ? 4'b0000 : 4'b0010;
							assign node26621 = (inp[1]) ? node26947 : node26622;
								assign node26622 = (inp[9]) ? node26808 : node26623;
									assign node26623 = (inp[4]) ? node26731 : node26624;
										assign node26624 = (inp[12]) ? node26680 : node26625;
											assign node26625 = (inp[10]) ? node26657 : node26626;
												assign node26626 = (inp[2]) ? node26648 : node26627;
													assign node26627 = (inp[0]) ? node26637 : node26628;
														assign node26628 = (inp[5]) ? node26630 : 4'b0100;
															assign node26630 = (inp[3]) ? node26634 : node26631;
																assign node26631 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node26634 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node26637 = (inp[15]) ? node26643 : node26638;
															assign node26638 = (inp[3]) ? node26640 : 4'b0100;
																assign node26640 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node26643 = (inp[3]) ? node26645 : 4'b0110;
																assign node26645 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node26648 = (inp[15]) ? 4'b0110 : node26649;
														assign node26649 = (inp[0]) ? 4'b0100 : node26650;
															assign node26650 = (inp[3]) ? node26652 : 4'b0110;
																assign node26652 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node26657 = (inp[3]) ? node26673 : node26658;
													assign node26658 = (inp[5]) ? node26668 : node26659;
														assign node26659 = (inp[2]) ? node26665 : node26660;
															assign node26660 = (inp[0]) ? node26662 : 4'b0110;
																assign node26662 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node26665 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node26668 = (inp[15]) ? node26670 : 4'b0100;
															assign node26670 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node26673 = (inp[15]) ? node26675 : 4'b0100;
														assign node26675 = (inp[0]) ? 4'b0100 : node26676;
															assign node26676 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node26680 = (inp[10]) ? node26704 : node26681;
												assign node26681 = (inp[5]) ? node26691 : node26682;
													assign node26682 = (inp[2]) ? node26684 : 4'b0100;
														assign node26684 = (inp[3]) ? node26686 : 4'b0110;
															assign node26686 = (inp[15]) ? 4'b0100 : node26687;
																assign node26687 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node26691 = (inp[15]) ? node26699 : node26692;
														assign node26692 = (inp[2]) ? node26696 : node26693;
															assign node26693 = (inp[3]) ? 4'b0110 : 4'b0100;
															assign node26696 = (inp[3]) ? 4'b0100 : 4'b0110;
														assign node26699 = (inp[0]) ? node26701 : 4'b0110;
															assign node26701 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node26704 = (inp[3]) ? node26714 : node26705;
													assign node26705 = (inp[5]) ? 4'b0010 : node26706;
														assign node26706 = (inp[0]) ? node26710 : node26707;
															assign node26707 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node26710 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26714 = (inp[2]) ? node26724 : node26715;
														assign node26715 = (inp[15]) ? node26717 : 4'b0010;
															assign node26717 = (inp[5]) ? node26721 : node26718;
																assign node26718 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node26721 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node26724 = (inp[15]) ? 4'b0000 : node26725;
															assign node26725 = (inp[5]) ? 4'b0000 : node26726;
																assign node26726 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node26731 = (inp[10]) ? node26771 : node26732;
											assign node26732 = (inp[2]) ? node26754 : node26733;
												assign node26733 = (inp[12]) ? node26745 : node26734;
													assign node26734 = (inp[0]) ? node26738 : node26735;
														assign node26735 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node26738 = (inp[15]) ? 4'b0010 : node26739;
															assign node26739 = (inp[5]) ? node26741 : 4'b0000;
																assign node26741 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node26745 = (inp[0]) ? node26751 : node26746;
														assign node26746 = (inp[15]) ? node26748 : 4'b0010;
															assign node26748 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node26751 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node26754 = (inp[0]) ? node26762 : node26755;
													assign node26755 = (inp[3]) ? node26757 : 4'b0000;
														assign node26757 = (inp[5]) ? node26759 : 4'b0000;
															assign node26759 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node26762 = (inp[5]) ? node26766 : node26763;
														assign node26763 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node26766 = (inp[15]) ? 4'b0000 : node26767;
															assign node26767 = (inp[3]) ? 4'b0010 : 4'b0000;
											assign node26771 = (inp[12]) ? node26787 : node26772;
												assign node26772 = (inp[15]) ? node26780 : node26773;
													assign node26773 = (inp[3]) ? node26775 : 4'b0000;
														assign node26775 = (inp[5]) ? node26777 : 4'b0000;
															assign node26777 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node26780 = (inp[0]) ? 4'b0010 : node26781;
														assign node26781 = (inp[3]) ? node26783 : 4'b0000;
															assign node26783 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node26787 = (inp[5]) ? node26797 : node26788;
													assign node26788 = (inp[0]) ? 4'b0100 : node26789;
														assign node26789 = (inp[15]) ? node26793 : node26790;
															assign node26790 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node26793 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node26797 = (inp[3]) ? 4'b0110 : node26798;
														assign node26798 = (inp[2]) ? node26800 : 4'b0100;
															assign node26800 = (inp[0]) ? node26804 : node26801;
																assign node26801 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node26804 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node26808 = (inp[4]) ? node26866 : node26809;
										assign node26809 = (inp[10]) ? node26833 : node26810;
											assign node26810 = (inp[0]) ? node26822 : node26811;
												assign node26811 = (inp[15]) ? node26817 : node26812;
													assign node26812 = (inp[5]) ? node26814 : 4'b0010;
														assign node26814 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node26817 = (inp[5]) ? node26819 : 4'b0000;
														assign node26819 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node26822 = (inp[15]) ? node26828 : node26823;
													assign node26823 = (inp[5]) ? node26825 : 4'b0000;
														assign node26825 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node26828 = (inp[3]) ? node26830 : 4'b0010;
														assign node26830 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node26833 = (inp[12]) ? node26851 : node26834;
												assign node26834 = (inp[15]) ? node26840 : node26835;
													assign node26835 = (inp[2]) ? node26837 : 4'b0010;
														assign node26837 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node26840 = (inp[0]) ? node26846 : node26841;
														assign node26841 = (inp[3]) ? node26843 : 4'b0000;
															assign node26843 = (inp[2]) ? 4'b0010 : 4'b0000;
														assign node26846 = (inp[3]) ? node26848 : 4'b0010;
															assign node26848 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node26851 = (inp[5]) ? node26859 : node26852;
													assign node26852 = (inp[3]) ? 4'b0110 : node26853;
														assign node26853 = (inp[15]) ? 4'b0100 : node26854;
															assign node26854 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node26859 = (inp[3]) ? 4'b0100 : node26860;
														assign node26860 = (inp[15]) ? 4'b0110 : node26861;
															assign node26861 = (inp[0]) ? 4'b0110 : 4'b0100;
										assign node26866 = (inp[10]) ? node26900 : node26867;
											assign node26867 = (inp[3]) ? node26887 : node26868;
												assign node26868 = (inp[5]) ? node26880 : node26869;
													assign node26869 = (inp[12]) ? node26871 : 4'b0110;
														assign node26871 = (inp[2]) ? 4'b0110 : node26872;
															assign node26872 = (inp[15]) ? node26876 : node26873;
																assign node26873 = (inp[0]) ? 4'b0100 : 4'b0110;
																assign node26876 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node26880 = (inp[15]) ? node26884 : node26881;
														assign node26881 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node26884 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node26887 = (inp[5]) ? node26895 : node26888;
													assign node26888 = (inp[15]) ? node26892 : node26889;
														assign node26889 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node26892 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node26895 = (inp[0]) ? node26897 : 4'b0110;
														assign node26897 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node26900 = (inp[12]) ? node26922 : node26901;
												assign node26901 = (inp[3]) ? node26907 : node26902;
													assign node26902 = (inp[2]) ? 4'b0110 : node26903;
														assign node26903 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node26907 = (inp[2]) ? node26913 : node26908;
														assign node26908 = (inp[0]) ? node26910 : 4'b0110;
															assign node26910 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node26913 = (inp[5]) ? node26915 : 4'b0100;
															assign node26915 = (inp[0]) ? node26919 : node26916;
																assign node26916 = (inp[15]) ? 4'b0110 : 4'b0100;
																assign node26919 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node26922 = (inp[2]) ? node26936 : node26923;
													assign node26923 = (inp[3]) ? node26931 : node26924;
														assign node26924 = (inp[5]) ? 4'b0000 : node26925;
															assign node26925 = (inp[0]) ? node26927 : 4'b0000;
																assign node26927 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node26931 = (inp[0]) ? 4'b0010 : node26932;
															assign node26932 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node26936 = (inp[3]) ? 4'b0000 : node26937;
														assign node26937 = (inp[15]) ? 4'b0000 : node26938;
															assign node26938 = (inp[0]) ? node26942 : node26939;
																assign node26939 = (inp[5]) ? 4'b0000 : 4'b0010;
																assign node26942 = (inp[5]) ? 4'b0010 : 4'b0000;
								assign node26947 = (inp[15]) ? node27085 : node26948;
									assign node26948 = (inp[0]) ? node27002 : node26949;
										assign node26949 = (inp[3]) ? node26983 : node26950;
											assign node26950 = (inp[5]) ? node26968 : node26951;
												assign node26951 = (inp[4]) ? node26959 : node26952;
													assign node26952 = (inp[12]) ? 4'b1110 : node26953;
														assign node26953 = (inp[2]) ? 4'b1010 : node26954;
															assign node26954 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node26959 = (inp[2]) ? node26965 : node26960;
														assign node26960 = (inp[10]) ? 4'b1010 : node26961;
															assign node26961 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node26965 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node26968 = (inp[9]) ? node26978 : node26969;
													assign node26969 = (inp[10]) ? node26975 : node26970;
														assign node26970 = (inp[4]) ? 4'b1010 : node26971;
															assign node26971 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node26975 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node26978 = (inp[4]) ? node26980 : 4'b1100;
														assign node26980 = (inp[10]) ? 4'b1000 : 4'b1100;
											assign node26983 = (inp[4]) ? node26991 : node26984;
												assign node26984 = (inp[9]) ? node26988 : node26985;
													assign node26985 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node26988 = (inp[10]) ? 4'b1100 : 4'b1000;
												assign node26991 = (inp[9]) ? node26997 : node26992;
													assign node26992 = (inp[12]) ? 4'b1100 : node26993;
														assign node26993 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node26997 = (inp[12]) ? 4'b1000 : node26998;
														assign node26998 = (inp[10]) ? 4'b1000 : 4'b1100;
										assign node27002 = (inp[3]) ? node27034 : node27003;
											assign node27003 = (inp[5]) ? node27017 : node27004;
												assign node27004 = (inp[12]) ? node27012 : node27005;
													assign node27005 = (inp[4]) ? 4'b1100 : node27006;
														assign node27006 = (inp[10]) ? node27008 : 4'b1000;
															assign node27008 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node27012 = (inp[9]) ? 4'b1000 : node27013;
														assign node27013 = (inp[4]) ? 4'b1100 : 4'b1000;
												assign node27017 = (inp[4]) ? node27027 : node27018;
													assign node27018 = (inp[9]) ? node27024 : node27019;
														assign node27019 = (inp[10]) ? 4'b1000 : node27020;
															assign node27020 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node27024 = (inp[12]) ? 4'b1110 : 4'b1000;
													assign node27027 = (inp[9]) ? 4'b1010 : node27028;
														assign node27028 = (inp[12]) ? 4'b1110 : node27029;
															assign node27029 = (inp[10]) ? 4'b1110 : 4'b1000;
											assign node27034 = (inp[2]) ? node27056 : node27035;
												assign node27035 = (inp[12]) ? node27043 : node27036;
													assign node27036 = (inp[10]) ? 4'b1110 : node27037;
														assign node27037 = (inp[9]) ? 4'b1110 : node27038;
															assign node27038 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node27043 = (inp[10]) ? node27049 : node27044;
														assign node27044 = (inp[9]) ? node27046 : 4'b1000;
															assign node27046 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node27049 = (inp[4]) ? node27053 : node27050;
															assign node27050 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node27053 = (inp[9]) ? 4'b1010 : 4'b1110;
												assign node27056 = (inp[5]) ? node27066 : node27057;
													assign node27057 = (inp[4]) ? node27059 : 4'b1000;
														assign node27059 = (inp[9]) ? 4'b1010 : node27060;
															assign node27060 = (inp[12]) ? 4'b1110 : node27061;
																assign node27061 = (inp[10]) ? 4'b1110 : 4'b1000;
													assign node27066 = (inp[4]) ? node27076 : node27067;
														assign node27067 = (inp[9]) ? node27071 : node27068;
															assign node27068 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node27071 = (inp[12]) ? 4'b1110 : node27072;
																assign node27072 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node27076 = (inp[9]) ? node27080 : node27077;
															assign node27077 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node27080 = (inp[10]) ? 4'b1010 : node27081;
																assign node27081 = (inp[12]) ? 4'b1010 : 4'b1110;
									assign node27085 = (inp[4]) ? node27143 : node27086;
										assign node27086 = (inp[9]) ? node27116 : node27087;
											assign node27087 = (inp[10]) ? node27105 : node27088;
												assign node27088 = (inp[12]) ? node27100 : node27089;
													assign node27089 = (inp[0]) ? node27095 : node27090;
														assign node27090 = (inp[3]) ? node27092 : 4'b1100;
															assign node27092 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node27095 = (inp[3]) ? node27097 : 4'b1110;
															assign node27097 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node27100 = (inp[5]) ? 4'b1000 : node27101;
														assign node27101 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node27105 = (inp[0]) ? node27111 : node27106;
													assign node27106 = (inp[3]) ? node27108 : 4'b1000;
														assign node27108 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node27111 = (inp[5]) ? node27113 : 4'b1010;
														assign node27113 = (inp[3]) ? 4'b1000 : 4'b1010;
											assign node27116 = (inp[0]) ? node27130 : node27117;
												assign node27117 = (inp[3]) ? node27125 : node27118;
													assign node27118 = (inp[5]) ? node27120 : 4'b1100;
														assign node27120 = (inp[12]) ? 4'b1110 : node27121;
															assign node27121 = (inp[10]) ? 4'b1110 : 4'b1000;
													assign node27125 = (inp[12]) ? 4'b1110 : node27126;
														assign node27126 = (inp[10]) ? 4'b1110 : 4'b1000;
												assign node27130 = (inp[5]) ? node27138 : node27131;
													assign node27131 = (inp[3]) ? node27133 : 4'b1110;
														assign node27133 = (inp[10]) ? 4'b1100 : node27134;
															assign node27134 = (inp[12]) ? 4'b1100 : 4'b1010;
													assign node27138 = (inp[12]) ? 4'b1100 : node27139;
														assign node27139 = (inp[10]) ? 4'b1100 : 4'b1000;
										assign node27143 = (inp[9]) ? node27173 : node27144;
											assign node27144 = (inp[12]) ? node27162 : node27145;
												assign node27145 = (inp[10]) ? node27155 : node27146;
													assign node27146 = (inp[2]) ? node27148 : 4'b1000;
														assign node27148 = (inp[3]) ? node27150 : 4'b1000;
															assign node27150 = (inp[5]) ? node27152 : 4'b1010;
																assign node27152 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node27155 = (inp[0]) ? 4'b1100 : node27156;
														assign node27156 = (inp[3]) ? 4'b1110 : node27157;
															assign node27157 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node27162 = (inp[0]) ? node27168 : node27163;
													assign node27163 = (inp[5]) ? 4'b1110 : node27164;
														assign node27164 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node27168 = (inp[3]) ? 4'b1100 : node27169;
														assign node27169 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node27173 = (inp[0]) ? node27181 : node27174;
												assign node27174 = (inp[5]) ? 4'b1010 : node27175;
													assign node27175 = (inp[3]) ? node27177 : 4'b1000;
														assign node27177 = (inp[12]) ? 4'b1010 : 4'b1110;
												assign node27181 = (inp[10]) ? node27193 : node27182;
													assign node27182 = (inp[12]) ? node27188 : node27183;
														assign node27183 = (inp[2]) ? 4'b1100 : node27184;
															assign node27184 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node27188 = (inp[5]) ? 4'b1000 : node27189;
															assign node27189 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node27193 = (inp[5]) ? 4'b1000 : node27194;
														assign node27194 = (inp[3]) ? 4'b1000 : 4'b1010;
					assign node27198 = (inp[11]) ? node28138 : node27199;
						assign node27199 = (inp[1]) ? node27581 : node27200;
							assign node27200 = (inp[4]) ? node27392 : node27201;
								assign node27201 = (inp[9]) ? node27287 : node27202;
									assign node27202 = (inp[12]) ? node27226 : node27203;
										assign node27203 = (inp[15]) ? node27215 : node27204;
											assign node27204 = (inp[0]) ? node27210 : node27205;
												assign node27205 = (inp[5]) ? node27207 : 4'b0110;
													assign node27207 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node27210 = (inp[5]) ? node27212 : 4'b0100;
													assign node27212 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node27215 = (inp[0]) ? node27221 : node27216;
												assign node27216 = (inp[3]) ? node27218 : 4'b0100;
													assign node27218 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node27221 = (inp[3]) ? node27223 : 4'b0110;
													assign node27223 = (inp[5]) ? 4'b0100 : 4'b0110;
										assign node27226 = (inp[10]) ? node27248 : node27227;
											assign node27227 = (inp[0]) ? node27239 : node27228;
												assign node27228 = (inp[15]) ? node27234 : node27229;
													assign node27229 = (inp[3]) ? node27231 : 4'b0110;
														assign node27231 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node27234 = (inp[5]) ? node27236 : 4'b0100;
														assign node27236 = (inp[3]) ? 4'b0110 : 4'b0100;
												assign node27239 = (inp[15]) ? node27245 : node27240;
													assign node27240 = (inp[3]) ? node27242 : 4'b0100;
														assign node27242 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node27245 = (inp[3]) ? 4'b0100 : 4'b0110;
											assign node27248 = (inp[2]) ? node27272 : node27249;
												assign node27249 = (inp[5]) ? node27261 : node27250;
													assign node27250 = (inp[13]) ? node27256 : node27251;
														assign node27251 = (inp[0]) ? 4'b0000 : node27252;
															assign node27252 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node27256 = (inp[15]) ? 4'b0010 : node27257;
															assign node27257 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node27261 = (inp[3]) ? 4'b0000 : node27262;
														assign node27262 = (inp[13]) ? 4'b0000 : node27263;
															assign node27263 = (inp[0]) ? node27267 : node27264;
																assign node27264 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node27267 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node27272 = (inp[15]) ? node27278 : node27273;
													assign node27273 = (inp[0]) ? node27275 : 4'b0010;
														assign node27275 = (inp[3]) ? 4'b0010 : 4'b0000;
													assign node27278 = (inp[0]) ? node27282 : node27279;
														assign node27279 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node27282 = (inp[13]) ? 4'b0010 : node27283;
															assign node27283 = (inp[3]) ? 4'b0000 : 4'b0010;
									assign node27287 = (inp[10]) ? node27311 : node27288;
										assign node27288 = (inp[0]) ? node27300 : node27289;
											assign node27289 = (inp[15]) ? node27295 : node27290;
												assign node27290 = (inp[3]) ? node27292 : 4'b0010;
													assign node27292 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node27295 = (inp[3]) ? node27297 : 4'b0000;
													assign node27297 = (inp[5]) ? 4'b0010 : 4'b0000;
											assign node27300 = (inp[15]) ? node27306 : node27301;
												assign node27301 = (inp[5]) ? node27303 : 4'b0000;
													assign node27303 = (inp[3]) ? 4'b0010 : 4'b0000;
												assign node27306 = (inp[5]) ? node27308 : 4'b0010;
													assign node27308 = (inp[3]) ? 4'b0000 : 4'b0010;
										assign node27311 = (inp[12]) ? node27357 : node27312;
											assign node27312 = (inp[13]) ? node27328 : node27313;
												assign node27313 = (inp[15]) ? node27323 : node27314;
													assign node27314 = (inp[3]) ? node27316 : 4'b0000;
														assign node27316 = (inp[2]) ? 4'b0010 : node27317;
															assign node27317 = (inp[5]) ? node27319 : 4'b0000;
																assign node27319 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node27323 = (inp[0]) ? node27325 : 4'b0000;
														assign node27325 = (inp[3]) ? 4'b0000 : 4'b0010;
												assign node27328 = (inp[2]) ? node27342 : node27329;
													assign node27329 = (inp[3]) ? node27331 : 4'b0000;
														assign node27331 = (inp[0]) ? node27337 : node27332;
															assign node27332 = (inp[5]) ? 4'b0010 : node27333;
																assign node27333 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node27337 = (inp[5]) ? 4'b0000 : node27338;
																assign node27338 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node27342 = (inp[15]) ? node27352 : node27343;
														assign node27343 = (inp[5]) ? node27347 : node27344;
															assign node27344 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node27347 = (inp[0]) ? 4'b0010 : node27348;
																assign node27348 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node27352 = (inp[0]) ? 4'b0010 : node27353;
															assign node27353 = (inp[5]) ? 4'b0010 : 4'b0000;
											assign node27357 = (inp[5]) ? node27375 : node27358;
												assign node27358 = (inp[15]) ? node27366 : node27359;
													assign node27359 = (inp[3]) ? node27363 : node27360;
														assign node27360 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node27363 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node27366 = (inp[2]) ? node27368 : 4'b0110;
														assign node27368 = (inp[3]) ? node27372 : node27369;
															assign node27369 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node27372 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node27375 = (inp[13]) ? node27383 : node27376;
													assign node27376 = (inp[3]) ? node27378 : 4'b0110;
														assign node27378 = (inp[0]) ? node27380 : 4'b0100;
															assign node27380 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node27383 = (inp[2]) ? 4'b0100 : node27384;
														assign node27384 = (inp[0]) ? node27388 : node27385;
															assign node27385 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node27388 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node27392 = (inp[9]) ? node27482 : node27393;
									assign node27393 = (inp[12]) ? node27443 : node27394;
										assign node27394 = (inp[2]) ? node27414 : node27395;
											assign node27395 = (inp[0]) ? node27405 : node27396;
												assign node27396 = (inp[15]) ? node27400 : node27397;
													assign node27397 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node27400 = (inp[13]) ? 4'b0000 : node27401;
														assign node27401 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node27405 = (inp[15]) ? node27409 : node27406;
													assign node27406 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node27409 = (inp[3]) ? node27411 : 4'b0010;
														assign node27411 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node27414 = (inp[10]) ? node27428 : node27415;
												assign node27415 = (inp[15]) ? node27423 : node27416;
													assign node27416 = (inp[0]) ? 4'b0000 : node27417;
														assign node27417 = (inp[5]) ? node27419 : 4'b0010;
															assign node27419 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node27423 = (inp[0]) ? node27425 : 4'b0000;
														assign node27425 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node27428 = (inp[0]) ? node27438 : node27429;
													assign node27429 = (inp[15]) ? node27435 : node27430;
														assign node27430 = (inp[5]) ? node27432 : 4'b0010;
															assign node27432 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node27435 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node27438 = (inp[15]) ? 4'b0010 : node27439;
														assign node27439 = (inp[3]) ? 4'b0010 : 4'b0000;
										assign node27443 = (inp[10]) ? node27461 : node27444;
											assign node27444 = (inp[0]) ? node27450 : node27445;
												assign node27445 = (inp[15]) ? node27447 : 4'b0010;
													assign node27447 = (inp[13]) ? 4'b0000 : 4'b0010;
												assign node27450 = (inp[15]) ? node27456 : node27451;
													assign node27451 = (inp[3]) ? node27453 : 4'b0000;
														assign node27453 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node27456 = (inp[3]) ? node27458 : 4'b0010;
														assign node27458 = (inp[5]) ? 4'b0000 : 4'b0010;
											assign node27461 = (inp[15]) ? node27473 : node27462;
												assign node27462 = (inp[0]) ? node27468 : node27463;
													assign node27463 = (inp[5]) ? 4'b0100 : node27464;
														assign node27464 = (inp[3]) ? 4'b0100 : 4'b0110;
													assign node27468 = (inp[3]) ? 4'b0110 : node27469;
														assign node27469 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node27473 = (inp[0]) ? node27479 : node27474;
													assign node27474 = (inp[5]) ? 4'b0110 : node27475;
														assign node27475 = (inp[2]) ? 4'b0100 : 4'b0110;
													assign node27479 = (inp[3]) ? 4'b0100 : 4'b0110;
									assign node27482 = (inp[12]) ? node27506 : node27483;
										assign node27483 = (inp[0]) ? node27495 : node27484;
											assign node27484 = (inp[15]) ? node27490 : node27485;
												assign node27485 = (inp[3]) ? 4'b0100 : node27486;
													assign node27486 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node27490 = (inp[5]) ? 4'b0110 : node27491;
													assign node27491 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node27495 = (inp[15]) ? node27501 : node27496;
												assign node27496 = (inp[3]) ? 4'b0110 : node27497;
													assign node27497 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node27501 = (inp[3]) ? 4'b0100 : node27502;
													assign node27502 = (inp[5]) ? 4'b0100 : 4'b0110;
										assign node27506 = (inp[10]) ? node27542 : node27507;
											assign node27507 = (inp[5]) ? node27523 : node27508;
												assign node27508 = (inp[0]) ? node27518 : node27509;
													assign node27509 = (inp[2]) ? node27511 : 4'b0100;
														assign node27511 = (inp[3]) ? node27515 : node27512;
															assign node27512 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node27515 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node27518 = (inp[15]) ? node27520 : 4'b0100;
														assign node27520 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node27523 = (inp[2]) ? node27531 : node27524;
													assign node27524 = (inp[15]) ? node27528 : node27525;
														assign node27525 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node27528 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node27531 = (inp[3]) ? node27533 : 4'b0100;
														assign node27533 = (inp[13]) ? 4'b0110 : node27534;
															assign node27534 = (inp[15]) ? node27538 : node27535;
																assign node27535 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node27538 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node27542 = (inp[2]) ? node27566 : node27543;
												assign node27543 = (inp[3]) ? node27561 : node27544;
													assign node27544 = (inp[15]) ? node27550 : node27545;
														assign node27545 = (inp[5]) ? node27547 : 4'b0000;
															assign node27547 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node27550 = (inp[13]) ? node27556 : node27551;
															assign node27551 = (inp[5]) ? 4'b0010 : node27552;
																assign node27552 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node27556 = (inp[5]) ? node27558 : 4'b0010;
																assign node27558 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node27561 = (inp[13]) ? 4'b0000 : node27562;
														assign node27562 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node27566 = (inp[13]) ? 4'b0010 : node27567;
													assign node27567 = (inp[15]) ? node27571 : node27568;
														assign node27568 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node27571 = (inp[0]) ? node27575 : node27572;
															assign node27572 = (inp[3]) ? 4'b0010 : 4'b0000;
															assign node27575 = (inp[3]) ? 4'b0000 : node27576;
																assign node27576 = (inp[5]) ? 4'b0000 : 4'b0010;
							assign node27581 = (inp[13]) ? node27861 : node27582;
								assign node27582 = (inp[3]) ? node27728 : node27583;
									assign node27583 = (inp[15]) ? node27665 : node27584;
										assign node27584 = (inp[0]) ? node27620 : node27585;
											assign node27585 = (inp[5]) ? node27599 : node27586;
												assign node27586 = (inp[12]) ? node27594 : node27587;
													assign node27587 = (inp[4]) ? node27591 : node27588;
														assign node27588 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node27591 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node27594 = (inp[2]) ? node27596 : 4'b0110;
														assign node27596 = (inp[10]) ? 4'b0010 : 4'b0110;
												assign node27599 = (inp[4]) ? node27611 : node27600;
													assign node27600 = (inp[9]) ? node27606 : node27601;
														assign node27601 = (inp[12]) ? node27603 : 4'b0110;
															assign node27603 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node27606 = (inp[10]) ? node27608 : 4'b0010;
															assign node27608 = (inp[12]) ? 4'b0100 : 4'b0010;
													assign node27611 = (inp[12]) ? node27615 : node27612;
														assign node27612 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node27615 = (inp[9]) ? node27617 : 4'b0100;
															assign node27617 = (inp[10]) ? 4'b0000 : 4'b0100;
											assign node27620 = (inp[5]) ? node27650 : node27621;
												assign node27621 = (inp[12]) ? node27631 : node27622;
													assign node27622 = (inp[2]) ? 4'b0000 : node27623;
														assign node27623 = (inp[4]) ? node27627 : node27624;
															assign node27624 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node27627 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node27631 = (inp[10]) ? node27641 : node27632;
														assign node27632 = (inp[2]) ? node27638 : node27633;
															assign node27633 = (inp[4]) ? 4'b0000 : node27634;
																assign node27634 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node27638 = (inp[9]) ? 4'b0100 : 4'b0000;
														assign node27641 = (inp[2]) ? node27643 : 4'b0100;
															assign node27643 = (inp[4]) ? node27647 : node27644;
																assign node27644 = (inp[9]) ? 4'b0100 : 4'b0000;
																assign node27647 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node27650 = (inp[4]) ? node27654 : node27651;
													assign node27651 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node27654 = (inp[9]) ? node27660 : node27655;
														assign node27655 = (inp[2]) ? node27657 : 4'b0000;
															assign node27657 = (inp[10]) ? 4'b0110 : 4'b0000;
														assign node27660 = (inp[10]) ? node27662 : 4'b0110;
															assign node27662 = (inp[2]) ? 4'b0110 : 4'b0010;
										assign node27665 = (inp[0]) ? node27697 : node27666;
											assign node27666 = (inp[5]) ? node27680 : node27667;
												assign node27667 = (inp[10]) ? node27673 : node27668;
													assign node27668 = (inp[4]) ? 4'b0100 : node27669;
														assign node27669 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node27673 = (inp[4]) ? 4'b0000 : node27674;
														assign node27674 = (inp[2]) ? 4'b0100 : node27675;
															assign node27675 = (inp[9]) ? 4'b0000 : 4'b0100;
												assign node27680 = (inp[9]) ? node27688 : node27681;
													assign node27681 = (inp[2]) ? node27685 : node27682;
														assign node27682 = (inp[10]) ? 4'b0110 : 4'b0100;
														assign node27685 = (inp[10]) ? 4'b0000 : 4'b0100;
													assign node27688 = (inp[2]) ? node27690 : 4'b0110;
														assign node27690 = (inp[12]) ? node27692 : 4'b0110;
															assign node27692 = (inp[10]) ? node27694 : 4'b0000;
																assign node27694 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node27697 = (inp[5]) ? node27717 : node27698;
												assign node27698 = (inp[12]) ? node27700 : 4'b0110;
													assign node27700 = (inp[2]) ? node27708 : node27701;
														assign node27701 = (inp[10]) ? 4'b0110 : node27702;
															assign node27702 = (inp[4]) ? node27704 : 4'b0110;
																assign node27704 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node27708 = (inp[4]) ? node27710 : 4'b0010;
															assign node27710 = (inp[10]) ? node27714 : node27711;
																assign node27711 = (inp[9]) ? 4'b0110 : 4'b0010;
																assign node27714 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node27717 = (inp[9]) ? 4'b0010 : node27718;
													assign node27718 = (inp[10]) ? node27722 : node27719;
														assign node27719 = (inp[4]) ? 4'b0010 : 4'b0110;
														assign node27722 = (inp[4]) ? node27724 : 4'b0010;
															assign node27724 = (inp[12]) ? 4'b0100 : 4'b0010;
									assign node27728 = (inp[10]) ? node27790 : node27729;
										assign node27729 = (inp[4]) ? node27759 : node27730;
											assign node27730 = (inp[9]) ? node27744 : node27731;
												assign node27731 = (inp[15]) ? node27739 : node27732;
													assign node27732 = (inp[0]) ? node27736 : node27733;
														assign node27733 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node27736 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node27739 = (inp[5]) ? node27741 : 4'b0110;
														assign node27741 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node27744 = (inp[5]) ? node27752 : node27745;
													assign node27745 = (inp[15]) ? node27749 : node27746;
														assign node27746 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node27749 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node27752 = (inp[2]) ? node27754 : 4'b0000;
														assign node27754 = (inp[15]) ? 4'b0000 : node27755;
															assign node27755 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node27759 = (inp[9]) ? node27775 : node27760;
												assign node27760 = (inp[15]) ? node27768 : node27761;
													assign node27761 = (inp[0]) ? node27765 : node27762;
														assign node27762 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node27765 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node27768 = (inp[0]) ? node27772 : node27769;
														assign node27769 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node27772 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node27775 = (inp[2]) ? node27787 : node27776;
													assign node27776 = (inp[12]) ? node27782 : node27777;
														assign node27777 = (inp[0]) ? node27779 : 4'b0100;
															assign node27779 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node27782 = (inp[5]) ? 4'b0110 : node27783;
															assign node27783 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node27787 = (inp[12]) ? 4'b0100 : 4'b0110;
										assign node27790 = (inp[9]) ? node27828 : node27791;
											assign node27791 = (inp[12]) ? node27811 : node27792;
												assign node27792 = (inp[4]) ? 4'b0010 : node27793;
													assign node27793 = (inp[2]) ? node27799 : node27794;
														assign node27794 = (inp[5]) ? 4'b0110 : node27795;
															assign node27795 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node27799 = (inp[5]) ? node27805 : node27800;
															assign node27800 = (inp[0]) ? node27802 : 4'b0110;
																assign node27802 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node27805 = (inp[0]) ? node27807 : 4'b0100;
																assign node27807 = (inp[15]) ? 4'b0100 : 4'b0110;
												assign node27811 = (inp[4]) ? node27823 : node27812;
													assign node27812 = (inp[15]) ? node27814 : 4'b0000;
														assign node27814 = (inp[2]) ? node27818 : node27815;
															assign node27815 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node27818 = (inp[5]) ? 4'b0010 : node27819;
																assign node27819 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node27823 = (inp[0]) ? 4'b0100 : node27824;
														assign node27824 = (inp[2]) ? 4'b0100 : 4'b0110;
											assign node27828 = (inp[15]) ? node27844 : node27829;
												assign node27829 = (inp[0]) ? node27835 : node27830;
													assign node27830 = (inp[12]) ? 4'b0000 : node27831;
														assign node27831 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node27835 = (inp[12]) ? node27841 : node27836;
														assign node27836 = (inp[4]) ? 4'b0110 : node27837;
															assign node27837 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node27841 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node27844 = (inp[0]) ? node27852 : node27845;
													assign node27845 = (inp[12]) ? 4'b0110 : node27846;
														assign node27846 = (inp[4]) ? 4'b0110 : node27847;
															assign node27847 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node27852 = (inp[12]) ? node27858 : node27853;
														assign node27853 = (inp[4]) ? 4'b0100 : node27854;
															assign node27854 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node27858 = (inp[4]) ? 4'b0000 : 4'b0100;
								assign node27861 = (inp[4]) ? node28015 : node27862;
									assign node27862 = (inp[9]) ? node27934 : node27863;
										assign node27863 = (inp[12]) ? node27913 : node27864;
											assign node27864 = (inp[10]) ? node27888 : node27865;
												assign node27865 = (inp[3]) ? node27873 : node27866;
													assign node27866 = (inp[5]) ? 4'b1100 : node27867;
														assign node27867 = (inp[0]) ? 4'b1100 : node27868;
															assign node27868 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node27873 = (inp[5]) ? node27877 : node27874;
														assign node27874 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node27877 = (inp[2]) ? node27883 : node27878;
															assign node27878 = (inp[15]) ? node27880 : 4'b1110;
																assign node27880 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node27883 = (inp[0]) ? 4'b1100 : node27884;
																assign node27884 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node27888 = (inp[5]) ? node27904 : node27889;
													assign node27889 = (inp[2]) ? node27895 : node27890;
														assign node27890 = (inp[0]) ? node27892 : 4'b1010;
															assign node27892 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node27895 = (inp[3]) ? 4'b1000 : node27896;
															assign node27896 = (inp[15]) ? node27900 : node27897;
																assign node27897 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node27900 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node27904 = (inp[2]) ? node27906 : 4'b1000;
														assign node27906 = (inp[0]) ? node27908 : 4'b1000;
															assign node27908 = (inp[3]) ? node27910 : 4'b1010;
																assign node27910 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node27913 = (inp[15]) ? node27925 : node27914;
												assign node27914 = (inp[0]) ? node27920 : node27915;
													assign node27915 = (inp[3]) ? node27917 : 4'b1010;
														assign node27917 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node27920 = (inp[3]) ? node27922 : 4'b1000;
														assign node27922 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node27925 = (inp[5]) ? node27927 : 4'b1010;
													assign node27927 = (inp[3]) ? node27931 : node27928;
														assign node27928 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node27931 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node27934 = (inp[12]) ? node27982 : node27935;
											assign node27935 = (inp[10]) ? node27949 : node27936;
												assign node27936 = (inp[15]) ? node27944 : node27937;
													assign node27937 = (inp[0]) ? node27941 : node27938;
														assign node27938 = (inp[3]) ? 4'b1000 : 4'b1010;
														assign node27941 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node27944 = (inp[0]) ? node27946 : 4'b1000;
														assign node27946 = (inp[3]) ? 4'b1000 : 4'b1010;
												assign node27949 = (inp[5]) ? node27963 : node27950;
													assign node27950 = (inp[3]) ? node27958 : node27951;
														assign node27951 = (inp[0]) ? node27955 : node27952;
															assign node27952 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node27955 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node27958 = (inp[15]) ? 4'b1100 : node27959;
															assign node27959 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node27963 = (inp[2]) ? node27971 : node27964;
														assign node27964 = (inp[0]) ? node27968 : node27965;
															assign node27965 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node27968 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node27971 = (inp[3]) ? node27977 : node27972;
															assign node27972 = (inp[0]) ? 4'b1110 : node27973;
																assign node27973 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node27977 = (inp[15]) ? node27979 : 4'b1110;
																assign node27979 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node27982 = (inp[2]) ? node27996 : node27983;
												assign node27983 = (inp[0]) ? node27985 : 4'b1110;
													assign node27985 = (inp[15]) ? node27991 : node27986;
														assign node27986 = (inp[3]) ? 4'b1110 : node27987;
															assign node27987 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node27991 = (inp[3]) ? 4'b1100 : node27992;
															assign node27992 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node27996 = (inp[15]) ? node28006 : node27997;
													assign node27997 = (inp[3]) ? 4'b1100 : node27998;
														assign node27998 = (inp[5]) ? node28002 : node27999;
															assign node27999 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node28002 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node28006 = (inp[0]) ? node28012 : node28007;
														assign node28007 = (inp[5]) ? 4'b1110 : node28008;
															assign node28008 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node28012 = (inp[3]) ? 4'b1100 : 4'b1110;
									assign node28015 = (inp[9]) ? node28077 : node28016;
										assign node28016 = (inp[10]) ? node28054 : node28017;
											assign node28017 = (inp[12]) ? node28035 : node28018;
												assign node28018 = (inp[5]) ? node28026 : node28019;
													assign node28019 = (inp[15]) ? node28023 : node28020;
														assign node28020 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node28023 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node28026 = (inp[15]) ? 4'b1010 : node28027;
														assign node28027 = (inp[2]) ? node28029 : 4'b1000;
															assign node28029 = (inp[3]) ? 4'b1010 : node28030;
																assign node28030 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node28035 = (inp[2]) ? node28045 : node28036;
													assign node28036 = (inp[5]) ? node28038 : 4'b1100;
														assign node28038 = (inp[15]) ? node28042 : node28039;
															assign node28039 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node28042 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node28045 = (inp[0]) ? node28047 : 4'b1110;
														assign node28047 = (inp[15]) ? node28051 : node28048;
															assign node28048 = (inp[5]) ? 4'b1110 : 4'b1100;
															assign node28051 = (inp[5]) ? 4'b1100 : 4'b1110;
											assign node28054 = (inp[15]) ? node28066 : node28055;
												assign node28055 = (inp[0]) ? node28061 : node28056;
													assign node28056 = (inp[5]) ? 4'b1100 : node28057;
														assign node28057 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node28061 = (inp[5]) ? 4'b1110 : node28062;
														assign node28062 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node28066 = (inp[0]) ? node28072 : node28067;
													assign node28067 = (inp[5]) ? 4'b1110 : node28068;
														assign node28068 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node28072 = (inp[3]) ? 4'b1100 : node28073;
														assign node28073 = (inp[12]) ? 4'b1100 : 4'b1110;
										assign node28077 = (inp[10]) ? node28115 : node28078;
											assign node28078 = (inp[12]) ? node28094 : node28079;
												assign node28079 = (inp[15]) ? node28083 : node28080;
													assign node28080 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node28083 = (inp[0]) ? node28089 : node28084;
														assign node28084 = (inp[3]) ? 4'b1110 : node28085;
															assign node28085 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node28089 = (inp[3]) ? 4'b1100 : node28090;
															assign node28090 = (inp[2]) ? 4'b1110 : 4'b1100;
												assign node28094 = (inp[0]) ? node28104 : node28095;
													assign node28095 = (inp[15]) ? node28101 : node28096;
														assign node28096 = (inp[3]) ? 4'b1000 : node28097;
															assign node28097 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node28101 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node28104 = (inp[3]) ? 4'b1010 : node28105;
														assign node28105 = (inp[2]) ? node28111 : node28106;
															assign node28106 = (inp[15]) ? 4'b1010 : node28107;
																assign node28107 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node28111 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node28115 = (inp[0]) ? node28127 : node28116;
												assign node28116 = (inp[15]) ? node28122 : node28117;
													assign node28117 = (inp[5]) ? 4'b1000 : node28118;
														assign node28118 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node28122 = (inp[5]) ? 4'b1010 : node28123;
														assign node28123 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node28127 = (inp[15]) ? node28133 : node28128;
													assign node28128 = (inp[5]) ? 4'b1010 : node28129;
														assign node28129 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node28133 = (inp[3]) ? 4'b1000 : node28134;
														assign node28134 = (inp[5]) ? 4'b1000 : 4'b1010;
						assign node28138 = (inp[1]) ? node28708 : node28139;
							assign node28139 = (inp[9]) ? node28463 : node28140;
								assign node28140 = (inp[4]) ? node28298 : node28141;
									assign node28141 = (inp[12]) ? node28235 : node28142;
										assign node28142 = (inp[10]) ? node28192 : node28143;
											assign node28143 = (inp[3]) ? node28173 : node28144;
												assign node28144 = (inp[2]) ? node28160 : node28145;
													assign node28145 = (inp[13]) ? node28153 : node28146;
														assign node28146 = (inp[0]) ? node28150 : node28147;
															assign node28147 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node28150 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node28153 = (inp[5]) ? node28155 : 4'b1100;
															assign node28155 = (inp[15]) ? 4'b1100 : node28156;
																assign node28156 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node28160 = (inp[13]) ? node28166 : node28161;
														assign node28161 = (inp[0]) ? 4'b1100 : node28162;
															assign node28162 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node28166 = (inp[5]) ? 4'b1110 : node28167;
															assign node28167 = (inp[15]) ? 4'b1110 : node28168;
																assign node28168 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node28173 = (inp[5]) ? node28179 : node28174;
													assign node28174 = (inp[15]) ? node28176 : 4'b1110;
														assign node28176 = (inp[2]) ? 4'b1100 : 4'b1110;
													assign node28179 = (inp[13]) ? node28185 : node28180;
														assign node28180 = (inp[15]) ? node28182 : 4'b1110;
															assign node28182 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node28185 = (inp[0]) ? node28189 : node28186;
															assign node28186 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node28189 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node28192 = (inp[2]) ? node28208 : node28193;
												assign node28193 = (inp[0]) ? node28199 : node28194;
													assign node28194 = (inp[15]) ? node28196 : 4'b1010;
														assign node28196 = (inp[13]) ? 4'b1000 : 4'b1010;
													assign node28199 = (inp[3]) ? node28201 : 4'b1000;
														assign node28201 = (inp[15]) ? node28205 : node28202;
															assign node28202 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node28205 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node28208 = (inp[5]) ? node28226 : node28209;
													assign node28209 = (inp[13]) ? node28217 : node28210;
														assign node28210 = (inp[15]) ? node28214 : node28211;
															assign node28211 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node28214 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node28217 = (inp[3]) ? node28219 : 4'b1000;
															assign node28219 = (inp[0]) ? node28223 : node28220;
																assign node28220 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node28223 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node28226 = (inp[0]) ? node28228 : 4'b1000;
														assign node28228 = (inp[13]) ? node28230 : 4'b1000;
															assign node28230 = (inp[15]) ? 4'b1010 : node28231;
																assign node28231 = (inp[3]) ? 4'b1010 : 4'b1000;
										assign node28235 = (inp[13]) ? node28275 : node28236;
											assign node28236 = (inp[5]) ? node28260 : node28237;
												assign node28237 = (inp[2]) ? node28247 : node28238;
													assign node28238 = (inp[10]) ? 4'b1010 : node28239;
														assign node28239 = (inp[0]) ? node28243 : node28240;
															assign node28240 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node28243 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node28247 = (inp[3]) ? node28253 : node28248;
														assign node28248 = (inp[15]) ? 4'b1000 : node28249;
															assign node28249 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node28253 = (inp[10]) ? node28255 : 4'b1010;
															assign node28255 = (inp[0]) ? node28257 : 4'b1000;
																assign node28257 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node28260 = (inp[2]) ? node28270 : node28261;
													assign node28261 = (inp[3]) ? 4'b1010 : node28262;
														assign node28262 = (inp[0]) ? node28266 : node28263;
															assign node28263 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node28266 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node28270 = (inp[3]) ? node28272 : 4'b1010;
														assign node28272 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node28275 = (inp[0]) ? node28287 : node28276;
												assign node28276 = (inp[15]) ? node28282 : node28277;
													assign node28277 = (inp[3]) ? node28279 : 4'b1010;
														assign node28279 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node28282 = (inp[3]) ? node28284 : 4'b1000;
														assign node28284 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node28287 = (inp[15]) ? node28293 : node28288;
													assign node28288 = (inp[3]) ? node28290 : 4'b1000;
														assign node28290 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node28293 = (inp[3]) ? node28295 : 4'b1010;
														assign node28295 = (inp[5]) ? 4'b1000 : 4'b1010;
									assign node28298 = (inp[12]) ? node28362 : node28299;
										assign node28299 = (inp[10]) ? node28339 : node28300;
											assign node28300 = (inp[13]) ? node28316 : node28301;
												assign node28301 = (inp[0]) ? node28307 : node28302;
													assign node28302 = (inp[15]) ? 4'b1000 : node28303;
														assign node28303 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node28307 = (inp[5]) ? node28311 : node28308;
														assign node28308 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28311 = (inp[3]) ? node28313 : 4'b1000;
															assign node28313 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node28316 = (inp[2]) ? node28334 : node28317;
													assign node28317 = (inp[5]) ? node28325 : node28318;
														assign node28318 = (inp[0]) ? node28322 : node28319;
															assign node28319 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node28322 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28325 = (inp[15]) ? 4'b1000 : node28326;
															assign node28326 = (inp[0]) ? node28330 : node28327;
																assign node28327 = (inp[3]) ? 4'b1000 : 4'b1010;
																assign node28330 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node28334 = (inp[15]) ? 4'b1010 : node28335;
														assign node28335 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node28339 = (inp[15]) ? node28351 : node28340;
												assign node28340 = (inp[0]) ? node28346 : node28341;
													assign node28341 = (inp[5]) ? 4'b1100 : node28342;
														assign node28342 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node28346 = (inp[3]) ? 4'b1110 : node28347;
														assign node28347 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node28351 = (inp[0]) ? node28357 : node28352;
													assign node28352 = (inp[5]) ? 4'b1110 : node28353;
														assign node28353 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node28357 = (inp[5]) ? 4'b1100 : node28358;
														assign node28358 = (inp[3]) ? 4'b1100 : 4'b1110;
										assign node28362 = (inp[5]) ? node28426 : node28363;
											assign node28363 = (inp[2]) ? node28399 : node28364;
												assign node28364 = (inp[15]) ? node28378 : node28365;
													assign node28365 = (inp[10]) ? node28373 : node28366;
														assign node28366 = (inp[3]) ? node28370 : node28367;
															assign node28367 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node28370 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node28373 = (inp[0]) ? 4'b1100 : node28374;
															assign node28374 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node28378 = (inp[10]) ? node28384 : node28379;
														assign node28379 = (inp[3]) ? 4'b1100 : node28380;
															assign node28380 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node28384 = (inp[13]) ? node28392 : node28385;
															assign node28385 = (inp[3]) ? node28389 : node28386;
																assign node28386 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node28389 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node28392 = (inp[0]) ? node28396 : node28393;
																assign node28393 = (inp[3]) ? 4'b1110 : 4'b1100;
																assign node28396 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node28399 = (inp[3]) ? node28413 : node28400;
													assign node28400 = (inp[10]) ? node28402 : 4'b1100;
														assign node28402 = (inp[13]) ? node28408 : node28403;
															assign node28403 = (inp[0]) ? node28405 : 4'b1110;
																assign node28405 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node28408 = (inp[0]) ? 4'b1110 : node28409;
																assign node28409 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node28413 = (inp[10]) ? node28419 : node28414;
														assign node28414 = (inp[0]) ? node28416 : 4'b1110;
															assign node28416 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node28419 = (inp[13]) ? 4'b1110 : node28420;
															assign node28420 = (inp[0]) ? 4'b1100 : node28421;
																assign node28421 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node28426 = (inp[3]) ? node28450 : node28427;
												assign node28427 = (inp[10]) ? node28443 : node28428;
													assign node28428 = (inp[13]) ? node28436 : node28429;
														assign node28429 = (inp[0]) ? node28433 : node28430;
															assign node28430 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node28433 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node28436 = (inp[0]) ? node28440 : node28437;
															assign node28437 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node28440 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node28443 = (inp[15]) ? node28447 : node28444;
														assign node28444 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node28447 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node28450 = (inp[10]) ? node28456 : node28451;
													assign node28451 = (inp[15]) ? 4'b1100 : node28452;
														assign node28452 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node28456 = (inp[0]) ? node28460 : node28457;
														assign node28457 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node28460 = (inp[15]) ? 4'b1100 : 4'b1110;
								assign node28463 = (inp[4]) ? node28591 : node28464;
									assign node28464 = (inp[12]) ? node28522 : node28465;
										assign node28465 = (inp[10]) ? node28489 : node28466;
											assign node28466 = (inp[15]) ? node28478 : node28467;
												assign node28467 = (inp[0]) ? node28473 : node28468;
													assign node28468 = (inp[5]) ? node28470 : 4'b1010;
														assign node28470 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node28473 = (inp[3]) ? node28475 : 4'b1000;
														assign node28475 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node28478 = (inp[0]) ? node28484 : node28479;
													assign node28479 = (inp[5]) ? node28481 : 4'b1000;
														assign node28481 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node28484 = (inp[3]) ? node28486 : 4'b1010;
														assign node28486 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node28489 = (inp[5]) ? node28507 : node28490;
												assign node28490 = (inp[15]) ? node28492 : 4'b1100;
													assign node28492 = (inp[13]) ? node28502 : node28493;
														assign node28493 = (inp[2]) ? node28495 : 4'b1110;
															assign node28495 = (inp[3]) ? node28499 : node28496;
																assign node28496 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node28499 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node28502 = (inp[0]) ? 4'b1100 : node28503;
															assign node28503 = (inp[3]) ? 4'b1110 : 4'b1100;
												assign node28507 = (inp[2]) ? node28515 : node28508;
													assign node28508 = (inp[13]) ? 4'b1110 : node28509;
														assign node28509 = (inp[0]) ? 4'b1110 : node28510;
															assign node28510 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node28515 = (inp[0]) ? node28519 : node28516;
														assign node28516 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node28519 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node28522 = (inp[2]) ? node28566 : node28523;
											assign node28523 = (inp[13]) ? node28543 : node28524;
												assign node28524 = (inp[15]) ? node28536 : node28525;
													assign node28525 = (inp[3]) ? node28533 : node28526;
														assign node28526 = (inp[0]) ? node28530 : node28527;
															assign node28527 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node28530 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node28533 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node28536 = (inp[3]) ? 4'b1110 : node28537;
														assign node28537 = (inp[5]) ? node28539 : 4'b1100;
															assign node28539 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node28543 = (inp[5]) ? node28555 : node28544;
													assign node28544 = (inp[0]) ? 4'b1110 : node28545;
														assign node28545 = (inp[10]) ? node28549 : node28546;
															assign node28546 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node28549 = (inp[15]) ? 4'b1110 : node28550;
																assign node28550 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node28555 = (inp[10]) ? node28561 : node28556;
														assign node28556 = (inp[15]) ? node28558 : 4'b1110;
															assign node28558 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node28561 = (inp[15]) ? 4'b1110 : node28562;
															assign node28562 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node28566 = (inp[5]) ? node28582 : node28567;
												assign node28567 = (inp[15]) ? node28575 : node28568;
													assign node28568 = (inp[3]) ? node28572 : node28569;
														assign node28569 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node28572 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node28575 = (inp[0]) ? node28579 : node28576;
														assign node28576 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node28579 = (inp[3]) ? 4'b1100 : 4'b1110;
												assign node28582 = (inp[13]) ? node28584 : 4'b1100;
													assign node28584 = (inp[15]) ? node28588 : node28585;
														assign node28585 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node28588 = (inp[0]) ? 4'b1100 : 4'b1110;
									assign node28591 = (inp[12]) ? node28663 : node28592;
										assign node28592 = (inp[10]) ? node28640 : node28593;
											assign node28593 = (inp[2]) ? node28617 : node28594;
												assign node28594 = (inp[0]) ? node28606 : node28595;
													assign node28595 = (inp[13]) ? 4'b1100 : node28596;
														assign node28596 = (inp[5]) ? 4'b1100 : node28597;
															assign node28597 = (inp[15]) ? node28601 : node28598;
																assign node28598 = (inp[3]) ? 4'b1100 : 4'b1110;
																assign node28601 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node28606 = (inp[15]) ? node28612 : node28607;
														assign node28607 = (inp[5]) ? 4'b1110 : node28608;
															assign node28608 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node28612 = (inp[5]) ? 4'b1100 : node28613;
															assign node28613 = (inp[13]) ? 4'b1110 : 4'b1100;
												assign node28617 = (inp[13]) ? node28633 : node28618;
													assign node28618 = (inp[15]) ? node28624 : node28619;
														assign node28619 = (inp[5]) ? node28621 : 4'b1100;
															assign node28621 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node28624 = (inp[0]) ? node28630 : node28625;
															assign node28625 = (inp[5]) ? 4'b1110 : node28626;
																assign node28626 = (inp[3]) ? 4'b1110 : 4'b1100;
															assign node28630 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node28633 = (inp[15]) ? 4'b1110 : node28634;
														assign node28634 = (inp[0]) ? 4'b1110 : node28635;
															assign node28635 = (inp[3]) ? 4'b1100 : 4'b1110;
											assign node28640 = (inp[0]) ? node28652 : node28641;
												assign node28641 = (inp[15]) ? node28647 : node28642;
													assign node28642 = (inp[3]) ? 4'b1000 : node28643;
														assign node28643 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node28647 = (inp[5]) ? 4'b1010 : node28648;
														assign node28648 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node28652 = (inp[15]) ? node28658 : node28653;
													assign node28653 = (inp[2]) ? 4'b1010 : node28654;
														assign node28654 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node28658 = (inp[5]) ? 4'b1000 : node28659;
														assign node28659 = (inp[3]) ? 4'b1000 : 4'b1010;
										assign node28663 = (inp[2]) ? node28687 : node28664;
											assign node28664 = (inp[15]) ? node28676 : node28665;
												assign node28665 = (inp[0]) ? node28671 : node28666;
													assign node28666 = (inp[5]) ? 4'b1000 : node28667;
														assign node28667 = (inp[3]) ? 4'b1000 : 4'b1010;
													assign node28671 = (inp[5]) ? 4'b1010 : node28672;
														assign node28672 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node28676 = (inp[0]) ? node28682 : node28677;
													assign node28677 = (inp[3]) ? 4'b1010 : node28678;
														assign node28678 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node28682 = (inp[3]) ? 4'b1000 : node28683;
														assign node28683 = (inp[5]) ? 4'b1000 : 4'b1010;
											assign node28687 = (inp[15]) ? node28699 : node28688;
												assign node28688 = (inp[0]) ? node28694 : node28689;
													assign node28689 = (inp[3]) ? 4'b1000 : node28690;
														assign node28690 = (inp[13]) ? 4'b1010 : 4'b1000;
													assign node28694 = (inp[5]) ? 4'b1010 : node28695;
														assign node28695 = (inp[3]) ? 4'b1010 : 4'b1000;
												assign node28699 = (inp[0]) ? node28703 : node28700;
													assign node28700 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node28703 = (inp[5]) ? 4'b1000 : node28704;
														assign node28704 = (inp[3]) ? 4'b1000 : 4'b1010;
							assign node28708 = (inp[13]) ? node29072 : node28709;
								assign node28709 = (inp[5]) ? node28877 : node28710;
									assign node28710 = (inp[10]) ? node28796 : node28711;
										assign node28711 = (inp[4]) ? node28753 : node28712;
											assign node28712 = (inp[2]) ? node28738 : node28713;
												assign node28713 = (inp[15]) ? node28721 : node28714;
													assign node28714 = (inp[0]) ? node28716 : 4'b1010;
														assign node28716 = (inp[12]) ? 4'b1000 : node28717;
															assign node28717 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node28721 = (inp[0]) ? node28731 : node28722;
														assign node28722 = (inp[9]) ? node28726 : node28723;
															assign node28723 = (inp[12]) ? 4'b1000 : 4'b1100;
															assign node28726 = (inp[12]) ? node28728 : 4'b1000;
																assign node28728 = (inp[3]) ? 4'b1110 : 4'b1100;
														assign node28731 = (inp[12]) ? node28735 : node28732;
															assign node28732 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node28735 = (inp[9]) ? 4'b1110 : 4'b1010;
												assign node28738 = (inp[12]) ? node28742 : node28739;
													assign node28739 = (inp[9]) ? 4'b1010 : 4'b1110;
													assign node28742 = (inp[9]) ? node28744 : 4'b1010;
														assign node28744 = (inp[0]) ? node28746 : 4'b1110;
															assign node28746 = (inp[3]) ? node28750 : node28747;
																assign node28747 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node28750 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node28753 = (inp[9]) ? node28771 : node28754;
												assign node28754 = (inp[12]) ? node28764 : node28755;
													assign node28755 = (inp[2]) ? node28757 : 4'b1010;
														assign node28757 = (inp[15]) ? node28761 : node28758;
															assign node28758 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node28761 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node28764 = (inp[15]) ? node28766 : 4'b1100;
														assign node28766 = (inp[2]) ? 4'b1110 : node28767;
															assign node28767 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node28771 = (inp[12]) ? node28783 : node28772;
													assign node28772 = (inp[15]) ? node28778 : node28773;
														assign node28773 = (inp[3]) ? 4'b1100 : node28774;
															assign node28774 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node28778 = (inp[0]) ? 4'b1110 : node28779;
															assign node28779 = (inp[3]) ? 4'b1110 : 4'b1100;
													assign node28783 = (inp[0]) ? node28791 : node28784;
														assign node28784 = (inp[3]) ? node28788 : node28785;
															assign node28785 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node28788 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28791 = (inp[3]) ? node28793 : 4'b1000;
															assign node28793 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node28796 = (inp[15]) ? node28834 : node28797;
											assign node28797 = (inp[4]) ? node28811 : node28798;
												assign node28798 = (inp[9]) ? node28802 : node28799;
													assign node28799 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node28802 = (inp[12]) ? 4'b1110 : node28803;
														assign node28803 = (inp[2]) ? node28805 : 4'b1110;
															assign node28805 = (inp[3]) ? node28807 : 4'b1100;
																assign node28807 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node28811 = (inp[9]) ? node28831 : node28812;
													assign node28812 = (inp[2]) ? node28820 : node28813;
														assign node28813 = (inp[3]) ? node28817 : node28814;
															assign node28814 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node28817 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node28820 = (inp[12]) ? node28826 : node28821;
															assign node28821 = (inp[3]) ? 4'b1110 : node28822;
																assign node28822 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node28826 = (inp[0]) ? 4'b1110 : node28827;
																assign node28827 = (inp[3]) ? 4'b1100 : 4'b1110;
													assign node28831 = (inp[12]) ? 4'b1010 : 4'b1000;
											assign node28834 = (inp[0]) ? node28856 : node28835;
												assign node28835 = (inp[3]) ? node28849 : node28836;
													assign node28836 = (inp[2]) ? node28842 : node28837;
														assign node28837 = (inp[12]) ? 4'b1000 : node28838;
															assign node28838 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node28842 = (inp[12]) ? 4'b1100 : node28843;
															assign node28843 = (inp[9]) ? node28845 : 4'b1000;
																assign node28845 = (inp[4]) ? 4'b1000 : 4'b1100;
													assign node28849 = (inp[9]) ? node28853 : node28850;
														assign node28850 = (inp[4]) ? 4'b1110 : 4'b1000;
														assign node28853 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node28856 = (inp[3]) ? node28870 : node28857;
													assign node28857 = (inp[12]) ? node28865 : node28858;
														assign node28858 = (inp[4]) ? node28862 : node28859;
															assign node28859 = (inp[9]) ? 4'b1110 : 4'b1010;
															assign node28862 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node28865 = (inp[2]) ? 4'b1010 : node28866;
															assign node28866 = (inp[4]) ? 4'b1110 : 4'b1010;
													assign node28870 = (inp[4]) ? node28874 : node28871;
														assign node28871 = (inp[9]) ? 4'b1100 : 4'b1010;
														assign node28874 = (inp[9]) ? 4'b1000 : 4'b1100;
									assign node28877 = (inp[12]) ? node28975 : node28878;
										assign node28878 = (inp[10]) ? node28926 : node28879;
											assign node28879 = (inp[0]) ? node28901 : node28880;
												assign node28880 = (inp[9]) ? node28892 : node28881;
													assign node28881 = (inp[4]) ? node28887 : node28882;
														assign node28882 = (inp[15]) ? 4'b1110 : node28883;
															assign node28883 = (inp[3]) ? 4'b1100 : 4'b1110;
														assign node28887 = (inp[3]) ? node28889 : 4'b1010;
															assign node28889 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node28892 = (inp[4]) ? node28898 : node28893;
														assign node28893 = (inp[3]) ? node28895 : 4'b1000;
															assign node28895 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28898 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node28901 = (inp[3]) ? node28917 : node28902;
													assign node28902 = (inp[2]) ? node28908 : node28903;
														assign node28903 = (inp[4]) ? node28905 : 4'b1000;
															assign node28905 = (inp[15]) ? 4'b1010 : 4'b1110;
														assign node28908 = (inp[15]) ? node28914 : node28909;
															assign node28909 = (inp[4]) ? 4'b1000 : node28910;
																assign node28910 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node28914 = (inp[4]) ? 4'b1100 : 4'b1010;
													assign node28917 = (inp[15]) ? node28919 : 4'b1110;
														assign node28919 = (inp[9]) ? node28923 : node28920;
															assign node28920 = (inp[4]) ? 4'b1000 : 4'b1100;
															assign node28923 = (inp[4]) ? 4'b1100 : 4'b1000;
											assign node28926 = (inp[3]) ? node28948 : node28927;
												assign node28927 = (inp[0]) ? node28939 : node28928;
													assign node28928 = (inp[4]) ? node28934 : node28929;
														assign node28929 = (inp[9]) ? 4'b1110 : node28930;
															assign node28930 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node28934 = (inp[9]) ? node28936 : 4'b1100;
															assign node28936 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node28939 = (inp[4]) ? node28945 : node28940;
														assign node28940 = (inp[9]) ? 4'b1100 : node28941;
															assign node28941 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node28945 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node28948 = (inp[0]) ? node28964 : node28949;
													assign node28949 = (inp[15]) ? node28957 : node28950;
														assign node28950 = (inp[4]) ? node28954 : node28951;
															assign node28951 = (inp[2]) ? 4'b1100 : 4'b1000;
															assign node28954 = (inp[9]) ? 4'b1000 : 4'b1100;
														assign node28957 = (inp[9]) ? node28961 : node28958;
															assign node28958 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node28961 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node28964 = (inp[15]) ? node28970 : node28965;
														assign node28965 = (inp[4]) ? node28967 : 4'b1010;
															assign node28967 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node28970 = (inp[9]) ? 4'b1000 : node28971;
															assign node28971 = (inp[2]) ? 4'b1000 : 4'b1100;
										assign node28975 = (inp[10]) ? node29015 : node28976;
											assign node28976 = (inp[4]) ? node28996 : node28977;
												assign node28977 = (inp[9]) ? node28991 : node28978;
													assign node28978 = (inp[0]) ? node28986 : node28979;
														assign node28979 = (inp[15]) ? node28983 : node28980;
															assign node28980 = (inp[3]) ? 4'b1000 : 4'b1010;
															assign node28983 = (inp[3]) ? 4'b1010 : 4'b1000;
														assign node28986 = (inp[15]) ? 4'b1010 : node28987;
															assign node28987 = (inp[3]) ? 4'b1010 : 4'b1000;
													assign node28991 = (inp[15]) ? 4'b1100 : node28992;
														assign node28992 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node28996 = (inp[9]) ? node29004 : node28997;
													assign node28997 = (inp[15]) ? node29001 : node28998;
														assign node28998 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node29001 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node29004 = (inp[2]) ? node29010 : node29005;
														assign node29005 = (inp[3]) ? 4'b1010 : node29006;
															assign node29006 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node29010 = (inp[0]) ? node29012 : 4'b1010;
															assign node29012 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node29015 = (inp[2]) ? node29037 : node29016;
												assign node29016 = (inp[0]) ? node29024 : node29017;
													assign node29017 = (inp[15]) ? node29019 : 4'b1100;
														assign node29019 = (inp[4]) ? 4'b1110 : node29020;
															assign node29020 = (inp[9]) ? 4'b1110 : 4'b1000;
													assign node29024 = (inp[15]) ? node29032 : node29025;
														assign node29025 = (inp[3]) ? node29027 : 4'b1110;
															assign node29027 = (inp[9]) ? node29029 : 4'b1010;
																assign node29029 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node29032 = (inp[4]) ? node29034 : 4'b1100;
															assign node29034 = (inp[9]) ? 4'b1000 : 4'b1100;
												assign node29037 = (inp[3]) ? node29057 : node29038;
													assign node29038 = (inp[9]) ? node29048 : node29039;
														assign node29039 = (inp[4]) ? node29041 : 4'b1010;
															assign node29041 = (inp[15]) ? node29045 : node29042;
																assign node29042 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node29045 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node29048 = (inp[4]) ? node29052 : node29049;
															assign node29049 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node29052 = (inp[0]) ? node29054 : 4'b1000;
																assign node29054 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node29057 = (inp[9]) ? node29065 : node29058;
														assign node29058 = (inp[4]) ? 4'b1100 : node29059;
															assign node29059 = (inp[0]) ? node29061 : 4'b1000;
																assign node29061 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node29065 = (inp[4]) ? node29067 : 4'b1110;
															assign node29067 = (inp[0]) ? node29069 : 4'b1010;
																assign node29069 = (inp[15]) ? 4'b1000 : 4'b1010;
								assign node29072 = (inp[4]) ? node29200 : node29073;
									assign node29073 = (inp[9]) ? node29137 : node29074;
										assign node29074 = (inp[12]) ? node29100 : node29075;
											assign node29075 = (inp[10]) ? node29091 : node29076;
												assign node29076 = (inp[2]) ? 4'b0110 : node29077;
													assign node29077 = (inp[3]) ? node29083 : node29078;
														assign node29078 = (inp[0]) ? 4'b0110 : node29079;
															assign node29079 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node29083 = (inp[15]) ? 4'b0100 : node29084;
															assign node29084 = (inp[0]) ? 4'b0100 : node29085;
																assign node29085 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node29091 = (inp[0]) ? node29095 : node29092;
													assign node29092 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node29095 = (inp[15]) ? 4'b0010 : node29096;
														assign node29096 = (inp[3]) ? 4'b0010 : 4'b0000;
											assign node29100 = (inp[3]) ? node29114 : node29101;
												assign node29101 = (inp[5]) ? node29107 : node29102;
													assign node29102 = (inp[2]) ? 4'b0010 : node29103;
														assign node29103 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node29107 = (inp[15]) ? node29111 : node29108;
														assign node29108 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node29111 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node29114 = (inp[10]) ? node29130 : node29115;
													assign node29115 = (inp[5]) ? node29123 : node29116;
														assign node29116 = (inp[15]) ? node29120 : node29117;
															assign node29117 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node29120 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node29123 = (inp[2]) ? node29125 : 4'b0000;
															assign node29125 = (inp[15]) ? node29127 : 4'b0000;
																assign node29127 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node29130 = (inp[5]) ? 4'b0010 : node29131;
														assign node29131 = (inp[15]) ? 4'b0000 : node29132;
															assign node29132 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node29137 = (inp[12]) ? node29167 : node29138;
											assign node29138 = (inp[10]) ? node29156 : node29139;
												assign node29139 = (inp[0]) ? node29147 : node29140;
													assign node29140 = (inp[15]) ? 4'b0000 : node29141;
														assign node29141 = (inp[5]) ? node29143 : 4'b0010;
															assign node29143 = (inp[2]) ? 4'b0000 : 4'b0010;
													assign node29147 = (inp[15]) ? node29153 : node29148;
														assign node29148 = (inp[5]) ? node29150 : 4'b0000;
															assign node29150 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node29153 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node29156 = (inp[2]) ? node29162 : node29157;
													assign node29157 = (inp[15]) ? node29159 : 4'b0100;
														assign node29159 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node29162 = (inp[15]) ? node29164 : 4'b0110;
														assign node29164 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node29167 = (inp[3]) ? node29193 : node29168;
												assign node29168 = (inp[15]) ? node29174 : node29169;
													assign node29169 = (inp[0]) ? node29171 : 4'b0110;
														assign node29171 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node29174 = (inp[10]) ? node29182 : node29175;
														assign node29175 = (inp[0]) ? node29179 : node29176;
															assign node29176 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node29179 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node29182 = (inp[2]) ? node29188 : node29183;
															assign node29183 = (inp[5]) ? node29185 : 4'b0110;
																assign node29185 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node29188 = (inp[5]) ? 4'b0110 : node29189;
																assign node29189 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node29193 = (inp[0]) ? node29197 : node29194;
													assign node29194 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node29197 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node29200 = (inp[9]) ? node29272 : node29201;
										assign node29201 = (inp[12]) ? node29231 : node29202;
											assign node29202 = (inp[10]) ? node29218 : node29203;
												assign node29203 = (inp[0]) ? node29209 : node29204;
													assign node29204 = (inp[15]) ? 4'b0000 : node29205;
														assign node29205 = (inp[5]) ? 4'b0000 : 4'b0010;
													assign node29209 = (inp[15]) ? node29215 : node29210;
														assign node29210 = (inp[5]) ? node29212 : 4'b0000;
															assign node29212 = (inp[3]) ? 4'b0010 : 4'b0000;
														assign node29215 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node29218 = (inp[15]) ? node29226 : node29219;
													assign node29219 = (inp[0]) ? node29221 : 4'b0100;
														assign node29221 = (inp[5]) ? 4'b0110 : node29222;
															assign node29222 = (inp[3]) ? 4'b0110 : 4'b0100;
													assign node29226 = (inp[0]) ? 4'b0100 : node29227;
														assign node29227 = (inp[3]) ? 4'b0110 : 4'b0100;
											assign node29231 = (inp[10]) ? node29255 : node29232;
												assign node29232 = (inp[2]) ? node29246 : node29233;
													assign node29233 = (inp[15]) ? node29241 : node29234;
														assign node29234 = (inp[0]) ? node29238 : node29235;
															assign node29235 = (inp[3]) ? 4'b0100 : 4'b0110;
															assign node29238 = (inp[3]) ? 4'b0110 : 4'b0100;
														assign node29241 = (inp[5]) ? node29243 : 4'b0100;
															assign node29243 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node29246 = (inp[5]) ? node29248 : 4'b0110;
														assign node29248 = (inp[15]) ? node29252 : node29249;
															assign node29249 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node29252 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node29255 = (inp[5]) ? node29265 : node29256;
													assign node29256 = (inp[15]) ? 4'b0100 : node29257;
														assign node29257 = (inp[3]) ? node29261 : node29258;
															assign node29258 = (inp[0]) ? 4'b0100 : 4'b0110;
															assign node29261 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node29265 = (inp[0]) ? node29269 : node29266;
														assign node29266 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node29269 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node29272 = (inp[12]) ? node29306 : node29273;
											assign node29273 = (inp[10]) ? node29289 : node29274;
												assign node29274 = (inp[0]) ? node29280 : node29275;
													assign node29275 = (inp[5]) ? node29277 : 4'b0100;
														assign node29277 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node29280 = (inp[15]) ? node29286 : node29281;
														assign node29281 = (inp[3]) ? 4'b0110 : node29282;
															assign node29282 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node29286 = (inp[3]) ? 4'b0100 : 4'b0110;
												assign node29289 = (inp[15]) ? node29299 : node29290;
													assign node29290 = (inp[0]) ? node29296 : node29291;
														assign node29291 = (inp[2]) ? node29293 : 4'b0000;
															assign node29293 = (inp[3]) ? 4'b0000 : 4'b0010;
														assign node29296 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node29299 = (inp[0]) ? node29301 : 4'b0010;
														assign node29301 = (inp[5]) ? 4'b0000 : node29302;
															assign node29302 = (inp[3]) ? 4'b0000 : 4'b0010;
											assign node29306 = (inp[0]) ? node29318 : node29307;
												assign node29307 = (inp[15]) ? node29313 : node29308;
													assign node29308 = (inp[5]) ? 4'b0000 : node29309;
														assign node29309 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node29313 = (inp[3]) ? 4'b0010 : node29314;
														assign node29314 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node29318 = (inp[5]) ? node29324 : node29319;
													assign node29319 = (inp[15]) ? node29321 : 4'b0000;
														assign node29321 = (inp[3]) ? 4'b0000 : 4'b0010;
													assign node29324 = (inp[15]) ? 4'b0000 : 4'b0010;
				assign node29327 = (inp[11]) ? node31351 : node29328;
					assign node29328 = (inp[6]) ? node30356 : node29329;
						assign node29329 = (inp[13]) ? node29925 : node29330;
							assign node29330 = (inp[1]) ? node29610 : node29331;
								assign node29331 = (inp[15]) ? node29465 : node29332;
									assign node29332 = (inp[0]) ? node29390 : node29333;
										assign node29333 = (inp[5]) ? node29357 : node29334;
											assign node29334 = (inp[4]) ? node29346 : node29335;
												assign node29335 = (inp[9]) ? node29341 : node29336;
													assign node29336 = (inp[10]) ? node29338 : 4'b1111;
														assign node29338 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node29341 = (inp[10]) ? node29343 : 4'b1011;
														assign node29343 = (inp[12]) ? 4'b1111 : 4'b1011;
												assign node29346 = (inp[9]) ? node29354 : node29347;
													assign node29347 = (inp[12]) ? node29349 : 4'b1011;
														assign node29349 = (inp[10]) ? node29351 : 4'b1011;
															assign node29351 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node29354 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node29357 = (inp[3]) ? node29375 : node29358;
												assign node29358 = (inp[9]) ? node29368 : node29359;
													assign node29359 = (inp[4]) ? node29365 : node29360;
														assign node29360 = (inp[2]) ? 4'b1111 : node29361;
															assign node29361 = (inp[10]) ? 4'b1011 : 4'b1111;
														assign node29365 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node29368 = (inp[10]) ? node29370 : 4'b1101;
														assign node29370 = (inp[4]) ? node29372 : 4'b1101;
															assign node29372 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node29375 = (inp[12]) ? node29383 : node29376;
													assign node29376 = (inp[9]) ? node29380 : node29377;
														assign node29377 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node29380 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node29383 = (inp[10]) ? 4'b1101 : node29384;
														assign node29384 = (inp[4]) ? node29386 : 4'b1101;
															assign node29386 = (inp[9]) ? 4'b1101 : 4'b1001;
										assign node29390 = (inp[5]) ? node29434 : node29391;
											assign node29391 = (inp[3]) ? node29415 : node29392;
												assign node29392 = (inp[12]) ? node29400 : node29393;
													assign node29393 = (inp[4]) ? node29397 : node29394;
														assign node29394 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node29397 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node29400 = (inp[4]) ? 4'b1001 : node29401;
														assign node29401 = (inp[2]) ? node29409 : node29402;
															assign node29402 = (inp[10]) ? node29406 : node29403;
																assign node29403 = (inp[9]) ? 4'b1001 : 4'b1101;
																assign node29406 = (inp[9]) ? 4'b1101 : 4'b1001;
															assign node29409 = (inp[9]) ? node29411 : 4'b1001;
																assign node29411 = (inp[10]) ? 4'b1101 : 4'b1001;
												assign node29415 = (inp[9]) ? node29423 : node29416;
													assign node29416 = (inp[4]) ? 4'b1001 : node29417;
														assign node29417 = (inp[12]) ? node29419 : 4'b1101;
															assign node29419 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node29423 = (inp[4]) ? node29427 : node29424;
														assign node29424 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node29427 = (inp[2]) ? 4'b1111 : node29428;
															assign node29428 = (inp[12]) ? node29430 : 4'b1111;
																assign node29430 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node29434 = (inp[3]) ? node29450 : node29435;
												assign node29435 = (inp[12]) ? node29441 : node29436;
													assign node29436 = (inp[4]) ? 4'b1001 : node29437;
														assign node29437 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node29441 = (inp[4]) ? node29447 : node29442;
														assign node29442 = (inp[10]) ? 4'b1111 : node29443;
															assign node29443 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node29447 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node29450 = (inp[9]) ? node29454 : node29451;
													assign node29451 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node29454 = (inp[4]) ? node29460 : node29455;
														assign node29455 = (inp[10]) ? node29457 : 4'b1011;
															assign node29457 = (inp[12]) ? 4'b1111 : 4'b1011;
														assign node29460 = (inp[10]) ? node29462 : 4'b1111;
															assign node29462 = (inp[2]) ? 4'b1011 : 4'b1111;
									assign node29465 = (inp[0]) ? node29537 : node29466;
										assign node29466 = (inp[5]) ? node29502 : node29467;
											assign node29467 = (inp[3]) ? node29487 : node29468;
												assign node29468 = (inp[9]) ? node29478 : node29469;
													assign node29469 = (inp[10]) ? node29473 : node29470;
														assign node29470 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node29473 = (inp[12]) ? node29475 : 4'b1001;
															assign node29475 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node29478 = (inp[4]) ? node29482 : node29479;
														assign node29479 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node29482 = (inp[12]) ? node29484 : 4'b1101;
															assign node29484 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node29487 = (inp[4]) ? node29497 : node29488;
													assign node29488 = (inp[9]) ? node29492 : node29489;
														assign node29489 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node29492 = (inp[12]) ? node29494 : 4'b1001;
															assign node29494 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node29497 = (inp[9]) ? node29499 : 4'b1001;
														assign node29499 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node29502 = (inp[3]) ? node29522 : node29503;
												assign node29503 = (inp[9]) ? node29513 : node29504;
													assign node29504 = (inp[4]) ? node29508 : node29505;
														assign node29505 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node29508 = (inp[12]) ? node29510 : 4'b1001;
															assign node29510 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node29513 = (inp[4]) ? node29517 : node29514;
														assign node29514 = (inp[12]) ? 4'b1111 : 4'b1001;
														assign node29517 = (inp[10]) ? node29519 : 4'b1111;
															assign node29519 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node29522 = (inp[2]) ? node29524 : 4'b1011;
													assign node29524 = (inp[10]) ? node29532 : node29525;
														assign node29525 = (inp[4]) ? node29529 : node29526;
															assign node29526 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node29529 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node29532 = (inp[4]) ? node29534 : 4'b1111;
															assign node29534 = (inp[9]) ? 4'b1111 : 4'b1011;
										assign node29537 = (inp[3]) ? node29577 : node29538;
											assign node29538 = (inp[5]) ? node29564 : node29539;
												assign node29539 = (inp[10]) ? node29549 : node29540;
													assign node29540 = (inp[2]) ? 4'b1011 : node29541;
														assign node29541 = (inp[4]) ? node29545 : node29542;
															assign node29542 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node29545 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node29549 = (inp[2]) ? node29551 : 4'b1111;
														assign node29551 = (inp[4]) ? node29559 : node29552;
															assign node29552 = (inp[12]) ? node29556 : node29553;
																assign node29553 = (inp[9]) ? 4'b1011 : 4'b1111;
																assign node29556 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node29559 = (inp[12]) ? 4'b1111 : node29560;
																assign node29560 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node29564 = (inp[12]) ? node29570 : node29565;
													assign node29565 = (inp[2]) ? 4'b1011 : node29566;
														assign node29566 = (inp[10]) ? 4'b1011 : 4'b1111;
													assign node29570 = (inp[9]) ? 4'b1101 : node29571;
														assign node29571 = (inp[2]) ? 4'b1011 : node29572;
															assign node29572 = (inp[10]) ? 4'b1101 : 4'b1011;
											assign node29577 = (inp[5]) ? node29593 : node29578;
												assign node29578 = (inp[4]) ? node29586 : node29579;
													assign node29579 = (inp[12]) ? node29583 : node29580;
														assign node29580 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node29583 = (inp[9]) ? 4'b1101 : 4'b1111;
													assign node29586 = (inp[9]) ? node29590 : node29587;
														assign node29587 = (inp[2]) ? 4'b1011 : 4'b1101;
														assign node29590 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node29593 = (inp[12]) ? node29599 : node29594;
													assign node29594 = (inp[9]) ? node29596 : 4'b1101;
														assign node29596 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node29599 = (inp[2]) ? node29601 : 4'b1001;
														assign node29601 = (inp[9]) ? node29603 : 4'b1001;
															assign node29603 = (inp[10]) ? node29607 : node29604;
																assign node29604 = (inp[4]) ? 4'b1101 : 4'b1001;
																assign node29607 = (inp[4]) ? 4'b1001 : 4'b1101;
								assign node29610 = (inp[2]) ? node29760 : node29611;
									assign node29611 = (inp[5]) ? node29687 : node29612;
										assign node29612 = (inp[15]) ? node29642 : node29613;
											assign node29613 = (inp[0]) ? node29635 : node29614;
												assign node29614 = (inp[12]) ? node29624 : node29615;
													assign node29615 = (inp[10]) ? 4'b0011 : node29616;
														assign node29616 = (inp[9]) ? node29620 : node29617;
															assign node29617 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node29620 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node29624 = (inp[3]) ? 4'b0101 : node29625;
														assign node29625 = (inp[10]) ? node29627 : 4'b0011;
															assign node29627 = (inp[9]) ? node29631 : node29628;
																assign node29628 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node29631 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node29635 = (inp[12]) ? 4'b0001 : node29636;
													assign node29636 = (inp[4]) ? 4'b0101 : node29637;
														assign node29637 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node29642 = (inp[0]) ? node29658 : node29643;
												assign node29643 = (inp[3]) ? node29645 : 4'b0001;
													assign node29645 = (inp[9]) ? node29653 : node29646;
														assign node29646 = (inp[12]) ? node29648 : 4'b0101;
															assign node29648 = (inp[4]) ? 4'b0001 : node29649;
																assign node29649 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node29653 = (inp[4]) ? 4'b0111 : node29654;
															assign node29654 = (inp[12]) ? 4'b0111 : 4'b0001;
												assign node29658 = (inp[3]) ? node29672 : node29659;
													assign node29659 = (inp[4]) ? node29667 : node29660;
														assign node29660 = (inp[10]) ? node29662 : 4'b0011;
															assign node29662 = (inp[12]) ? 4'b0111 : node29663;
																assign node29663 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node29667 = (inp[9]) ? node29669 : 4'b0011;
															assign node29669 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node29672 = (inp[9]) ? node29682 : node29673;
														assign node29673 = (inp[4]) ? node29677 : node29674;
															assign node29674 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node29677 = (inp[10]) ? node29679 : 4'b0011;
																assign node29679 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node29682 = (inp[12]) ? 4'b0101 : node29683;
															assign node29683 = (inp[4]) ? 4'b0101 : 4'b0011;
										assign node29687 = (inp[9]) ? node29721 : node29688;
											assign node29688 = (inp[4]) ? node29706 : node29689;
												assign node29689 = (inp[10]) ? node29697 : node29690;
													assign node29690 = (inp[15]) ? 4'b0101 : node29691;
														assign node29691 = (inp[0]) ? 4'b0101 : node29692;
															assign node29692 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node29697 = (inp[12]) ? node29699 : 4'b0101;
														assign node29699 = (inp[3]) ? 4'b0011 : node29700;
															assign node29700 = (inp[0]) ? node29702 : 4'b0001;
																assign node29702 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node29706 = (inp[12]) ? node29712 : node29707;
													assign node29707 = (inp[15]) ? node29709 : 4'b0001;
														assign node29709 = (inp[10]) ? 4'b0011 : 4'b0001;
													assign node29712 = (inp[15]) ? node29718 : node29713;
														assign node29713 = (inp[0]) ? 4'b0011 : node29714;
															assign node29714 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node29718 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node29721 = (inp[4]) ? node29749 : node29722;
												assign node29722 = (inp[12]) ? node29742 : node29723;
													assign node29723 = (inp[10]) ? node29737 : node29724;
														assign node29724 = (inp[15]) ? node29730 : node29725;
															assign node29725 = (inp[3]) ? node29727 : 4'b0011;
																assign node29727 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node29730 = (inp[0]) ? node29734 : node29731;
																assign node29731 = (inp[3]) ? 4'b0011 : 4'b0001;
																assign node29734 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node29737 = (inp[0]) ? 4'b0001 : node29738;
															assign node29738 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node29742 = (inp[10]) ? node29746 : node29743;
														assign node29743 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node29746 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node29749 = (inp[10]) ? node29757 : node29750;
													assign node29750 = (inp[3]) ? 4'b0111 : node29751;
														assign node29751 = (inp[0]) ? 4'b0101 : node29752;
															assign node29752 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node29757 = (inp[15]) ? 4'b0001 : 4'b0011;
									assign node29760 = (inp[9]) ? node29846 : node29761;
										assign node29761 = (inp[4]) ? node29811 : node29762;
											assign node29762 = (inp[10]) ? node29784 : node29763;
												assign node29763 = (inp[3]) ? node29781 : node29764;
													assign node29764 = (inp[12]) ? node29774 : node29765;
														assign node29765 = (inp[5]) ? node29767 : 4'b0111;
															assign node29767 = (inp[0]) ? node29771 : node29768;
																assign node29768 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node29771 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node29774 = (inp[5]) ? 4'b0111 : node29775;
															assign node29775 = (inp[0]) ? node29777 : 4'b0101;
																assign node29777 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node29781 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node29784 = (inp[12]) ? node29794 : node29785;
													assign node29785 = (inp[15]) ? node29791 : node29786;
														assign node29786 = (inp[5]) ? 4'b0101 : node29787;
															assign node29787 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node29791 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node29794 = (inp[5]) ? node29802 : node29795;
														assign node29795 = (inp[15]) ? node29799 : node29796;
															assign node29796 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node29799 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node29802 = (inp[3]) ? node29804 : 4'b0011;
															assign node29804 = (inp[0]) ? node29808 : node29805;
																assign node29805 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node29808 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node29811 = (inp[10]) ? node29831 : node29812;
												assign node29812 = (inp[15]) ? node29824 : node29813;
													assign node29813 = (inp[0]) ? node29819 : node29814;
														assign node29814 = (inp[3]) ? node29816 : 4'b0011;
															assign node29816 = (inp[5]) ? 4'b0001 : 4'b0011;
														assign node29819 = (inp[5]) ? node29821 : 4'b0001;
															assign node29821 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node29824 = (inp[0]) ? node29826 : 4'b0001;
														assign node29826 = (inp[3]) ? node29828 : 4'b0011;
															assign node29828 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node29831 = (inp[12]) ? node29837 : node29832;
													assign node29832 = (inp[15]) ? 4'b0001 : node29833;
														assign node29833 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node29837 = (inp[5]) ? 4'b0101 : node29838;
														assign node29838 = (inp[15]) ? 4'b0111 : node29839;
															assign node29839 = (inp[3]) ? 4'b0101 : node29840;
																assign node29840 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node29846 = (inp[4]) ? node29888 : node29847;
											assign node29847 = (inp[10]) ? node29865 : node29848;
												assign node29848 = (inp[0]) ? node29860 : node29849;
													assign node29849 = (inp[12]) ? node29855 : node29850;
														assign node29850 = (inp[15]) ? node29852 : 4'b0011;
															assign node29852 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node29855 = (inp[15]) ? 4'b0001 : node29856;
															assign node29856 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node29860 = (inp[15]) ? 4'b0011 : node29861;
														assign node29861 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node29865 = (inp[12]) ? node29875 : node29866;
													assign node29866 = (inp[5]) ? node29872 : node29867;
														assign node29867 = (inp[15]) ? node29869 : 4'b0001;
															assign node29869 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node29872 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node29875 = (inp[15]) ? node29879 : node29876;
														assign node29876 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node29879 = (inp[0]) ? node29885 : node29880;
															assign node29880 = (inp[5]) ? 4'b0111 : node29881;
																assign node29881 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node29885 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node29888 = (inp[12]) ? node29910 : node29889;
												assign node29889 = (inp[5]) ? node29903 : node29890;
													assign node29890 = (inp[15]) ? 4'b0111 : node29891;
														assign node29891 = (inp[10]) ? node29897 : node29892;
															assign node29892 = (inp[0]) ? 4'b0111 : node29893;
																assign node29893 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node29897 = (inp[0]) ? 4'b0101 : node29898;
																assign node29898 = (inp[3]) ? 4'b0101 : 4'b0111;
													assign node29903 = (inp[15]) ? node29907 : node29904;
														assign node29904 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node29907 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node29910 = (inp[10]) ? node29920 : node29911;
													assign node29911 = (inp[15]) ? 4'b0111 : node29912;
														assign node29912 = (inp[0]) ? 4'b0101 : node29913;
															assign node29913 = (inp[3]) ? 4'b0101 : node29914;
																assign node29914 = (inp[5]) ? 4'b0101 : 4'b0111;
													assign node29920 = (inp[3]) ? 4'b0001 : node29921;
														assign node29921 = (inp[5]) ? 4'b0001 : 4'b0011;
							assign node29925 = (inp[0]) ? node30121 : node29926;
								assign node29926 = (inp[15]) ? node30018 : node29927;
									assign node29927 = (inp[3]) ? node29963 : node29928;
										assign node29928 = (inp[4]) ? node29942 : node29929;
											assign node29929 = (inp[9]) ? node29935 : node29930;
												assign node29930 = (inp[12]) ? node29932 : 4'b0111;
													assign node29932 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node29935 = (inp[10]) ? node29937 : 4'b0011;
													assign node29937 = (inp[12]) ? node29939 : 4'b0011;
														assign node29939 = (inp[2]) ? 4'b0101 : 4'b0111;
											assign node29942 = (inp[5]) ? node29952 : node29943;
												assign node29943 = (inp[1]) ? node29945 : 4'b0111;
													assign node29945 = (inp[9]) ? node29947 : 4'b0011;
														assign node29947 = (inp[10]) ? node29949 : 4'b0111;
															assign node29949 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node29952 = (inp[9]) ? node29958 : node29953;
													assign node29953 = (inp[12]) ? node29955 : 4'b0011;
														assign node29955 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node29958 = (inp[10]) ? node29960 : 4'b0101;
														assign node29960 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node29963 = (inp[5]) ? node29987 : node29964;
											assign node29964 = (inp[9]) ? node29976 : node29965;
												assign node29965 = (inp[4]) ? node29971 : node29966;
													assign node29966 = (inp[12]) ? node29968 : 4'b0111;
														assign node29968 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node29971 = (inp[12]) ? node29973 : 4'b0011;
														assign node29973 = (inp[10]) ? 4'b0101 : 4'b0011;
												assign node29976 = (inp[4]) ? node29982 : node29977;
													assign node29977 = (inp[12]) ? node29979 : 4'b0011;
														assign node29979 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node29982 = (inp[12]) ? node29984 : 4'b0101;
														assign node29984 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node29987 = (inp[1]) ? node30007 : node29988;
												assign node29988 = (inp[10]) ? node29994 : node29989;
													assign node29989 = (inp[9]) ? node29991 : 4'b0001;
														assign node29991 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node29994 = (inp[9]) ? node30000 : node29995;
														assign node29995 = (inp[12]) ? 4'b0101 : node29996;
															assign node29996 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node30000 = (inp[4]) ? node30004 : node30001;
															assign node30001 = (inp[12]) ? 4'b0101 : 4'b0001;
															assign node30004 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node30007 = (inp[9]) ? node30013 : node30008;
													assign node30008 = (inp[12]) ? 4'b0001 : node30009;
														assign node30009 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node30013 = (inp[2]) ? 4'b0001 : node30014;
														assign node30014 = (inp[10]) ? 4'b0001 : 4'b0101;
									assign node30018 = (inp[3]) ? node30068 : node30019;
										assign node30019 = (inp[5]) ? node30051 : node30020;
											assign node30020 = (inp[9]) ? node30040 : node30021;
												assign node30021 = (inp[12]) ? node30025 : node30022;
													assign node30022 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node30025 = (inp[2]) ? node30035 : node30026;
														assign node30026 = (inp[1]) ? 4'b0101 : node30027;
															assign node30027 = (inp[10]) ? node30031 : node30028;
																assign node30028 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node30031 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node30035 = (inp[1]) ? node30037 : 4'b0001;
															assign node30037 = (inp[10]) ? 4'b0101 : 4'b0001;
												assign node30040 = (inp[4]) ? node30046 : node30041;
													assign node30041 = (inp[12]) ? node30043 : 4'b0001;
														assign node30043 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node30046 = (inp[12]) ? node30048 : 4'b0101;
														assign node30048 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node30051 = (inp[4]) ? node30059 : node30052;
												assign node30052 = (inp[9]) ? 4'b0001 : node30053;
													assign node30053 = (inp[10]) ? node30055 : 4'b0101;
														assign node30055 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node30059 = (inp[9]) ? node30065 : node30060;
													assign node30060 = (inp[12]) ? node30062 : 4'b0001;
														assign node30062 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node30065 = (inp[10]) ? 4'b0011 : 4'b0111;
										assign node30068 = (inp[5]) ? node30088 : node30069;
											assign node30069 = (inp[9]) ? node30081 : node30070;
												assign node30070 = (inp[4]) ? node30076 : node30071;
													assign node30071 = (inp[12]) ? node30073 : 4'b0101;
														assign node30073 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node30076 = (inp[12]) ? node30078 : 4'b0001;
														assign node30078 = (inp[1]) ? 4'b0111 : 4'b0001;
												assign node30081 = (inp[4]) ? 4'b0111 : node30082;
													assign node30082 = (inp[10]) ? node30084 : 4'b0001;
														assign node30084 = (inp[12]) ? 4'b0111 : 4'b0001;
											assign node30088 = (inp[1]) ? node30104 : node30089;
												assign node30089 = (inp[4]) ? node30095 : node30090;
													assign node30090 = (inp[9]) ? 4'b0011 : node30091;
														assign node30091 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node30095 = (inp[9]) ? node30099 : node30096;
														assign node30096 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node30099 = (inp[10]) ? node30101 : 4'b0111;
															assign node30101 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node30104 = (inp[9]) ? node30116 : node30105;
													assign node30105 = (inp[4]) ? node30111 : node30106;
														assign node30106 = (inp[12]) ? node30108 : 4'b0111;
															assign node30108 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node30111 = (inp[12]) ? node30113 : 4'b0011;
															assign node30113 = (inp[2]) ? 4'b0111 : 4'b0011;
													assign node30116 = (inp[4]) ? 4'b0111 : node30117;
														assign node30117 = (inp[10]) ? 4'b0111 : 4'b0011;
								assign node30121 = (inp[15]) ? node30237 : node30122;
									assign node30122 = (inp[3]) ? node30182 : node30123;
										assign node30123 = (inp[5]) ? node30165 : node30124;
											assign node30124 = (inp[1]) ? node30148 : node30125;
												assign node30125 = (inp[12]) ? node30135 : node30126;
													assign node30126 = (inp[10]) ? node30132 : node30127;
														assign node30127 = (inp[4]) ? 4'b0001 : node30128;
															assign node30128 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node30132 = (inp[2]) ? 4'b0001 : 4'b0101;
													assign node30135 = (inp[9]) ? node30141 : node30136;
														assign node30136 = (inp[10]) ? 4'b0001 : node30137;
															assign node30137 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node30141 = (inp[10]) ? node30145 : node30142;
															assign node30142 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node30145 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node30148 = (inp[9]) ? node30160 : node30149;
													assign node30149 = (inp[4]) ? node30155 : node30150;
														assign node30150 = (inp[10]) ? node30152 : 4'b0101;
															assign node30152 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node30155 = (inp[12]) ? node30157 : 4'b0001;
															assign node30157 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node30160 = (inp[12]) ? node30162 : 4'b0101;
														assign node30162 = (inp[10]) ? 4'b0101 : 4'b0001;
											assign node30165 = (inp[4]) ? node30173 : node30166;
												assign node30166 = (inp[9]) ? node30168 : 4'b0101;
													assign node30168 = (inp[10]) ? node30170 : 4'b0001;
														assign node30170 = (inp[12]) ? 4'b0111 : 4'b0001;
												assign node30173 = (inp[9]) ? node30177 : node30174;
													assign node30174 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node30177 = (inp[12]) ? node30179 : 4'b0111;
														assign node30179 = (inp[10]) ? 4'b0011 : 4'b0111;
										assign node30182 = (inp[5]) ? node30204 : node30183;
											assign node30183 = (inp[9]) ? node30193 : node30184;
												assign node30184 = (inp[4]) ? node30188 : node30185;
													assign node30185 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node30188 = (inp[12]) ? node30190 : 4'b0001;
														assign node30190 = (inp[10]) ? 4'b0111 : 4'b0001;
												assign node30193 = (inp[4]) ? node30199 : node30194;
													assign node30194 = (inp[10]) ? node30196 : 4'b0001;
														assign node30196 = (inp[12]) ? 4'b0111 : 4'b0001;
													assign node30199 = (inp[10]) ? node30201 : 4'b0111;
														assign node30201 = (inp[12]) ? 4'b0011 : 4'b0111;
											assign node30204 = (inp[12]) ? node30228 : node30205;
												assign node30205 = (inp[1]) ? node30221 : node30206;
													assign node30206 = (inp[10]) ? node30216 : node30207;
														assign node30207 = (inp[2]) ? node30213 : node30208;
															assign node30208 = (inp[9]) ? 4'b0011 : node30209;
																assign node30209 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node30213 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node30216 = (inp[4]) ? 4'b0111 : node30217;
															assign node30217 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node30221 = (inp[9]) ? node30225 : node30222;
														assign node30222 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node30225 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node30228 = (inp[2]) ? node30232 : node30229;
													assign node30229 = (inp[9]) ? 4'b0111 : 4'b0011;
													assign node30232 = (inp[9]) ? node30234 : 4'b0111;
														assign node30234 = (inp[10]) ? 4'b0111 : 4'b0011;
									assign node30237 = (inp[5]) ? node30283 : node30238;
										assign node30238 = (inp[3]) ? node30260 : node30239;
											assign node30239 = (inp[9]) ? node30249 : node30240;
												assign node30240 = (inp[10]) ? node30242 : 4'b0111;
													assign node30242 = (inp[12]) ? node30246 : node30243;
														assign node30243 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node30246 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node30249 = (inp[4]) ? node30255 : node30250;
													assign node30250 = (inp[10]) ? node30252 : 4'b0011;
														assign node30252 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node30255 = (inp[12]) ? node30257 : 4'b0111;
														assign node30257 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node30260 = (inp[9]) ? node30272 : node30261;
												assign node30261 = (inp[4]) ? node30267 : node30262;
													assign node30262 = (inp[12]) ? node30264 : 4'b0111;
														assign node30264 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node30267 = (inp[12]) ? node30269 : 4'b0011;
														assign node30269 = (inp[10]) ? 4'b0101 : 4'b0011;
												assign node30272 = (inp[4]) ? node30278 : node30273;
													assign node30273 = (inp[12]) ? node30275 : 4'b0011;
														assign node30275 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node30278 = (inp[12]) ? node30280 : 4'b0101;
														assign node30280 = (inp[10]) ? 4'b0001 : 4'b0101;
										assign node30283 = (inp[3]) ? node30301 : node30284;
											assign node30284 = (inp[4]) ? node30290 : node30285;
												assign node30285 = (inp[9]) ? 4'b0011 : node30286;
													assign node30286 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node30290 = (inp[9]) ? node30296 : node30291;
													assign node30291 = (inp[12]) ? node30293 : 4'b0011;
														assign node30293 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node30296 = (inp[12]) ? node30298 : 4'b0101;
														assign node30298 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node30301 = (inp[2]) ? node30325 : node30302;
												assign node30302 = (inp[9]) ? node30314 : node30303;
													assign node30303 = (inp[4]) ? node30309 : node30304;
														assign node30304 = (inp[12]) ? node30306 : 4'b0101;
															assign node30306 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node30309 = (inp[12]) ? node30311 : 4'b0001;
															assign node30311 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node30314 = (inp[4]) ? node30320 : node30315;
														assign node30315 = (inp[12]) ? node30317 : 4'b0001;
															assign node30317 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node30320 = (inp[10]) ? node30322 : 4'b0101;
															assign node30322 = (inp[12]) ? 4'b0001 : 4'b0101;
												assign node30325 = (inp[12]) ? node30341 : node30326;
													assign node30326 = (inp[1]) ? node30332 : node30327;
														assign node30327 = (inp[4]) ? 4'b0101 : node30328;
															assign node30328 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node30332 = (inp[10]) ? node30334 : 4'b0001;
															assign node30334 = (inp[9]) ? node30338 : node30335;
																assign node30335 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node30338 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node30341 = (inp[9]) ? node30347 : node30342;
														assign node30342 = (inp[1]) ? 4'b0001 : node30343;
															assign node30343 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node30347 = (inp[1]) ? node30349 : 4'b0001;
															assign node30349 = (inp[10]) ? node30353 : node30350;
																assign node30350 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node30353 = (inp[4]) ? 4'b0001 : 4'b0101;
						assign node30356 = (inp[1]) ? node31018 : node30357;
							assign node30357 = (inp[13]) ? node30729 : node30358;
								assign node30358 = (inp[12]) ? node30526 : node30359;
									assign node30359 = (inp[5]) ? node30465 : node30360;
										assign node30360 = (inp[2]) ? node30408 : node30361;
											assign node30361 = (inp[9]) ? node30381 : node30362;
												assign node30362 = (inp[4]) ? node30368 : node30363;
													assign node30363 = (inp[15]) ? node30365 : 4'b0101;
														assign node30365 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node30368 = (inp[3]) ? node30370 : 4'b0001;
														assign node30370 = (inp[10]) ? node30376 : node30371;
															assign node30371 = (inp[0]) ? 4'b0001 : node30372;
																assign node30372 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node30376 = (inp[0]) ? node30378 : 4'b0001;
																assign node30378 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node30381 = (inp[4]) ? node30395 : node30382;
													assign node30382 = (inp[3]) ? node30388 : node30383;
														assign node30383 = (inp[15]) ? node30385 : 4'b0011;
															assign node30385 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node30388 = (inp[15]) ? node30392 : node30389;
															assign node30389 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node30392 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node30395 = (inp[3]) ? node30403 : node30396;
														assign node30396 = (inp[10]) ? node30398 : 4'b0111;
															assign node30398 = (inp[0]) ? node30400 : 4'b0101;
																assign node30400 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node30403 = (inp[10]) ? 4'b0111 : node30404;
															assign node30404 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node30408 = (inp[3]) ? node30444 : node30409;
												assign node30409 = (inp[9]) ? node30423 : node30410;
													assign node30410 = (inp[4]) ? node30416 : node30411;
														assign node30411 = (inp[0]) ? node30413 : 4'b0111;
															assign node30413 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node30416 = (inp[15]) ? node30420 : node30417;
															assign node30417 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node30420 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node30423 = (inp[4]) ? node30429 : node30424;
														assign node30424 = (inp[15]) ? node30426 : 4'b0001;
															assign node30426 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node30429 = (inp[10]) ? node30437 : node30430;
															assign node30430 = (inp[15]) ? node30434 : node30431;
																assign node30431 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node30434 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node30437 = (inp[0]) ? node30441 : node30438;
																assign node30438 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node30441 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node30444 = (inp[4]) ? node30458 : node30445;
													assign node30445 = (inp[9]) ? node30451 : node30446;
														assign node30446 = (inp[15]) ? node30448 : 4'b0111;
															assign node30448 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node30451 = (inp[15]) ? node30455 : node30452;
															assign node30452 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node30455 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node30458 = (inp[9]) ? node30460 : 4'b0011;
														assign node30460 = (inp[0]) ? node30462 : 4'b0111;
															assign node30462 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node30465 = (inp[0]) ? node30499 : node30466;
											assign node30466 = (inp[15]) ? node30486 : node30467;
												assign node30467 = (inp[3]) ? node30475 : node30468;
													assign node30468 = (inp[10]) ? 4'b0011 : node30469;
														assign node30469 = (inp[9]) ? 4'b0101 : node30470;
															assign node30470 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node30475 = (inp[10]) ? node30481 : node30476;
														assign node30476 = (inp[4]) ? node30478 : 4'b0001;
															assign node30478 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node30481 = (inp[4]) ? node30483 : 4'b0101;
															assign node30483 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node30486 = (inp[3]) ? node30492 : node30487;
													assign node30487 = (inp[9]) ? 4'b0001 : node30488;
														assign node30488 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node30492 = (inp[4]) ? node30496 : node30493;
														assign node30493 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node30496 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node30499 = (inp[15]) ? node30513 : node30500;
												assign node30500 = (inp[3]) ? node30508 : node30501;
													assign node30501 = (inp[4]) ? node30505 : node30502;
														assign node30502 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node30505 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node30508 = (inp[4]) ? node30510 : 4'b0111;
														assign node30510 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node30513 = (inp[3]) ? node30519 : node30514;
													assign node30514 = (inp[9]) ? 4'b0101 : node30515;
														assign node30515 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node30519 = (inp[9]) ? node30523 : node30520;
														assign node30520 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node30523 = (inp[4]) ? 4'b0101 : 4'b0001;
									assign node30526 = (inp[9]) ? node30608 : node30527;
										assign node30527 = (inp[3]) ? node30567 : node30528;
											assign node30528 = (inp[4]) ? node30544 : node30529;
												assign node30529 = (inp[10]) ? node30537 : node30530;
													assign node30530 = (inp[5]) ? node30532 : 4'b0101;
														assign node30532 = (inp[15]) ? 4'b0111 : node30533;
															assign node30533 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node30537 = (inp[15]) ? node30541 : node30538;
														assign node30538 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node30541 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node30544 = (inp[10]) ? node30552 : node30545;
													assign node30545 = (inp[2]) ? 4'b0011 : node30546;
														assign node30546 = (inp[0]) ? node30548 : 4'b0011;
															assign node30548 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node30552 = (inp[5]) ? node30560 : node30553;
														assign node30553 = (inp[0]) ? node30557 : node30554;
															assign node30554 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node30557 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node30560 = (inp[15]) ? node30564 : node30561;
															assign node30561 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node30564 = (inp[0]) ? 4'b0101 : 4'b0111;
											assign node30567 = (inp[5]) ? node30589 : node30568;
												assign node30568 = (inp[10]) ? node30576 : node30569;
													assign node30569 = (inp[15]) ? node30573 : node30570;
														assign node30570 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node30573 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node30576 = (inp[4]) ? node30582 : node30577;
														assign node30577 = (inp[15]) ? 4'b0011 : node30578;
															assign node30578 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node30582 = (inp[2]) ? node30586 : node30583;
															assign node30583 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node30586 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node30589 = (inp[15]) ? node30601 : node30590;
													assign node30590 = (inp[0]) ? node30598 : node30591;
														assign node30591 = (inp[4]) ? node30595 : node30592;
															assign node30592 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node30595 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node30598 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node30601 = (inp[0]) ? node30603 : 4'b0111;
														assign node30603 = (inp[2]) ? 4'b0101 : node30604;
															assign node30604 = (inp[10]) ? 4'b0101 : 4'b0001;
										assign node30608 = (inp[2]) ? node30660 : node30609;
											assign node30609 = (inp[5]) ? node30647 : node30610;
												assign node30610 = (inp[0]) ? node30630 : node30611;
													assign node30611 = (inp[3]) ? node30621 : node30612;
														assign node30612 = (inp[15]) ? node30614 : 4'b0011;
															assign node30614 = (inp[10]) ? node30618 : node30615;
																assign node30615 = (inp[4]) ? 4'b0101 : 4'b0001;
																assign node30618 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node30621 = (inp[15]) ? node30627 : node30622;
															assign node30622 = (inp[4]) ? node30624 : 4'b0101;
																assign node30624 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node30627 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node30630 = (inp[15]) ? node30640 : node30631;
														assign node30631 = (inp[3]) ? node30635 : node30632;
															assign node30632 = (inp[10]) ? 4'b0001 : 4'b0101;
															assign node30635 = (inp[4]) ? node30637 : 4'b0111;
																assign node30637 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node30640 = (inp[10]) ? node30642 : 4'b0011;
															assign node30642 = (inp[3]) ? node30644 : 4'b0011;
																assign node30644 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node30647 = (inp[0]) ? node30653 : node30648;
													assign node30648 = (inp[15]) ? node30650 : 4'b0001;
														assign node30650 = (inp[3]) ? 4'b0011 : 4'b0111;
													assign node30653 = (inp[15]) ? 4'b0101 : node30654;
														assign node30654 = (inp[3]) ? node30656 : 4'b0111;
															assign node30656 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node30660 = (inp[5]) ? node30698 : node30661;
												assign node30661 = (inp[0]) ? node30685 : node30662;
													assign node30662 = (inp[4]) ? node30672 : node30663;
														assign node30663 = (inp[10]) ? node30667 : node30664;
															assign node30664 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node30667 = (inp[15]) ? node30669 : 4'b0101;
																assign node30669 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node30672 = (inp[10]) ? node30680 : node30673;
															assign node30673 = (inp[3]) ? node30677 : node30674;
																assign node30674 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node30677 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node30680 = (inp[15]) ? 4'b0011 : node30681;
																assign node30681 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node30685 = (inp[4]) ? node30693 : node30686;
														assign node30686 = (inp[15]) ? node30690 : node30687;
															assign node30687 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node30690 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node30693 = (inp[10]) ? 4'b0001 : node30694;
															assign node30694 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node30698 = (inp[3]) ? node30712 : node30699;
													assign node30699 = (inp[0]) ? node30705 : node30700;
														assign node30700 = (inp[4]) ? 4'b0111 : node30701;
															assign node30701 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node30705 = (inp[15]) ? node30707 : 4'b0001;
															assign node30707 = (inp[4]) ? node30709 : 4'b0101;
																assign node30709 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node30712 = (inp[4]) ? node30722 : node30713;
														assign node30713 = (inp[10]) ? node30719 : node30714;
															assign node30714 = (inp[15]) ? node30716 : 4'b0011;
																assign node30716 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node30719 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node30722 = (inp[10]) ? node30724 : 4'b0101;
															assign node30724 = (inp[15]) ? 4'b0001 : node30725;
																assign node30725 = (inp[0]) ? 4'b0011 : 4'b0001;
								assign node30729 = (inp[3]) ? node30853 : node30730;
									assign node30730 = (inp[0]) ? node30778 : node30731;
										assign node30731 = (inp[15]) ? node30759 : node30732;
											assign node30732 = (inp[5]) ? node30746 : node30733;
												assign node30733 = (inp[2]) ? node30739 : node30734;
													assign node30734 = (inp[4]) ? 4'b1011 : node30735;
														assign node30735 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node30739 = (inp[12]) ? node30741 : 4'b1011;
														assign node30741 = (inp[4]) ? 4'b1111 : node30742;
															assign node30742 = (inp[9]) ? 4'b1111 : 4'b1011;
												assign node30746 = (inp[9]) ? node30754 : node30747;
													assign node30747 = (inp[10]) ? 4'b1011 : node30748;
														assign node30748 = (inp[12]) ? 4'b1101 : node30749;
															assign node30749 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node30754 = (inp[4]) ? 4'b1001 : node30755;
														assign node30755 = (inp[10]) ? 4'b1101 : 4'b1011;
											assign node30759 = (inp[4]) ? node30767 : node30760;
												assign node30760 = (inp[10]) ? 4'b1001 : node30761;
													assign node30761 = (inp[2]) ? 4'b1001 : node30762;
														assign node30762 = (inp[12]) ? 4'b1001 : 4'b1101;
												assign node30767 = (inp[5]) ? node30769 : 4'b1001;
													assign node30769 = (inp[9]) ? node30773 : node30770;
														assign node30770 = (inp[10]) ? 4'b1111 : 4'b1001;
														assign node30773 = (inp[10]) ? 4'b1011 : node30774;
															assign node30774 = (inp[2]) ? 4'b1111 : 4'b1011;
										assign node30778 = (inp[15]) ? node30822 : node30779;
											assign node30779 = (inp[5]) ? node30803 : node30780;
												assign node30780 = (inp[12]) ? node30796 : node30781;
													assign node30781 = (inp[9]) ? node30791 : node30782;
														assign node30782 = (inp[2]) ? 4'b1001 : node30783;
															assign node30783 = (inp[4]) ? node30787 : node30784;
																assign node30784 = (inp[10]) ? 4'b1001 : 4'b1101;
																assign node30787 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node30791 = (inp[10]) ? 4'b1101 : node30792;
															assign node30792 = (inp[4]) ? 4'b1101 : 4'b1001;
													assign node30796 = (inp[9]) ? node30800 : node30797;
														assign node30797 = (inp[4]) ? 4'b1101 : 4'b1001;
														assign node30800 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node30803 = (inp[4]) ? node30815 : node30804;
													assign node30804 = (inp[12]) ? node30812 : node30805;
														assign node30805 = (inp[2]) ? 4'b1001 : node30806;
															assign node30806 = (inp[10]) ? 4'b1001 : node30807;
																assign node30807 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node30812 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node30815 = (inp[9]) ? 4'b1011 : node30816;
														assign node30816 = (inp[12]) ? 4'b1111 : node30817;
															assign node30817 = (inp[10]) ? 4'b1111 : 4'b1001;
											assign node30822 = (inp[5]) ? node30842 : node30823;
												assign node30823 = (inp[4]) ? node30837 : node30824;
													assign node30824 = (inp[2]) ? node30830 : node30825;
														assign node30825 = (inp[9]) ? node30827 : 4'b1011;
															assign node30827 = (inp[10]) ? 4'b1111 : 4'b1011;
														assign node30830 = (inp[10]) ? 4'b1011 : node30831;
															assign node30831 = (inp[9]) ? node30833 : 4'b1111;
																assign node30833 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node30837 = (inp[10]) ? node30839 : 4'b1111;
														assign node30839 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node30842 = (inp[4]) ? node30848 : node30843;
													assign node30843 = (inp[2]) ? node30845 : 4'b1011;
														assign node30845 = (inp[9]) ? 4'b1101 : 4'b1011;
													assign node30848 = (inp[10]) ? node30850 : 4'b1101;
														assign node30850 = (inp[9]) ? 4'b1001 : 4'b1101;
									assign node30853 = (inp[4]) ? node30933 : node30854;
										assign node30854 = (inp[9]) ? node30900 : node30855;
											assign node30855 = (inp[12]) ? node30875 : node30856;
												assign node30856 = (inp[10]) ? node30866 : node30857;
													assign node30857 = (inp[15]) ? node30859 : 4'b1101;
														assign node30859 = (inp[0]) ? node30863 : node30860;
															assign node30860 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node30863 = (inp[5]) ? 4'b1101 : 4'b1111;
													assign node30866 = (inp[5]) ? node30868 : 4'b1001;
														assign node30868 = (inp[2]) ? node30870 : 4'b1011;
															assign node30870 = (inp[0]) ? node30872 : 4'b1001;
																assign node30872 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node30875 = (inp[10]) ? node30893 : node30876;
													assign node30876 = (inp[2]) ? node30878 : 4'b1001;
														assign node30878 = (inp[0]) ? node30886 : node30879;
															assign node30879 = (inp[15]) ? node30883 : node30880;
																assign node30880 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node30883 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node30886 = (inp[15]) ? node30890 : node30887;
																assign node30887 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node30890 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node30893 = (inp[5]) ? node30895 : 4'b1001;
														assign node30895 = (inp[15]) ? node30897 : 4'b1001;
															assign node30897 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node30900 = (inp[10]) ? node30926 : node30901;
												assign node30901 = (inp[12]) ? node30913 : node30902;
													assign node30902 = (inp[15]) ? node30904 : 4'b1001;
														assign node30904 = (inp[2]) ? node30908 : node30905;
															assign node30905 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node30908 = (inp[0]) ? 4'b1001 : node30909;
																assign node30909 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node30913 = (inp[2]) ? node30919 : node30914;
														assign node30914 = (inp[15]) ? 4'b1101 : node30915;
															assign node30915 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node30919 = (inp[0]) ? node30923 : node30920;
															assign node30920 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node30923 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node30926 = (inp[0]) ? node30930 : node30927;
													assign node30927 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node30930 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node30933 = (inp[9]) ? node30973 : node30934;
											assign node30934 = (inp[12]) ? node30954 : node30935;
												assign node30935 = (inp[10]) ? node30947 : node30936;
													assign node30936 = (inp[15]) ? node30942 : node30937;
														assign node30937 = (inp[0]) ? 4'b1001 : node30938;
															assign node30938 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node30942 = (inp[0]) ? 4'b1011 : node30943;
															assign node30943 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node30947 = (inp[5]) ? node30949 : 4'b1111;
														assign node30949 = (inp[0]) ? 4'b1101 : node30950;
															assign node30950 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node30954 = (inp[2]) ? node30960 : node30955;
													assign node30955 = (inp[5]) ? node30957 : 4'b1111;
														assign node30957 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node30960 = (inp[5]) ? node30966 : node30961;
														assign node30961 = (inp[10]) ? node30963 : 4'b1101;
															assign node30963 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node30966 = (inp[0]) ? node30970 : node30967;
															assign node30967 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node30970 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node30973 = (inp[10]) ? node30995 : node30974;
												assign node30974 = (inp[12]) ? node30982 : node30975;
													assign node30975 = (inp[2]) ? node30977 : 4'b1101;
														assign node30977 = (inp[15]) ? 4'b1111 : node30978;
															assign node30978 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node30982 = (inp[5]) ? node30990 : node30983;
														assign node30983 = (inp[2]) ? node30985 : 4'b1001;
															assign node30985 = (inp[0]) ? 4'b1011 : node30986;
																assign node30986 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node30990 = (inp[0]) ? 4'b1001 : node30991;
															assign node30991 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node30995 = (inp[12]) ? node31003 : node30996;
													assign node30996 = (inp[15]) ? node31000 : node30997;
														assign node30997 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node31000 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node31003 = (inp[2]) ? node31011 : node31004;
														assign node31004 = (inp[0]) ? node31008 : node31005;
															assign node31005 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node31008 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node31011 = (inp[15]) ? node31015 : node31012;
															assign node31012 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node31015 = (inp[0]) ? 4'b1001 : 4'b1011;
							assign node31018 = (inp[0]) ? node31202 : node31019;
								assign node31019 = (inp[15]) ? node31109 : node31020;
									assign node31020 = (inp[5]) ? node31064 : node31021;
										assign node31021 = (inp[3]) ? node31045 : node31022;
											assign node31022 = (inp[4]) ? node31034 : node31023;
												assign node31023 = (inp[2]) ? 4'b1011 : node31024;
													assign node31024 = (inp[9]) ? node31030 : node31025;
														assign node31025 = (inp[10]) ? 4'b1011 : node31026;
															assign node31026 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node31030 = (inp[10]) ? 4'b1111 : 4'b1011;
												assign node31034 = (inp[9]) ? node31040 : node31035;
													assign node31035 = (inp[12]) ? 4'b1111 : node31036;
														assign node31036 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node31040 = (inp[10]) ? 4'b1011 : node31041;
														assign node31041 = (inp[12]) ? 4'b1011 : 4'b1111;
											assign node31045 = (inp[9]) ? node31057 : node31046;
												assign node31046 = (inp[4]) ? node31052 : node31047;
													assign node31047 = (inp[10]) ? 4'b1011 : node31048;
														assign node31048 = (inp[12]) ? 4'b1011 : 4'b1111;
													assign node31052 = (inp[10]) ? 4'b1101 : node31053;
														assign node31053 = (inp[12]) ? 4'b1101 : 4'b1011;
												assign node31057 = (inp[4]) ? node31059 : 4'b1101;
													assign node31059 = (inp[10]) ? 4'b1001 : node31060;
														assign node31060 = (inp[12]) ? 4'b1001 : 4'b1101;
										assign node31064 = (inp[3]) ? node31086 : node31065;
											assign node31065 = (inp[9]) ? node31077 : node31066;
												assign node31066 = (inp[4]) ? node31072 : node31067;
													assign node31067 = (inp[12]) ? 4'b1011 : node31068;
														assign node31068 = (inp[2]) ? 4'b1011 : 4'b1111;
													assign node31072 = (inp[2]) ? 4'b1101 : node31073;
														assign node31073 = (inp[13]) ? 4'b1101 : 4'b1011;
												assign node31077 = (inp[4]) ? node31083 : node31078;
													assign node31078 = (inp[10]) ? 4'b1101 : node31079;
														assign node31079 = (inp[12]) ? 4'b1101 : 4'b1011;
													assign node31083 = (inp[10]) ? 4'b1001 : 4'b1101;
											assign node31086 = (inp[9]) ? node31098 : node31087;
												assign node31087 = (inp[4]) ? node31093 : node31088;
													assign node31088 = (inp[10]) ? 4'b1001 : node31089;
														assign node31089 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node31093 = (inp[10]) ? 4'b1101 : node31094;
														assign node31094 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node31098 = (inp[4]) ? node31104 : node31099;
													assign node31099 = (inp[10]) ? 4'b1101 : node31100;
														assign node31100 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node31104 = (inp[13]) ? node31106 : 4'b1001;
														assign node31106 = (inp[2]) ? 4'b1101 : 4'b1001;
									assign node31109 = (inp[5]) ? node31155 : node31110;
										assign node31110 = (inp[3]) ? node31132 : node31111;
											assign node31111 = (inp[9]) ? node31123 : node31112;
												assign node31112 = (inp[4]) ? node31118 : node31113;
													assign node31113 = (inp[12]) ? 4'b1001 : node31114;
														assign node31114 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node31118 = (inp[10]) ? 4'b1101 : node31119;
														assign node31119 = (inp[12]) ? 4'b1101 : 4'b1001;
												assign node31123 = (inp[4]) ? node31129 : node31124;
													assign node31124 = (inp[12]) ? 4'b1101 : node31125;
														assign node31125 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node31129 = (inp[10]) ? 4'b1001 : 4'b1101;
											assign node31132 = (inp[4]) ? node31144 : node31133;
												assign node31133 = (inp[9]) ? node31139 : node31134;
													assign node31134 = (inp[10]) ? 4'b1001 : node31135;
														assign node31135 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node31139 = (inp[10]) ? 4'b1111 : node31140;
														assign node31140 = (inp[13]) ? 4'b1001 : 4'b1111;
												assign node31144 = (inp[9]) ? node31150 : node31145;
													assign node31145 = (inp[12]) ? 4'b1111 : node31146;
														assign node31146 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node31150 = (inp[12]) ? 4'b1011 : node31151;
														assign node31151 = (inp[2]) ? 4'b1011 : 4'b1111;
										assign node31155 = (inp[3]) ? node31175 : node31156;
											assign node31156 = (inp[4]) ? node31168 : node31157;
												assign node31157 = (inp[9]) ? node31163 : node31158;
													assign node31158 = (inp[12]) ? 4'b1001 : node31159;
														assign node31159 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node31163 = (inp[10]) ? 4'b1111 : node31164;
														assign node31164 = (inp[12]) ? 4'b1111 : 4'b1001;
												assign node31168 = (inp[9]) ? 4'b1011 : node31169;
													assign node31169 = (inp[10]) ? 4'b1111 : node31170;
														assign node31170 = (inp[13]) ? 4'b1001 : 4'b1111;
											assign node31175 = (inp[2]) ? node31189 : node31176;
												assign node31176 = (inp[4]) ? node31184 : node31177;
													assign node31177 = (inp[9]) ? node31179 : 4'b1011;
														assign node31179 = (inp[12]) ? 4'b1111 : node31180;
															assign node31180 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node31184 = (inp[10]) ? node31186 : 4'b1111;
														assign node31186 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node31189 = (inp[9]) ? node31195 : node31190;
													assign node31190 = (inp[4]) ? node31192 : 4'b1011;
														assign node31192 = (inp[12]) ? 4'b1111 : 4'b1011;
													assign node31195 = (inp[4]) ? 4'b1011 : node31196;
														assign node31196 = (inp[10]) ? 4'b1111 : node31197;
															assign node31197 = (inp[12]) ? 4'b1111 : 4'b1011;
								assign node31202 = (inp[4]) ? node31272 : node31203;
									assign node31203 = (inp[9]) ? node31237 : node31204;
										assign node31204 = (inp[15]) ? node31224 : node31205;
											assign node31205 = (inp[3]) ? node31213 : node31206;
												assign node31206 = (inp[5]) ? 4'b1001 : node31207;
													assign node31207 = (inp[2]) ? node31209 : 4'b1001;
														assign node31209 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node31213 = (inp[5]) ? node31219 : node31214;
													assign node31214 = (inp[2]) ? node31216 : 4'b1001;
														assign node31216 = (inp[13]) ? 4'b1101 : 4'b1001;
													assign node31219 = (inp[2]) ? 4'b1011 : node31220;
														assign node31220 = (inp[13]) ? 4'b1111 : 4'b1011;
											assign node31224 = (inp[10]) ? node31232 : node31225;
												assign node31225 = (inp[12]) ? 4'b1011 : node31226;
													assign node31226 = (inp[3]) ? node31228 : 4'b1111;
														assign node31228 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node31232 = (inp[5]) ? node31234 : 4'b1011;
													assign node31234 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node31237 = (inp[10]) ? node31261 : node31238;
											assign node31238 = (inp[12]) ? node31250 : node31239;
												assign node31239 = (inp[15]) ? node31245 : node31240;
													assign node31240 = (inp[3]) ? node31242 : 4'b1001;
														assign node31242 = (inp[13]) ? 4'b1001 : 4'b1011;
													assign node31245 = (inp[5]) ? node31247 : 4'b1011;
														assign node31247 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node31250 = (inp[15]) ? node31256 : node31251;
													assign node31251 = (inp[3]) ? 4'b1111 : node31252;
														assign node31252 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node31256 = (inp[5]) ? 4'b1101 : node31257;
														assign node31257 = (inp[2]) ? 4'b1101 : 4'b1111;
											assign node31261 = (inp[15]) ? node31267 : node31262;
												assign node31262 = (inp[5]) ? 4'b1111 : node31263;
													assign node31263 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node31267 = (inp[3]) ? 4'b1101 : node31268;
													assign node31268 = (inp[5]) ? 4'b1101 : 4'b1111;
									assign node31272 = (inp[9]) ? node31320 : node31273;
										assign node31273 = (inp[10]) ? node31309 : node31274;
											assign node31274 = (inp[12]) ? node31286 : node31275;
												assign node31275 = (inp[15]) ? node31281 : node31276;
													assign node31276 = (inp[13]) ? 4'b1001 : node31277;
														assign node31277 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node31281 = (inp[3]) ? node31283 : 4'b1011;
														assign node31283 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node31286 = (inp[5]) ? 4'b1111 : node31287;
													assign node31287 = (inp[2]) ? node31293 : node31288;
														assign node31288 = (inp[13]) ? node31290 : 4'b1101;
															assign node31290 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node31293 = (inp[13]) ? node31301 : node31294;
															assign node31294 = (inp[3]) ? node31298 : node31295;
																assign node31295 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node31298 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node31301 = (inp[3]) ? node31305 : node31302;
																assign node31302 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node31305 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node31309 = (inp[15]) ? node31315 : node31310;
												assign node31310 = (inp[3]) ? 4'b1111 : node31311;
													assign node31311 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node31315 = (inp[12]) ? node31317 : 4'b1101;
													assign node31317 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node31320 = (inp[15]) ? node31338 : node31321;
											assign node31321 = (inp[5]) ? node31333 : node31322;
												assign node31322 = (inp[3]) ? node31328 : node31323;
													assign node31323 = (inp[12]) ? 4'b1001 : node31324;
														assign node31324 = (inp[10]) ? 4'b1001 : 4'b1101;
													assign node31328 = (inp[10]) ? 4'b1011 : node31329;
														assign node31329 = (inp[12]) ? 4'b1011 : 4'b1111;
												assign node31333 = (inp[12]) ? 4'b1011 : node31334;
													assign node31334 = (inp[10]) ? 4'b1011 : 4'b1111;
											assign node31338 = (inp[5]) ? node31346 : node31339;
												assign node31339 = (inp[3]) ? node31341 : 4'b1011;
													assign node31341 = (inp[10]) ? 4'b1001 : node31342;
														assign node31342 = (inp[2]) ? 4'b1001 : 4'b1101;
												assign node31346 = (inp[10]) ? 4'b1001 : node31347;
													assign node31347 = (inp[12]) ? 4'b1001 : 4'b1101;
					assign node31351 = (inp[6]) ? node32467 : node31352;
						assign node31352 = (inp[13]) ? node31930 : node31353;
							assign node31353 = (inp[1]) ? node31653 : node31354;
								assign node31354 = (inp[3]) ? node31500 : node31355;
									assign node31355 = (inp[15]) ? node31431 : node31356;
										assign node31356 = (inp[0]) ? node31398 : node31357;
											assign node31357 = (inp[5]) ? node31377 : node31358;
												assign node31358 = (inp[12]) ? node31366 : node31359;
													assign node31359 = (inp[9]) ? node31363 : node31360;
														assign node31360 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node31363 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node31366 = (inp[4]) ? node31372 : node31367;
														assign node31367 = (inp[9]) ? node31369 : 4'b0111;
															assign node31369 = (inp[10]) ? 4'b0111 : 4'b0011;
														assign node31372 = (inp[2]) ? 4'b0011 : node31373;
															assign node31373 = (inp[9]) ? 4'b0111 : 4'b0011;
												assign node31377 = (inp[9]) ? node31387 : node31378;
													assign node31378 = (inp[4]) ? node31384 : node31379;
														assign node31379 = (inp[12]) ? node31381 : 4'b0111;
															assign node31381 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node31384 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node31387 = (inp[4]) ? node31393 : node31388;
														assign node31388 = (inp[10]) ? node31390 : 4'b0011;
															assign node31390 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node31393 = (inp[10]) ? node31395 : 4'b0101;
															assign node31395 = (inp[2]) ? 4'b0101 : 4'b0001;
											assign node31398 = (inp[5]) ? node31416 : node31399;
												assign node31399 = (inp[9]) ? node31409 : node31400;
													assign node31400 = (inp[10]) ? node31402 : 4'b0101;
														assign node31402 = (inp[12]) ? node31406 : node31403;
															assign node31403 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node31406 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node31409 = (inp[4]) ? 4'b0101 : node31410;
														assign node31410 = (inp[10]) ? node31412 : 4'b0001;
															assign node31412 = (inp[2]) ? 4'b0101 : 4'b0001;
												assign node31416 = (inp[12]) ? node31424 : node31417;
													assign node31417 = (inp[9]) ? node31421 : node31418;
														assign node31418 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node31421 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node31424 = (inp[2]) ? 4'b0111 : node31425;
														assign node31425 = (inp[10]) ? node31427 : 4'b0001;
															assign node31427 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node31431 = (inp[0]) ? node31465 : node31432;
											assign node31432 = (inp[5]) ? node31450 : node31433;
												assign node31433 = (inp[9]) ? node31443 : node31434;
													assign node31434 = (inp[4]) ? node31438 : node31435;
														assign node31435 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node31438 = (inp[12]) ? node31440 : 4'b0001;
															assign node31440 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node31443 = (inp[4]) ? 4'b0101 : node31444;
														assign node31444 = (inp[10]) ? node31446 : 4'b0001;
															assign node31446 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node31450 = (inp[10]) ? 4'b0001 : node31451;
													assign node31451 = (inp[12]) ? node31459 : node31452;
														assign node31452 = (inp[4]) ? node31456 : node31453;
															assign node31453 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node31456 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node31459 = (inp[9]) ? 4'b0001 : node31460;
															assign node31460 = (inp[2]) ? 4'b0101 : 4'b0001;
											assign node31465 = (inp[5]) ? node31481 : node31466;
												assign node31466 = (inp[9]) ? node31476 : node31467;
													assign node31467 = (inp[4]) ? node31471 : node31468;
														assign node31468 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node31471 = (inp[12]) ? node31473 : 4'b0011;
															assign node31473 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node31476 = (inp[4]) ? 4'b0111 : node31477;
														assign node31477 = (inp[10]) ? 4'b0111 : 4'b0011;
												assign node31481 = (inp[9]) ? node31491 : node31482;
													assign node31482 = (inp[2]) ? node31484 : 4'b0011;
														assign node31484 = (inp[4]) ? node31488 : node31485;
															assign node31485 = (inp[12]) ? 4'b0011 : 4'b0111;
															assign node31488 = (inp[12]) ? 4'b0101 : 4'b0011;
													assign node31491 = (inp[10]) ? node31495 : node31492;
														assign node31492 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node31495 = (inp[4]) ? node31497 : 4'b0101;
															assign node31497 = (inp[12]) ? 4'b0001 : 4'b0101;
									assign node31500 = (inp[0]) ? node31578 : node31501;
										assign node31501 = (inp[15]) ? node31537 : node31502;
											assign node31502 = (inp[5]) ? node31520 : node31503;
												assign node31503 = (inp[4]) ? node31511 : node31504;
													assign node31504 = (inp[9]) ? 4'b0011 : node31505;
														assign node31505 = (inp[10]) ? node31507 : 4'b0111;
															assign node31507 = (inp[12]) ? 4'b0011 : 4'b0111;
													assign node31511 = (inp[9]) ? node31517 : node31512;
														assign node31512 = (inp[10]) ? node31514 : 4'b0011;
															assign node31514 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node31517 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node31520 = (inp[9]) ? node31532 : node31521;
													assign node31521 = (inp[4]) ? node31527 : node31522;
														assign node31522 = (inp[12]) ? node31524 : 4'b0101;
															assign node31524 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node31527 = (inp[12]) ? node31529 : 4'b0001;
															assign node31529 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node31532 = (inp[4]) ? node31534 : 4'b0001;
														assign node31534 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node31537 = (inp[5]) ? node31557 : node31538;
												assign node31538 = (inp[9]) ? node31548 : node31539;
													assign node31539 = (inp[12]) ? node31543 : node31540;
														assign node31540 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node31543 = (inp[4]) ? node31545 : 4'b0001;
															assign node31545 = (inp[10]) ? 4'b0111 : 4'b0001;
													assign node31548 = (inp[4]) ? node31552 : node31549;
														assign node31549 = (inp[12]) ? 4'b0111 : 4'b0001;
														assign node31552 = (inp[10]) ? node31554 : 4'b0111;
															assign node31554 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node31557 = (inp[2]) ? node31567 : node31558;
													assign node31558 = (inp[12]) ? 4'b0111 : node31559;
														assign node31559 = (inp[9]) ? node31563 : node31560;
															assign node31560 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node31563 = (inp[4]) ? 4'b0111 : 4'b0011;
													assign node31567 = (inp[9]) ? node31575 : node31568;
														assign node31568 = (inp[4]) ? node31570 : 4'b0111;
															assign node31570 = (inp[10]) ? node31572 : 4'b0011;
																assign node31572 = (inp[12]) ? 4'b0111 : 4'b0011;
														assign node31575 = (inp[4]) ? 4'b0111 : 4'b0011;
										assign node31578 = (inp[15]) ? node31622 : node31579;
											assign node31579 = (inp[5]) ? node31597 : node31580;
												assign node31580 = (inp[9]) ? node31588 : node31581;
													assign node31581 = (inp[4]) ? 4'b0001 : node31582;
														assign node31582 = (inp[12]) ? node31584 : 4'b0101;
															assign node31584 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node31588 = (inp[10]) ? node31590 : 4'b0111;
														assign node31590 = (inp[4]) ? node31594 : node31591;
															assign node31591 = (inp[12]) ? 4'b0111 : 4'b0001;
															assign node31594 = (inp[12]) ? 4'b0011 : 4'b0111;
												assign node31597 = (inp[2]) ? node31609 : node31598;
													assign node31598 = (inp[12]) ? node31604 : node31599;
														assign node31599 = (inp[9]) ? node31601 : 4'b0111;
															assign node31601 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node31604 = (inp[9]) ? 4'b0111 : node31605;
															assign node31605 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node31609 = (inp[10]) ? node31615 : node31610;
														assign node31610 = (inp[4]) ? 4'b0011 : node31611;
															assign node31611 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node31615 = (inp[4]) ? node31617 : 4'b0011;
															assign node31617 = (inp[12]) ? 4'b0111 : node31618;
																assign node31618 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node31622 = (inp[5]) ? node31642 : node31623;
												assign node31623 = (inp[9]) ? node31633 : node31624;
													assign node31624 = (inp[12]) ? node31628 : node31625;
														assign node31625 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node31628 = (inp[4]) ? node31630 : 4'b0011;
															assign node31630 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node31633 = (inp[4]) ? node31637 : node31634;
														assign node31634 = (inp[12]) ? 4'b0101 : 4'b0011;
														assign node31637 = (inp[12]) ? node31639 : 4'b0101;
															assign node31639 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node31642 = (inp[9]) ? node31646 : node31643;
													assign node31643 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node31646 = (inp[2]) ? 4'b0001 : node31647;
														assign node31647 = (inp[10]) ? 4'b0101 : node31648;
															assign node31648 = (inp[4]) ? 4'b0101 : 4'b0001;
								assign node31653 = (inp[9]) ? node31795 : node31654;
									assign node31654 = (inp[4]) ? node31722 : node31655;
										assign node31655 = (inp[10]) ? node31691 : node31656;
											assign node31656 = (inp[12]) ? node31680 : node31657;
												assign node31657 = (inp[3]) ? node31665 : node31658;
													assign node31658 = (inp[15]) ? node31662 : node31659;
														assign node31659 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node31662 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node31665 = (inp[15]) ? 4'b1111 : node31666;
														assign node31666 = (inp[2]) ? node31672 : node31667;
															assign node31667 = (inp[0]) ? 4'b1111 : node31668;
																assign node31668 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node31672 = (inp[5]) ? node31676 : node31673;
																assign node31673 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node31676 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node31680 = (inp[0]) ? node31688 : node31681;
													assign node31681 = (inp[15]) ? node31683 : 4'b1011;
														assign node31683 = (inp[5]) ? node31685 : 4'b1001;
															assign node31685 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node31688 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node31691 = (inp[5]) ? node31699 : node31692;
												assign node31692 = (inp[0]) ? node31696 : node31693;
													assign node31693 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node31696 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node31699 = (inp[12]) ? node31715 : node31700;
													assign node31700 = (inp[0]) ? node31706 : node31701;
														assign node31701 = (inp[15]) ? node31703 : 4'b1001;
															assign node31703 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node31706 = (inp[2]) ? node31708 : 4'b1011;
															assign node31708 = (inp[3]) ? node31712 : node31709;
																assign node31709 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node31712 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node31715 = (inp[0]) ? 4'b1001 : node31716;
														assign node31716 = (inp[2]) ? node31718 : 4'b1001;
															assign node31718 = (inp[3]) ? 4'b1001 : 4'b1011;
										assign node31722 = (inp[10]) ? node31752 : node31723;
											assign node31723 = (inp[12]) ? node31735 : node31724;
												assign node31724 = (inp[3]) ? node31728 : node31725;
													assign node31725 = (inp[2]) ? 4'b1001 : 4'b1011;
													assign node31728 = (inp[2]) ? node31730 : 4'b1001;
														assign node31730 = (inp[5]) ? node31732 : 4'b1001;
															assign node31732 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node31735 = (inp[15]) ? node31745 : node31736;
													assign node31736 = (inp[3]) ? 4'b1101 : node31737;
														assign node31737 = (inp[2]) ? 4'b1101 : node31738;
															assign node31738 = (inp[5]) ? node31740 : 4'b1111;
																assign node31740 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node31745 = (inp[0]) ? node31747 : 4'b1111;
														assign node31747 = (inp[5]) ? 4'b1101 : node31748;
															assign node31748 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node31752 = (inp[2]) ? node31778 : node31753;
												assign node31753 = (inp[5]) ? node31769 : node31754;
													assign node31754 = (inp[3]) ? node31762 : node31755;
														assign node31755 = (inp[0]) ? node31759 : node31756;
															assign node31756 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node31759 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node31762 = (inp[0]) ? node31766 : node31763;
															assign node31763 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node31766 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node31769 = (inp[12]) ? node31771 : 4'b1101;
														assign node31771 = (inp[0]) ? node31775 : node31772;
															assign node31772 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node31775 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node31778 = (inp[12]) ? node31780 : 4'b1111;
													assign node31780 = (inp[15]) ? node31790 : node31781;
														assign node31781 = (inp[0]) ? node31787 : node31782;
															assign node31782 = (inp[5]) ? 4'b1101 : node31783;
																assign node31783 = (inp[3]) ? 4'b1101 : 4'b1111;
															assign node31787 = (inp[3]) ? 4'b1111 : 4'b1101;
														assign node31790 = (inp[3]) ? node31792 : 4'b1111;
															assign node31792 = (inp[0]) ? 4'b1101 : 4'b1111;
									assign node31795 = (inp[4]) ? node31863 : node31796;
										assign node31796 = (inp[10]) ? node31826 : node31797;
											assign node31797 = (inp[12]) ? node31809 : node31798;
												assign node31798 = (inp[0]) ? node31804 : node31799;
													assign node31799 = (inp[15]) ? 4'b1001 : node31800;
														assign node31800 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node31804 = (inp[15]) ? 4'b1011 : node31805;
														assign node31805 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node31809 = (inp[5]) ? node31821 : node31810;
													assign node31810 = (inp[3]) ? node31816 : node31811;
														assign node31811 = (inp[15]) ? node31813 : 4'b1101;
															assign node31813 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node31816 = (inp[0]) ? node31818 : 4'b1111;
															assign node31818 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node31821 = (inp[2]) ? 4'b1111 : node31822;
														assign node31822 = (inp[3]) ? 4'b1111 : 4'b1101;
											assign node31826 = (inp[12]) ? node31844 : node31827;
												assign node31827 = (inp[15]) ? node31839 : node31828;
													assign node31828 = (inp[0]) ? node31834 : node31829;
														assign node31829 = (inp[5]) ? 4'b1101 : node31830;
															assign node31830 = (inp[2]) ? 4'b1111 : 4'b1101;
														assign node31834 = (inp[3]) ? 4'b1111 : node31835;
															assign node31835 = (inp[2]) ? 4'b1101 : 4'b1111;
													assign node31839 = (inp[0]) ? node31841 : 4'b1111;
														assign node31841 = (inp[5]) ? 4'b1101 : 4'b1111;
												assign node31844 = (inp[15]) ? node31854 : node31845;
													assign node31845 = (inp[0]) ? node31849 : node31846;
														assign node31846 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node31849 = (inp[2]) ? 4'b1111 : node31850;
															assign node31850 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node31854 = (inp[5]) ? 4'b1101 : node31855;
														assign node31855 = (inp[3]) ? node31859 : node31856;
															assign node31856 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node31859 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node31863 = (inp[10]) ? node31897 : node31864;
											assign node31864 = (inp[12]) ? node31876 : node31865;
												assign node31865 = (inp[0]) ? node31871 : node31866;
													assign node31866 = (inp[15]) ? node31868 : 4'b1101;
														assign node31868 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node31871 = (inp[15]) ? node31873 : 4'b1111;
														assign node31873 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node31876 = (inp[5]) ? node31890 : node31877;
													assign node31877 = (inp[15]) ? node31885 : node31878;
														assign node31878 = (inp[3]) ? node31882 : node31879;
															assign node31879 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node31882 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node31885 = (inp[3]) ? node31887 : 4'b1001;
															assign node31887 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node31890 = (inp[15]) ? node31894 : node31891;
														assign node31891 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node31894 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node31897 = (inp[12]) ? node31917 : node31898;
												assign node31898 = (inp[15]) ? node31908 : node31899;
													assign node31899 = (inp[0]) ? node31903 : node31900;
														assign node31900 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node31903 = (inp[3]) ? 4'b1011 : node31904;
															assign node31904 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node31908 = (inp[0]) ? node31912 : node31909;
														assign node31909 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node31912 = (inp[3]) ? 4'b1001 : node31913;
															assign node31913 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node31917 = (inp[3]) ? node31925 : node31918;
													assign node31918 = (inp[0]) ? 4'b1011 : node31919;
														assign node31919 = (inp[5]) ? node31921 : 4'b1011;
															assign node31921 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node31925 = (inp[0]) ? 4'b1001 : node31926;
														assign node31926 = (inp[15]) ? 4'b1011 : 4'b1001;
							assign node31930 = (inp[12]) ? node32224 : node31931;
								assign node31931 = (inp[4]) ? node32077 : node31932;
									assign node31932 = (inp[1]) ? node32002 : node31933;
										assign node31933 = (inp[15]) ? node31969 : node31934;
											assign node31934 = (inp[9]) ? node31952 : node31935;
												assign node31935 = (inp[10]) ? node31945 : node31936;
													assign node31936 = (inp[0]) ? node31940 : node31937;
														assign node31937 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node31940 = (inp[5]) ? node31942 : 4'b1101;
															assign node31942 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node31945 = (inp[5]) ? node31947 : 4'b1011;
														assign node31947 = (inp[2]) ? node31949 : 4'b1001;
															assign node31949 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node31952 = (inp[10]) ? node31964 : node31953;
													assign node31953 = (inp[0]) ? node31959 : node31954;
														assign node31954 = (inp[3]) ? node31956 : 4'b1011;
															assign node31956 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node31959 = (inp[5]) ? node31961 : 4'b1001;
															assign node31961 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node31964 = (inp[5]) ? node31966 : 4'b1101;
														assign node31966 = (inp[2]) ? 4'b1111 : 4'b1101;
											assign node31969 = (inp[0]) ? node31987 : node31970;
												assign node31970 = (inp[3]) ? node31976 : node31971;
													assign node31971 = (inp[9]) ? node31973 : 4'b1001;
														assign node31973 = (inp[10]) ? 4'b1111 : 4'b1001;
													assign node31976 = (inp[5]) ? node31982 : node31977;
														assign node31977 = (inp[9]) ? 4'b1111 : node31978;
															assign node31978 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node31982 = (inp[2]) ? node31984 : 4'b1011;
															assign node31984 = (inp[10]) ? 4'b1011 : 4'b1111;
												assign node31987 = (inp[5]) ? node31995 : node31988;
													assign node31988 = (inp[3]) ? 4'b1011 : node31989;
														assign node31989 = (inp[10]) ? node31991 : 4'b1011;
															assign node31991 = (inp[9]) ? 4'b1111 : 4'b1011;
													assign node31995 = (inp[2]) ? node31997 : 4'b1011;
														assign node31997 = (inp[3]) ? 4'b1001 : node31998;
															assign node31998 = (inp[9]) ? 4'b1101 : 4'b1111;
										assign node32002 = (inp[10]) ? node32038 : node32003;
											assign node32003 = (inp[9]) ? node32023 : node32004;
												assign node32004 = (inp[0]) ? node32012 : node32005;
													assign node32005 = (inp[15]) ? node32007 : 4'b1111;
														assign node32007 = (inp[3]) ? node32009 : 4'b1101;
															assign node32009 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node32012 = (inp[2]) ? node32014 : 4'b1101;
														assign node32014 = (inp[5]) ? node32018 : node32015;
															assign node32015 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node32018 = (inp[15]) ? 4'b1101 : node32019;
																assign node32019 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node32023 = (inp[3]) ? node32035 : node32024;
													assign node32024 = (inp[2]) ? node32030 : node32025;
														assign node32025 = (inp[15]) ? node32027 : 4'b1011;
															assign node32027 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node32030 = (inp[0]) ? node32032 : 4'b1001;
															assign node32032 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node32035 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node32038 = (inp[9]) ? node32060 : node32039;
												assign node32039 = (inp[2]) ? node32047 : node32040;
													assign node32040 = (inp[5]) ? 4'b1011 : node32041;
														assign node32041 = (inp[0]) ? 4'b1011 : node32042;
															assign node32042 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node32047 = (inp[3]) ? node32053 : node32048;
														assign node32048 = (inp[0]) ? node32050 : 4'b1011;
															assign node32050 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node32053 = (inp[0]) ? node32055 : 4'b1001;
															assign node32055 = (inp[15]) ? 4'b1011 : node32056;
																assign node32056 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node32060 = (inp[5]) ? node32070 : node32061;
													assign node32061 = (inp[0]) ? 4'b1111 : node32062;
														assign node32062 = (inp[2]) ? node32066 : node32063;
															assign node32063 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node32066 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node32070 = (inp[0]) ? node32074 : node32071;
														assign node32071 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node32074 = (inp[15]) ? 4'b1101 : 4'b1111;
									assign node32077 = (inp[10]) ? node32143 : node32078;
										assign node32078 = (inp[9]) ? node32124 : node32079;
											assign node32079 = (inp[1]) ? node32107 : node32080;
												assign node32080 = (inp[2]) ? node32090 : node32081;
													assign node32081 = (inp[15]) ? 4'b1001 : node32082;
														assign node32082 = (inp[3]) ? node32084 : 4'b1001;
															assign node32084 = (inp[0]) ? 4'b1011 : node32085;
																assign node32085 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node32090 = (inp[3]) ? node32096 : node32091;
														assign node32091 = (inp[15]) ? 4'b1011 : node32092;
															assign node32092 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node32096 = (inp[0]) ? node32102 : node32097;
															assign node32097 = (inp[5]) ? node32099 : 4'b1001;
																assign node32099 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node32102 = (inp[5]) ? node32104 : 4'b1011;
																assign node32104 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node32107 = (inp[0]) ? node32119 : node32108;
													assign node32108 = (inp[15]) ? node32114 : node32109;
														assign node32109 = (inp[3]) ? node32111 : 4'b1011;
															assign node32111 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node32114 = (inp[3]) ? node32116 : 4'b1001;
															assign node32116 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node32119 = (inp[15]) ? 4'b1011 : node32120;
														assign node32120 = (inp[3]) ? 4'b1011 : 4'b1001;
											assign node32124 = (inp[0]) ? node32134 : node32125;
												assign node32125 = (inp[15]) ? node32129 : node32126;
													assign node32126 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node32129 = (inp[3]) ? 4'b1111 : node32130;
														assign node32130 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node32134 = (inp[15]) ? node32140 : node32135;
													assign node32135 = (inp[5]) ? 4'b1111 : node32136;
														assign node32136 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node32140 = (inp[5]) ? 4'b1101 : 4'b1111;
										assign node32143 = (inp[9]) ? node32185 : node32144;
											assign node32144 = (inp[3]) ? node32168 : node32145;
												assign node32145 = (inp[0]) ? node32155 : node32146;
													assign node32146 = (inp[1]) ? node32148 : 4'b1111;
														assign node32148 = (inp[15]) ? node32152 : node32149;
															assign node32149 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node32152 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node32155 = (inp[1]) ? node32163 : node32156;
														assign node32156 = (inp[15]) ? node32160 : node32157;
															assign node32157 = (inp[5]) ? 4'b1111 : 4'b1101;
															assign node32160 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node32163 = (inp[5]) ? 4'b1101 : node32164;
															assign node32164 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node32168 = (inp[2]) ? node32178 : node32169;
													assign node32169 = (inp[5]) ? node32171 : 4'b1101;
														assign node32171 = (inp[15]) ? node32175 : node32172;
															assign node32172 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node32175 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node32178 = (inp[15]) ? node32182 : node32179;
														assign node32179 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node32182 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node32185 = (inp[1]) ? node32213 : node32186;
												assign node32186 = (inp[5]) ? node32206 : node32187;
													assign node32187 = (inp[2]) ? node32197 : node32188;
														assign node32188 = (inp[3]) ? node32190 : 4'b1001;
															assign node32190 = (inp[15]) ? node32194 : node32191;
																assign node32191 = (inp[0]) ? 4'b1011 : 4'b1001;
																assign node32194 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node32197 = (inp[3]) ? 4'b1011 : node32198;
															assign node32198 = (inp[0]) ? node32202 : node32199;
																assign node32199 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node32202 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node32206 = (inp[15]) ? node32210 : node32207;
														assign node32207 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node32210 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node32213 = (inp[0]) ? node32219 : node32214;
													assign node32214 = (inp[15]) ? node32216 : 4'b1001;
														assign node32216 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node32219 = (inp[15]) ? 4'b1001 : node32220;
														assign node32220 = (inp[3]) ? 4'b1011 : 4'b1001;
								assign node32224 = (inp[9]) ? node32352 : node32225;
									assign node32225 = (inp[4]) ? node32297 : node32226;
										assign node32226 = (inp[5]) ? node32254 : node32227;
											assign node32227 = (inp[3]) ? node32235 : node32228;
												assign node32228 = (inp[2]) ? 4'b1001 : node32229;
													assign node32229 = (inp[1]) ? node32231 : 4'b1001;
														assign node32231 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node32235 = (inp[1]) ? node32249 : node32236;
													assign node32236 = (inp[10]) ? 4'b1001 : node32237;
														assign node32237 = (inp[2]) ? node32243 : node32238;
															assign node32238 = (inp[0]) ? node32240 : 4'b1001;
																assign node32240 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node32243 = (inp[15]) ? node32245 : 4'b1011;
																assign node32245 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node32249 = (inp[15]) ? node32251 : 4'b1011;
														assign node32251 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node32254 = (inp[10]) ? node32278 : node32255;
												assign node32255 = (inp[3]) ? node32269 : node32256;
													assign node32256 = (inp[2]) ? node32262 : node32257;
														assign node32257 = (inp[15]) ? 4'b1001 : node32258;
															assign node32258 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node32262 = (inp[15]) ? node32266 : node32263;
															assign node32263 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node32266 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node32269 = (inp[1]) ? node32273 : node32270;
														assign node32270 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node32273 = (inp[15]) ? 4'b1011 : node32274;
															assign node32274 = (inp[0]) ? 4'b1011 : 4'b1001;
												assign node32278 = (inp[15]) ? node32292 : node32279;
													assign node32279 = (inp[2]) ? node32287 : node32280;
														assign node32280 = (inp[0]) ? node32284 : node32281;
															assign node32281 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node32284 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node32287 = (inp[3]) ? 4'b1001 : node32288;
															assign node32288 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node32292 = (inp[3]) ? node32294 : 4'b1011;
														assign node32294 = (inp[0]) ? 4'b1001 : 4'b1011;
										assign node32297 = (inp[3]) ? node32345 : node32298;
											assign node32298 = (inp[0]) ? node32326 : node32299;
												assign node32299 = (inp[2]) ? node32305 : node32300;
													assign node32300 = (inp[10]) ? 4'b1111 : node32301;
														assign node32301 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node32305 = (inp[10]) ? node32313 : node32306;
														assign node32306 = (inp[5]) ? node32310 : node32307;
															assign node32307 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node32310 = (inp[1]) ? 4'b1101 : 4'b1111;
														assign node32313 = (inp[1]) ? node32319 : node32314;
															assign node32314 = (inp[5]) ? node32316 : 4'b1101;
																assign node32316 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node32319 = (inp[15]) ? node32323 : node32320;
																assign node32320 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node32323 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node32326 = (inp[10]) ? node32334 : node32327;
													assign node32327 = (inp[5]) ? node32331 : node32328;
														assign node32328 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node32331 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node32334 = (inp[1]) ? node32340 : node32335;
														assign node32335 = (inp[5]) ? 4'b1101 : node32336;
															assign node32336 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node32340 = (inp[15]) ? 4'b1111 : node32341;
															assign node32341 = (inp[5]) ? 4'b1111 : 4'b1101;
											assign node32345 = (inp[0]) ? node32349 : node32346;
												assign node32346 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node32349 = (inp[15]) ? 4'b1101 : 4'b1111;
									assign node32352 = (inp[4]) ? node32412 : node32353;
										assign node32353 = (inp[5]) ? node32405 : node32354;
											assign node32354 = (inp[1]) ? node32372 : node32355;
												assign node32355 = (inp[10]) ? node32363 : node32356;
													assign node32356 = (inp[3]) ? 4'b1111 : node32357;
														assign node32357 = (inp[0]) ? node32359 : 4'b1111;
															assign node32359 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node32363 = (inp[0]) ? 4'b1111 : node32364;
														assign node32364 = (inp[15]) ? node32368 : node32365;
															assign node32365 = (inp[2]) ? 4'b1101 : 4'b1111;
															assign node32368 = (inp[3]) ? 4'b1111 : 4'b1101;
												assign node32372 = (inp[3]) ? node32388 : node32373;
													assign node32373 = (inp[10]) ? node32381 : node32374;
														assign node32374 = (inp[15]) ? node32378 : node32375;
															assign node32375 = (inp[2]) ? 4'b1111 : 4'b1101;
															assign node32378 = (inp[2]) ? 4'b1101 : 4'b1111;
														assign node32381 = (inp[0]) ? node32385 : node32382;
															assign node32382 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node32385 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node32388 = (inp[10]) ? node32400 : node32389;
														assign node32389 = (inp[2]) ? node32395 : node32390;
															assign node32390 = (inp[0]) ? 4'b1111 : node32391;
																assign node32391 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node32395 = (inp[0]) ? node32397 : 4'b1101;
																assign node32397 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node32400 = (inp[0]) ? 4'b1101 : node32401;
															assign node32401 = (inp[15]) ? 4'b1111 : 4'b1101;
											assign node32405 = (inp[15]) ? node32409 : node32406;
												assign node32406 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node32409 = (inp[0]) ? 4'b1101 : 4'b1111;
										assign node32412 = (inp[3]) ? node32440 : node32413;
											assign node32413 = (inp[15]) ? node32427 : node32414;
												assign node32414 = (inp[2]) ? node32422 : node32415;
													assign node32415 = (inp[0]) ? node32419 : node32416;
														assign node32416 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node32419 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node32422 = (inp[5]) ? 4'b1011 : node32423;
														assign node32423 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node32427 = (inp[2]) ? node32435 : node32428;
													assign node32428 = (inp[0]) ? node32432 : node32429;
														assign node32429 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node32432 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node32435 = (inp[0]) ? node32437 : 4'b1001;
														assign node32437 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node32440 = (inp[1]) ? node32448 : node32441;
												assign node32441 = (inp[15]) ? node32445 : node32442;
													assign node32442 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node32445 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node32448 = (inp[2]) ? node32460 : node32449;
													assign node32449 = (inp[5]) ? node32457 : node32450;
														assign node32450 = (inp[10]) ? node32452 : 4'b1011;
															assign node32452 = (inp[0]) ? node32454 : 4'b1011;
																assign node32454 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node32457 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node32460 = (inp[10]) ? 4'b1011 : node32461;
														assign node32461 = (inp[0]) ? node32463 : 4'b1011;
															assign node32463 = (inp[15]) ? 4'b1001 : 4'b1011;
						assign node32467 = (inp[1]) ? node33007 : node32468;
							assign node32468 = (inp[13]) ? node32738 : node32469;
								assign node32469 = (inp[4]) ? node32613 : node32470;
									assign node32470 = (inp[9]) ? node32542 : node32471;
										assign node32471 = (inp[10]) ? node32505 : node32472;
											assign node32472 = (inp[12]) ? node32496 : node32473;
												assign node32473 = (inp[15]) ? node32487 : node32474;
													assign node32474 = (inp[3]) ? node32478 : node32475;
														assign node32475 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node32478 = (inp[2]) ? node32484 : node32479;
															assign node32479 = (inp[0]) ? 4'b1111 : node32480;
																assign node32480 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node32484 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node32487 = (inp[3]) ? node32489 : 4'b1111;
														assign node32489 = (inp[5]) ? node32493 : node32490;
															assign node32490 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node32493 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node32496 = (inp[0]) ? 4'b1011 : node32497;
													assign node32497 = (inp[15]) ? node32501 : node32498;
														assign node32498 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node32501 = (inp[5]) ? 4'b1011 : 4'b1001;
											assign node32505 = (inp[2]) ? node32529 : node32506;
												assign node32506 = (inp[5]) ? node32516 : node32507;
													assign node32507 = (inp[12]) ? node32513 : node32508;
														assign node32508 = (inp[0]) ? 4'b1001 : node32509;
															assign node32509 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node32513 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node32516 = (inp[3]) ? node32522 : node32517;
														assign node32517 = (inp[0]) ? 4'b1011 : node32518;
															assign node32518 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node32522 = (inp[15]) ? node32526 : node32523;
															assign node32523 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node32526 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node32529 = (inp[0]) ? 4'b1001 : node32530;
													assign node32530 = (inp[15]) ? node32534 : node32531;
														assign node32531 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node32534 = (inp[12]) ? 4'b1001 : node32535;
															assign node32535 = (inp[5]) ? node32537 : 4'b1001;
																assign node32537 = (inp[3]) ? 4'b1011 : 4'b1001;
										assign node32542 = (inp[12]) ? node32576 : node32543;
											assign node32543 = (inp[10]) ? node32561 : node32544;
												assign node32544 = (inp[5]) ? node32550 : node32545;
													assign node32545 = (inp[0]) ? node32547 : 4'b1001;
														assign node32547 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node32550 = (inp[15]) ? node32556 : node32551;
														assign node32551 = (inp[3]) ? node32553 : 4'b1011;
															assign node32553 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node32556 = (inp[0]) ? node32558 : 4'b1001;
															assign node32558 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node32561 = (inp[5]) ? node32567 : node32562;
													assign node32562 = (inp[0]) ? node32564 : 4'b1111;
														assign node32564 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node32567 = (inp[3]) ? node32569 : 4'b1101;
														assign node32569 = (inp[15]) ? node32573 : node32570;
															assign node32570 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node32573 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node32576 = (inp[3]) ? node32600 : node32577;
												assign node32577 = (inp[10]) ? node32591 : node32578;
													assign node32578 = (inp[15]) ? node32586 : node32579;
														assign node32579 = (inp[0]) ? node32583 : node32580;
															assign node32580 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node32583 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node32586 = (inp[2]) ? 4'b1101 : node32587;
															assign node32587 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node32591 = (inp[5]) ? node32593 : 4'b1111;
														assign node32593 = (inp[2]) ? node32595 : 4'b1101;
															assign node32595 = (inp[15]) ? node32597 : 4'b1111;
																assign node32597 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node32600 = (inp[5]) ? node32608 : node32601;
													assign node32601 = (inp[15]) ? node32605 : node32602;
														assign node32602 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node32605 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node32608 = (inp[0]) ? 4'b1101 : node32609;
														assign node32609 = (inp[15]) ? 4'b1111 : 4'b1101;
									assign node32613 = (inp[9]) ? node32669 : node32614;
										assign node32614 = (inp[12]) ? node32654 : node32615;
											assign node32615 = (inp[10]) ? node32643 : node32616;
												assign node32616 = (inp[5]) ? node32630 : node32617;
													assign node32617 = (inp[2]) ? node32623 : node32618;
														assign node32618 = (inp[15]) ? 4'b1011 : node32619;
															assign node32619 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node32623 = (inp[0]) ? node32627 : node32624;
															assign node32624 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node32627 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node32630 = (inp[0]) ? node32636 : node32631;
														assign node32631 = (inp[15]) ? 4'b1001 : node32632;
															assign node32632 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node32636 = (inp[15]) ? node32640 : node32637;
															assign node32637 = (inp[3]) ? 4'b1011 : 4'b1001;
															assign node32640 = (inp[3]) ? 4'b1001 : 4'b1011;
												assign node32643 = (inp[5]) ? node32649 : node32644;
													assign node32644 = (inp[0]) ? 4'b1111 : node32645;
														assign node32645 = (inp[2]) ? 4'b1111 : 4'b1101;
													assign node32649 = (inp[15]) ? node32651 : 4'b1101;
														assign node32651 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node32654 = (inp[15]) ? node32662 : node32655;
												assign node32655 = (inp[0]) ? node32657 : 4'b1101;
													assign node32657 = (inp[5]) ? 4'b1111 : node32658;
														assign node32658 = (inp[2]) ? 4'b1111 : 4'b1101;
												assign node32662 = (inp[0]) ? node32664 : 4'b1111;
													assign node32664 = (inp[5]) ? 4'b1101 : node32665;
														assign node32665 = (inp[3]) ? 4'b1101 : 4'b1111;
										assign node32669 = (inp[12]) ? node32711 : node32670;
											assign node32670 = (inp[10]) ? node32690 : node32671;
												assign node32671 = (inp[0]) ? node32685 : node32672;
													assign node32672 = (inp[2]) ? node32678 : node32673;
														assign node32673 = (inp[3]) ? node32675 : 4'b1111;
															assign node32675 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node32678 = (inp[5]) ? 4'b1101 : node32679;
															assign node32679 = (inp[3]) ? 4'b1101 : node32680;
																assign node32680 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node32685 = (inp[15]) ? node32687 : 4'b1111;
														assign node32687 = (inp[3]) ? 4'b1101 : 4'b1111;
												assign node32690 = (inp[2]) ? node32696 : node32691;
													assign node32691 = (inp[3]) ? node32693 : 4'b1001;
														assign node32693 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node32696 = (inp[3]) ? node32704 : node32697;
														assign node32697 = (inp[15]) ? node32699 : 4'b1011;
															assign node32699 = (inp[5]) ? 4'b1011 : node32700;
																assign node32700 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node32704 = (inp[0]) ? node32708 : node32705;
															assign node32705 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node32708 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node32711 = (inp[5]) ? node32731 : node32712;
												assign node32712 = (inp[15]) ? node32720 : node32713;
													assign node32713 = (inp[2]) ? node32715 : 4'b1001;
														assign node32715 = (inp[3]) ? node32717 : 4'b1011;
															assign node32717 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node32720 = (inp[2]) ? node32722 : 4'b1011;
														assign node32722 = (inp[10]) ? node32728 : node32723;
															assign node32723 = (inp[3]) ? node32725 : 4'b1011;
																assign node32725 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node32728 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node32731 = (inp[15]) ? node32735 : node32732;
													assign node32732 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node32735 = (inp[0]) ? 4'b1001 : 4'b1011;
								assign node32738 = (inp[9]) ? node32886 : node32739;
									assign node32739 = (inp[4]) ? node32823 : node32740;
										assign node32740 = (inp[10]) ? node32790 : node32741;
											assign node32741 = (inp[12]) ? node32771 : node32742;
												assign node32742 = (inp[2]) ? node32758 : node32743;
													assign node32743 = (inp[0]) ? node32751 : node32744;
														assign node32744 = (inp[3]) ? node32746 : 4'b0111;
															assign node32746 = (inp[15]) ? 4'b0111 : node32747;
																assign node32747 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node32751 = (inp[3]) ? node32755 : node32752;
															assign node32752 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node32755 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node32758 = (inp[15]) ? node32766 : node32759;
														assign node32759 = (inp[0]) ? node32763 : node32760;
															assign node32760 = (inp[3]) ? 4'b0101 : 4'b0111;
															assign node32763 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node32766 = (inp[0]) ? node32768 : 4'b0101;
															assign node32768 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node32771 = (inp[2]) ? node32781 : node32772;
													assign node32772 = (inp[0]) ? node32776 : node32773;
														assign node32773 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node32776 = (inp[15]) ? node32778 : 4'b0001;
															assign node32778 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node32781 = (inp[15]) ? 4'b0011 : node32782;
														assign node32782 = (inp[5]) ? node32784 : 4'b0011;
															assign node32784 = (inp[3]) ? node32786 : 4'b0001;
																assign node32786 = (inp[0]) ? 4'b0011 : 4'b0001;
											assign node32790 = (inp[5]) ? node32798 : node32791;
												assign node32791 = (inp[15]) ? node32795 : node32792;
													assign node32792 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node32795 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node32798 = (inp[0]) ? node32814 : node32799;
													assign node32799 = (inp[2]) ? node32805 : node32800;
														assign node32800 = (inp[3]) ? node32802 : 4'b0011;
															assign node32802 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node32805 = (inp[12]) ? node32809 : node32806;
															assign node32806 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node32809 = (inp[15]) ? 4'b0001 : node32810;
																assign node32810 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node32814 = (inp[12]) ? 4'b0011 : node32815;
														assign node32815 = (inp[15]) ? node32819 : node32816;
															assign node32816 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node32819 = (inp[2]) ? 4'b0011 : 4'b0001;
										assign node32823 = (inp[10]) ? node32857 : node32824;
											assign node32824 = (inp[12]) ? node32844 : node32825;
												assign node32825 = (inp[3]) ? node32831 : node32826;
													assign node32826 = (inp[0]) ? node32828 : 4'b0001;
														assign node32828 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node32831 = (inp[5]) ? node32839 : node32832;
														assign node32832 = (inp[0]) ? node32836 : node32833;
															assign node32833 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node32836 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node32839 = (inp[0]) ? 4'b0011 : node32840;
															assign node32840 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node32844 = (inp[0]) ? node32854 : node32845;
													assign node32845 = (inp[15]) ? node32849 : node32846;
														assign node32846 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node32849 = (inp[5]) ? 4'b0111 : node32850;
															assign node32850 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node32854 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node32857 = (inp[12]) ? node32871 : node32858;
												assign node32858 = (inp[5]) ? node32864 : node32859;
													assign node32859 = (inp[3]) ? 4'b0101 : node32860;
														assign node32860 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node32864 = (inp[15]) ? node32868 : node32865;
														assign node32865 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node32868 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node32871 = (inp[15]) ? node32875 : node32872;
													assign node32872 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node32875 = (inp[0]) ? node32881 : node32876;
														assign node32876 = (inp[5]) ? 4'b0111 : node32877;
															assign node32877 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node32881 = (inp[5]) ? 4'b0101 : node32882;
															assign node32882 = (inp[3]) ? 4'b0101 : 4'b0111;
									assign node32886 = (inp[4]) ? node32960 : node32887;
										assign node32887 = (inp[10]) ? node32927 : node32888;
											assign node32888 = (inp[12]) ? node32908 : node32889;
												assign node32889 = (inp[5]) ? node32895 : node32890;
													assign node32890 = (inp[0]) ? node32892 : 4'b0011;
														assign node32892 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node32895 = (inp[2]) ? 4'b0001 : node32896;
														assign node32896 = (inp[3]) ? node32902 : node32897;
															assign node32897 = (inp[0]) ? node32899 : 4'b0001;
																assign node32899 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node32902 = (inp[15]) ? node32904 : 4'b0011;
																assign node32904 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node32908 = (inp[0]) ? node32920 : node32909;
													assign node32909 = (inp[15]) ? node32915 : node32910;
														assign node32910 = (inp[5]) ? 4'b0101 : node32911;
															assign node32911 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node32915 = (inp[5]) ? 4'b0111 : node32916;
															assign node32916 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node32920 = (inp[15]) ? node32922 : 4'b0111;
														assign node32922 = (inp[5]) ? 4'b0101 : node32923;
															assign node32923 = (inp[3]) ? 4'b0101 : 4'b0111;
											assign node32927 = (inp[2]) ? node32941 : node32928;
												assign node32928 = (inp[15]) ? node32932 : node32929;
													assign node32929 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node32932 = (inp[0]) ? node32936 : node32933;
														assign node32933 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node32936 = (inp[5]) ? 4'b0101 : node32937;
															assign node32937 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node32941 = (inp[0]) ? node32951 : node32942;
													assign node32942 = (inp[5]) ? node32948 : node32943;
														assign node32943 = (inp[12]) ? 4'b0111 : node32944;
															assign node32944 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node32948 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node32951 = (inp[15]) ? node32955 : node32952;
														assign node32952 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node32955 = (inp[5]) ? 4'b0101 : node32956;
															assign node32956 = (inp[3]) ? 4'b0101 : 4'b0111;
										assign node32960 = (inp[10]) ? node32990 : node32961;
											assign node32961 = (inp[12]) ? node32973 : node32962;
												assign node32962 = (inp[0]) ? node32968 : node32963;
													assign node32963 = (inp[5]) ? node32965 : 4'b0101;
														assign node32965 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node32968 = (inp[15]) ? node32970 : 4'b0111;
														assign node32970 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node32973 = (inp[3]) ? node32985 : node32974;
													assign node32974 = (inp[0]) ? node32980 : node32975;
														assign node32975 = (inp[5]) ? node32977 : 4'b0001;
															assign node32977 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node32980 = (inp[15]) ? node32982 : 4'b0011;
															assign node32982 = (inp[5]) ? 4'b0001 : 4'b0011;
													assign node32985 = (inp[15]) ? node32987 : 4'b0001;
														assign node32987 = (inp[5]) ? 4'b0001 : 4'b0011;
											assign node32990 = (inp[15]) ? node32996 : node32991;
												assign node32991 = (inp[0]) ? node32993 : 4'b0001;
													assign node32993 = (inp[5]) ? 4'b0011 : 4'b0001;
												assign node32996 = (inp[0]) ? node33002 : node32997;
													assign node32997 = (inp[3]) ? 4'b0011 : node32998;
														assign node32998 = (inp[5]) ? 4'b0011 : 4'b0001;
													assign node33002 = (inp[3]) ? 4'b0001 : node33003;
														assign node33003 = (inp[5]) ? 4'b0001 : 4'b0011;
							assign node33007 = (inp[5]) ? node33305 : node33008;
								assign node33008 = (inp[12]) ? node33220 : node33009;
									assign node33009 = (inp[13]) ? node33107 : node33010;
										assign node33010 = (inp[9]) ? node33062 : node33011;
											assign node33011 = (inp[3]) ? node33039 : node33012;
												assign node33012 = (inp[15]) ? node33032 : node33013;
													assign node33013 = (inp[0]) ? node33025 : node33014;
														assign node33014 = (inp[2]) ? node33020 : node33015;
															assign node33015 = (inp[4]) ? node33017 : 4'b0111;
																assign node33017 = (inp[10]) ? 4'b0111 : 4'b0011;
															assign node33020 = (inp[4]) ? 4'b0111 : node33021;
																assign node33021 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node33025 = (inp[10]) ? node33029 : node33026;
															assign node33026 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node33029 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node33032 = (inp[0]) ? 4'b0111 : node33033;
														assign node33033 = (inp[10]) ? node33035 : 4'b0101;
															assign node33035 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node33039 = (inp[10]) ? node33051 : node33040;
													assign node33040 = (inp[4]) ? node33046 : node33041;
														assign node33041 = (inp[15]) ? 4'b0101 : node33042;
															assign node33042 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node33046 = (inp[15]) ? 4'b0011 : node33047;
															assign node33047 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node33051 = (inp[4]) ? node33057 : node33052;
														assign node33052 = (inp[15]) ? node33054 : 4'b0011;
															assign node33054 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node33057 = (inp[0]) ? 4'b0111 : node33058;
															assign node33058 = (inp[15]) ? 4'b0111 : 4'b0101;
											assign node33062 = (inp[15]) ? node33086 : node33063;
												assign node33063 = (inp[0]) ? node33071 : node33064;
													assign node33064 = (inp[4]) ? node33066 : 4'b0011;
														assign node33066 = (inp[2]) ? node33068 : 4'b0101;
															assign node33068 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node33071 = (inp[3]) ? node33079 : node33072;
														assign node33072 = (inp[2]) ? node33074 : 4'b0101;
															assign node33074 = (inp[10]) ? 4'b0001 : node33075;
																assign node33075 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node33079 = (inp[4]) ? node33083 : node33080;
															assign node33080 = (inp[10]) ? 4'b0111 : 4'b0001;
															assign node33083 = (inp[10]) ? 4'b0011 : 4'b0111;
												assign node33086 = (inp[0]) ? node33096 : node33087;
													assign node33087 = (inp[10]) ? node33089 : 4'b0001;
														assign node33089 = (inp[3]) ? node33093 : node33090;
															assign node33090 = (inp[2]) ? 4'b0101 : 4'b0001;
															assign node33093 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node33096 = (inp[3]) ? node33104 : node33097;
														assign node33097 = (inp[10]) ? node33101 : node33098;
															assign node33098 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node33101 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node33104 = (inp[10]) ? 4'b0001 : 4'b0011;
										assign node33107 = (inp[2]) ? node33165 : node33108;
											assign node33108 = (inp[3]) ? node33138 : node33109;
												assign node33109 = (inp[4]) ? node33123 : node33110;
													assign node33110 = (inp[9]) ? node33116 : node33111;
														assign node33111 = (inp[15]) ? node33113 : 4'b0001;
															assign node33113 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node33116 = (inp[10]) ? 4'b0101 : node33117;
															assign node33117 = (inp[0]) ? 4'b0001 : node33118;
																assign node33118 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node33123 = (inp[10]) ? node33129 : node33124;
														assign node33124 = (inp[0]) ? 4'b0011 : node33125;
															assign node33125 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node33129 = (inp[9]) ? node33131 : 4'b0101;
															assign node33131 = (inp[0]) ? node33135 : node33132;
																assign node33132 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node33135 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node33138 = (inp[4]) ? node33152 : node33139;
													assign node33139 = (inp[0]) ? node33143 : node33140;
														assign node33140 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node33143 = (inp[15]) ? node33147 : node33144;
															assign node33144 = (inp[9]) ? 4'b0111 : 4'b0101;
															assign node33147 = (inp[10]) ? 4'b0011 : node33148;
																assign node33148 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node33152 = (inp[0]) ? node33158 : node33153;
														assign node33153 = (inp[10]) ? node33155 : 4'b0011;
															assign node33155 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node33158 = (inp[15]) ? node33160 : 4'b0011;
															assign node33160 = (inp[9]) ? node33162 : 4'b0011;
																assign node33162 = (inp[10]) ? 4'b0001 : 4'b0101;
											assign node33165 = (inp[10]) ? node33201 : node33166;
												assign node33166 = (inp[4]) ? node33180 : node33167;
													assign node33167 = (inp[9]) ? node33177 : node33168;
														assign node33168 = (inp[3]) ? 4'b0111 : node33169;
															assign node33169 = (inp[0]) ? node33173 : node33170;
																assign node33170 = (inp[15]) ? 4'b0101 : 4'b0111;
																assign node33173 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node33177 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node33180 = (inp[9]) ? node33194 : node33181;
														assign node33181 = (inp[3]) ? node33189 : node33182;
															assign node33182 = (inp[0]) ? node33186 : node33183;
																assign node33183 = (inp[15]) ? 4'b0001 : 4'b0011;
																assign node33186 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node33189 = (inp[0]) ? 4'b0001 : node33190;
																assign node33190 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node33194 = (inp[3]) ? node33198 : node33195;
															assign node33195 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node33198 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node33201 = (inp[3]) ? node33215 : node33202;
													assign node33202 = (inp[9]) ? node33210 : node33203;
														assign node33203 = (inp[4]) ? 4'b0101 : node33204;
															assign node33204 = (inp[0]) ? node33206 : 4'b0001;
																assign node33206 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node33210 = (inp[0]) ? 4'b0111 : node33211;
															assign node33211 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node33215 = (inp[4]) ? 4'b0111 : node33216;
														assign node33216 = (inp[9]) ? 4'b0101 : 4'b0001;
									assign node33220 = (inp[0]) ? node33264 : node33221;
										assign node33221 = (inp[15]) ? node33249 : node33222;
											assign node33222 = (inp[3]) ? node33242 : node33223;
												assign node33223 = (inp[2]) ? node33231 : node33224;
													assign node33224 = (inp[4]) ? node33228 : node33225;
														assign node33225 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node33228 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node33231 = (inp[10]) ? 4'b0011 : node33232;
														assign node33232 = (inp[13]) ? node33236 : node33233;
															assign node33233 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node33236 = (inp[4]) ? node33238 : 4'b0011;
																assign node33238 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node33242 = (inp[9]) ? node33246 : node33243;
													assign node33243 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node33246 = (inp[4]) ? 4'b0001 : 4'b0101;
											assign node33249 = (inp[3]) ? node33257 : node33250;
												assign node33250 = (inp[9]) ? node33254 : node33251;
													assign node33251 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node33254 = (inp[4]) ? 4'b0001 : 4'b0101;
												assign node33257 = (inp[4]) ? node33261 : node33258;
													assign node33258 = (inp[9]) ? 4'b0111 : 4'b0001;
													assign node33261 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node33264 = (inp[15]) ? node33282 : node33265;
											assign node33265 = (inp[3]) ? node33273 : node33266;
												assign node33266 = (inp[4]) ? node33270 : node33267;
													assign node33267 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node33270 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node33273 = (inp[10]) ? 4'b0111 : node33274;
													assign node33274 = (inp[9]) ? node33278 : node33275;
														assign node33275 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node33278 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node33282 = (inp[3]) ? node33298 : node33283;
												assign node33283 = (inp[10]) ? node33291 : node33284;
													assign node33284 = (inp[2]) ? node33286 : 4'b0111;
														assign node33286 = (inp[9]) ? node33288 : 4'b0011;
															assign node33288 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node33291 = (inp[9]) ? node33295 : node33292;
														assign node33292 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node33295 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node33298 = (inp[4]) ? node33302 : node33299;
													assign node33299 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node33302 = (inp[9]) ? 4'b0001 : 4'b0101;
								assign node33305 = (inp[12]) ? node33489 : node33306;
									assign node33306 = (inp[13]) ? node33408 : node33307;
										assign node33307 = (inp[0]) ? node33357 : node33308;
											assign node33308 = (inp[15]) ? node33330 : node33309;
												assign node33309 = (inp[3]) ? node33321 : node33310;
													assign node33310 = (inp[9]) ? node33316 : node33311;
														assign node33311 = (inp[4]) ? 4'b0011 : node33312;
															assign node33312 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node33316 = (inp[10]) ? node33318 : 4'b0011;
															assign node33318 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node33321 = (inp[2]) ? 4'b0001 : node33322;
														assign node33322 = (inp[4]) ? 4'b0101 : node33323;
															assign node33323 = (inp[10]) ? node33325 : 4'b0101;
																assign node33325 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node33330 = (inp[3]) ? node33346 : node33331;
													assign node33331 = (inp[9]) ? node33341 : node33332;
														assign node33332 = (inp[2]) ? 4'b0111 : node33333;
															assign node33333 = (inp[4]) ? node33337 : node33334;
																assign node33334 = (inp[10]) ? 4'b0001 : 4'b0101;
																assign node33337 = (inp[10]) ? 4'b0111 : 4'b0001;
														assign node33341 = (inp[4]) ? node33343 : 4'b0111;
															assign node33343 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node33346 = (inp[2]) ? node33348 : 4'b0111;
														assign node33348 = (inp[10]) ? node33350 : 4'b0011;
															assign node33350 = (inp[9]) ? node33354 : node33351;
																assign node33351 = (inp[4]) ? 4'b0111 : 4'b0011;
																assign node33354 = (inp[4]) ? 4'b0011 : 4'b0111;
											assign node33357 = (inp[15]) ? node33387 : node33358;
												assign node33358 = (inp[3]) ? node33370 : node33359;
													assign node33359 = (inp[10]) ? node33365 : node33360;
														assign node33360 = (inp[4]) ? 4'b0001 : node33361;
															assign node33361 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node33365 = (inp[2]) ? node33367 : 4'b0111;
															assign node33367 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node33370 = (inp[9]) ? node33378 : node33371;
														assign node33371 = (inp[2]) ? 4'b0011 : node33372;
															assign node33372 = (inp[4]) ? 4'b0011 : node33373;
																assign node33373 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node33378 = (inp[2]) ? node33384 : node33379;
															assign node33379 = (inp[4]) ? node33381 : 4'b0111;
																assign node33381 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node33384 = (inp[4]) ? 4'b0111 : 4'b0011;
												assign node33387 = (inp[3]) ? node33395 : node33388;
													assign node33388 = (inp[4]) ? node33390 : 4'b0111;
														assign node33390 = (inp[9]) ? 4'b0101 : node33391;
															assign node33391 = (inp[10]) ? 4'b0101 : 4'b0011;
													assign node33395 = (inp[10]) ? node33401 : node33396;
														assign node33396 = (inp[4]) ? node33398 : 4'b0001;
															assign node33398 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node33401 = (inp[9]) ? node33405 : node33402;
															assign node33402 = (inp[4]) ? 4'b0101 : 4'b0001;
															assign node33405 = (inp[4]) ? 4'b0001 : 4'b0101;
										assign node33408 = (inp[4]) ? node33452 : node33409;
											assign node33409 = (inp[0]) ? node33433 : node33410;
												assign node33410 = (inp[9]) ? node33424 : node33411;
													assign node33411 = (inp[10]) ? node33417 : node33412;
														assign node33412 = (inp[2]) ? node33414 : 4'b0111;
															assign node33414 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node33417 = (inp[3]) ? node33421 : node33418;
															assign node33418 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node33421 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node33424 = (inp[10]) ? node33430 : node33425;
														assign node33425 = (inp[15]) ? 4'b0001 : node33426;
															assign node33426 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node33430 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node33433 = (inp[9]) ? node33443 : node33434;
													assign node33434 = (inp[2]) ? 4'b0101 : node33435;
														assign node33435 = (inp[3]) ? node33439 : node33436;
															assign node33436 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node33439 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node33443 = (inp[10]) ? node33449 : node33444;
														assign node33444 = (inp[2]) ? 4'b0011 : node33445;
															assign node33445 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node33449 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node33452 = (inp[2]) ? node33466 : node33453;
												assign node33453 = (inp[15]) ? node33455 : 4'b0001;
													assign node33455 = (inp[0]) ? node33459 : node33456;
														assign node33456 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node33459 = (inp[10]) ? node33463 : node33460;
															assign node33460 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node33463 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node33466 = (inp[0]) ? node33476 : node33467;
													assign node33467 = (inp[15]) ? node33473 : node33468;
														assign node33468 = (inp[9]) ? node33470 : 4'b0001;
															assign node33470 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node33473 = (inp[9]) ? 4'b0011 : 4'b0001;
													assign node33476 = (inp[15]) ? node33484 : node33477;
														assign node33477 = (inp[3]) ? node33479 : 4'b0111;
															assign node33479 = (inp[10]) ? node33481 : 4'b0011;
																assign node33481 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node33484 = (inp[10]) ? 4'b0001 : node33485;
															assign node33485 = (inp[3]) ? 4'b0001 : 4'b0011;
									assign node33489 = (inp[13]) ? node33561 : node33490;
										assign node33490 = (inp[10]) ? node33524 : node33491;
											assign node33491 = (inp[4]) ? node33505 : node33492;
												assign node33492 = (inp[9]) ? node33500 : node33493;
													assign node33493 = (inp[3]) ? node33495 : 4'b0011;
														assign node33495 = (inp[0]) ? 4'b0011 : node33496;
															assign node33496 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node33500 = (inp[15]) ? 4'b0101 : node33501;
														assign node33501 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node33505 = (inp[9]) ? node33519 : node33506;
													assign node33506 = (inp[3]) ? node33514 : node33507;
														assign node33507 = (inp[15]) ? node33511 : node33508;
															assign node33508 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node33511 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node33514 = (inp[15]) ? node33516 : 4'b0111;
															assign node33516 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node33519 = (inp[15]) ? node33521 : 4'b0011;
														assign node33521 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node33524 = (inp[9]) ? node33546 : node33525;
												assign node33525 = (inp[4]) ? node33541 : node33526;
													assign node33526 = (inp[2]) ? node33538 : node33527;
														assign node33527 = (inp[15]) ? node33533 : node33528;
															assign node33528 = (inp[0]) ? 4'b0011 : node33529;
																assign node33529 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node33533 = (inp[0]) ? node33535 : 4'b0001;
																assign node33535 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node33538 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node33541 = (inp[0]) ? 4'b0101 : node33542;
														assign node33542 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node33546 = (inp[4]) ? node33554 : node33547;
													assign node33547 = (inp[0]) ? node33551 : node33548;
														assign node33548 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node33551 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node33554 = (inp[15]) ? node33558 : node33555;
														assign node33555 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node33558 = (inp[0]) ? 4'b0001 : 4'b0011;
										assign node33561 = (inp[4]) ? node33579 : node33562;
											assign node33562 = (inp[9]) ? node33572 : node33563;
												assign node33563 = (inp[15]) ? node33565 : 4'b0011;
													assign node33565 = (inp[3]) ? node33569 : node33566;
														assign node33566 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node33569 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node33572 = (inp[0]) ? node33576 : node33573;
													assign node33573 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node33576 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node33579 = (inp[9]) ? node33601 : node33580;
												assign node33580 = (inp[2]) ? node33588 : node33581;
													assign node33581 = (inp[15]) ? node33585 : node33582;
														assign node33582 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node33585 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node33588 = (inp[10]) ? node33596 : node33589;
														assign node33589 = (inp[0]) ? node33593 : node33590;
															assign node33590 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node33593 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node33596 = (inp[0]) ? node33598 : 4'b0111;
															assign node33598 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node33601 = (inp[3]) ? node33607 : node33602;
													assign node33602 = (inp[15]) ? node33604 : 4'b0011;
														assign node33604 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node33607 = (inp[15]) ? 4'b0011 : node33608;
														assign node33608 = (inp[0]) ? 4'b0011 : 4'b0001;
			assign node33612 = (inp[7]) ? node38970 : node33613;
				assign node33613 = (inp[13]) ? node36467 : node33614;
					assign node33614 = (inp[4]) ? node35028 : node33615;
						assign node33615 = (inp[5]) ? node34271 : node33616;
							assign node33616 = (inp[15]) ? node33966 : node33617;
								assign node33617 = (inp[0]) ? node33791 : node33618;
									assign node33618 = (inp[9]) ? node33702 : node33619;
										assign node33619 = (inp[10]) ? node33651 : node33620;
											assign node33620 = (inp[12]) ? node33640 : node33621;
												assign node33621 = (inp[3]) ? node33627 : node33622;
													assign node33622 = (inp[11]) ? 4'b1111 : node33623;
														assign node33623 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node33627 = (inp[2]) ? node33633 : node33628;
														assign node33628 = (inp[11]) ? node33630 : 4'b1111;
															assign node33630 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node33633 = (inp[11]) ? node33635 : 4'b0111;
															assign node33635 = (inp[1]) ? 4'b0111 : node33636;
																assign node33636 = (inp[6]) ? 4'b1111 : 4'b0111;
												assign node33640 = (inp[11]) ? node33648 : node33641;
													assign node33641 = (inp[6]) ? node33645 : node33642;
														assign node33642 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node33645 = (inp[1]) ? 4'b1011 : 4'b0111;
													assign node33648 = (inp[2]) ? 4'b1011 : 4'b0011;
											assign node33651 = (inp[12]) ? node33669 : node33652;
												assign node33652 = (inp[1]) ? node33660 : node33653;
													assign node33653 = (inp[6]) ? node33657 : node33654;
														assign node33654 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node33657 = (inp[11]) ? 4'b1011 : 4'b0111;
													assign node33660 = (inp[3]) ? 4'b1011 : node33661;
														assign node33661 = (inp[2]) ? 4'b1011 : node33662;
															assign node33662 = (inp[11]) ? node33664 : 4'b0111;
																assign node33664 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node33669 = (inp[6]) ? node33685 : node33670;
													assign node33670 = (inp[3]) ? 4'b1011 : node33671;
														assign node33671 = (inp[2]) ? node33679 : node33672;
															assign node33672 = (inp[11]) ? node33676 : node33673;
																assign node33673 = (inp[1]) ? 4'b0011 : 4'b1011;
																assign node33676 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node33679 = (inp[11]) ? node33681 : 4'b1011;
																assign node33681 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node33685 = (inp[2]) ? node33695 : node33686;
														assign node33686 = (inp[3]) ? node33688 : 4'b0011;
															assign node33688 = (inp[1]) ? node33692 : node33689;
																assign node33689 = (inp[11]) ? 4'b1011 : 4'b0011;
																assign node33692 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node33695 = (inp[11]) ? node33699 : node33696;
															assign node33696 = (inp[3]) ? 4'b0011 : 4'b1011;
															assign node33699 = (inp[1]) ? 4'b0011 : 4'b1011;
										assign node33702 = (inp[12]) ? node33746 : node33703;
											assign node33703 = (inp[10]) ? node33729 : node33704;
												assign node33704 = (inp[6]) ? node33716 : node33705;
													assign node33705 = (inp[2]) ? node33711 : node33706;
														assign node33706 = (inp[1]) ? node33708 : 4'b1011;
															assign node33708 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node33711 = (inp[1]) ? node33713 : 4'b0011;
															assign node33713 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node33716 = (inp[2]) ? node33722 : node33717;
														assign node33717 = (inp[3]) ? 4'b0011 : node33718;
															assign node33718 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node33722 = (inp[11]) ? node33726 : node33723;
															assign node33723 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node33726 = (inp[1]) ? 4'b0011 : 4'b1011;
												assign node33729 = (inp[6]) ? node33739 : node33730;
													assign node33730 = (inp[11]) ? node33734 : node33731;
														assign node33731 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node33734 = (inp[1]) ? node33736 : 4'b0011;
															assign node33736 = (inp[3]) ? 4'b1101 : 4'b1111;
													assign node33739 = (inp[11]) ? node33743 : node33740;
														assign node33740 = (inp[1]) ? 4'b1101 : 4'b0011;
														assign node33743 = (inp[1]) ? 4'b0101 : 4'b1101;
											assign node33746 = (inp[3]) ? node33770 : node33747;
												assign node33747 = (inp[10]) ? node33761 : node33748;
													assign node33748 = (inp[1]) ? node33754 : node33749;
														assign node33749 = (inp[11]) ? 4'b0011 : node33750;
															assign node33750 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node33754 = (inp[2]) ? node33756 : 4'b1111;
															assign node33756 = (inp[6]) ? node33758 : 4'b0011;
																assign node33758 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node33761 = (inp[11]) ? 4'b0111 : node33762;
														assign node33762 = (inp[6]) ? node33766 : node33763;
															assign node33763 = (inp[1]) ? 4'b0111 : 4'b1111;
															assign node33766 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node33770 = (inp[10]) ? node33780 : node33771;
													assign node33771 = (inp[6]) ? node33775 : node33772;
														assign node33772 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node33775 = (inp[1]) ? node33777 : 4'b1101;
															assign node33777 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node33780 = (inp[2]) ? node33784 : node33781;
														assign node33781 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node33784 = (inp[1]) ? node33786 : 4'b0101;
															assign node33786 = (inp[11]) ? 4'b1101 : node33787;
																assign node33787 = (inp[6]) ? 4'b1101 : 4'b0101;
									assign node33791 = (inp[3]) ? node33869 : node33792;
										assign node33792 = (inp[1]) ? node33832 : node33793;
											assign node33793 = (inp[9]) ? node33817 : node33794;
												assign node33794 = (inp[12]) ? node33800 : node33795;
													assign node33795 = (inp[11]) ? 4'b0101 : node33796;
														assign node33796 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node33800 = (inp[10]) ? node33808 : node33801;
														assign node33801 = (inp[11]) ? node33805 : node33802;
															assign node33802 = (inp[2]) ? 4'b0101 : 4'b1101;
															assign node33805 = (inp[6]) ? 4'b1001 : 4'b0101;
														assign node33808 = (inp[2]) ? node33810 : 4'b0001;
															assign node33810 = (inp[11]) ? node33814 : node33811;
																assign node33811 = (inp[6]) ? 4'b0001 : 4'b1001;
																assign node33814 = (inp[6]) ? 4'b1001 : 4'b0001;
												assign node33817 = (inp[11]) ? node33821 : node33818;
													assign node33818 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node33821 = (inp[6]) ? node33827 : node33822;
														assign node33822 = (inp[2]) ? node33824 : 4'b0001;
															assign node33824 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node33827 = (inp[10]) ? 4'b1101 : node33828;
															assign node33828 = (inp[12]) ? 4'b1101 : 4'b1001;
											assign node33832 = (inp[9]) ? node33852 : node33833;
												assign node33833 = (inp[11]) ? node33845 : node33834;
													assign node33834 = (inp[6]) ? node33840 : node33835;
														assign node33835 = (inp[10]) ? node33837 : 4'b0101;
															assign node33837 = (inp[12]) ? 4'b0001 : 4'b0101;
														assign node33840 = (inp[12]) ? 4'b1001 : node33841;
															assign node33841 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node33845 = (inp[6]) ? 4'b0001 : node33846;
														assign node33846 = (inp[2]) ? 4'b1001 : node33847;
															assign node33847 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node33852 = (inp[11]) ? node33860 : node33853;
													assign node33853 = (inp[6]) ? node33855 : 4'b0001;
														assign node33855 = (inp[10]) ? 4'b1101 : node33856;
															assign node33856 = (inp[12]) ? 4'b1101 : 4'b1001;
													assign node33860 = (inp[6]) ? node33862 : 4'b1101;
														assign node33862 = (inp[2]) ? node33864 : 4'b0101;
															assign node33864 = (inp[12]) ? 4'b0101 : node33865;
																assign node33865 = (inp[10]) ? 4'b0101 : 4'b0001;
										assign node33869 = (inp[9]) ? node33925 : node33870;
											assign node33870 = (inp[10]) ? node33892 : node33871;
												assign node33871 = (inp[11]) ? node33885 : node33872;
													assign node33872 = (inp[12]) ? node33878 : node33873;
														assign node33873 = (inp[1]) ? 4'b1101 : node33874;
															assign node33874 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node33878 = (inp[1]) ? node33882 : node33879;
															assign node33879 = (inp[6]) ? 4'b0101 : 4'b1101;
															assign node33882 = (inp[6]) ? 4'b1001 : 4'b0101;
													assign node33885 = (inp[12]) ? node33889 : node33886;
														assign node33886 = (inp[6]) ? 4'b1101 : 4'b0101;
														assign node33889 = (inp[2]) ? 4'b1001 : 4'b0001;
												assign node33892 = (inp[12]) ? node33910 : node33893;
													assign node33893 = (inp[1]) ? node33901 : node33894;
														assign node33894 = (inp[2]) ? node33896 : 4'b1101;
															assign node33896 = (inp[11]) ? 4'b0101 : node33897;
																assign node33897 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node33901 = (inp[2]) ? node33903 : 4'b1001;
															assign node33903 = (inp[11]) ? node33907 : node33904;
																assign node33904 = (inp[6]) ? 4'b1001 : 4'b0101;
																assign node33907 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node33910 = (inp[6]) ? node33916 : node33911;
														assign node33911 = (inp[11]) ? 4'b0001 : node33912;
															assign node33912 = (inp[2]) ? 4'b0001 : 4'b1001;
														assign node33916 = (inp[2]) ? 4'b1001 : node33917;
															assign node33917 = (inp[1]) ? node33921 : node33918;
																assign node33918 = (inp[11]) ? 4'b1001 : 4'b0001;
																assign node33921 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node33925 = (inp[10]) ? node33943 : node33926;
												assign node33926 = (inp[11]) ? node33934 : node33927;
													assign node33927 = (inp[6]) ? node33931 : node33928;
														assign node33928 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node33931 = (inp[1]) ? 4'b1001 : 4'b0001;
													assign node33934 = (inp[12]) ? node33940 : node33935;
														assign node33935 = (inp[6]) ? 4'b0001 : node33936;
															assign node33936 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node33940 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node33943 = (inp[12]) ? node33955 : node33944;
													assign node33944 = (inp[11]) ? node33950 : node33945;
														assign node33945 = (inp[6]) ? 4'b0001 : node33946;
															assign node33946 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node33950 = (inp[2]) ? node33952 : 4'b1111;
															assign node33952 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node33955 = (inp[2]) ? 4'b1111 : node33956;
														assign node33956 = (inp[1]) ? node33958 : 4'b0111;
															assign node33958 = (inp[11]) ? node33962 : node33959;
																assign node33959 = (inp[6]) ? 4'b1111 : 4'b0111;
																assign node33962 = (inp[6]) ? 4'b0111 : 4'b1111;
								assign node33966 = (inp[0]) ? node34122 : node33967;
									assign node33967 = (inp[3]) ? node34043 : node33968;
										assign node33968 = (inp[1]) ? node34012 : node33969;
											assign node33969 = (inp[12]) ? node33987 : node33970;
												assign node33970 = (inp[10]) ? node33980 : node33971;
													assign node33971 = (inp[9]) ? node33973 : 4'b1101;
														assign node33973 = (inp[11]) ? node33977 : node33974;
															assign node33974 = (inp[6]) ? 4'b0001 : 4'b1001;
															assign node33977 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node33980 = (inp[11]) ? node33982 : 4'b1001;
														assign node33982 = (inp[6]) ? node33984 : 4'b0101;
															assign node33984 = (inp[9]) ? 4'b1101 : 4'b1001;
												assign node33987 = (inp[9]) ? node33997 : node33988;
													assign node33988 = (inp[11]) ? node33992 : node33989;
														assign node33989 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node33992 = (inp[6]) ? 4'b1001 : node33993;
															assign node33993 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node33997 = (inp[10]) ? node34005 : node33998;
														assign node33998 = (inp[6]) ? node34002 : node33999;
															assign node33999 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node34002 = (inp[11]) ? 4'b1101 : 4'b0001;
														assign node34005 = (inp[11]) ? node34009 : node34006;
															assign node34006 = (inp[6]) ? 4'b0101 : 4'b1101;
															assign node34009 = (inp[6]) ? 4'b1101 : 4'b0101;
											assign node34012 = (inp[9]) ? node34032 : node34013;
												assign node34013 = (inp[12]) ? node34023 : node34014;
													assign node34014 = (inp[6]) ? node34016 : 4'b0101;
														assign node34016 = (inp[11]) ? node34020 : node34017;
															assign node34017 = (inp[10]) ? 4'b1001 : 4'b1101;
															assign node34020 = (inp[2]) ? 4'b0101 : 4'b0001;
													assign node34023 = (inp[11]) ? node34029 : node34024;
														assign node34024 = (inp[6]) ? 4'b1001 : node34025;
															assign node34025 = (inp[10]) ? 4'b0001 : 4'b0101;
														assign node34029 = (inp[6]) ? 4'b0001 : 4'b1001;
												assign node34032 = (inp[11]) ? node34036 : node34033;
													assign node34033 = (inp[10]) ? 4'b0101 : 4'b0001;
													assign node34036 = (inp[6]) ? node34038 : 4'b1101;
														assign node34038 = (inp[12]) ? 4'b0101 : node34039;
															assign node34039 = (inp[10]) ? 4'b0101 : 4'b0001;
										assign node34043 = (inp[9]) ? node34081 : node34044;
											assign node34044 = (inp[10]) ? node34062 : node34045;
												assign node34045 = (inp[1]) ? node34053 : node34046;
													assign node34046 = (inp[11]) ? node34050 : node34047;
														assign node34047 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node34050 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node34053 = (inp[6]) ? node34057 : node34054;
														assign node34054 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node34057 = (inp[12]) ? node34059 : 4'b0101;
															assign node34059 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node34062 = (inp[12]) ? node34072 : node34063;
													assign node34063 = (inp[1]) ? node34065 : 4'b0101;
														assign node34065 = (inp[6]) ? node34069 : node34066;
															assign node34066 = (inp[11]) ? 4'b1001 : 4'b0101;
															assign node34069 = (inp[11]) ? 4'b0001 : 4'b1001;
													assign node34072 = (inp[6]) ? 4'b0001 : node34073;
														assign node34073 = (inp[1]) ? node34077 : node34074;
															assign node34074 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node34077 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node34081 = (inp[12]) ? node34099 : node34082;
												assign node34082 = (inp[1]) ? node34088 : node34083;
													assign node34083 = (inp[11]) ? 4'b0001 : node34084;
														assign node34084 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node34088 = (inp[10]) ? node34094 : node34089;
														assign node34089 = (inp[6]) ? 4'b1001 : node34090;
															assign node34090 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node34094 = (inp[2]) ? 4'b1111 : node34095;
															assign node34095 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node34099 = (inp[10]) ? node34107 : node34100;
													assign node34100 = (inp[6]) ? node34104 : node34101;
														assign node34101 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node34104 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node34107 = (inp[2]) ? node34119 : node34108;
														assign node34108 = (inp[11]) ? node34114 : node34109;
															assign node34109 = (inp[6]) ? 4'b1111 : node34110;
																assign node34110 = (inp[1]) ? 4'b0111 : 4'b1111;
															assign node34114 = (inp[1]) ? 4'b0111 : node34115;
																assign node34115 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node34119 = (inp[11]) ? 4'b1111 : 4'b0111;
									assign node34122 = (inp[3]) ? node34204 : node34123;
										assign node34123 = (inp[6]) ? node34163 : node34124;
											assign node34124 = (inp[10]) ? node34134 : node34125;
												assign node34125 = (inp[9]) ? node34127 : 4'b0111;
													assign node34127 = (inp[11]) ? node34131 : node34128;
														assign node34128 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node34131 = (inp[12]) ? 4'b0011 : 4'b1011;
												assign node34134 = (inp[2]) ? node34150 : node34135;
													assign node34135 = (inp[9]) ? node34145 : node34136;
														assign node34136 = (inp[12]) ? node34140 : node34137;
															assign node34137 = (inp[11]) ? 4'b1011 : 4'b0111;
															assign node34140 = (inp[11]) ? 4'b0011 : node34141;
																assign node34141 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node34145 = (inp[12]) ? node34147 : 4'b0011;
															assign node34147 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node34150 = (inp[11]) ? node34154 : node34151;
														assign node34151 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node34154 = (inp[1]) ? node34160 : node34155;
															assign node34155 = (inp[12]) ? 4'b0111 : node34156;
																assign node34156 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node34160 = (inp[9]) ? 4'b1111 : 4'b1011;
											assign node34163 = (inp[10]) ? node34189 : node34164;
												assign node34164 = (inp[9]) ? node34180 : node34165;
													assign node34165 = (inp[12]) ? node34173 : node34166;
														assign node34166 = (inp[1]) ? node34170 : node34167;
															assign node34167 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node34170 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node34173 = (inp[11]) ? node34177 : node34174;
															assign node34174 = (inp[1]) ? 4'b1011 : 4'b0111;
															assign node34177 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node34180 = (inp[12]) ? node34184 : node34181;
														assign node34181 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node34184 = (inp[11]) ? node34186 : 4'b0011;
															assign node34186 = (inp[2]) ? 4'b0111 : 4'b1111;
												assign node34189 = (inp[9]) ? node34197 : node34190;
													assign node34190 = (inp[11]) ? node34194 : node34191;
														assign node34191 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node34194 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node34197 = (inp[1]) ? node34201 : node34198;
														assign node34198 = (inp[11]) ? 4'b1111 : 4'b0011;
														assign node34201 = (inp[11]) ? 4'b0111 : 4'b1111;
										assign node34204 = (inp[9]) ? node34256 : node34205;
											assign node34205 = (inp[10]) ? node34227 : node34206;
												assign node34206 = (inp[6]) ? node34222 : node34207;
													assign node34207 = (inp[2]) ? node34213 : node34208;
														assign node34208 = (inp[11]) ? 4'b0111 : node34209;
															assign node34209 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node34213 = (inp[12]) ? node34217 : node34214;
															assign node34214 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node34217 = (inp[1]) ? 4'b1011 : node34218;
																assign node34218 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node34222 = (inp[12]) ? 4'b1011 : node34223;
														assign node34223 = (inp[11]) ? 4'b1111 : 4'b0111;
												assign node34227 = (inp[12]) ? node34235 : node34228;
													assign node34228 = (inp[1]) ? node34230 : 4'b0111;
														assign node34230 = (inp[11]) ? node34232 : 4'b1011;
															assign node34232 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node34235 = (inp[2]) ? node34243 : node34236;
														assign node34236 = (inp[1]) ? 4'b0011 : node34237;
															assign node34237 = (inp[6]) ? node34239 : 4'b0011;
																assign node34239 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node34243 = (inp[1]) ? node34249 : node34244;
															assign node34244 = (inp[11]) ? node34246 : 4'b1011;
																assign node34246 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node34249 = (inp[11]) ? node34253 : node34250;
																assign node34250 = (inp[6]) ? 4'b1011 : 4'b0011;
																assign node34253 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node34256 = (inp[1]) ? node34262 : node34257;
												assign node34257 = (inp[6]) ? 4'b0011 : node34258;
													assign node34258 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node34262 = (inp[11]) ? node34268 : node34263;
													assign node34263 = (inp[6]) ? node34265 : 4'b0011;
														assign node34265 = (inp[2]) ? 4'b1011 : 4'b1101;
													assign node34268 = (inp[6]) ? 4'b0101 : 4'b1101;
							assign node34271 = (inp[9]) ? node34653 : node34272;
								assign node34272 = (inp[12]) ? node34452 : node34273;
									assign node34273 = (inp[10]) ? node34385 : node34274;
										assign node34274 = (inp[1]) ? node34332 : node34275;
											assign node34275 = (inp[6]) ? node34299 : node34276;
												assign node34276 = (inp[11]) ? node34288 : node34277;
													assign node34277 = (inp[2]) ? node34283 : node34278;
														assign node34278 = (inp[0]) ? node34280 : 4'b1101;
															assign node34280 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node34283 = (inp[15]) ? node34285 : 4'b1111;
															assign node34285 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node34288 = (inp[2]) ? node34292 : node34289;
														assign node34289 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node34292 = (inp[0]) ? 4'b0111 : node34293;
															assign node34293 = (inp[15]) ? 4'b0101 : node34294;
																assign node34294 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node34299 = (inp[11]) ? node34311 : node34300;
													assign node34300 = (inp[3]) ? node34306 : node34301;
														assign node34301 = (inp[2]) ? 4'b0111 : node34302;
															assign node34302 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node34306 = (inp[0]) ? node34308 : 4'b0101;
															assign node34308 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node34311 = (inp[2]) ? node34319 : node34312;
														assign node34312 = (inp[3]) ? node34314 : 4'b1111;
															assign node34314 = (inp[15]) ? 4'b1111 : node34315;
																assign node34315 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node34319 = (inp[3]) ? node34327 : node34320;
															assign node34320 = (inp[15]) ? node34324 : node34321;
																assign node34321 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node34324 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node34327 = (inp[15]) ? node34329 : 4'b1101;
																assign node34329 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node34332 = (inp[11]) ? node34364 : node34333;
												assign node34333 = (inp[6]) ? node34357 : node34334;
													assign node34334 = (inp[15]) ? node34344 : node34335;
														assign node34335 = (inp[2]) ? node34337 : 4'b0101;
															assign node34337 = (inp[3]) ? node34341 : node34338;
																assign node34338 = (inp[0]) ? 4'b0101 : 4'b0111;
																assign node34341 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node34344 = (inp[2]) ? node34350 : node34345;
															assign node34345 = (inp[0]) ? 4'b0111 : node34346;
																assign node34346 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node34350 = (inp[3]) ? node34354 : node34351;
																assign node34351 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node34354 = (inp[0]) ? 4'b0101 : 4'b0111;
													assign node34357 = (inp[3]) ? 4'b1101 : node34358;
														assign node34358 = (inp[15]) ? 4'b1111 : node34359;
															assign node34359 = (inp[2]) ? 4'b1101 : 4'b1111;
												assign node34364 = (inp[6]) ? node34376 : node34365;
													assign node34365 = (inp[2]) ? node34371 : node34366;
														assign node34366 = (inp[15]) ? 4'b1101 : node34367;
															assign node34367 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node34371 = (inp[15]) ? 4'b1111 : node34372;
															assign node34372 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node34376 = (inp[3]) ? 4'b0101 : node34377;
														assign node34377 = (inp[2]) ? 4'b0101 : node34378;
															assign node34378 = (inp[15]) ? 4'b0111 : node34379;
																assign node34379 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node34385 = (inp[1]) ? node34413 : node34386;
											assign node34386 = (inp[6]) ? node34402 : node34387;
												assign node34387 = (inp[11]) ? node34393 : node34388;
													assign node34388 = (inp[2]) ? node34390 : 4'b1101;
														assign node34390 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node34393 = (inp[3]) ? 4'b0101 : node34394;
														assign node34394 = (inp[15]) ? node34398 : node34395;
															assign node34395 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node34398 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node34402 = (inp[11]) ? 4'b1001 : node34403;
													assign node34403 = (inp[2]) ? node34405 : 4'b0101;
														assign node34405 = (inp[0]) ? node34407 : 4'b0101;
															assign node34407 = (inp[15]) ? 4'b0111 : node34408;
																assign node34408 = (inp[3]) ? 4'b0111 : 4'b0101;
											assign node34413 = (inp[11]) ? node34437 : node34414;
												assign node34414 = (inp[6]) ? node34430 : node34415;
													assign node34415 = (inp[3]) ? node34423 : node34416;
														assign node34416 = (inp[0]) ? node34420 : node34417;
															assign node34417 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node34420 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node34423 = (inp[0]) ? node34427 : node34424;
															assign node34424 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node34427 = (inp[2]) ? 4'b0101 : 4'b0111;
													assign node34430 = (inp[15]) ? node34432 : 4'b1011;
														assign node34432 = (inp[0]) ? 4'b1011 : node34433;
															assign node34433 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node34437 = (inp[6]) ? node34445 : node34438;
													assign node34438 = (inp[15]) ? 4'b1011 : node34439;
														assign node34439 = (inp[0]) ? 4'b1001 : node34440;
															assign node34440 = (inp[3]) ? 4'b1001 : 4'b1011;
													assign node34445 = (inp[0]) ? 4'b0001 : node34446;
														assign node34446 = (inp[3]) ? node34448 : 4'b0011;
															assign node34448 = (inp[15]) ? 4'b0011 : 4'b0001;
									assign node34452 = (inp[10]) ? node34542 : node34453;
										assign node34453 = (inp[6]) ? node34493 : node34454;
											assign node34454 = (inp[11]) ? node34478 : node34455;
												assign node34455 = (inp[1]) ? node34469 : node34456;
													assign node34456 = (inp[3]) ? node34462 : node34457;
														assign node34457 = (inp[0]) ? node34459 : 4'b1101;
															assign node34459 = (inp[2]) ? 4'b1101 : 4'b1111;
														assign node34462 = (inp[0]) ? node34466 : node34463;
															assign node34463 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node34466 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node34469 = (inp[0]) ? 4'b0111 : node34470;
														assign node34470 = (inp[15]) ? node34474 : node34471;
															assign node34471 = (inp[2]) ? 4'b0111 : 4'b0101;
															assign node34474 = (inp[3]) ? 4'b0111 : 4'b0101;
												assign node34478 = (inp[1]) ? node34486 : node34479;
													assign node34479 = (inp[15]) ? node34481 : 4'b0111;
														assign node34481 = (inp[3]) ? 4'b0101 : node34482;
															assign node34482 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node34486 = (inp[2]) ? node34488 : 4'b1001;
														assign node34488 = (inp[3]) ? 4'b1001 : node34489;
															assign node34489 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node34493 = (inp[1]) ? node34515 : node34494;
												assign node34494 = (inp[11]) ? node34502 : node34495;
													assign node34495 = (inp[0]) ? 4'b0111 : node34496;
														assign node34496 = (inp[3]) ? 4'b0101 : node34497;
															assign node34497 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node34502 = (inp[0]) ? node34510 : node34503;
														assign node34503 = (inp[2]) ? node34507 : node34504;
															assign node34504 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node34507 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node34510 = (inp[15]) ? node34512 : 4'b1001;
															assign node34512 = (inp[2]) ? 4'b1001 : 4'b1011;
												assign node34515 = (inp[11]) ? node34529 : node34516;
													assign node34516 = (inp[3]) ? node34522 : node34517;
														assign node34517 = (inp[15]) ? 4'b1011 : node34518;
															assign node34518 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node34522 = (inp[15]) ? node34526 : node34523;
															assign node34523 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node34526 = (inp[0]) ? 4'b1001 : 4'b1011;
													assign node34529 = (inp[0]) ? node34535 : node34530;
														assign node34530 = (inp[2]) ? 4'b0011 : node34531;
															assign node34531 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node34535 = (inp[3]) ? node34539 : node34536;
															assign node34536 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node34539 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node34542 = (inp[15]) ? node34600 : node34543;
											assign node34543 = (inp[11]) ? node34575 : node34544;
												assign node34544 = (inp[1]) ? node34562 : node34545;
													assign node34545 = (inp[6]) ? node34555 : node34546;
														assign node34546 = (inp[2]) ? node34548 : 4'b1001;
															assign node34548 = (inp[0]) ? node34552 : node34549;
																assign node34549 = (inp[3]) ? 4'b1001 : 4'b1011;
																assign node34552 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node34555 = (inp[3]) ? node34559 : node34556;
															assign node34556 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node34559 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node34562 = (inp[6]) ? node34568 : node34563;
														assign node34563 = (inp[2]) ? node34565 : 4'b0001;
															assign node34565 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node34568 = (inp[0]) ? node34572 : node34569;
															assign node34569 = (inp[3]) ? 4'b1001 : 4'b1011;
															assign node34572 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node34575 = (inp[2]) ? node34581 : node34576;
													assign node34576 = (inp[1]) ? 4'b1011 : node34577;
														assign node34577 = (inp[6]) ? 4'b1011 : 4'b0001;
													assign node34581 = (inp[6]) ? node34589 : node34582;
														assign node34582 = (inp[1]) ? 4'b1011 : node34583;
															assign node34583 = (inp[0]) ? 4'b0011 : node34584;
																assign node34584 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node34589 = (inp[1]) ? node34595 : node34590;
															assign node34590 = (inp[3]) ? node34592 : 4'b1001;
																assign node34592 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node34595 = (inp[0]) ? 4'b0001 : node34596;
																assign node34596 = (inp[3]) ? 4'b0001 : 4'b0011;
											assign node34600 = (inp[2]) ? node34624 : node34601;
												assign node34601 = (inp[0]) ? node34611 : node34602;
													assign node34602 = (inp[3]) ? node34604 : 4'b0001;
														assign node34604 = (inp[11]) ? 4'b0011 : node34605;
															assign node34605 = (inp[6]) ? node34607 : 4'b0011;
																assign node34607 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node34611 = (inp[3]) ? node34617 : node34612;
														assign node34612 = (inp[11]) ? 4'b1011 : node34613;
															assign node34613 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node34617 = (inp[6]) ? 4'b0001 : node34618;
															assign node34618 = (inp[1]) ? node34620 : 4'b0001;
																assign node34620 = (inp[11]) ? 4'b1001 : 4'b0001;
												assign node34624 = (inp[11]) ? node34636 : node34625;
													assign node34625 = (inp[0]) ? node34631 : node34626;
														assign node34626 = (inp[6]) ? 4'b1001 : node34627;
															assign node34627 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node34631 = (inp[3]) ? node34633 : 4'b0011;
															assign node34633 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node34636 = (inp[1]) ? node34646 : node34637;
														assign node34637 = (inp[6]) ? node34643 : node34638;
															assign node34638 = (inp[0]) ? 4'b0001 : node34639;
																assign node34639 = (inp[3]) ? 4'b0011 : 4'b0001;
															assign node34643 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node34646 = (inp[6]) ? 4'b0011 : node34647;
															assign node34647 = (inp[0]) ? 4'b1011 : node34648;
																assign node34648 = (inp[3]) ? 4'b1011 : 4'b1001;
								assign node34653 = (inp[10]) ? node34851 : node34654;
									assign node34654 = (inp[12]) ? node34754 : node34655;
										assign node34655 = (inp[3]) ? node34715 : node34656;
											assign node34656 = (inp[11]) ? node34694 : node34657;
												assign node34657 = (inp[2]) ? node34671 : node34658;
													assign node34658 = (inp[1]) ? node34664 : node34659;
														assign node34659 = (inp[6]) ? node34661 : 4'b1001;
															assign node34661 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node34664 = (inp[6]) ? node34666 : 4'b0011;
															assign node34666 = (inp[0]) ? node34668 : 4'b1011;
																assign node34668 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node34671 = (inp[1]) ? node34685 : node34672;
														assign node34672 = (inp[6]) ? node34680 : node34673;
															assign node34673 = (inp[0]) ? node34677 : node34674;
																assign node34674 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node34677 = (inp[15]) ? 4'b1011 : 4'b1001;
															assign node34680 = (inp[0]) ? node34682 : 4'b0001;
																assign node34682 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34685 = (inp[6]) ? 4'b1001 : node34686;
															assign node34686 = (inp[15]) ? node34690 : node34687;
																assign node34687 = (inp[0]) ? 4'b0001 : 4'b0011;
																assign node34690 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node34694 = (inp[0]) ? node34704 : node34695;
													assign node34695 = (inp[15]) ? node34697 : 4'b0011;
														assign node34697 = (inp[1]) ? node34701 : node34698;
															assign node34698 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node34701 = (inp[2]) ? 4'b0001 : 4'b1001;
													assign node34704 = (inp[15]) ? node34710 : node34705;
														assign node34705 = (inp[6]) ? node34707 : 4'b0001;
															assign node34707 = (inp[1]) ? 4'b0001 : 4'b1001;
														assign node34710 = (inp[6]) ? 4'b0011 : node34711;
															assign node34711 = (inp[1]) ? 4'b1011 : 4'b0011;
											assign node34715 = (inp[11]) ? node34733 : node34716;
												assign node34716 = (inp[15]) ? node34724 : node34717;
													assign node34717 = (inp[0]) ? 4'b0011 : node34718;
														assign node34718 = (inp[2]) ? 4'b0001 : node34719;
															assign node34719 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node34724 = (inp[0]) ? 4'b0001 : node34725;
														assign node34725 = (inp[2]) ? 4'b1011 : node34726;
															assign node34726 = (inp[6]) ? node34728 : 4'b0011;
																assign node34728 = (inp[1]) ? 4'b1011 : 4'b0011;
												assign node34733 = (inp[15]) ? node34743 : node34734;
													assign node34734 = (inp[0]) ? node34736 : 4'b1001;
														assign node34736 = (inp[1]) ? node34740 : node34737;
															assign node34737 = (inp[6]) ? 4'b1011 : 4'b0011;
															assign node34740 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node34743 = (inp[0]) ? node34751 : node34744;
														assign node34744 = (inp[6]) ? node34748 : node34745;
															assign node34745 = (inp[2]) ? 4'b0011 : 4'b1011;
															assign node34748 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node34751 = (inp[1]) ? 4'b0001 : 4'b1001;
										assign node34754 = (inp[6]) ? node34804 : node34755;
											assign node34755 = (inp[1]) ? node34779 : node34756;
												assign node34756 = (inp[11]) ? node34760 : node34757;
													assign node34757 = (inp[2]) ? 4'b1001 : 4'b1011;
													assign node34760 = (inp[2]) ? node34774 : node34761;
														assign node34761 = (inp[0]) ? node34767 : node34762;
															assign node34762 = (inp[3]) ? node34764 : 4'b0001;
																assign node34764 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node34767 = (inp[3]) ? node34771 : node34768;
																assign node34768 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node34771 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node34774 = (inp[3]) ? 4'b0011 : node34775;
															assign node34775 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node34779 = (inp[11]) ? node34793 : node34780;
													assign node34780 = (inp[0]) ? node34788 : node34781;
														assign node34781 = (inp[3]) ? node34785 : node34782;
															assign node34782 = (inp[15]) ? 4'b0001 : 4'b0011;
															assign node34785 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34788 = (inp[15]) ? 4'b0001 : node34789;
															assign node34789 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node34793 = (inp[3]) ? node34799 : node34794;
														assign node34794 = (inp[15]) ? node34796 : 4'b1101;
															assign node34796 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node34799 = (inp[15]) ? 4'b1101 : node34800;
															assign node34800 = (inp[0]) ? 4'b1111 : 4'b1101;
											assign node34804 = (inp[1]) ? node34836 : node34805;
												assign node34805 = (inp[11]) ? node34823 : node34806;
													assign node34806 = (inp[0]) ? node34814 : node34807;
														assign node34807 = (inp[2]) ? 4'b0011 : node34808;
															assign node34808 = (inp[3]) ? node34810 : 4'b0001;
																assign node34810 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34814 = (inp[2]) ? node34818 : node34815;
															assign node34815 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node34818 = (inp[15]) ? 4'b0001 : node34819;
																assign node34819 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node34823 = (inp[2]) ? node34831 : node34824;
														assign node34824 = (inp[3]) ? 4'b1101 : node34825;
															assign node34825 = (inp[0]) ? 4'b1111 : node34826;
																assign node34826 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node34831 = (inp[15]) ? 4'b1111 : node34832;
															assign node34832 = (inp[0]) ? 4'b1111 : 4'b1101;
												assign node34836 = (inp[11]) ? node34844 : node34837;
													assign node34837 = (inp[0]) ? node34841 : node34838;
														assign node34838 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node34841 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node34844 = (inp[0]) ? node34848 : node34845;
														assign node34845 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node34848 = (inp[15]) ? 4'b0101 : 4'b0111;
									assign node34851 = (inp[12]) ? node34929 : node34852;
										assign node34852 = (inp[6]) ? node34896 : node34853;
											assign node34853 = (inp[1]) ? node34875 : node34854;
												assign node34854 = (inp[11]) ? node34862 : node34855;
													assign node34855 = (inp[0]) ? 4'b1001 : node34856;
														assign node34856 = (inp[3]) ? node34858 : 4'b1011;
															assign node34858 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node34862 = (inp[0]) ? node34870 : node34863;
														assign node34863 = (inp[15]) ? node34867 : node34864;
															assign node34864 = (inp[3]) ? 4'b0001 : 4'b0011;
															assign node34867 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node34870 = (inp[2]) ? node34872 : 4'b0001;
															assign node34872 = (inp[15]) ? 4'b0011 : 4'b0001;
												assign node34875 = (inp[11]) ? node34887 : node34876;
													assign node34876 = (inp[3]) ? node34882 : node34877;
														assign node34877 = (inp[2]) ? 4'b0001 : node34878;
															assign node34878 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node34882 = (inp[0]) ? node34884 : 4'b0011;
															assign node34884 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node34887 = (inp[3]) ? node34893 : node34888;
														assign node34888 = (inp[15]) ? 4'b1111 : node34889;
															assign node34889 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node34893 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node34896 = (inp[1]) ? node34908 : node34897;
												assign node34897 = (inp[11]) ? node34903 : node34898;
													assign node34898 = (inp[0]) ? node34900 : 4'b0001;
														assign node34900 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node34903 = (inp[0]) ? 4'b1101 : node34904;
														assign node34904 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node34908 = (inp[11]) ? node34924 : node34909;
													assign node34909 = (inp[3]) ? node34915 : node34910;
														assign node34910 = (inp[0]) ? node34912 : 4'b1101;
															assign node34912 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node34915 = (inp[2]) ? node34919 : node34916;
															assign node34916 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node34919 = (inp[15]) ? node34921 : 4'b1101;
																assign node34921 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node34924 = (inp[0]) ? node34926 : 4'b0111;
														assign node34926 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node34929 = (inp[6]) ? node34963 : node34930;
											assign node34930 = (inp[0]) ? node34948 : node34931;
												assign node34931 = (inp[15]) ? node34939 : node34932;
													assign node34932 = (inp[1]) ? node34936 : node34933;
														assign node34933 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node34936 = (inp[3]) ? 4'b0101 : 4'b1101;
													assign node34939 = (inp[2]) ? node34945 : node34940;
														assign node34940 = (inp[3]) ? 4'b1111 : node34941;
															assign node34941 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node34945 = (inp[3]) ? 4'b0111 : 4'b1111;
												assign node34948 = (inp[15]) ? node34956 : node34949;
													assign node34949 = (inp[11]) ? node34953 : node34950;
														assign node34950 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node34953 = (inp[1]) ? 4'b1111 : 4'b0111;
													assign node34956 = (inp[2]) ? node34958 : 4'b0101;
														assign node34958 = (inp[11]) ? node34960 : 4'b0101;
															assign node34960 = (inp[1]) ? 4'b1101 : 4'b0101;
											assign node34963 = (inp[3]) ? node35005 : node34964;
												assign node34964 = (inp[1]) ? node34976 : node34965;
													assign node34965 = (inp[11]) ? node34971 : node34966;
														assign node34966 = (inp[0]) ? 4'b0111 : node34967;
															assign node34967 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node34971 = (inp[0]) ? node34973 : 4'b1111;
															assign node34973 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node34976 = (inp[11]) ? node34990 : node34977;
														assign node34977 = (inp[2]) ? node34983 : node34978;
															assign node34978 = (inp[0]) ? node34980 : 4'b1111;
																assign node34980 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node34983 = (inp[15]) ? node34987 : node34984;
																assign node34984 = (inp[0]) ? 4'b1111 : 4'b1101;
																assign node34987 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node34990 = (inp[2]) ? node34998 : node34991;
															assign node34991 = (inp[0]) ? node34995 : node34992;
																assign node34992 = (inp[15]) ? 4'b0111 : 4'b0101;
																assign node34995 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node34998 = (inp[15]) ? node35002 : node34999;
																assign node34999 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node35002 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node35005 = (inp[15]) ? node35023 : node35006;
													assign node35006 = (inp[0]) ? node35014 : node35007;
														assign node35007 = (inp[1]) ? node35011 : node35008;
															assign node35008 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node35011 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node35014 = (inp[2]) ? 4'b0111 : node35015;
															assign node35015 = (inp[1]) ? node35019 : node35016;
																assign node35016 = (inp[11]) ? 4'b1111 : 4'b0111;
																assign node35019 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node35023 = (inp[0]) ? node35025 : 4'b0111;
														assign node35025 = (inp[1]) ? 4'b0101 : 4'b1101;
						assign node35028 = (inp[15]) ? node35752 : node35029;
							assign node35029 = (inp[0]) ? node35431 : node35030;
								assign node35030 = (inp[3]) ? node35224 : node35031;
									assign node35031 = (inp[5]) ? node35125 : node35032;
										assign node35032 = (inp[10]) ? node35082 : node35033;
											assign node35033 = (inp[9]) ? node35055 : node35034;
												assign node35034 = (inp[12]) ? node35046 : node35035;
													assign node35035 = (inp[11]) ? node35041 : node35036;
														assign node35036 = (inp[2]) ? 4'b1011 : node35037;
															assign node35037 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node35041 = (inp[6]) ? node35043 : 4'b0011;
															assign node35043 = (inp[1]) ? 4'b0011 : 4'b1011;
													assign node35046 = (inp[11]) ? node35048 : 4'b0011;
														assign node35048 = (inp[2]) ? 4'b1111 : node35049;
															assign node35049 = (inp[1]) ? node35051 : 4'b0011;
																assign node35051 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node35055 = (inp[12]) ? node35071 : node35056;
													assign node35056 = (inp[11]) ? node35066 : node35057;
														assign node35057 = (inp[2]) ? node35061 : node35058;
															assign node35058 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node35061 = (inp[1]) ? node35063 : 4'b1111;
																assign node35063 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node35066 = (inp[1]) ? node35068 : 4'b1111;
															assign node35068 = (inp[2]) ? 4'b0111 : 4'b1111;
													assign node35071 = (inp[1]) ? node35077 : node35072;
														assign node35072 = (inp[11]) ? 4'b0111 : node35073;
															assign node35073 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node35077 = (inp[11]) ? node35079 : 4'b1011;
															assign node35079 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node35082 = (inp[9]) ? node35102 : node35083;
												assign node35083 = (inp[12]) ? node35089 : node35084;
													assign node35084 = (inp[11]) ? node35086 : 4'b0011;
														assign node35086 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node35089 = (inp[1]) ? node35095 : node35090;
														assign node35090 = (inp[6]) ? 4'b0111 : node35091;
															assign node35091 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node35095 = (inp[6]) ? node35099 : node35096;
															assign node35096 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node35099 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node35102 = (inp[12]) ? node35114 : node35103;
													assign node35103 = (inp[11]) ? node35109 : node35104;
														assign node35104 = (inp[1]) ? 4'b0111 : node35105;
															assign node35105 = (inp[2]) ? 4'b1111 : 4'b0111;
														assign node35109 = (inp[6]) ? 4'b1011 : node35110;
															assign node35110 = (inp[1]) ? 4'b1011 : 4'b0111;
													assign node35114 = (inp[6]) ? node35120 : node35115;
														assign node35115 = (inp[11]) ? 4'b0011 : node35116;
															assign node35116 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node35120 = (inp[1]) ? node35122 : 4'b1011;
															assign node35122 = (inp[11]) ? 4'b0011 : 4'b1011;
										assign node35125 = (inp[9]) ? node35173 : node35126;
											assign node35126 = (inp[10]) ? node35154 : node35127;
												assign node35127 = (inp[12]) ? node35141 : node35128;
													assign node35128 = (inp[11]) ? node35136 : node35129;
														assign node35129 = (inp[6]) ? node35133 : node35130;
															assign node35130 = (inp[1]) ? 4'b0011 : 4'b1011;
															assign node35133 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node35136 = (inp[1]) ? 4'b1011 : node35137;
															assign node35137 = (inp[2]) ? 4'b0011 : 4'b1011;
													assign node35141 = (inp[6]) ? node35149 : node35142;
														assign node35142 = (inp[1]) ? node35146 : node35143;
															assign node35143 = (inp[11]) ? 4'b0011 : 4'b1011;
															assign node35146 = (inp[11]) ? 4'b1101 : 4'b0011;
														assign node35149 = (inp[1]) ? node35151 : 4'b1101;
															assign node35151 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node35154 = (inp[6]) ? node35168 : node35155;
													assign node35155 = (inp[12]) ? node35163 : node35156;
														assign node35156 = (inp[11]) ? node35160 : node35157;
															assign node35157 = (inp[1]) ? 4'b0011 : 4'b1011;
															assign node35160 = (inp[1]) ? 4'b1101 : 4'b0011;
														assign node35163 = (inp[2]) ? node35165 : 4'b0101;
															assign node35165 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node35168 = (inp[11]) ? node35170 : 4'b1101;
														assign node35170 = (inp[1]) ? 4'b0101 : 4'b1101;
											assign node35173 = (inp[12]) ? node35199 : node35174;
												assign node35174 = (inp[6]) ? node35188 : node35175;
													assign node35175 = (inp[2]) ? node35183 : node35176;
														assign node35176 = (inp[11]) ? node35180 : node35177;
															assign node35177 = (inp[1]) ? 4'b0101 : 4'b1101;
															assign node35180 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node35183 = (inp[11]) ? 4'b0101 : node35184;
															assign node35184 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node35188 = (inp[10]) ? node35196 : node35189;
														assign node35189 = (inp[11]) ? node35193 : node35190;
															assign node35190 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node35193 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node35196 = (inp[1]) ? 4'b0001 : 4'b0101;
												assign node35199 = (inp[10]) ? node35207 : node35200;
													assign node35200 = (inp[6]) ? node35202 : 4'b0101;
														assign node35202 = (inp[11]) ? node35204 : 4'b1001;
															assign node35204 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node35207 = (inp[6]) ? node35219 : node35208;
														assign node35208 = (inp[2]) ? node35214 : node35209;
															assign node35209 = (inp[1]) ? node35211 : 4'b0001;
																assign node35211 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node35214 = (inp[1]) ? 4'b1001 : node35215;
																assign node35215 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node35219 = (inp[2]) ? 4'b0001 : node35220;
															assign node35220 = (inp[1]) ? 4'b0001 : 4'b1001;
									assign node35224 = (inp[5]) ? node35320 : node35225;
										assign node35225 = (inp[9]) ? node35281 : node35226;
											assign node35226 = (inp[12]) ? node35252 : node35227;
												assign node35227 = (inp[10]) ? node35243 : node35228;
													assign node35228 = (inp[6]) ? node35238 : node35229;
														assign node35229 = (inp[2]) ? node35233 : node35230;
															assign node35230 = (inp[1]) ? 4'b1011 : 4'b0011;
															assign node35233 = (inp[1]) ? node35235 : 4'b1011;
																assign node35235 = (inp[11]) ? 4'b1011 : 4'b0011;
														assign node35238 = (inp[11]) ? 4'b0011 : node35239;
															assign node35239 = (inp[2]) ? 4'b0011 : 4'b1011;
													assign node35243 = (inp[1]) ? node35249 : node35244;
														assign node35244 = (inp[11]) ? 4'b1101 : node35245;
															assign node35245 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node35249 = (inp[2]) ? 4'b1101 : 4'b0101;
												assign node35252 = (inp[10]) ? node35264 : node35253;
													assign node35253 = (inp[6]) ? node35259 : node35254;
														assign node35254 = (inp[1]) ? 4'b1101 : node35255;
															assign node35255 = (inp[2]) ? 4'b0011 : 4'b1011;
														assign node35259 = (inp[11]) ? node35261 : 4'b1101;
															assign node35261 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node35264 = (inp[11]) ? node35272 : node35265;
														assign node35265 = (inp[6]) ? node35269 : node35266;
															assign node35266 = (inp[1]) ? 4'b0101 : 4'b1101;
															assign node35269 = (inp[1]) ? 4'b1101 : 4'b0101;
														assign node35272 = (inp[2]) ? node35274 : 4'b0101;
															assign node35274 = (inp[1]) ? node35278 : node35275;
																assign node35275 = (inp[6]) ? 4'b1101 : 4'b0101;
																assign node35278 = (inp[6]) ? 4'b0101 : 4'b1101;
											assign node35281 = (inp[10]) ? node35299 : node35282;
												assign node35282 = (inp[11]) ? node35288 : node35283;
													assign node35283 = (inp[6]) ? 4'b0101 : node35284;
														assign node35284 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node35288 = (inp[2]) ? node35294 : node35289;
														assign node35289 = (inp[1]) ? node35291 : 4'b0101;
															assign node35291 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node35294 = (inp[1]) ? 4'b1001 : node35295;
															assign node35295 = (inp[6]) ? 4'b1101 : 4'b0101;
												assign node35299 = (inp[12]) ? node35311 : node35300;
													assign node35300 = (inp[1]) ? node35306 : node35301;
														assign node35301 = (inp[2]) ? node35303 : 4'b0101;
															assign node35303 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node35306 = (inp[2]) ? node35308 : 4'b1001;
															assign node35308 = (inp[6]) ? 4'b1001 : 4'b0101;
													assign node35311 = (inp[1]) ? 4'b0001 : node35312;
														assign node35312 = (inp[11]) ? node35316 : node35313;
															assign node35313 = (inp[6]) ? 4'b0001 : 4'b1001;
															assign node35316 = (inp[6]) ? 4'b1001 : 4'b0001;
										assign node35320 = (inp[2]) ? node35380 : node35321;
											assign node35321 = (inp[1]) ? node35347 : node35322;
												assign node35322 = (inp[12]) ? node35336 : node35323;
													assign node35323 = (inp[9]) ? node35329 : node35324;
														assign node35324 = (inp[11]) ? 4'b1101 : node35325;
															assign node35325 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node35329 = (inp[6]) ? node35333 : node35330;
															assign node35330 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node35333 = (inp[11]) ? 4'b1001 : 4'b0101;
													assign node35336 = (inp[9]) ? node35344 : node35337;
														assign node35337 = (inp[6]) ? node35341 : node35338;
															assign node35338 = (inp[10]) ? 4'b1101 : 4'b1001;
															assign node35341 = (inp[10]) ? 4'b0101 : 4'b1101;
														assign node35344 = (inp[10]) ? 4'b1001 : 4'b1101;
												assign node35347 = (inp[9]) ? node35369 : node35348;
													assign node35348 = (inp[10]) ? node35362 : node35349;
														assign node35349 = (inp[12]) ? node35357 : node35350;
															assign node35350 = (inp[11]) ? node35354 : node35351;
																assign node35351 = (inp[6]) ? 4'b1001 : 4'b0001;
																assign node35354 = (inp[6]) ? 4'b0001 : 4'b1001;
															assign node35357 = (inp[11]) ? 4'b1101 : node35358;
																assign node35358 = (inp[6]) ? 4'b1101 : 4'b0001;
														assign node35362 = (inp[12]) ? node35364 : 4'b1101;
															assign node35364 = (inp[11]) ? 4'b0101 : node35365;
																assign node35365 = (inp[6]) ? 4'b1101 : 4'b0101;
													assign node35369 = (inp[10]) ? node35375 : node35370;
														assign node35370 = (inp[6]) ? 4'b1001 : node35371;
															assign node35371 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node35375 = (inp[6]) ? node35377 : 4'b1001;
															assign node35377 = (inp[11]) ? 4'b0001 : 4'b1001;
											assign node35380 = (inp[12]) ? node35412 : node35381;
												assign node35381 = (inp[1]) ? node35393 : node35382;
													assign node35382 = (inp[6]) ? node35386 : node35383;
														assign node35383 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node35386 = (inp[11]) ? node35388 : 4'b0101;
															assign node35388 = (inp[10]) ? node35390 : 4'b1001;
																assign node35390 = (inp[9]) ? 4'b1001 : 4'b1101;
													assign node35393 = (inp[6]) ? node35401 : node35394;
														assign node35394 = (inp[9]) ? node35398 : node35395;
															assign node35395 = (inp[10]) ? 4'b1101 : 4'b1001;
															assign node35398 = (inp[10]) ? 4'b1001 : 4'b1101;
														assign node35401 = (inp[11]) ? node35409 : node35402;
															assign node35402 = (inp[10]) ? node35406 : node35403;
																assign node35403 = (inp[9]) ? 4'b1101 : 4'b1001;
																assign node35406 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node35409 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node35412 = (inp[9]) ? node35420 : node35413;
													assign node35413 = (inp[10]) ? node35417 : node35414;
														assign node35414 = (inp[11]) ? 4'b0101 : 4'b0001;
														assign node35417 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node35420 = (inp[1]) ? node35424 : node35421;
														assign node35421 = (inp[11]) ? 4'b0101 : 4'b0001;
														assign node35424 = (inp[10]) ? 4'b0001 : node35425;
															assign node35425 = (inp[6]) ? node35427 : 4'b1001;
																assign node35427 = (inp[11]) ? 4'b0001 : 4'b1001;
								assign node35431 = (inp[3]) ? node35581 : node35432;
									assign node35432 = (inp[5]) ? node35494 : node35433;
										assign node35433 = (inp[6]) ? node35461 : node35434;
											assign node35434 = (inp[1]) ? node35448 : node35435;
												assign node35435 = (inp[11]) ? node35441 : node35436;
													assign node35436 = (inp[10]) ? 4'b1101 : node35437;
														assign node35437 = (inp[9]) ? 4'b1101 : 4'b1001;
													assign node35441 = (inp[2]) ? 4'b0101 : node35442;
														assign node35442 = (inp[9]) ? node35444 : 4'b0101;
															assign node35444 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node35448 = (inp[11]) ? node35452 : node35449;
													assign node35449 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node35452 = (inp[9]) ? node35456 : node35453;
														assign node35453 = (inp[12]) ? 4'b1101 : 4'b1001;
														assign node35456 = (inp[12]) ? 4'b1001 : node35457;
															assign node35457 = (inp[10]) ? 4'b1001 : 4'b1101;
											assign node35461 = (inp[9]) ? node35481 : node35462;
												assign node35462 = (inp[11]) ? node35474 : node35463;
													assign node35463 = (inp[1]) ? node35469 : node35464;
														assign node35464 = (inp[10]) ? node35466 : 4'b0001;
															assign node35466 = (inp[12]) ? 4'b0101 : 4'b0001;
														assign node35469 = (inp[12]) ? 4'b1101 : node35470;
															assign node35470 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node35474 = (inp[1]) ? node35476 : 4'b1101;
														assign node35476 = (inp[10]) ? 4'b0101 : node35477;
															assign node35477 = (inp[12]) ? 4'b0101 : 4'b0001;
												assign node35481 = (inp[11]) ? node35487 : node35482;
													assign node35482 = (inp[10]) ? node35484 : 4'b0101;
														assign node35484 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node35487 = (inp[1]) ? node35489 : 4'b1001;
														assign node35489 = (inp[2]) ? 4'b0001 : node35490;
															assign node35490 = (inp[12]) ? 4'b0001 : 4'b0101;
										assign node35494 = (inp[9]) ? node35544 : node35495;
											assign node35495 = (inp[12]) ? node35517 : node35496;
												assign node35496 = (inp[10]) ? node35506 : node35497;
													assign node35497 = (inp[2]) ? 4'b1001 : node35498;
														assign node35498 = (inp[11]) ? 4'b1001 : node35499;
															assign node35499 = (inp[1]) ? 4'b1001 : node35500;
																assign node35500 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node35506 = (inp[1]) ? node35512 : node35507;
														assign node35507 = (inp[6]) ? node35509 : 4'b0001;
															assign node35509 = (inp[11]) ? 4'b1111 : 4'b0001;
														assign node35512 = (inp[6]) ? 4'b1111 : node35513;
															assign node35513 = (inp[11]) ? 4'b1111 : 4'b0001;
												assign node35517 = (inp[10]) ? node35529 : node35518;
													assign node35518 = (inp[1]) ? node35524 : node35519;
														assign node35519 = (inp[11]) ? 4'b1111 : node35520;
															assign node35520 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node35524 = (inp[6]) ? node35526 : 4'b1111;
															assign node35526 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node35529 = (inp[6]) ? node35537 : node35530;
														assign node35530 = (inp[1]) ? node35534 : node35531;
															assign node35531 = (inp[11]) ? 4'b0111 : 4'b1111;
															assign node35534 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node35537 = (inp[1]) ? node35541 : node35538;
															assign node35538 = (inp[2]) ? 4'b0111 : 4'b1111;
															assign node35541 = (inp[11]) ? 4'b0111 : 4'b1111;
											assign node35544 = (inp[10]) ? node35564 : node35545;
												assign node35545 = (inp[2]) ? 4'b0111 : node35546;
													assign node35546 = (inp[11]) ? node35554 : node35547;
														assign node35547 = (inp[1]) ? node35551 : node35548;
															assign node35548 = (inp[6]) ? 4'b0111 : 4'b1111;
															assign node35551 = (inp[12]) ? 4'b1011 : 4'b1111;
														assign node35554 = (inp[12]) ? 4'b0111 : node35555;
															assign node35555 = (inp[6]) ? node35559 : node35556;
																assign node35556 = (inp[1]) ? 4'b1111 : 4'b0111;
																assign node35559 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node35564 = (inp[12]) ? node35574 : node35565;
													assign node35565 = (inp[11]) ? 4'b1011 : node35566;
														assign node35566 = (inp[1]) ? node35570 : node35567;
															assign node35567 = (inp[2]) ? 4'b0111 : 4'b1111;
															assign node35570 = (inp[6]) ? 4'b1011 : 4'b0111;
													assign node35574 = (inp[1]) ? 4'b1011 : node35575;
														assign node35575 = (inp[6]) ? node35577 : 4'b0011;
															assign node35577 = (inp[11]) ? 4'b1011 : 4'b0011;
									assign node35581 = (inp[5]) ? node35657 : node35582;
										assign node35582 = (inp[9]) ? node35620 : node35583;
											assign node35583 = (inp[10]) ? node35599 : node35584;
												assign node35584 = (inp[11]) ? node35594 : node35585;
													assign node35585 = (inp[2]) ? node35591 : node35586;
														assign node35586 = (inp[1]) ? node35588 : 4'b0001;
															assign node35588 = (inp[12]) ? 4'b0001 : 4'b1001;
														assign node35591 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node35594 = (inp[12]) ? node35596 : 4'b0001;
														assign node35596 = (inp[2]) ? 4'b0111 : 4'b1111;
												assign node35599 = (inp[6]) ? node35613 : node35600;
													assign node35600 = (inp[12]) ? node35608 : node35601;
														assign node35601 = (inp[2]) ? 4'b1111 : node35602;
															assign node35602 = (inp[1]) ? 4'b0001 : node35603;
																assign node35603 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node35608 = (inp[11]) ? 4'b1111 : node35609;
															assign node35609 = (inp[1]) ? 4'b0111 : 4'b1111;
													assign node35613 = (inp[1]) ? node35617 : node35614;
														assign node35614 = (inp[11]) ? 4'b1111 : 4'b0111;
														assign node35617 = (inp[11]) ? 4'b0111 : 4'b1111;
											assign node35620 = (inp[10]) ? node35644 : node35621;
												assign node35621 = (inp[12]) ? node35629 : node35622;
													assign node35622 = (inp[1]) ? node35624 : 4'b1111;
														assign node35624 = (inp[11]) ? node35626 : 4'b0111;
															assign node35626 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node35629 = (inp[6]) ? node35639 : node35630;
														assign node35630 = (inp[2]) ? node35632 : 4'b0111;
															assign node35632 = (inp[1]) ? node35636 : node35633;
																assign node35633 = (inp[11]) ? 4'b0111 : 4'b1111;
																assign node35636 = (inp[11]) ? 4'b1011 : 4'b0111;
														assign node35639 = (inp[1]) ? 4'b1011 : node35640;
															assign node35640 = (inp[11]) ? 4'b1011 : 4'b0111;
												assign node35644 = (inp[12]) ? node35652 : node35645;
													assign node35645 = (inp[11]) ? node35647 : 4'b0111;
														assign node35647 = (inp[2]) ? node35649 : 4'b1011;
															assign node35649 = (inp[1]) ? 4'b0011 : 4'b0111;
													assign node35652 = (inp[2]) ? 4'b0011 : node35653;
														assign node35653 = (inp[6]) ? 4'b1011 : 4'b0011;
										assign node35657 = (inp[10]) ? node35707 : node35658;
											assign node35658 = (inp[9]) ? node35686 : node35659;
												assign node35659 = (inp[12]) ? node35671 : node35660;
													assign node35660 = (inp[6]) ? node35666 : node35661;
														assign node35661 = (inp[11]) ? 4'b1011 : node35662;
															assign node35662 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node35666 = (inp[1]) ? node35668 : 4'b0011;
															assign node35668 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node35671 = (inp[11]) ? node35679 : node35672;
														assign node35672 = (inp[2]) ? 4'b0011 : node35673;
															assign node35673 = (inp[1]) ? node35675 : 4'b0011;
																assign node35675 = (inp[6]) ? 4'b1111 : 4'b0011;
														assign node35679 = (inp[6]) ? node35683 : node35680;
															assign node35680 = (inp[1]) ? 4'b1111 : 4'b0011;
															assign node35683 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node35686 = (inp[11]) ? node35698 : node35687;
													assign node35687 = (inp[12]) ? 4'b0111 : node35688;
														assign node35688 = (inp[2]) ? node35694 : node35689;
															assign node35689 = (inp[6]) ? node35691 : 4'b0111;
																assign node35691 = (inp[1]) ? 4'b1111 : 4'b0111;
															assign node35694 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node35698 = (inp[12]) ? node35702 : node35699;
														assign node35699 = (inp[2]) ? 4'b0111 : 4'b1111;
														assign node35702 = (inp[6]) ? node35704 : 4'b1011;
															assign node35704 = (inp[1]) ? 4'b0011 : 4'b1011;
											assign node35707 = (inp[9]) ? node35731 : node35708;
												assign node35708 = (inp[12]) ? node35718 : node35709;
													assign node35709 = (inp[1]) ? node35711 : 4'b0011;
														assign node35711 = (inp[6]) ? node35715 : node35712;
															assign node35712 = (inp[2]) ? 4'b1111 : 4'b0011;
															assign node35715 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node35718 = (inp[11]) ? node35724 : node35719;
														assign node35719 = (inp[6]) ? node35721 : 4'b1111;
															assign node35721 = (inp[1]) ? 4'b1111 : 4'b0111;
														assign node35724 = (inp[1]) ? node35728 : node35725;
															assign node35725 = (inp[6]) ? 4'b1111 : 4'b0111;
															assign node35728 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node35731 = (inp[12]) ? node35743 : node35732;
													assign node35732 = (inp[6]) ? node35738 : node35733;
														assign node35733 = (inp[1]) ? 4'b0111 : node35734;
															assign node35734 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node35738 = (inp[2]) ? 4'b0111 : node35739;
															assign node35739 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node35743 = (inp[11]) ? node35745 : 4'b0011;
														assign node35745 = (inp[2]) ? 4'b1011 : node35746;
															assign node35746 = (inp[1]) ? 4'b0011 : node35747;
																assign node35747 = (inp[6]) ? 4'b1011 : 4'b0011;
							assign node35752 = (inp[0]) ? node36090 : node35753;
								assign node35753 = (inp[5]) ? node35951 : node35754;
									assign node35754 = (inp[3]) ? node35846 : node35755;
										assign node35755 = (inp[6]) ? node35801 : node35756;
											assign node35756 = (inp[9]) ? node35786 : node35757;
												assign node35757 = (inp[12]) ? node35767 : node35758;
													assign node35758 = (inp[1]) ? node35762 : node35759;
														assign node35759 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node35762 = (inp[11]) ? node35764 : 4'b0001;
															assign node35764 = (inp[10]) ? 4'b1101 : 4'b1001;
													assign node35767 = (inp[10]) ? node35775 : node35768;
														assign node35768 = (inp[11]) ? node35772 : node35769;
															assign node35769 = (inp[1]) ? 4'b0001 : 4'b1001;
															assign node35772 = (inp[1]) ? 4'b1101 : 4'b0001;
														assign node35775 = (inp[2]) ? node35781 : node35776;
															assign node35776 = (inp[11]) ? node35778 : 4'b1101;
																assign node35778 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node35781 = (inp[1]) ? node35783 : 4'b1101;
																assign node35783 = (inp[11]) ? 4'b1101 : 4'b0101;
												assign node35786 = (inp[12]) ? node35792 : node35787;
													assign node35787 = (inp[10]) ? node35789 : 4'b1101;
														assign node35789 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node35792 = (inp[10]) ? node35796 : node35793;
														assign node35793 = (inp[1]) ? 4'b0101 : 4'b1101;
														assign node35796 = (inp[1]) ? node35798 : 4'b1001;
															assign node35798 = (inp[11]) ? 4'b1001 : 4'b0001;
											assign node35801 = (inp[11]) ? node35823 : node35802;
												assign node35802 = (inp[1]) ? node35814 : node35803;
													assign node35803 = (inp[9]) ? node35809 : node35804;
														assign node35804 = (inp[12]) ? node35806 : 4'b0001;
															assign node35806 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node35809 = (inp[10]) ? node35811 : 4'b0101;
															assign node35811 = (inp[12]) ? 4'b0001 : 4'b0101;
													assign node35814 = (inp[12]) ? node35820 : node35815;
														assign node35815 = (inp[2]) ? node35817 : 4'b1001;
															assign node35817 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node35820 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node35823 = (inp[1]) ? node35835 : node35824;
													assign node35824 = (inp[9]) ? node35830 : node35825;
														assign node35825 = (inp[12]) ? 4'b1101 : node35826;
															assign node35826 = (inp[10]) ? 4'b1101 : 4'b1001;
														assign node35830 = (inp[10]) ? 4'b1001 : node35831;
															assign node35831 = (inp[12]) ? 4'b1001 : 4'b1101;
													assign node35835 = (inp[9]) ? node35841 : node35836;
														assign node35836 = (inp[12]) ? 4'b0101 : node35837;
															assign node35837 = (inp[10]) ? 4'b0101 : 4'b0001;
														assign node35841 = (inp[12]) ? 4'b0001 : node35842;
															assign node35842 = (inp[2]) ? 4'b0001 : 4'b0101;
										assign node35846 = (inp[9]) ? node35906 : node35847;
											assign node35847 = (inp[12]) ? node35885 : node35848;
												assign node35848 = (inp[10]) ? node35866 : node35849;
													assign node35849 = (inp[2]) ? node35861 : node35850;
														assign node35850 = (inp[1]) ? node35856 : node35851;
															assign node35851 = (inp[6]) ? node35853 : 4'b1001;
																assign node35853 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node35856 = (inp[6]) ? 4'b0001 : node35857;
																assign node35857 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node35861 = (inp[11]) ? 4'b0001 : node35862;
															assign node35862 = (inp[6]) ? 4'b1001 : 4'b0001;
													assign node35866 = (inp[11]) ? node35876 : node35867;
														assign node35867 = (inp[2]) ? node35869 : 4'b0001;
															assign node35869 = (inp[6]) ? node35873 : node35870;
																assign node35870 = (inp[1]) ? 4'b0001 : 4'b1001;
																assign node35873 = (inp[1]) ? 4'b1111 : 4'b0001;
														assign node35876 = (inp[2]) ? 4'b0001 : node35877;
															assign node35877 = (inp[1]) ? node35881 : node35878;
																assign node35878 = (inp[6]) ? 4'b1111 : 4'b0001;
																assign node35881 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node35885 = (inp[10]) ? node35895 : node35886;
													assign node35886 = (inp[11]) ? node35888 : 4'b0001;
														assign node35888 = (inp[1]) ? node35892 : node35889;
															assign node35889 = (inp[6]) ? 4'b1111 : 4'b0001;
															assign node35892 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node35895 = (inp[2]) ? node35899 : node35896;
														assign node35896 = (inp[6]) ? 4'b1111 : 4'b0111;
														assign node35899 = (inp[1]) ? node35901 : 4'b1111;
															assign node35901 = (inp[6]) ? node35903 : 4'b1111;
																assign node35903 = (inp[11]) ? 4'b0111 : 4'b1111;
											assign node35906 = (inp[10]) ? node35930 : node35907;
												assign node35907 = (inp[12]) ? node35921 : node35908;
													assign node35908 = (inp[1]) ? node35910 : 4'b1111;
														assign node35910 = (inp[2]) ? node35916 : node35911;
															assign node35911 = (inp[11]) ? node35913 : 4'b0111;
																assign node35913 = (inp[6]) ? 4'b0111 : 4'b1111;
															assign node35916 = (inp[6]) ? node35918 : 4'b1111;
																assign node35918 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node35921 = (inp[11]) ? 4'b1011 : node35922;
														assign node35922 = (inp[2]) ? 4'b0111 : node35923;
															assign node35923 = (inp[1]) ? 4'b1011 : node35924;
																assign node35924 = (inp[6]) ? 4'b0111 : 4'b1111;
												assign node35930 = (inp[11]) ? node35942 : node35931;
													assign node35931 = (inp[12]) ? node35935 : node35932;
														assign node35932 = (inp[1]) ? 4'b1011 : 4'b0111;
														assign node35935 = (inp[2]) ? node35937 : 4'b0011;
															assign node35937 = (inp[1]) ? 4'b0011 : node35938;
																assign node35938 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node35942 = (inp[1]) ? node35948 : node35943;
														assign node35943 = (inp[6]) ? 4'b1011 : node35944;
															assign node35944 = (inp[12]) ? 4'b0011 : 4'b0111;
														assign node35948 = (inp[6]) ? 4'b0011 : 4'b1011;
									assign node35951 = (inp[9]) ? node36029 : node35952;
										assign node35952 = (inp[10]) ? node35994 : node35953;
											assign node35953 = (inp[3]) ? node35979 : node35954;
												assign node35954 = (inp[12]) ? node35972 : node35955;
													assign node35955 = (inp[2]) ? node35967 : node35956;
														assign node35956 = (inp[6]) ? node35962 : node35957;
															assign node35957 = (inp[1]) ? 4'b0001 : node35958;
																assign node35958 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node35962 = (inp[1]) ? 4'b1001 : node35963;
																assign node35963 = (inp[11]) ? 4'b1001 : 4'b0001;
														assign node35967 = (inp[6]) ? node35969 : 4'b1001;
															assign node35969 = (inp[1]) ? 4'b0001 : 4'b1001;
													assign node35972 = (inp[2]) ? node35976 : node35973;
														assign node35973 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node35976 = (inp[1]) ? 4'b0111 : 4'b0001;
												assign node35979 = (inp[11]) ? node35985 : node35980;
													assign node35980 = (inp[6]) ? node35982 : 4'b1011;
														assign node35982 = (inp[1]) ? 4'b1011 : 4'b0011;
													assign node35985 = (inp[1]) ? node35987 : 4'b0011;
														assign node35987 = (inp[12]) ? node35991 : node35988;
															assign node35988 = (inp[6]) ? 4'b0011 : 4'b1011;
															assign node35991 = (inp[2]) ? 4'b1111 : 4'b0111;
											assign node35994 = (inp[12]) ? node36016 : node35995;
												assign node35995 = (inp[1]) ? node36009 : node35996;
													assign node35996 = (inp[3]) ? node36004 : node35997;
														assign node35997 = (inp[11]) ? node36001 : node35998;
															assign node35998 = (inp[6]) ? 4'b0001 : 4'b1001;
															assign node36001 = (inp[6]) ? 4'b1111 : 4'b0001;
														assign node36004 = (inp[6]) ? 4'b1111 : node36005;
															assign node36005 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node36009 = (inp[6]) ? node36013 : node36010;
														assign node36010 = (inp[11]) ? 4'b1111 : 4'b0001;
														assign node36013 = (inp[11]) ? 4'b0111 : 4'b1111;
												assign node36016 = (inp[1]) ? node36024 : node36017;
													assign node36017 = (inp[6]) ? node36021 : node36018;
														assign node36018 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node36021 = (inp[11]) ? 4'b1111 : 4'b0111;
													assign node36024 = (inp[6]) ? 4'b1111 : node36025;
														assign node36025 = (inp[11]) ? 4'b1111 : 4'b0111;
										assign node36029 = (inp[12]) ? node36063 : node36030;
											assign node36030 = (inp[6]) ? node36046 : node36031;
												assign node36031 = (inp[3]) ? node36041 : node36032;
													assign node36032 = (inp[11]) ? node36036 : node36033;
														assign node36033 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node36036 = (inp[1]) ? node36038 : 4'b0111;
															assign node36038 = (inp[2]) ? 4'b1111 : 4'b1011;
													assign node36041 = (inp[11]) ? 4'b0111 : node36042;
														assign node36042 = (inp[1]) ? 4'b0111 : 4'b1111;
												assign node36046 = (inp[10]) ? node36056 : node36047;
													assign node36047 = (inp[2]) ? node36049 : 4'b1111;
														assign node36049 = (inp[1]) ? node36053 : node36050;
															assign node36050 = (inp[11]) ? 4'b1111 : 4'b0111;
															assign node36053 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node36056 = (inp[11]) ? node36060 : node36057;
														assign node36057 = (inp[1]) ? 4'b1011 : 4'b0111;
														assign node36060 = (inp[1]) ? 4'b0011 : 4'b1011;
											assign node36063 = (inp[10]) ? node36077 : node36064;
												assign node36064 = (inp[1]) ? node36070 : node36065;
													assign node36065 = (inp[6]) ? 4'b0111 : node36066;
														assign node36066 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node36070 = (inp[6]) ? node36074 : node36071;
														assign node36071 = (inp[11]) ? 4'b1011 : 4'b0111;
														assign node36074 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node36077 = (inp[6]) ? node36085 : node36078;
													assign node36078 = (inp[1]) ? node36082 : node36079;
														assign node36079 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node36082 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node36085 = (inp[11]) ? node36087 : 4'b0011;
														assign node36087 = (inp[1]) ? 4'b0011 : 4'b1011;
								assign node36090 = (inp[5]) ? node36288 : node36091;
									assign node36091 = (inp[3]) ? node36193 : node36092;
										assign node36092 = (inp[11]) ? node36136 : node36093;
											assign node36093 = (inp[12]) ? node36111 : node36094;
												assign node36094 = (inp[9]) ? node36104 : node36095;
													assign node36095 = (inp[6]) ? node36099 : node36096;
														assign node36096 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node36099 = (inp[1]) ? node36101 : 4'b0011;
															assign node36101 = (inp[10]) ? 4'b1111 : 4'b1011;
													assign node36104 = (inp[10]) ? node36106 : 4'b1111;
														assign node36106 = (inp[6]) ? node36108 : 4'b0111;
															assign node36108 = (inp[1]) ? 4'b1011 : 4'b0111;
												assign node36111 = (inp[9]) ? node36123 : node36112;
													assign node36112 = (inp[10]) ? node36116 : node36113;
														assign node36113 = (inp[2]) ? 4'b1111 : 4'b1011;
														assign node36116 = (inp[1]) ? node36120 : node36117;
															assign node36117 = (inp[6]) ? 4'b0111 : 4'b1111;
															assign node36120 = (inp[6]) ? 4'b1111 : 4'b0111;
													assign node36123 = (inp[10]) ? node36131 : node36124;
														assign node36124 = (inp[2]) ? 4'b1011 : node36125;
															assign node36125 = (inp[6]) ? 4'b0111 : node36126;
																assign node36126 = (inp[1]) ? 4'b0111 : 4'b1111;
														assign node36131 = (inp[1]) ? 4'b1011 : node36132;
															assign node36132 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node36136 = (inp[9]) ? node36158 : node36137;
												assign node36137 = (inp[10]) ? node36145 : node36138;
													assign node36138 = (inp[6]) ? node36142 : node36139;
														assign node36139 = (inp[1]) ? 4'b1011 : 4'b0011;
														assign node36142 = (inp[12]) ? 4'b0111 : 4'b0011;
													assign node36145 = (inp[2]) ? node36153 : node36146;
														assign node36146 = (inp[1]) ? node36150 : node36147;
															assign node36147 = (inp[6]) ? 4'b1111 : 4'b0011;
															assign node36150 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node36153 = (inp[6]) ? 4'b0111 : node36154;
															assign node36154 = (inp[1]) ? 4'b1111 : 4'b0111;
												assign node36158 = (inp[10]) ? node36170 : node36159;
													assign node36159 = (inp[12]) ? node36167 : node36160;
														assign node36160 = (inp[2]) ? 4'b0111 : node36161;
															assign node36161 = (inp[1]) ? node36163 : 4'b1111;
																assign node36163 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node36167 = (inp[1]) ? 4'b1011 : 4'b0111;
													assign node36170 = (inp[2]) ? node36180 : node36171;
														assign node36171 = (inp[12]) ? node36173 : 4'b1011;
															assign node36173 = (inp[1]) ? node36177 : node36174;
																assign node36174 = (inp[6]) ? 4'b1011 : 4'b0011;
																assign node36177 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node36180 = (inp[12]) ? node36186 : node36181;
															assign node36181 = (inp[6]) ? node36183 : 4'b0111;
																assign node36183 = (inp[1]) ? 4'b0011 : 4'b1011;
															assign node36186 = (inp[6]) ? node36190 : node36187;
																assign node36187 = (inp[1]) ? 4'b1011 : 4'b0011;
																assign node36190 = (inp[1]) ? 4'b0011 : 4'b1011;
										assign node36193 = (inp[9]) ? node36243 : node36194;
											assign node36194 = (inp[12]) ? node36220 : node36195;
												assign node36195 = (inp[10]) ? node36209 : node36196;
													assign node36196 = (inp[2]) ? node36202 : node36197;
														assign node36197 = (inp[11]) ? node36199 : 4'b0011;
															assign node36199 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node36202 = (inp[6]) ? node36204 : 4'b1011;
															assign node36204 = (inp[1]) ? node36206 : 4'b0011;
																assign node36206 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node36209 = (inp[1]) ? node36215 : node36210;
														assign node36210 = (inp[11]) ? 4'b0011 : node36211;
															assign node36211 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node36215 = (inp[6]) ? node36217 : 4'b0011;
															assign node36217 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node36220 = (inp[10]) ? node36232 : node36221;
													assign node36221 = (inp[1]) ? node36225 : node36222;
														assign node36222 = (inp[2]) ? 4'b0011 : 4'b1101;
														assign node36225 = (inp[6]) ? node36229 : node36226;
															assign node36226 = (inp[11]) ? 4'b1101 : 4'b0011;
															assign node36229 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node36232 = (inp[1]) ? 4'b1101 : node36233;
														assign node36233 = (inp[2]) ? 4'b0101 : node36234;
															assign node36234 = (inp[6]) ? node36238 : node36235;
																assign node36235 = (inp[11]) ? 4'b0101 : 4'b1101;
																assign node36238 = (inp[11]) ? 4'b1101 : 4'b0101;
											assign node36243 = (inp[10]) ? node36265 : node36244;
												assign node36244 = (inp[1]) ? node36252 : node36245;
													assign node36245 = (inp[6]) ? node36249 : node36246;
														assign node36246 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node36249 = (inp[11]) ? 4'b1101 : 4'b0101;
													assign node36252 = (inp[12]) ? node36258 : node36253;
														assign node36253 = (inp[6]) ? 4'b1101 : node36254;
															assign node36254 = (inp[2]) ? 4'b1101 : 4'b0101;
														assign node36258 = (inp[6]) ? node36262 : node36259;
															assign node36259 = (inp[2]) ? 4'b1001 : 4'b0101;
															assign node36262 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node36265 = (inp[12]) ? node36275 : node36266;
													assign node36266 = (inp[11]) ? 4'b1001 : node36267;
														assign node36267 = (inp[6]) ? node36271 : node36268;
															assign node36268 = (inp[1]) ? 4'b0101 : 4'b1101;
															assign node36271 = (inp[1]) ? 4'b1001 : 4'b0101;
													assign node36275 = (inp[1]) ? node36281 : node36276;
														assign node36276 = (inp[11]) ? node36278 : 4'b0001;
															assign node36278 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node36281 = (inp[6]) ? node36285 : node36282;
															assign node36282 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node36285 = (inp[11]) ? 4'b0001 : 4'b1001;
									assign node36288 = (inp[9]) ? node36380 : node36289;
										assign node36289 = (inp[12]) ? node36335 : node36290;
											assign node36290 = (inp[3]) ? node36312 : node36291;
												assign node36291 = (inp[6]) ? node36305 : node36292;
													assign node36292 = (inp[2]) ? node36300 : node36293;
														assign node36293 = (inp[10]) ? 4'b0011 : node36294;
															assign node36294 = (inp[11]) ? 4'b1011 : node36295;
																assign node36295 = (inp[1]) ? 4'b0011 : 4'b1011;
														assign node36300 = (inp[11]) ? 4'b0011 : node36301;
															assign node36301 = (inp[10]) ? 4'b1011 : 4'b0011;
													assign node36305 = (inp[10]) ? node36307 : 4'b1011;
														assign node36307 = (inp[11]) ? node36309 : 4'b0011;
															assign node36309 = (inp[1]) ? 4'b0101 : 4'b1101;
												assign node36312 = (inp[10]) ? node36322 : node36313;
													assign node36313 = (inp[1]) ? 4'b1001 : node36314;
														assign node36314 = (inp[2]) ? node36316 : 4'b0001;
															assign node36316 = (inp[6]) ? node36318 : 4'b1001;
																assign node36318 = (inp[11]) ? 4'b1001 : 4'b0001;
													assign node36322 = (inp[1]) ? node36330 : node36323;
														assign node36323 = (inp[2]) ? 4'b1001 : node36324;
															assign node36324 = (inp[6]) ? node36326 : 4'b0001;
																assign node36326 = (inp[11]) ? 4'b1101 : 4'b0001;
														assign node36330 = (inp[11]) ? node36332 : 4'b1101;
															assign node36332 = (inp[6]) ? 4'b0101 : 4'b1101;
											assign node36335 = (inp[10]) ? node36351 : node36336;
												assign node36336 = (inp[1]) ? node36346 : node36337;
													assign node36337 = (inp[3]) ? node36343 : node36338;
														assign node36338 = (inp[11]) ? node36340 : 4'b0011;
															assign node36340 = (inp[6]) ? 4'b1101 : 4'b0011;
														assign node36343 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node36346 = (inp[11]) ? node36348 : 4'b1101;
														assign node36348 = (inp[6]) ? 4'b0101 : 4'b1101;
												assign node36351 = (inp[2]) ? node36363 : node36352;
													assign node36352 = (inp[1]) ? node36358 : node36353;
														assign node36353 = (inp[6]) ? node36355 : 4'b1101;
															assign node36355 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node36358 = (inp[6]) ? node36360 : 4'b0101;
															assign node36360 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node36363 = (inp[3]) ? node36371 : node36364;
														assign node36364 = (inp[11]) ? node36366 : 4'b1101;
															assign node36366 = (inp[1]) ? node36368 : 4'b1101;
																assign node36368 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node36371 = (inp[6]) ? 4'b0101 : node36372;
															assign node36372 = (inp[1]) ? node36376 : node36373;
																assign node36373 = (inp[11]) ? 4'b0101 : 4'b1101;
																assign node36376 = (inp[11]) ? 4'b1101 : 4'b0101;
										assign node36380 = (inp[12]) ? node36430 : node36381;
											assign node36381 = (inp[10]) ? node36411 : node36382;
												assign node36382 = (inp[2]) ? node36396 : node36383;
													assign node36383 = (inp[3]) ? node36385 : 4'b0101;
														assign node36385 = (inp[11]) ? node36391 : node36386;
															assign node36386 = (inp[6]) ? node36388 : 4'b0101;
																assign node36388 = (inp[1]) ? 4'b1101 : 4'b0101;
															assign node36391 = (inp[6]) ? node36393 : 4'b1101;
																assign node36393 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node36396 = (inp[1]) ? node36404 : node36397;
														assign node36397 = (inp[6]) ? node36401 : node36398;
															assign node36398 = (inp[11]) ? 4'b0101 : 4'b1101;
															assign node36401 = (inp[11]) ? 4'b1101 : 4'b0101;
														assign node36404 = (inp[6]) ? node36408 : node36405;
															assign node36405 = (inp[11]) ? 4'b1101 : 4'b0101;
															assign node36408 = (inp[11]) ? 4'b0101 : 4'b1101;
												assign node36411 = (inp[11]) ? node36423 : node36412;
													assign node36412 = (inp[2]) ? node36418 : node36413;
														assign node36413 = (inp[1]) ? 4'b1001 : node36414;
															assign node36414 = (inp[6]) ? 4'b0101 : 4'b1101;
														assign node36418 = (inp[1]) ? 4'b0101 : node36419;
															assign node36419 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node36423 = (inp[1]) ? node36427 : node36424;
														assign node36424 = (inp[6]) ? 4'b1001 : 4'b0101;
														assign node36427 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node36430 = (inp[10]) ? node36446 : node36431;
												assign node36431 = (inp[6]) ? node36439 : node36432;
													assign node36432 = (inp[2]) ? node36434 : 4'b0101;
														assign node36434 = (inp[11]) ? 4'b1001 : node36435;
															assign node36435 = (inp[1]) ? 4'b0101 : 4'b1101;
													assign node36439 = (inp[11]) ? node36443 : node36440;
														assign node36440 = (inp[1]) ? 4'b1001 : 4'b0101;
														assign node36443 = (inp[1]) ? 4'b0001 : 4'b1001;
												assign node36446 = (inp[2]) ? node36458 : node36447;
													assign node36447 = (inp[11]) ? node36453 : node36448;
														assign node36448 = (inp[1]) ? node36450 : 4'b0001;
															assign node36450 = (inp[6]) ? 4'b1001 : 4'b0001;
														assign node36453 = (inp[1]) ? node36455 : 4'b1001;
															assign node36455 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node36458 = (inp[11]) ? node36460 : 4'b1001;
														assign node36460 = (inp[1]) ? node36464 : node36461;
															assign node36461 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node36464 = (inp[6]) ? 4'b0001 : 4'b1001;
					assign node36467 = (inp[12]) ? node37719 : node36468;
						assign node36468 = (inp[10]) ? node37074 : node36469;
							assign node36469 = (inp[3]) ? node36761 : node36470;
								assign node36470 = (inp[11]) ? node36614 : node36471;
									assign node36471 = (inp[6]) ? node36553 : node36472;
										assign node36472 = (inp[2]) ? node36518 : node36473;
											assign node36473 = (inp[0]) ? node36495 : node36474;
												assign node36474 = (inp[15]) ? node36486 : node36475;
													assign node36475 = (inp[5]) ? node36483 : node36476;
														assign node36476 = (inp[4]) ? node36480 : node36477;
															assign node36477 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node36480 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node36483 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node36486 = (inp[9]) ? node36490 : node36487;
														assign node36487 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node36490 = (inp[4]) ? node36492 : 4'b0001;
															assign node36492 = (inp[5]) ? 4'b0111 : 4'b0101;
												assign node36495 = (inp[15]) ? node36505 : node36496;
													assign node36496 = (inp[4]) ? node36500 : node36497;
														assign node36497 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node36500 = (inp[9]) ? node36502 : 4'b0001;
															assign node36502 = (inp[1]) ? 4'b0111 : 4'b0101;
													assign node36505 = (inp[5]) ? node36511 : node36506;
														assign node36506 = (inp[9]) ? 4'b0111 : node36507;
															assign node36507 = (inp[4]) ? 4'b0011 : 4'b0111;
														assign node36511 = (inp[9]) ? node36515 : node36512;
															assign node36512 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node36515 = (inp[4]) ? 4'b0101 : 4'b0011;
											assign node36518 = (inp[0]) ? node36538 : node36519;
												assign node36519 = (inp[15]) ? node36533 : node36520;
													assign node36520 = (inp[1]) ? node36528 : node36521;
														assign node36521 = (inp[4]) ? node36525 : node36522;
															assign node36522 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node36525 = (inp[9]) ? 4'b0111 : 4'b0011;
														assign node36528 = (inp[9]) ? node36530 : 4'b0011;
															assign node36530 = (inp[4]) ? 4'b0101 : 4'b0011;
													assign node36533 = (inp[4]) ? 4'b0001 : node36534;
														assign node36534 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node36538 = (inp[15]) ? node36546 : node36539;
													assign node36539 = (inp[9]) ? node36543 : node36540;
														assign node36540 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node36543 = (inp[4]) ? 4'b0101 : 4'b0001;
													assign node36546 = (inp[4]) ? node36550 : node36547;
														assign node36547 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node36550 = (inp[9]) ? 4'b0101 : 4'b0011;
										assign node36553 = (inp[4]) ? node36579 : node36554;
											assign node36554 = (inp[9]) ? node36570 : node36555;
												assign node36555 = (inp[2]) ? node36563 : node36556;
													assign node36556 = (inp[5]) ? 4'b1101 : node36557;
														assign node36557 = (inp[0]) ? node36559 : 4'b1111;
															assign node36559 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node36563 = (inp[0]) ? node36567 : node36564;
														assign node36564 = (inp[1]) ? 4'b1111 : 4'b1101;
														assign node36567 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node36570 = (inp[2]) ? 4'b1001 : node36571;
													assign node36571 = (inp[0]) ? node36575 : node36572;
														assign node36572 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node36575 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node36579 = (inp[9]) ? node36597 : node36580;
												assign node36580 = (inp[5]) ? node36592 : node36581;
													assign node36581 = (inp[1]) ? node36589 : node36582;
														assign node36582 = (inp[2]) ? 4'b1011 : node36583;
															assign node36583 = (inp[0]) ? 4'b1001 : node36584;
																assign node36584 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node36589 = (inp[2]) ? 4'b1001 : 4'b1011;
													assign node36592 = (inp[0]) ? node36594 : 4'b1011;
														assign node36594 = (inp[2]) ? 4'b1011 : 4'b1001;
												assign node36597 = (inp[15]) ? node36603 : node36598;
													assign node36598 = (inp[5]) ? node36600 : 4'b1111;
														assign node36600 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node36603 = (inp[1]) ? node36609 : node36604;
														assign node36604 = (inp[5]) ? node36606 : 4'b1111;
															assign node36606 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node36609 = (inp[0]) ? node36611 : 4'b1101;
															assign node36611 = (inp[5]) ? 4'b1101 : 4'b1111;
									assign node36614 = (inp[6]) ? node36714 : node36615;
										assign node36615 = (inp[1]) ? node36669 : node36616;
											assign node36616 = (inp[2]) ? node36642 : node36617;
												assign node36617 = (inp[15]) ? node36633 : node36618;
													assign node36618 = (inp[0]) ? node36624 : node36619;
														assign node36619 = (inp[9]) ? node36621 : 4'b1111;
															assign node36621 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node36624 = (inp[5]) ? node36626 : 4'b1101;
															assign node36626 = (inp[9]) ? node36630 : node36627;
																assign node36627 = (inp[4]) ? 4'b1001 : 4'b1101;
																assign node36630 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node36633 = (inp[0]) ? node36637 : node36634;
														assign node36634 = (inp[9]) ? 4'b1111 : 4'b1101;
														assign node36637 = (inp[4]) ? 4'b1011 : node36638;
															assign node36638 = (inp[9]) ? 4'b1011 : 4'b1111;
												assign node36642 = (inp[0]) ? node36656 : node36643;
													assign node36643 = (inp[15]) ? node36649 : node36644;
														assign node36644 = (inp[9]) ? 4'b1011 : node36645;
															assign node36645 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node36649 = (inp[5]) ? node36651 : 4'b1001;
															assign node36651 = (inp[4]) ? node36653 : 4'b1001;
																assign node36653 = (inp[9]) ? 4'b1111 : 4'b1001;
													assign node36656 = (inp[4]) ? node36662 : node36657;
														assign node36657 = (inp[9]) ? node36659 : 4'b1111;
															assign node36659 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node36662 = (inp[9]) ? node36664 : 4'b1011;
															assign node36664 = (inp[15]) ? node36666 : 4'b1111;
																assign node36666 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node36669 = (inp[15]) ? node36691 : node36670;
												assign node36670 = (inp[0]) ? node36674 : node36671;
													assign node36671 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node36674 = (inp[2]) ? node36684 : node36675;
														assign node36675 = (inp[5]) ? node36679 : node36676;
															assign node36676 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node36679 = (inp[9]) ? 4'b1001 : node36680;
																assign node36680 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node36684 = (inp[5]) ? 4'b1001 : node36685;
															assign node36685 = (inp[9]) ? 4'b1001 : node36686;
																assign node36686 = (inp[4]) ? 4'b1001 : 4'b1101;
												assign node36691 = (inp[0]) ? node36705 : node36692;
													assign node36692 = (inp[5]) ? node36694 : 4'b1101;
														assign node36694 = (inp[2]) ? node36700 : node36695;
															assign node36695 = (inp[4]) ? 4'b1001 : node36696;
																assign node36696 = (inp[9]) ? 4'b1001 : 4'b1101;
															assign node36700 = (inp[9]) ? node36702 : 4'b1001;
																assign node36702 = (inp[4]) ? 4'b1111 : 4'b1001;
													assign node36705 = (inp[4]) ? node36709 : node36706;
														assign node36706 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node36709 = (inp[5]) ? 4'b1101 : node36710;
															assign node36710 = (inp[9]) ? 4'b1111 : 4'b1011;
										assign node36714 = (inp[4]) ? node36740 : node36715;
											assign node36715 = (inp[9]) ? node36733 : node36716;
												assign node36716 = (inp[5]) ? node36724 : node36717;
													assign node36717 = (inp[2]) ? node36719 : 4'b0111;
														assign node36719 = (inp[15]) ? node36721 : 4'b0101;
															assign node36721 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node36724 = (inp[1]) ? node36726 : 4'b0101;
														assign node36726 = (inp[15]) ? node36730 : node36727;
															assign node36727 = (inp[0]) ? 4'b0101 : 4'b0111;
															assign node36730 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node36733 = (inp[0]) ? node36737 : node36734;
													assign node36734 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node36737 = (inp[15]) ? 4'b0011 : 4'b0001;
											assign node36740 = (inp[9]) ? node36748 : node36741;
												assign node36741 = (inp[15]) ? node36745 : node36742;
													assign node36742 = (inp[0]) ? 4'b0001 : 4'b0011;
													assign node36745 = (inp[0]) ? 4'b0011 : 4'b0001;
												assign node36748 = (inp[15]) ? node36756 : node36749;
													assign node36749 = (inp[0]) ? node36753 : node36750;
														assign node36750 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node36753 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node36756 = (inp[0]) ? 4'b0111 : node36757;
														assign node36757 = (inp[5]) ? 4'b0111 : 4'b0101;
								assign node36761 = (inp[6]) ? node36917 : node36762;
									assign node36762 = (inp[11]) ? node36852 : node36763;
										assign node36763 = (inp[4]) ? node36811 : node36764;
											assign node36764 = (inp[9]) ? node36792 : node36765;
												assign node36765 = (inp[5]) ? node36773 : node36766;
													assign node36766 = (inp[15]) ? node36770 : node36767;
														assign node36767 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node36770 = (inp[0]) ? 4'b0111 : 4'b0101;
													assign node36773 = (inp[2]) ? node36787 : node36774;
														assign node36774 = (inp[1]) ? node36780 : node36775;
															assign node36775 = (inp[0]) ? node36777 : 4'b0101;
																assign node36777 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node36780 = (inp[15]) ? node36784 : node36781;
																assign node36781 = (inp[0]) ? 4'b0111 : 4'b0101;
																assign node36784 = (inp[0]) ? 4'b0101 : 4'b0111;
														assign node36787 = (inp[15]) ? node36789 : 4'b0111;
															assign node36789 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node36792 = (inp[0]) ? node36804 : node36793;
													assign node36793 = (inp[2]) ? node36799 : node36794;
														assign node36794 = (inp[15]) ? node36796 : 4'b0011;
															assign node36796 = (inp[5]) ? 4'b0011 : 4'b0001;
														assign node36799 = (inp[5]) ? 4'b0001 : node36800;
															assign node36800 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node36804 = (inp[5]) ? node36808 : node36805;
														assign node36805 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node36808 = (inp[15]) ? 4'b0001 : 4'b0011;
											assign node36811 = (inp[9]) ? node36839 : node36812;
												assign node36812 = (inp[5]) ? node36820 : node36813;
													assign node36813 = (inp[15]) ? node36817 : node36814;
														assign node36814 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node36817 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node36820 = (inp[2]) ? node36826 : node36821;
														assign node36821 = (inp[15]) ? 4'b0001 : node36822;
															assign node36822 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node36826 = (inp[1]) ? node36832 : node36827;
															assign node36827 = (inp[15]) ? node36829 : 4'b0001;
																assign node36829 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node36832 = (inp[0]) ? node36836 : node36833;
																assign node36833 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node36836 = (inp[15]) ? 4'b0001 : 4'b0011;
												assign node36839 = (inp[5]) ? node36847 : node36840;
													assign node36840 = (inp[1]) ? 4'b0111 : node36841;
														assign node36841 = (inp[2]) ? node36843 : 4'b0101;
															assign node36843 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node36847 = (inp[0]) ? 4'b0101 : node36848;
														assign node36848 = (inp[15]) ? 4'b0111 : 4'b0101;
										assign node36852 = (inp[4]) ? node36884 : node36853;
											assign node36853 = (inp[9]) ? node36873 : node36854;
												assign node36854 = (inp[15]) ? node36868 : node36855;
													assign node36855 = (inp[1]) ? node36863 : node36856;
														assign node36856 = (inp[0]) ? node36860 : node36857;
															assign node36857 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node36860 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node36863 = (inp[5]) ? 4'b1101 : node36864;
															assign node36864 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node36868 = (inp[0]) ? 4'b1111 : node36869;
														assign node36869 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node36873 = (inp[0]) ? node36879 : node36874;
													assign node36874 = (inp[5]) ? node36876 : 4'b1011;
														assign node36876 = (inp[1]) ? 4'b1001 : 4'b1011;
													assign node36879 = (inp[5]) ? node36881 : 4'b1001;
														assign node36881 = (inp[15]) ? 4'b1001 : 4'b1011;
											assign node36884 = (inp[9]) ? node36910 : node36885;
												assign node36885 = (inp[15]) ? node36897 : node36886;
													assign node36886 = (inp[2]) ? 4'b1001 : node36887;
														assign node36887 = (inp[1]) ? node36889 : 4'b1001;
															assign node36889 = (inp[0]) ? node36893 : node36890;
																assign node36890 = (inp[5]) ? 4'b1001 : 4'b1011;
																assign node36893 = (inp[5]) ? 4'b1011 : 4'b1001;
													assign node36897 = (inp[2]) ? node36903 : node36898;
														assign node36898 = (inp[0]) ? node36900 : 4'b1011;
															assign node36900 = (inp[5]) ? 4'b1001 : 4'b1011;
														assign node36903 = (inp[1]) ? node36905 : 4'b1001;
															assign node36905 = (inp[0]) ? 4'b1011 : node36906;
																assign node36906 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node36910 = (inp[15]) ? node36914 : node36911;
													assign node36911 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node36914 = (inp[0]) ? 4'b1101 : 4'b1111;
									assign node36917 = (inp[11]) ? node37007 : node36918;
										assign node36918 = (inp[4]) ? node36960 : node36919;
											assign node36919 = (inp[9]) ? node36945 : node36920;
												assign node36920 = (inp[1]) ? node36932 : node36921;
													assign node36921 = (inp[5]) ? node36923 : 4'b1101;
														assign node36923 = (inp[2]) ? node36929 : node36924;
															assign node36924 = (inp[15]) ? 4'b1101 : node36925;
																assign node36925 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node36929 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node36932 = (inp[5]) ? node36940 : node36933;
														assign node36933 = (inp[15]) ? node36937 : node36934;
															assign node36934 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node36937 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node36940 = (inp[0]) ? node36942 : 4'b1101;
															assign node36942 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node36945 = (inp[0]) ? node36953 : node36946;
													assign node36946 = (inp[1]) ? 4'b1001 : node36947;
														assign node36947 = (inp[15]) ? 4'b1001 : node36948;
															assign node36948 = (inp[2]) ? 4'b1011 : 4'b1001;
													assign node36953 = (inp[15]) ? node36957 : node36954;
														assign node36954 = (inp[5]) ? 4'b1011 : 4'b1001;
														assign node36957 = (inp[5]) ? 4'b1001 : 4'b1011;
											assign node36960 = (inp[9]) ? node36994 : node36961;
												assign node36961 = (inp[2]) ? node36985 : node36962;
													assign node36962 = (inp[1]) ? node36972 : node36963;
														assign node36963 = (inp[5]) ? 4'b1001 : node36964;
															assign node36964 = (inp[0]) ? node36968 : node36965;
																assign node36965 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node36968 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node36972 = (inp[15]) ? node36978 : node36973;
															assign node36973 = (inp[0]) ? node36975 : 4'b1011;
																assign node36975 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node36978 = (inp[0]) ? node36982 : node36979;
																assign node36979 = (inp[5]) ? 4'b1011 : 4'b1001;
																assign node36982 = (inp[5]) ? 4'b1001 : 4'b1011;
													assign node36985 = (inp[15]) ? node36987 : 4'b1001;
														assign node36987 = (inp[0]) ? node36991 : node36988;
															assign node36988 = (inp[5]) ? 4'b1011 : 4'b1001;
															assign node36991 = (inp[5]) ? 4'b1001 : 4'b1011;
												assign node36994 = (inp[5]) ? node37002 : node36995;
													assign node36995 = (inp[0]) ? node36999 : node36996;
														assign node36996 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node36999 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node37002 = (inp[0]) ? 4'b1101 : node37003;
														assign node37003 = (inp[15]) ? 4'b1111 : 4'b1101;
										assign node37007 = (inp[0]) ? node37043 : node37008;
											assign node37008 = (inp[15]) ? node37028 : node37009;
												assign node37009 = (inp[5]) ? node37015 : node37010;
													assign node37010 = (inp[4]) ? 4'b0101 : node37011;
														assign node37011 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node37015 = (inp[1]) ? node37021 : node37016;
														assign node37016 = (inp[9]) ? node37018 : 4'b0101;
															assign node37018 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node37021 = (inp[4]) ? node37025 : node37022;
															assign node37022 = (inp[9]) ? 4'b0001 : 4'b0101;
															assign node37025 = (inp[9]) ? 4'b0101 : 4'b0001;
												assign node37028 = (inp[5]) ? node37036 : node37029;
													assign node37029 = (inp[9]) ? node37033 : node37030;
														assign node37030 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node37033 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node37036 = (inp[4]) ? node37040 : node37037;
														assign node37037 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node37040 = (inp[9]) ? 4'b0111 : 4'b0011;
											assign node37043 = (inp[15]) ? node37061 : node37044;
												assign node37044 = (inp[5]) ? node37050 : node37045;
													assign node37045 = (inp[2]) ? node37047 : 4'b0001;
														assign node37047 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node37050 = (inp[1]) ? node37054 : node37051;
														assign node37051 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node37054 = (inp[9]) ? node37058 : node37055;
															assign node37055 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37058 = (inp[2]) ? 4'b0011 : 4'b0111;
												assign node37061 = (inp[5]) ? node37067 : node37062;
													assign node37062 = (inp[4]) ? node37064 : 4'b0011;
														assign node37064 = (inp[9]) ? 4'b0101 : 4'b0011;
													assign node37067 = (inp[4]) ? node37071 : node37068;
														assign node37068 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node37071 = (inp[9]) ? 4'b0101 : 4'b0001;
							assign node37074 = (inp[1]) ? node37442 : node37075;
								assign node37075 = (inp[15]) ? node37275 : node37076;
									assign node37076 = (inp[0]) ? node37172 : node37077;
										assign node37077 = (inp[3]) ? node37129 : node37078;
											assign node37078 = (inp[5]) ? node37106 : node37079;
												assign node37079 = (inp[2]) ? node37097 : node37080;
													assign node37080 = (inp[9]) ? node37090 : node37081;
														assign node37081 = (inp[6]) ? node37087 : node37082;
															assign node37082 = (inp[11]) ? 4'b1011 : node37083;
																assign node37083 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37087 = (inp[4]) ? 4'b1111 : 4'b1011;
														assign node37090 = (inp[11]) ? node37094 : node37091;
															assign node37091 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node37094 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node37097 = (inp[9]) ? 4'b0011 : node37098;
														assign node37098 = (inp[11]) ? node37100 : 4'b0111;
															assign node37100 = (inp[4]) ? 4'b0111 : node37101;
																assign node37101 = (inp[6]) ? 4'b0011 : 4'b1011;
												assign node37106 = (inp[4]) ? node37120 : node37107;
													assign node37107 = (inp[9]) ? node37115 : node37108;
														assign node37108 = (inp[11]) ? node37112 : node37109;
															assign node37109 = (inp[6]) ? 4'b1011 : 4'b0111;
															assign node37112 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node37115 = (inp[6]) ? node37117 : 4'b0011;
															assign node37117 = (inp[11]) ? 4'b0101 : 4'b1101;
													assign node37120 = (inp[2]) ? node37126 : node37121;
														assign node37121 = (inp[6]) ? node37123 : 4'b1101;
															assign node37123 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node37126 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node37129 = (inp[9]) ? node37159 : node37130;
												assign node37130 = (inp[5]) ? node37146 : node37131;
													assign node37131 = (inp[4]) ? node37141 : node37132;
														assign node37132 = (inp[2]) ? node37138 : node37133;
															assign node37133 = (inp[6]) ? node37135 : 4'b1011;
																assign node37135 = (inp[11]) ? 4'b0011 : 4'b1011;
															assign node37138 = (inp[6]) ? 4'b0011 : 4'b0111;
														assign node37141 = (inp[6]) ? 4'b1101 : node37142;
															assign node37142 = (inp[11]) ? 4'b1101 : 4'b0011;
													assign node37146 = (inp[4]) ? node37154 : node37147;
														assign node37147 = (inp[11]) ? node37151 : node37148;
															assign node37148 = (inp[6]) ? 4'b1001 : 4'b0101;
															assign node37151 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node37154 = (inp[6]) ? node37156 : 4'b0001;
															assign node37156 = (inp[2]) ? 4'b0101 : 4'b1101;
												assign node37159 = (inp[4]) ? node37165 : node37160;
													assign node37160 = (inp[11]) ? node37162 : 4'b1101;
														assign node37162 = (inp[6]) ? 4'b0101 : 4'b1101;
													assign node37165 = (inp[6]) ? node37169 : node37166;
														assign node37166 = (inp[11]) ? 4'b1001 : 4'b0101;
														assign node37169 = (inp[11]) ? 4'b0001 : 4'b1001;
										assign node37172 = (inp[5]) ? node37218 : node37173;
											assign node37173 = (inp[3]) ? node37197 : node37174;
												assign node37174 = (inp[4]) ? node37184 : node37175;
													assign node37175 = (inp[9]) ? node37181 : node37176;
														assign node37176 = (inp[11]) ? node37178 : 4'b1001;
															assign node37178 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node37181 = (inp[6]) ? 4'b1101 : 4'b0001;
													assign node37184 = (inp[11]) ? node37190 : node37185;
														assign node37185 = (inp[6]) ? 4'b1001 : node37186;
															assign node37186 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node37190 = (inp[9]) ? node37194 : node37191;
															assign node37191 = (inp[6]) ? 4'b0101 : 4'b1101;
															assign node37194 = (inp[2]) ? 4'b0001 : 4'b1001;
												assign node37197 = (inp[9]) ? node37207 : node37198;
													assign node37198 = (inp[4]) ? node37202 : node37199;
														assign node37199 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node37202 = (inp[6]) ? node37204 : 4'b0001;
															assign node37204 = (inp[2]) ? 4'b0111 : 4'b1111;
													assign node37207 = (inp[6]) ? node37213 : node37208;
														assign node37208 = (inp[4]) ? node37210 : 4'b0001;
															assign node37210 = (inp[11]) ? 4'b1011 : 4'b0111;
														assign node37213 = (inp[11]) ? 4'b0111 : node37214;
															assign node37214 = (inp[4]) ? 4'b1011 : 4'b1111;
											assign node37218 = (inp[3]) ? node37246 : node37219;
												assign node37219 = (inp[4]) ? node37231 : node37220;
													assign node37220 = (inp[11]) ? node37224 : node37221;
														assign node37221 = (inp[9]) ? 4'b0001 : 4'b0101;
														assign node37224 = (inp[9]) ? node37228 : node37225;
															assign node37225 = (inp[6]) ? 4'b0001 : 4'b1001;
															assign node37228 = (inp[6]) ? 4'b0111 : 4'b1111;
													assign node37231 = (inp[9]) ? node37239 : node37232;
														assign node37232 = (inp[2]) ? 4'b1111 : node37233;
															assign node37233 = (inp[11]) ? node37235 : 4'b0001;
																assign node37235 = (inp[6]) ? 4'b0111 : 4'b1111;
														assign node37239 = (inp[6]) ? node37243 : node37240;
															assign node37240 = (inp[11]) ? 4'b1011 : 4'b0111;
															assign node37243 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node37246 = (inp[6]) ? node37262 : node37247;
													assign node37247 = (inp[11]) ? node37253 : node37248;
														assign node37248 = (inp[4]) ? 4'b0011 : node37249;
															assign node37249 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node37253 = (inp[2]) ? node37255 : 4'b1011;
															assign node37255 = (inp[4]) ? node37259 : node37256;
																assign node37256 = (inp[9]) ? 4'b1111 : 4'b1011;
																assign node37259 = (inp[9]) ? 4'b1011 : 4'b1111;
													assign node37262 = (inp[11]) ? node37268 : node37263;
														assign node37263 = (inp[4]) ? node37265 : 4'b1111;
															assign node37265 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node37268 = (inp[9]) ? node37272 : node37269;
															assign node37269 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node37272 = (inp[4]) ? 4'b0011 : 4'b0111;
									assign node37275 = (inp[0]) ? node37363 : node37276;
										assign node37276 = (inp[3]) ? node37312 : node37277;
											assign node37277 = (inp[5]) ? node37293 : node37278;
												assign node37278 = (inp[2]) ? node37288 : node37279;
													assign node37279 = (inp[9]) ? node37281 : 4'b0101;
														assign node37281 = (inp[4]) ? node37283 : 4'b1101;
															assign node37283 = (inp[6]) ? 4'b1001 : node37284;
																assign node37284 = (inp[11]) ? 4'b1001 : 4'b0101;
													assign node37288 = (inp[4]) ? node37290 : 4'b1001;
														assign node37290 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node37293 = (inp[9]) ? node37305 : node37294;
													assign node37294 = (inp[6]) ? node37298 : node37295;
														assign node37295 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node37298 = (inp[4]) ? node37302 : node37299;
															assign node37299 = (inp[11]) ? 4'b0001 : 4'b1001;
															assign node37302 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node37305 = (inp[4]) ? node37309 : node37306;
														assign node37306 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node37309 = (inp[6]) ? 4'b0011 : 4'b1011;
											assign node37312 = (inp[5]) ? node37328 : node37313;
												assign node37313 = (inp[4]) ? node37319 : node37314;
													assign node37314 = (inp[9]) ? node37316 : 4'b1001;
														assign node37316 = (inp[6]) ? 4'b1111 : 4'b0001;
													assign node37319 = (inp[9]) ? node37321 : 4'b1111;
														assign node37321 = (inp[6]) ? node37325 : node37322;
															assign node37322 = (inp[11]) ? 4'b1011 : 4'b0111;
															assign node37325 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node37328 = (inp[6]) ? node37350 : node37329;
													assign node37329 = (inp[11]) ? node37337 : node37330;
														assign node37330 = (inp[2]) ? 4'b0011 : node37331;
															assign node37331 = (inp[4]) ? 4'b0111 : node37332;
																assign node37332 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node37337 = (inp[2]) ? node37343 : node37338;
															assign node37338 = (inp[4]) ? 4'b1011 : node37339;
																assign node37339 = (inp[9]) ? 4'b1111 : 4'b1011;
															assign node37343 = (inp[9]) ? node37347 : node37344;
																assign node37344 = (inp[4]) ? 4'b1111 : 4'b1011;
																assign node37347 = (inp[4]) ? 4'b1011 : 4'b1111;
													assign node37350 = (inp[11]) ? node37354 : node37351;
														assign node37351 = (inp[9]) ? 4'b1011 : 4'b1111;
														assign node37354 = (inp[2]) ? node37356 : 4'b0011;
															assign node37356 = (inp[4]) ? node37360 : node37357;
																assign node37357 = (inp[9]) ? 4'b0111 : 4'b0011;
																assign node37360 = (inp[9]) ? 4'b0011 : 4'b0111;
										assign node37363 = (inp[5]) ? node37407 : node37364;
											assign node37364 = (inp[3]) ? node37386 : node37365;
												assign node37365 = (inp[9]) ? node37377 : node37366;
													assign node37366 = (inp[4]) ? node37368 : 4'b1011;
														assign node37368 = (inp[2]) ? 4'b1111 : node37369;
															assign node37369 = (inp[6]) ? node37373 : node37370;
																assign node37370 = (inp[11]) ? 4'b1111 : 4'b0011;
																assign node37373 = (inp[11]) ? 4'b0111 : 4'b1111;
													assign node37377 = (inp[11]) ? node37381 : node37378;
														assign node37378 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node37381 = (inp[6]) ? node37383 : 4'b1011;
															assign node37383 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node37386 = (inp[9]) ? node37396 : node37387;
													assign node37387 = (inp[4]) ? 4'b1101 : node37388;
														assign node37388 = (inp[11]) ? node37392 : node37389;
															assign node37389 = (inp[6]) ? 4'b1011 : 4'b0111;
															assign node37392 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node37396 = (inp[4]) ? node37402 : node37397;
														assign node37397 = (inp[6]) ? node37399 : 4'b1101;
															assign node37399 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node37402 = (inp[11]) ? node37404 : 4'b1001;
															assign node37404 = (inp[6]) ? 4'b0001 : 4'b1001;
											assign node37407 = (inp[4]) ? node37425 : node37408;
												assign node37408 = (inp[9]) ? node37418 : node37409;
													assign node37409 = (inp[3]) ? node37415 : node37410;
														assign node37410 = (inp[2]) ? 4'b1011 : node37411;
															assign node37411 = (inp[6]) ? 4'b0011 : 4'b1011;
														assign node37415 = (inp[6]) ? 4'b0001 : 4'b1001;
													assign node37418 = (inp[11]) ? 4'b1101 : node37419;
														assign node37419 = (inp[6]) ? 4'b1101 : node37420;
															assign node37420 = (inp[3]) ? 4'b0001 : 4'b0011;
												assign node37425 = (inp[11]) ? node37435 : node37426;
													assign node37426 = (inp[6]) ? node37432 : node37427;
														assign node37427 = (inp[9]) ? 4'b0101 : node37428;
															assign node37428 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node37432 = (inp[3]) ? 4'b1101 : 4'b1001;
													assign node37435 = (inp[6]) ? node37439 : node37436;
														assign node37436 = (inp[9]) ? 4'b1001 : 4'b1101;
														assign node37439 = (inp[9]) ? 4'b0001 : 4'b0101;
								assign node37442 = (inp[4]) ? node37578 : node37443;
									assign node37443 = (inp[9]) ? node37513 : node37444;
										assign node37444 = (inp[6]) ? node37480 : node37445;
											assign node37445 = (inp[11]) ? node37469 : node37446;
												assign node37446 = (inp[15]) ? node37458 : node37447;
													assign node37447 = (inp[0]) ? node37453 : node37448;
														assign node37448 = (inp[5]) ? node37450 : 4'b0111;
															assign node37450 = (inp[3]) ? 4'b0101 : 4'b0111;
														assign node37453 = (inp[3]) ? node37455 : 4'b0101;
															assign node37455 = (inp[5]) ? 4'b0111 : 4'b0101;
													assign node37458 = (inp[0]) ? node37464 : node37459;
														assign node37459 = (inp[5]) ? node37461 : 4'b0101;
															assign node37461 = (inp[3]) ? 4'b0111 : 4'b0101;
														assign node37464 = (inp[5]) ? node37466 : 4'b0111;
															assign node37466 = (inp[3]) ? 4'b0101 : 4'b0111;
												assign node37469 = (inp[15]) ? node37475 : node37470;
													assign node37470 = (inp[0]) ? node37472 : 4'b1011;
														assign node37472 = (inp[2]) ? 4'b1001 : 4'b1011;
													assign node37475 = (inp[5]) ? node37477 : 4'b1001;
														assign node37477 = (inp[2]) ? 4'b1011 : 4'b1001;
											assign node37480 = (inp[11]) ? node37494 : node37481;
												assign node37481 = (inp[0]) ? 4'b1011 : node37482;
													assign node37482 = (inp[15]) ? node37488 : node37483;
														assign node37483 = (inp[5]) ? node37485 : 4'b1011;
															assign node37485 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node37488 = (inp[3]) ? node37490 : 4'b1001;
															assign node37490 = (inp[5]) ? 4'b1011 : 4'b1001;
												assign node37494 = (inp[15]) ? node37508 : node37495;
													assign node37495 = (inp[0]) ? node37503 : node37496;
														assign node37496 = (inp[2]) ? node37498 : 4'b0011;
															assign node37498 = (inp[5]) ? node37500 : 4'b0011;
																assign node37500 = (inp[3]) ? 4'b0001 : 4'b0011;
														assign node37503 = (inp[5]) ? node37505 : 4'b0001;
															assign node37505 = (inp[3]) ? 4'b0011 : 4'b0001;
													assign node37508 = (inp[0]) ? 4'b0011 : node37509;
														assign node37509 = (inp[3]) ? 4'b0011 : 4'b0001;
										assign node37513 = (inp[6]) ? node37543 : node37514;
											assign node37514 = (inp[11]) ? node37530 : node37515;
												assign node37515 = (inp[15]) ? node37521 : node37516;
													assign node37516 = (inp[0]) ? 4'b0001 : node37517;
														assign node37517 = (inp[3]) ? 4'b0001 : 4'b0011;
													assign node37521 = (inp[0]) ? node37525 : node37522;
														assign node37522 = (inp[3]) ? 4'b0011 : 4'b0001;
														assign node37525 = (inp[3]) ? node37527 : 4'b0011;
															assign node37527 = (inp[5]) ? 4'b0001 : 4'b0011;
												assign node37530 = (inp[0]) ? node37534 : node37531;
													assign node37531 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node37534 = (inp[15]) ? node37540 : node37535;
														assign node37535 = (inp[5]) ? 4'b1111 : node37536;
															assign node37536 = (inp[2]) ? 4'b1101 : 4'b1111;
														assign node37540 = (inp[3]) ? 4'b1101 : 4'b1111;
											assign node37543 = (inp[11]) ? node37563 : node37544;
												assign node37544 = (inp[5]) ? node37556 : node37545;
													assign node37545 = (inp[3]) ? 4'b1111 : node37546;
														assign node37546 = (inp[2]) ? node37548 : 4'b1111;
															assign node37548 = (inp[15]) ? node37552 : node37549;
																assign node37549 = (inp[0]) ? 4'b1101 : 4'b1111;
																assign node37552 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node37556 = (inp[15]) ? node37560 : node37557;
														assign node37557 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node37560 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node37563 = (inp[5]) ? node37571 : node37564;
													assign node37564 = (inp[0]) ? 4'b0111 : node37565;
														assign node37565 = (inp[15]) ? node37567 : 4'b0111;
															assign node37567 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node37571 = (inp[15]) ? node37575 : node37572;
														assign node37572 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node37575 = (inp[0]) ? 4'b0101 : 4'b0111;
									assign node37578 = (inp[9]) ? node37660 : node37579;
										assign node37579 = (inp[11]) ? node37615 : node37580;
											assign node37580 = (inp[6]) ? node37594 : node37581;
												assign node37581 = (inp[0]) ? node37589 : node37582;
													assign node37582 = (inp[15]) ? 4'b0001 : node37583;
														assign node37583 = (inp[5]) ? node37585 : 4'b0011;
															assign node37585 = (inp[2]) ? 4'b0011 : 4'b0001;
													assign node37589 = (inp[15]) ? 4'b0011 : node37590;
														assign node37590 = (inp[3]) ? 4'b0011 : 4'b0001;
												assign node37594 = (inp[15]) ? node37604 : node37595;
													assign node37595 = (inp[2]) ? 4'b1111 : node37596;
														assign node37596 = (inp[3]) ? 4'b1101 : node37597;
															assign node37597 = (inp[0]) ? node37599 : 4'b1111;
																assign node37599 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node37604 = (inp[0]) ? node37610 : node37605;
														assign node37605 = (inp[5]) ? 4'b1111 : node37606;
															assign node37606 = (inp[2]) ? 4'b1101 : 4'b1111;
														assign node37610 = (inp[3]) ? 4'b1101 : node37611;
															assign node37611 = (inp[5]) ? 4'b1101 : 4'b1111;
											assign node37615 = (inp[6]) ? node37635 : node37616;
												assign node37616 = (inp[0]) ? node37628 : node37617;
													assign node37617 = (inp[15]) ? node37623 : node37618;
														assign node37618 = (inp[5]) ? 4'b1101 : node37619;
															assign node37619 = (inp[3]) ? 4'b1101 : 4'b1111;
														assign node37623 = (inp[5]) ? 4'b1111 : node37624;
															assign node37624 = (inp[3]) ? 4'b1111 : 4'b1101;
													assign node37628 = (inp[5]) ? 4'b1111 : node37629;
														assign node37629 = (inp[3]) ? 4'b1101 : node37630;
															assign node37630 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node37635 = (inp[2]) ? node37645 : node37636;
													assign node37636 = (inp[3]) ? 4'b0111 : node37637;
														assign node37637 = (inp[0]) ? node37639 : 4'b0111;
															assign node37639 = (inp[5]) ? 4'b0101 : node37640;
																assign node37640 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node37645 = (inp[0]) ? node37651 : node37646;
														assign node37646 = (inp[15]) ? node37648 : 4'b0101;
															assign node37648 = (inp[5]) ? 4'b0111 : 4'b0101;
														assign node37651 = (inp[5]) ? node37657 : node37652;
															assign node37652 = (inp[15]) ? 4'b0111 : node37653;
																assign node37653 = (inp[3]) ? 4'b0111 : 4'b0101;
															assign node37657 = (inp[15]) ? 4'b0101 : 4'b0111;
										assign node37660 = (inp[6]) ? node37686 : node37661;
											assign node37661 = (inp[11]) ? node37675 : node37662;
												assign node37662 = (inp[5]) ? node37666 : node37663;
													assign node37663 = (inp[3]) ? 4'b0111 : 4'b0101;
													assign node37666 = (inp[3]) ? 4'b0101 : node37667;
														assign node37667 = (inp[2]) ? node37669 : 4'b0111;
															assign node37669 = (inp[15]) ? 4'b0101 : node37670;
																assign node37670 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node37675 = (inp[0]) ? node37679 : node37676;
													assign node37676 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node37679 = (inp[15]) ? node37683 : node37680;
														assign node37680 = (inp[3]) ? 4'b1011 : 4'b1001;
														assign node37683 = (inp[3]) ? 4'b1001 : 4'b1011;
											assign node37686 = (inp[11]) ? node37704 : node37687;
												assign node37687 = (inp[0]) ? node37697 : node37688;
													assign node37688 = (inp[15]) ? node37694 : node37689;
														assign node37689 = (inp[5]) ? 4'b1001 : node37690;
															assign node37690 = (inp[3]) ? 4'b1001 : 4'b1011;
														assign node37694 = (inp[3]) ? 4'b1011 : 4'b1001;
													assign node37697 = (inp[15]) ? 4'b1001 : node37698;
														assign node37698 = (inp[5]) ? 4'b1011 : node37699;
															assign node37699 = (inp[3]) ? 4'b1011 : 4'b1001;
												assign node37704 = (inp[5]) ? node37714 : node37705;
													assign node37705 = (inp[3]) ? node37707 : 4'b0011;
														assign node37707 = (inp[0]) ? node37711 : node37708;
															assign node37708 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node37711 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node37714 = (inp[0]) ? node37716 : 4'b0001;
														assign node37716 = (inp[15]) ? 4'b0001 : 4'b0011;
						assign node37719 = (inp[3]) ? node38295 : node37720;
							assign node37720 = (inp[11]) ? node37990 : node37721;
								assign node37721 = (inp[6]) ? node37863 : node37722;
									assign node37722 = (inp[15]) ? node37796 : node37723;
										assign node37723 = (inp[0]) ? node37755 : node37724;
											assign node37724 = (inp[4]) ? node37742 : node37725;
												assign node37725 = (inp[5]) ? node37735 : node37726;
													assign node37726 = (inp[1]) ? 4'b0111 : node37727;
														assign node37727 = (inp[9]) ? node37731 : node37728;
															assign node37728 = (inp[10]) ? 4'b0011 : 4'b0111;
															assign node37731 = (inp[10]) ? 4'b0111 : 4'b0011;
													assign node37735 = (inp[9]) ? node37739 : node37736;
														assign node37736 = (inp[10]) ? 4'b0011 : 4'b0111;
														assign node37739 = (inp[10]) ? 4'b0101 : 4'b0011;
												assign node37742 = (inp[5]) ? node37750 : node37743;
													assign node37743 = (inp[1]) ? 4'b0111 : node37744;
														assign node37744 = (inp[9]) ? node37746 : 4'b0011;
															assign node37746 = (inp[10]) ? 4'b0011 : 4'b0111;
													assign node37750 = (inp[2]) ? node37752 : 4'b0101;
														assign node37752 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node37755 = (inp[5]) ? node37779 : node37756;
												assign node37756 = (inp[2]) ? node37772 : node37757;
													assign node37757 = (inp[10]) ? node37765 : node37758;
														assign node37758 = (inp[1]) ? 4'b0001 : node37759;
															assign node37759 = (inp[9]) ? node37761 : 4'b0101;
																assign node37761 = (inp[4]) ? 4'b0101 : 4'b0001;
														assign node37765 = (inp[4]) ? node37769 : node37766;
															assign node37766 = (inp[9]) ? 4'b0101 : 4'b0001;
															assign node37769 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node37772 = (inp[4]) ? node37774 : 4'b0001;
														assign node37774 = (inp[9]) ? node37776 : 4'b0101;
															assign node37776 = (inp[10]) ? 4'b0001 : 4'b0101;
												assign node37779 = (inp[4]) ? node37789 : node37780;
													assign node37780 = (inp[1]) ? node37784 : node37781;
														assign node37781 = (inp[2]) ? 4'b0111 : 4'b0001;
														assign node37784 = (inp[10]) ? 4'b0001 : node37785;
															assign node37785 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node37789 = (inp[9]) ? node37793 : node37790;
														assign node37790 = (inp[10]) ? 4'b0111 : 4'b0001;
														assign node37793 = (inp[10]) ? 4'b0011 : 4'b0111;
										assign node37796 = (inp[0]) ? node37822 : node37797;
											assign node37797 = (inp[5]) ? node37811 : node37798;
												assign node37798 = (inp[1]) ? 4'b0001 : node37799;
													assign node37799 = (inp[2]) ? node37801 : 4'b0001;
														assign node37801 = (inp[10]) ? 4'b0101 : node37802;
															assign node37802 = (inp[9]) ? node37806 : node37803;
																assign node37803 = (inp[4]) ? 4'b0001 : 4'b0101;
																assign node37806 = (inp[4]) ? 4'b0101 : 4'b0001;
												assign node37811 = (inp[9]) ? node37815 : node37812;
													assign node37812 = (inp[10]) ? 4'b0001 : 4'b0101;
													assign node37815 = (inp[1]) ? node37817 : 4'b0001;
														assign node37817 = (inp[4]) ? node37819 : 4'b0111;
															assign node37819 = (inp[10]) ? 4'b0011 : 4'b0111;
											assign node37822 = (inp[10]) ? node37854 : node37823;
												assign node37823 = (inp[5]) ? node37839 : node37824;
													assign node37824 = (inp[2]) ? node37832 : node37825;
														assign node37825 = (inp[1]) ? 4'b0111 : node37826;
															assign node37826 = (inp[9]) ? node37828 : 4'b0011;
																assign node37828 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node37832 = (inp[1]) ? 4'b0011 : node37833;
															assign node37833 = (inp[9]) ? 4'b0111 : node37834;
																assign node37834 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node37839 = (inp[2]) ? node37847 : node37840;
														assign node37840 = (inp[9]) ? node37844 : node37841;
															assign node37841 = (inp[4]) ? 4'b0011 : 4'b0111;
															assign node37844 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node37847 = (inp[1]) ? node37849 : 4'b0011;
															assign node37849 = (inp[9]) ? 4'b0011 : node37850;
																assign node37850 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node37854 = (inp[5]) ? node37856 : 4'b0011;
													assign node37856 = (inp[4]) ? node37860 : node37857;
														assign node37857 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node37860 = (inp[9]) ? 4'b0001 : 4'b0101;
									assign node37863 = (inp[9]) ? node37907 : node37864;
										assign node37864 = (inp[4]) ? node37872 : node37865;
											assign node37865 = (inp[15]) ? node37869 : node37866;
												assign node37866 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node37869 = (inp[0]) ? 4'b1011 : 4'b1001;
											assign node37872 = (inp[10]) ? node37894 : node37873;
												assign node37873 = (inp[0]) ? node37887 : node37874;
													assign node37874 = (inp[1]) ? node37880 : node37875;
														assign node37875 = (inp[5]) ? node37877 : 4'b1111;
															assign node37877 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node37880 = (inp[5]) ? node37884 : node37881;
															assign node37881 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node37884 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node37887 = (inp[5]) ? node37891 : node37888;
														assign node37888 = (inp[2]) ? 4'b1111 : 4'b1101;
														assign node37891 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node37894 = (inp[0]) ? node37900 : node37895;
													assign node37895 = (inp[5]) ? 4'b1101 : node37896;
														assign node37896 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node37900 = (inp[5]) ? node37904 : node37901;
														assign node37901 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node37904 = (inp[15]) ? 4'b1101 : 4'b1111;
										assign node37907 = (inp[4]) ? node37953 : node37908;
											assign node37908 = (inp[0]) ? node37934 : node37909;
												assign node37909 = (inp[2]) ? node37927 : node37910;
													assign node37910 = (inp[10]) ? node37920 : node37911;
														assign node37911 = (inp[1]) ? node37913 : 4'b1111;
															assign node37913 = (inp[15]) ? node37917 : node37914;
																assign node37914 = (inp[5]) ? 4'b1101 : 4'b1111;
																assign node37917 = (inp[5]) ? 4'b1111 : 4'b1101;
														assign node37920 = (inp[15]) ? node37924 : node37921;
															assign node37921 = (inp[5]) ? 4'b1101 : 4'b1111;
															assign node37924 = (inp[5]) ? 4'b1111 : 4'b1101;
													assign node37927 = (inp[15]) ? node37931 : node37928;
														assign node37928 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node37931 = (inp[5]) ? 4'b1111 : 4'b1101;
												assign node37934 = (inp[2]) ? node37946 : node37935;
													assign node37935 = (inp[1]) ? node37941 : node37936;
														assign node37936 = (inp[5]) ? node37938 : 4'b1111;
															assign node37938 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node37941 = (inp[5]) ? node37943 : 4'b1101;
															assign node37943 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node37946 = (inp[5]) ? node37950 : node37947;
														assign node37947 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node37950 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node37953 = (inp[5]) ? node37983 : node37954;
												assign node37954 = (inp[10]) ? node37972 : node37955;
													assign node37955 = (inp[2]) ? node37965 : node37956;
														assign node37956 = (inp[1]) ? node37958 : 4'b1011;
															assign node37958 = (inp[0]) ? node37962 : node37959;
																assign node37959 = (inp[15]) ? 4'b1001 : 4'b1011;
																assign node37962 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node37965 = (inp[0]) ? node37969 : node37966;
															assign node37966 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node37969 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node37972 = (inp[2]) ? node37978 : node37973;
														assign node37973 = (inp[15]) ? 4'b1001 : node37974;
															assign node37974 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node37978 = (inp[15]) ? 4'b1011 : node37979;
															assign node37979 = (inp[0]) ? 4'b1001 : 4'b1011;
												assign node37983 = (inp[15]) ? node37987 : node37984;
													assign node37984 = (inp[0]) ? 4'b1011 : 4'b1001;
													assign node37987 = (inp[0]) ? 4'b1001 : 4'b1011;
								assign node37990 = (inp[6]) ? node38168 : node37991;
									assign node37991 = (inp[10]) ? node38091 : node37992;
										assign node37992 = (inp[1]) ? node38036 : node37993;
											assign node37993 = (inp[9]) ? node38015 : node37994;
												assign node37994 = (inp[4]) ? node38002 : node37995;
													assign node37995 = (inp[0]) ? node37999 : node37996;
														assign node37996 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node37999 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node38002 = (inp[15]) ? node38008 : node38003;
														assign node38003 = (inp[0]) ? 4'b1101 : node38004;
															assign node38004 = (inp[5]) ? 4'b1101 : 4'b1111;
														assign node38008 = (inp[5]) ? node38012 : node38009;
															assign node38009 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node38012 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node38015 = (inp[4]) ? node38031 : node38016;
													assign node38016 = (inp[5]) ? node38022 : node38017;
														assign node38017 = (inp[0]) ? node38019 : 4'b1101;
															assign node38019 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node38022 = (inp[2]) ? node38028 : node38023;
															assign node38023 = (inp[15]) ? node38025 : 4'b1101;
																assign node38025 = (inp[0]) ? 4'b1101 : 4'b1111;
															assign node38028 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node38031 = (inp[15]) ? 4'b1001 : node38032;
														assign node38032 = (inp[2]) ? 4'b1001 : 4'b1011;
											assign node38036 = (inp[15]) ? node38068 : node38037;
												assign node38037 = (inp[0]) ? node38055 : node38038;
													assign node38038 = (inp[5]) ? node38050 : node38039;
														assign node38039 = (inp[2]) ? node38045 : node38040;
															assign node38040 = (inp[4]) ? node38042 : 4'b1011;
																assign node38042 = (inp[9]) ? 4'b1011 : 4'b1111;
															assign node38045 = (inp[9]) ? node38047 : 4'b1111;
																assign node38047 = (inp[4]) ? 4'b1011 : 4'b1111;
														assign node38050 = (inp[4]) ? node38052 : 4'b1011;
															assign node38052 = (inp[2]) ? 4'b1001 : 4'b1101;
													assign node38055 = (inp[5]) ? node38061 : node38056;
														assign node38056 = (inp[4]) ? 4'b1101 : node38057;
															assign node38057 = (inp[9]) ? 4'b1101 : 4'b1001;
														assign node38061 = (inp[2]) ? 4'b1111 : node38062;
															assign node38062 = (inp[9]) ? node38064 : 4'b1001;
																assign node38064 = (inp[4]) ? 4'b1011 : 4'b1111;
												assign node38068 = (inp[0]) ? node38080 : node38069;
													assign node38069 = (inp[5]) ? node38077 : node38070;
														assign node38070 = (inp[9]) ? node38074 : node38071;
															assign node38071 = (inp[4]) ? 4'b1101 : 4'b1001;
															assign node38074 = (inp[4]) ? 4'b1001 : 4'b1101;
														assign node38077 = (inp[9]) ? 4'b1011 : 4'b1001;
													assign node38080 = (inp[5]) ? node38086 : node38081;
														assign node38081 = (inp[4]) ? 4'b1011 : node38082;
															assign node38082 = (inp[9]) ? 4'b1111 : 4'b1011;
														assign node38086 = (inp[2]) ? node38088 : 4'b1011;
															assign node38088 = (inp[4]) ? 4'b1001 : 4'b1101;
										assign node38091 = (inp[4]) ? node38127 : node38092;
											assign node38092 = (inp[9]) ? node38102 : node38093;
												assign node38093 = (inp[1]) ? 4'b1011 : node38094;
													assign node38094 = (inp[0]) ? node38098 : node38095;
														assign node38095 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node38098 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node38102 = (inp[1]) ? node38110 : node38103;
													assign node38103 = (inp[0]) ? 4'b1111 : node38104;
														assign node38104 = (inp[2]) ? node38106 : 4'b1101;
															assign node38106 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node38110 = (inp[15]) ? node38116 : node38111;
														assign node38111 = (inp[5]) ? 4'b1101 : node38112;
															assign node38112 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node38116 = (inp[2]) ? node38122 : node38117;
															assign node38117 = (inp[5]) ? 4'b1111 : node38118;
																assign node38118 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node38122 = (inp[5]) ? node38124 : 4'b1111;
																assign node38124 = (inp[0]) ? 4'b1101 : 4'b1111;
											assign node38127 = (inp[9]) ? node38147 : node38128;
												assign node38128 = (inp[1]) ? node38138 : node38129;
													assign node38129 = (inp[0]) ? node38133 : node38130;
														assign node38130 = (inp[2]) ? 4'b1101 : 4'b1111;
														assign node38133 = (inp[5]) ? node38135 : 4'b1111;
															assign node38135 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node38138 = (inp[5]) ? node38140 : 4'b1111;
														assign node38140 = (inp[15]) ? node38144 : node38141;
															assign node38141 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node38144 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node38147 = (inp[5]) ? node38163 : node38148;
													assign node38148 = (inp[2]) ? node38152 : node38149;
														assign node38149 = (inp[1]) ? 4'b1011 : 4'b1001;
														assign node38152 = (inp[1]) ? node38158 : node38153;
															assign node38153 = (inp[15]) ? node38155 : 4'b1011;
																assign node38155 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node38158 = (inp[0]) ? 4'b1001 : node38159;
																assign node38159 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node38163 = (inp[0]) ? 4'b1001 : node38164;
														assign node38164 = (inp[15]) ? 4'b1011 : 4'b1001;
									assign node38168 = (inp[10]) ? node38234 : node38169;
										assign node38169 = (inp[15]) ? node38205 : node38170;
											assign node38170 = (inp[5]) ? node38190 : node38171;
												assign node38171 = (inp[0]) ? node38187 : node38172;
													assign node38172 = (inp[2]) ? node38180 : node38173;
														assign node38173 = (inp[4]) ? node38177 : node38174;
															assign node38174 = (inp[9]) ? 4'b0111 : 4'b0011;
															assign node38177 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node38180 = (inp[4]) ? node38184 : node38181;
															assign node38181 = (inp[1]) ? 4'b0111 : 4'b0011;
															assign node38184 = (inp[9]) ? 4'b0011 : 4'b0111;
													assign node38187 = (inp[1]) ? 4'b0101 : 4'b0001;
												assign node38190 = (inp[0]) ? node38198 : node38191;
													assign node38191 = (inp[9]) ? node38195 : node38192;
														assign node38192 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node38195 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node38198 = (inp[4]) ? node38202 : node38199;
														assign node38199 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node38202 = (inp[9]) ? 4'b0011 : 4'b0111;
											assign node38205 = (inp[4]) ? node38225 : node38206;
												assign node38206 = (inp[9]) ? node38210 : node38207;
													assign node38207 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node38210 = (inp[2]) ? node38218 : node38211;
														assign node38211 = (inp[0]) ? node38215 : node38212;
															assign node38212 = (inp[5]) ? 4'b0111 : 4'b0101;
															assign node38215 = (inp[5]) ? 4'b0101 : 4'b0111;
														assign node38218 = (inp[0]) ? node38222 : node38219;
															assign node38219 = (inp[1]) ? 4'b0111 : 4'b0101;
															assign node38222 = (inp[5]) ? 4'b0101 : 4'b0111;
												assign node38225 = (inp[9]) ? 4'b0011 : node38226;
													assign node38226 = (inp[5]) ? node38230 : node38227;
														assign node38227 = (inp[0]) ? 4'b0111 : 4'b0101;
														assign node38230 = (inp[0]) ? 4'b0101 : 4'b0111;
										assign node38234 = (inp[0]) ? node38262 : node38235;
											assign node38235 = (inp[15]) ? node38253 : node38236;
												assign node38236 = (inp[5]) ? node38246 : node38237;
													assign node38237 = (inp[1]) ? node38239 : 4'b0111;
														assign node38239 = (inp[9]) ? node38243 : node38240;
															assign node38240 = (inp[4]) ? 4'b0111 : 4'b0011;
															assign node38243 = (inp[2]) ? 4'b0011 : 4'b0111;
													assign node38246 = (inp[4]) ? node38250 : node38247;
														assign node38247 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node38250 = (inp[9]) ? 4'b0001 : 4'b0101;
												assign node38253 = (inp[4]) ? node38257 : node38254;
													assign node38254 = (inp[9]) ? 4'b0101 : 4'b0001;
													assign node38257 = (inp[5]) ? 4'b0111 : node38258;
														assign node38258 = (inp[9]) ? 4'b0001 : 4'b0101;
											assign node38262 = (inp[15]) ? node38278 : node38263;
												assign node38263 = (inp[5]) ? node38271 : node38264;
													assign node38264 = (inp[4]) ? node38268 : node38265;
														assign node38265 = (inp[9]) ? 4'b0101 : 4'b0001;
														assign node38268 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node38271 = (inp[9]) ? node38275 : node38272;
														assign node38272 = (inp[4]) ? 4'b0111 : 4'b0001;
														assign node38275 = (inp[4]) ? 4'b0011 : 4'b0111;
												assign node38278 = (inp[5]) ? node38286 : node38279;
													assign node38279 = (inp[9]) ? node38283 : node38280;
														assign node38280 = (inp[4]) ? 4'b0111 : 4'b0011;
														assign node38283 = (inp[4]) ? 4'b0011 : 4'b0111;
													assign node38286 = (inp[2]) ? node38288 : 4'b0011;
														assign node38288 = (inp[9]) ? node38292 : node38289;
															assign node38289 = (inp[4]) ? 4'b0101 : 4'b0011;
															assign node38292 = (inp[4]) ? 4'b0001 : 4'b0101;
							assign node38295 = (inp[5]) ? node38661 : node38296;
								assign node38296 = (inp[1]) ? node38502 : node38297;
									assign node38297 = (inp[10]) ? node38403 : node38298;
										assign node38298 = (inp[15]) ? node38348 : node38299;
											assign node38299 = (inp[6]) ? node38325 : node38300;
												assign node38300 = (inp[11]) ? node38316 : node38301;
													assign node38301 = (inp[0]) ? node38309 : node38302;
														assign node38302 = (inp[4]) ? node38306 : node38303;
															assign node38303 = (inp[9]) ? 4'b0011 : 4'b0111;
															assign node38306 = (inp[9]) ? 4'b0101 : 4'b0011;
														assign node38309 = (inp[9]) ? node38313 : node38310;
															assign node38310 = (inp[4]) ? 4'b0001 : 4'b0101;
															assign node38313 = (inp[4]) ? 4'b0111 : 4'b0001;
													assign node38316 = (inp[4]) ? node38322 : node38317;
														assign node38317 = (inp[9]) ? 4'b1111 : node38318;
															assign node38318 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node38322 = (inp[9]) ? 4'b1001 : 4'b1101;
												assign node38325 = (inp[11]) ? node38335 : node38326;
													assign node38326 = (inp[0]) ? node38332 : node38327;
														assign node38327 = (inp[9]) ? 4'b1101 : node38328;
															assign node38328 = (inp[4]) ? 4'b1101 : 4'b1011;
														assign node38332 = (inp[4]) ? 4'b1011 : 4'b1001;
													assign node38335 = (inp[0]) ? node38343 : node38336;
														assign node38336 = (inp[2]) ? node38338 : 4'b0101;
															assign node38338 = (inp[9]) ? node38340 : 4'b0101;
																assign node38340 = (inp[4]) ? 4'b0001 : 4'b0101;
														assign node38343 = (inp[2]) ? 4'b0111 : node38344;
															assign node38344 = (inp[9]) ? 4'b0111 : 4'b0001;
											assign node38348 = (inp[0]) ? node38374 : node38349;
												assign node38349 = (inp[9]) ? node38361 : node38350;
													assign node38350 = (inp[4]) ? node38356 : node38351;
														assign node38351 = (inp[6]) ? node38353 : 4'b0101;
															assign node38353 = (inp[11]) ? 4'b0001 : 4'b1001;
														assign node38356 = (inp[6]) ? 4'b1111 : node38357;
															assign node38357 = (inp[11]) ? 4'b1111 : 4'b0001;
													assign node38361 = (inp[4]) ? node38367 : node38362;
														assign node38362 = (inp[6]) ? node38364 : 4'b1111;
															assign node38364 = (inp[11]) ? 4'b0111 : 4'b1111;
														assign node38367 = (inp[6]) ? node38371 : node38368;
															assign node38368 = (inp[11]) ? 4'b1011 : 4'b0111;
															assign node38371 = (inp[11]) ? 4'b0011 : 4'b1011;
												assign node38374 = (inp[9]) ? node38388 : node38375;
													assign node38375 = (inp[4]) ? node38383 : node38376;
														assign node38376 = (inp[6]) ? node38380 : node38377;
															assign node38377 = (inp[11]) ? 4'b1011 : 4'b0111;
															assign node38380 = (inp[11]) ? 4'b0011 : 4'b1011;
														assign node38383 = (inp[11]) ? 4'b1101 : node38384;
															assign node38384 = (inp[6]) ? 4'b1101 : 4'b0011;
													assign node38388 = (inp[4]) ? node38396 : node38389;
														assign node38389 = (inp[2]) ? 4'b0101 : node38390;
															assign node38390 = (inp[6]) ? node38392 : 4'b1101;
																assign node38392 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node38396 = (inp[11]) ? node38400 : node38397;
															assign node38397 = (inp[2]) ? 4'b1001 : 4'b0101;
															assign node38400 = (inp[6]) ? 4'b0001 : 4'b1001;
										assign node38403 = (inp[9]) ? node38449 : node38404;
											assign node38404 = (inp[4]) ? node38422 : node38405;
												assign node38405 = (inp[15]) ? node38415 : node38406;
													assign node38406 = (inp[2]) ? 4'b0011 : node38407;
														assign node38407 = (inp[6]) ? node38411 : node38408;
															assign node38408 = (inp[11]) ? 4'b1011 : 4'b0011;
															assign node38411 = (inp[11]) ? 4'b0011 : 4'b1011;
													assign node38415 = (inp[0]) ? node38417 : 4'b1001;
														assign node38417 = (inp[6]) ? 4'b1011 : node38418;
															assign node38418 = (inp[11]) ? 4'b1011 : 4'b0011;
												assign node38422 = (inp[11]) ? node38438 : node38423;
													assign node38423 = (inp[6]) ? node38431 : node38424;
														assign node38424 = (inp[2]) ? 4'b0111 : node38425;
															assign node38425 = (inp[0]) ? 4'b0101 : node38426;
																assign node38426 = (inp[15]) ? 4'b0111 : 4'b0101;
														assign node38431 = (inp[15]) ? node38435 : node38432;
															assign node38432 = (inp[0]) ? 4'b1111 : 4'b1101;
															assign node38435 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node38438 = (inp[6]) ? node38440 : 4'b1111;
														assign node38440 = (inp[2]) ? node38446 : node38441;
															assign node38441 = (inp[15]) ? 4'b0111 : node38442;
																assign node38442 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node38446 = (inp[15]) ? 4'b0101 : 4'b0111;
											assign node38449 = (inp[4]) ? node38485 : node38450;
												assign node38450 = (inp[2]) ? node38476 : node38451;
													assign node38451 = (inp[11]) ? node38463 : node38452;
														assign node38452 = (inp[6]) ? node38458 : node38453;
															assign node38453 = (inp[15]) ? 4'b0111 : node38454;
																assign node38454 = (inp[0]) ? 4'b0111 : 4'b0101;
															assign node38458 = (inp[0]) ? 4'b1111 : node38459;
																assign node38459 = (inp[15]) ? 4'b1111 : 4'b1101;
														assign node38463 = (inp[6]) ? node38471 : node38464;
															assign node38464 = (inp[0]) ? node38468 : node38465;
																assign node38465 = (inp[15]) ? 4'b1111 : 4'b1101;
																assign node38468 = (inp[15]) ? 4'b1101 : 4'b1111;
															assign node38471 = (inp[0]) ? node38473 : 4'b0111;
																assign node38473 = (inp[15]) ? 4'b0101 : 4'b0111;
													assign node38476 = (inp[15]) ? node38482 : node38477;
														assign node38477 = (inp[6]) ? node38479 : 4'b0101;
															assign node38479 = (inp[11]) ? 4'b0101 : 4'b1101;
														assign node38482 = (inp[0]) ? 4'b0101 : 4'b0111;
												assign node38485 = (inp[15]) ? node38495 : node38486;
													assign node38486 = (inp[0]) ? node38490 : node38487;
														assign node38487 = (inp[2]) ? 4'b1001 : 4'b0001;
														assign node38490 = (inp[11]) ? node38492 : 4'b1011;
															assign node38492 = (inp[6]) ? 4'b0011 : 4'b1011;
													assign node38495 = (inp[0]) ? node38497 : 4'b1011;
														assign node38497 = (inp[11]) ? node38499 : 4'b1001;
															assign node38499 = (inp[6]) ? 4'b0001 : 4'b1001;
									assign node38502 = (inp[6]) ? node38594 : node38503;
										assign node38503 = (inp[11]) ? node38549 : node38504;
											assign node38504 = (inp[4]) ? node38528 : node38505;
												assign node38505 = (inp[10]) ? node38515 : node38506;
													assign node38506 = (inp[9]) ? node38508 : 4'b0111;
														assign node38508 = (inp[15]) ? node38512 : node38509;
															assign node38509 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node38512 = (inp[0]) ? 4'b0011 : 4'b0001;
													assign node38515 = (inp[9]) ? node38521 : node38516;
														assign node38516 = (inp[0]) ? 4'b0011 : node38517;
															assign node38517 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node38521 = (inp[0]) ? node38525 : node38522;
															assign node38522 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node38525 = (inp[15]) ? 4'b0101 : 4'b0111;
												assign node38528 = (inp[15]) ? node38544 : node38529;
													assign node38529 = (inp[2]) ? node38537 : node38530;
														assign node38530 = (inp[10]) ? node38534 : node38531;
															assign node38531 = (inp[0]) ? 4'b0001 : 4'b0101;
															assign node38534 = (inp[9]) ? 4'b0011 : 4'b0111;
														assign node38537 = (inp[10]) ? node38541 : node38538;
															assign node38538 = (inp[0]) ? 4'b0001 : 4'b0011;
															assign node38541 = (inp[9]) ? 4'b0001 : 4'b0101;
													assign node38544 = (inp[0]) ? 4'b0001 : node38545;
														assign node38545 = (inp[9]) ? 4'b0011 : 4'b0001;
											assign node38549 = (inp[9]) ? node38569 : node38550;
												assign node38550 = (inp[4]) ? node38558 : node38551;
													assign node38551 = (inp[0]) ? node38555 : node38552;
														assign node38552 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node38555 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node38558 = (inp[2]) ? node38564 : node38559;
														assign node38559 = (inp[10]) ? node38561 : 4'b1101;
															assign node38561 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node38564 = (inp[0]) ? 4'b1101 : node38565;
															assign node38565 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node38569 = (inp[4]) ? node38577 : node38570;
													assign node38570 = (inp[10]) ? node38574 : node38571;
														assign node38571 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node38574 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node38577 = (inp[10]) ? node38585 : node38578;
														assign node38578 = (inp[15]) ? node38582 : node38579;
															assign node38579 = (inp[0]) ? 4'b1011 : 4'b1001;
															assign node38582 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node38585 = (inp[2]) ? node38589 : node38586;
															assign node38586 = (inp[0]) ? 4'b1001 : 4'b1011;
															assign node38589 = (inp[0]) ? node38591 : 4'b1001;
																assign node38591 = (inp[15]) ? 4'b1001 : 4'b1011;
										assign node38594 = (inp[11]) ? node38632 : node38595;
											assign node38595 = (inp[4]) ? node38611 : node38596;
												assign node38596 = (inp[9]) ? node38604 : node38597;
													assign node38597 = (inp[0]) ? node38601 : node38598;
														assign node38598 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node38601 = (inp[15]) ? 4'b1011 : 4'b1001;
													assign node38604 = (inp[15]) ? node38608 : node38605;
														assign node38605 = (inp[0]) ? 4'b1111 : 4'b1101;
														assign node38608 = (inp[0]) ? 4'b1101 : 4'b1111;
												assign node38611 = (inp[9]) ? node38625 : node38612;
													assign node38612 = (inp[2]) ? node38618 : node38613;
														assign node38613 = (inp[0]) ? node38615 : 4'b1101;
															assign node38615 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node38618 = (inp[0]) ? node38622 : node38619;
															assign node38619 = (inp[15]) ? 4'b1111 : 4'b1101;
															assign node38622 = (inp[15]) ? 4'b1101 : 4'b1111;
													assign node38625 = (inp[2]) ? 4'b1011 : node38626;
														assign node38626 = (inp[0]) ? 4'b1001 : node38627;
															assign node38627 = (inp[15]) ? 4'b1011 : 4'b1001;
											assign node38632 = (inp[0]) ? node38648 : node38633;
												assign node38633 = (inp[15]) ? node38641 : node38634;
													assign node38634 = (inp[9]) ? node38638 : node38635;
														assign node38635 = (inp[4]) ? 4'b0101 : 4'b0011;
														assign node38638 = (inp[4]) ? 4'b0001 : 4'b0101;
													assign node38641 = (inp[4]) ? node38645 : node38642;
														assign node38642 = (inp[9]) ? 4'b0111 : 4'b0001;
														assign node38645 = (inp[9]) ? 4'b0011 : 4'b0111;
												assign node38648 = (inp[9]) ? node38654 : node38649;
													assign node38649 = (inp[4]) ? 4'b0101 : node38650;
														assign node38650 = (inp[15]) ? 4'b0011 : 4'b0001;
													assign node38654 = (inp[4]) ? node38658 : node38655;
														assign node38655 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node38658 = (inp[15]) ? 4'b0001 : 4'b0011;
								assign node38661 = (inp[4]) ? node38789 : node38662;
									assign node38662 = (inp[9]) ? node38718 : node38663;
										assign node38663 = (inp[6]) ? node38697 : node38664;
											assign node38664 = (inp[11]) ? node38678 : node38665;
												assign node38665 = (inp[10]) ? node38671 : node38666;
													assign node38666 = (inp[0]) ? 4'b0111 : node38667;
														assign node38667 = (inp[2]) ? 4'b0111 : 4'b0101;
													assign node38671 = (inp[15]) ? node38675 : node38672;
														assign node38672 = (inp[0]) ? 4'b0011 : 4'b0001;
														assign node38675 = (inp[0]) ? 4'b0001 : 4'b0011;
												assign node38678 = (inp[1]) ? node38690 : node38679;
													assign node38679 = (inp[10]) ? node38685 : node38680;
														assign node38680 = (inp[15]) ? node38682 : 4'b1001;
															assign node38682 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node38685 = (inp[0]) ? node38687 : 4'b1011;
															assign node38687 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node38690 = (inp[15]) ? node38694 : node38691;
														assign node38691 = (inp[0]) ? 4'b1011 : 4'b1001;
														assign node38694 = (inp[0]) ? 4'b1001 : 4'b1011;
											assign node38697 = (inp[11]) ? node38703 : node38698;
												assign node38698 = (inp[0]) ? 4'b1001 : node38699;
													assign node38699 = (inp[15]) ? 4'b1011 : 4'b1001;
												assign node38703 = (inp[1]) ? node38711 : node38704;
													assign node38704 = (inp[0]) ? node38708 : node38705;
														assign node38705 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node38708 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node38711 = (inp[0]) ? node38715 : node38712;
														assign node38712 = (inp[15]) ? 4'b0011 : 4'b0001;
														assign node38715 = (inp[15]) ? 4'b0001 : 4'b0011;
										assign node38718 = (inp[6]) ? node38762 : node38719;
											assign node38719 = (inp[11]) ? node38743 : node38720;
												assign node38720 = (inp[10]) ? node38738 : node38721;
													assign node38721 = (inp[1]) ? node38729 : node38722;
														assign node38722 = (inp[0]) ? node38726 : node38723;
															assign node38723 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node38726 = (inp[15]) ? 4'b0001 : 4'b0011;
														assign node38729 = (inp[2]) ? 4'b0011 : node38730;
															assign node38730 = (inp[0]) ? node38734 : node38731;
																assign node38731 = (inp[15]) ? 4'b0011 : 4'b0001;
																assign node38734 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node38738 = (inp[0]) ? 4'b0111 : node38739;
														assign node38739 = (inp[15]) ? 4'b0111 : 4'b0101;
												assign node38743 = (inp[1]) ? node38749 : node38744;
													assign node38744 = (inp[15]) ? node38746 : 4'b1111;
														assign node38746 = (inp[10]) ? 4'b1101 : 4'b1111;
													assign node38749 = (inp[10]) ? node38755 : node38750;
														assign node38750 = (inp[15]) ? node38752 : 4'b1101;
															assign node38752 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node38755 = (inp[2]) ? node38757 : 4'b1101;
															assign node38757 = (inp[0]) ? node38759 : 4'b1111;
																assign node38759 = (inp[15]) ? 4'b1101 : 4'b1111;
											assign node38762 = (inp[11]) ? node38770 : node38763;
												assign node38763 = (inp[0]) ? node38767 : node38764;
													assign node38764 = (inp[15]) ? 4'b1111 : 4'b1101;
													assign node38767 = (inp[15]) ? 4'b1101 : 4'b1111;
												assign node38770 = (inp[1]) ? node38776 : node38771;
													assign node38771 = (inp[0]) ? 4'b0101 : node38772;
														assign node38772 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node38776 = (inp[10]) ? node38784 : node38777;
														assign node38777 = (inp[0]) ? node38781 : node38778;
															assign node38778 = (inp[15]) ? 4'b0111 : 4'b0101;
															assign node38781 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node38784 = (inp[15]) ? node38786 : 4'b0111;
															assign node38786 = (inp[2]) ? 4'b0101 : 4'b0111;
									assign node38789 = (inp[9]) ? node38859 : node38790;
										assign node38790 = (inp[11]) ? node38824 : node38791;
											assign node38791 = (inp[6]) ? node38807 : node38792;
												assign node38792 = (inp[10]) ? node38804 : node38793;
													assign node38793 = (inp[1]) ? node38799 : node38794;
														assign node38794 = (inp[15]) ? node38796 : 4'b0001;
															assign node38796 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node38799 = (inp[0]) ? node38801 : 4'b0011;
															assign node38801 = (inp[15]) ? 4'b0001 : 4'b0011;
													assign node38804 = (inp[0]) ? 4'b0111 : 4'b0101;
												assign node38807 = (inp[10]) ? node38813 : node38808;
													assign node38808 = (inp[15]) ? node38810 : 4'b1111;
														assign node38810 = (inp[0]) ? 4'b1101 : 4'b1111;
													assign node38813 = (inp[1]) ? node38819 : node38814;
														assign node38814 = (inp[15]) ? node38816 : 4'b1101;
															assign node38816 = (inp[0]) ? 4'b1101 : 4'b1111;
														assign node38819 = (inp[0]) ? 4'b1111 : node38820;
															assign node38820 = (inp[15]) ? 4'b1111 : 4'b1101;
											assign node38824 = (inp[6]) ? node38844 : node38825;
												assign node38825 = (inp[1]) ? node38837 : node38826;
													assign node38826 = (inp[10]) ? node38832 : node38827;
														assign node38827 = (inp[0]) ? node38829 : 4'b1111;
															assign node38829 = (inp[15]) ? 4'b1101 : 4'b1111;
														assign node38832 = (inp[2]) ? 4'b1111 : node38833;
															assign node38833 = (inp[0]) ? 4'b1111 : 4'b1101;
													assign node38837 = (inp[10]) ? node38839 : 4'b1101;
														assign node38839 = (inp[2]) ? 4'b1101 : node38840;
															assign node38840 = (inp[15]) ? 4'b1111 : 4'b1101;
												assign node38844 = (inp[1]) ? node38846 : 4'b0101;
													assign node38846 = (inp[10]) ? node38848 : 4'b0101;
														assign node38848 = (inp[2]) ? node38854 : node38849;
															assign node38849 = (inp[0]) ? node38851 : 4'b0101;
																assign node38851 = (inp[15]) ? 4'b0101 : 4'b0111;
															assign node38854 = (inp[0]) ? 4'b0101 : node38855;
																assign node38855 = (inp[15]) ? 4'b0111 : 4'b0101;
										assign node38859 = (inp[10]) ? node38903 : node38860;
											assign node38860 = (inp[11]) ? node38886 : node38861;
												assign node38861 = (inp[6]) ? node38875 : node38862;
													assign node38862 = (inp[1]) ? node38870 : node38863;
														assign node38863 = (inp[2]) ? node38865 : 4'b0111;
															assign node38865 = (inp[0]) ? node38867 : 4'b0101;
																assign node38867 = (inp[15]) ? 4'b0101 : 4'b0111;
														assign node38870 = (inp[0]) ? 4'b0101 : node38871;
															assign node38871 = (inp[15]) ? 4'b0111 : 4'b0101;
													assign node38875 = (inp[2]) ? node38881 : node38876;
														assign node38876 = (inp[0]) ? node38878 : 4'b1001;
															assign node38878 = (inp[15]) ? 4'b1001 : 4'b1011;
														assign node38881 = (inp[0]) ? node38883 : 4'b1011;
															assign node38883 = (inp[15]) ? 4'b1001 : 4'b1011;
												assign node38886 = (inp[6]) ? node38894 : node38887;
													assign node38887 = (inp[0]) ? node38891 : node38888;
														assign node38888 = (inp[15]) ? 4'b1011 : 4'b1001;
														assign node38891 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node38894 = (inp[1]) ? node38896 : 4'b0011;
														assign node38896 = (inp[15]) ? node38900 : node38897;
															assign node38897 = (inp[0]) ? 4'b0011 : 4'b0001;
															assign node38900 = (inp[0]) ? 4'b0001 : 4'b0011;
											assign node38903 = (inp[1]) ? node38933 : node38904;
												assign node38904 = (inp[15]) ? node38920 : node38905;
													assign node38905 = (inp[0]) ? node38913 : node38906;
														assign node38906 = (inp[11]) ? node38910 : node38907;
															assign node38907 = (inp[6]) ? 4'b1001 : 4'b0001;
															assign node38910 = (inp[6]) ? 4'b0001 : 4'b1001;
														assign node38913 = (inp[2]) ? 4'b1011 : node38914;
															assign node38914 = (inp[6]) ? 4'b1011 : node38915;
																assign node38915 = (inp[11]) ? 4'b1011 : 4'b0011;
													assign node38920 = (inp[0]) ? node38926 : node38921;
														assign node38921 = (inp[11]) ? 4'b1011 : node38922;
															assign node38922 = (inp[6]) ? 4'b1011 : 4'b0011;
														assign node38926 = (inp[6]) ? node38930 : node38927;
															assign node38927 = (inp[11]) ? 4'b1001 : 4'b0001;
															assign node38930 = (inp[11]) ? 4'b0001 : 4'b1001;
												assign node38933 = (inp[11]) ? node38953 : node38934;
													assign node38934 = (inp[6]) ? node38944 : node38935;
														assign node38935 = (inp[2]) ? 4'b0011 : node38936;
															assign node38936 = (inp[15]) ? node38940 : node38937;
																assign node38937 = (inp[0]) ? 4'b0011 : 4'b0001;
																assign node38940 = (inp[0]) ? 4'b0001 : 4'b0011;
														assign node38944 = (inp[2]) ? 4'b1001 : node38945;
															assign node38945 = (inp[0]) ? node38949 : node38946;
																assign node38946 = (inp[15]) ? 4'b1011 : 4'b1001;
																assign node38949 = (inp[15]) ? 4'b1001 : 4'b1011;
													assign node38953 = (inp[6]) ? node38963 : node38954;
														assign node38954 = (inp[2]) ? node38960 : node38955;
															assign node38955 = (inp[0]) ? node38957 : 4'b1001;
																assign node38957 = (inp[15]) ? 4'b1001 : 4'b1011;
															assign node38960 = (inp[0]) ? 4'b1001 : 4'b1011;
														assign node38963 = (inp[0]) ? node38967 : node38964;
															assign node38964 = (inp[15]) ? 4'b0011 : 4'b0001;
															assign node38967 = (inp[15]) ? 4'b0001 : 4'b0011;
				assign node38970 = (inp[3]) ? node41496 : node38971;
					assign node38971 = (inp[9]) ? node40229 : node38972;
						assign node38972 = (inp[4]) ? node39538 : node38973;
							assign node38973 = (inp[10]) ? node39217 : node38974;
								assign node38974 = (inp[12]) ? node39094 : node38975;
									assign node38975 = (inp[6]) ? node39043 : node38976;
										assign node38976 = (inp[11]) ? node39006 : node38977;
											assign node38977 = (inp[13]) ? node38991 : node38978;
												assign node38978 = (inp[1]) ? node38984 : node38979;
													assign node38979 = (inp[0]) ? 4'b1110 : node38980;
														assign node38980 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node38984 = (inp[15]) ? node38988 : node38985;
														assign node38985 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node38988 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node38991 = (inp[5]) ? node39001 : node38992;
													assign node38992 = (inp[2]) ? node38994 : 4'b0110;
														assign node38994 = (inp[0]) ? node38998 : node38995;
															assign node38995 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node38998 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node39001 = (inp[0]) ? 4'b0100 : node39002;
														assign node39002 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node39006 = (inp[13]) ? node39024 : node39007;
												assign node39007 = (inp[1]) ? node39015 : node39008;
													assign node39008 = (inp[2]) ? 4'b0110 : node39009;
														assign node39009 = (inp[0]) ? 4'b0100 : node39010;
															assign node39010 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node39015 = (inp[5]) ? node39017 : 4'b1110;
														assign node39017 = (inp[0]) ? node39021 : node39018;
															assign node39018 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node39021 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node39024 = (inp[5]) ? node39030 : node39025;
													assign node39025 = (inp[0]) ? 4'b1100 : node39026;
														assign node39026 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node39030 = (inp[2]) ? node39038 : node39031;
														assign node39031 = (inp[1]) ? node39033 : 4'b1110;
															assign node39033 = (inp[15]) ? node39035 : 4'b1100;
																assign node39035 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node39038 = (inp[15]) ? node39040 : 4'b1100;
															assign node39040 = (inp[0]) ? 4'b1110 : 4'b1100;
										assign node39043 = (inp[11]) ? node39073 : node39044;
											assign node39044 = (inp[13]) ? node39060 : node39045;
												assign node39045 = (inp[1]) ? node39053 : node39046;
													assign node39046 = (inp[0]) ? node39050 : node39047;
														assign node39047 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node39050 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node39053 = (inp[0]) ? node39057 : node39054;
														assign node39054 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node39057 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node39060 = (inp[2]) ? node39066 : node39061;
													assign node39061 = (inp[15]) ? 4'b1110 : node39062;
														assign node39062 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node39066 = (inp[15]) ? node39070 : node39067;
														assign node39067 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node39070 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node39073 = (inp[1]) ? node39087 : node39074;
												assign node39074 = (inp[13]) ? node39082 : node39075;
													assign node39075 = (inp[5]) ? node39077 : 4'b1110;
														assign node39077 = (inp[15]) ? 4'b1100 : node39078;
															assign node39078 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node39082 = (inp[15]) ? node39084 : 4'b0100;
														assign node39084 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node39087 = (inp[15]) ? node39091 : node39088;
													assign node39088 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node39091 = (inp[0]) ? 4'b0110 : 4'b0100;
									assign node39094 = (inp[11]) ? node39168 : node39095;
										assign node39095 = (inp[6]) ? node39125 : node39096;
											assign node39096 = (inp[1]) ? node39108 : node39097;
												assign node39097 = (inp[13]) ? node39103 : node39098;
													assign node39098 = (inp[2]) ? node39100 : 4'b1110;
														assign node39100 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node39103 = (inp[0]) ? node39105 : 4'b0110;
														assign node39105 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node39108 = (inp[2]) ? node39116 : node39109;
													assign node39109 = (inp[0]) ? node39113 : node39110;
														assign node39110 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node39113 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node39116 = (inp[13]) ? node39122 : node39117;
														assign node39117 = (inp[15]) ? node39119 : 4'b0100;
															assign node39119 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node39122 = (inp[15]) ? 4'b0100 : 4'b0110;
											assign node39125 = (inp[13]) ? node39141 : node39126;
												assign node39126 = (inp[1]) ? node39134 : node39127;
													assign node39127 = (inp[0]) ? node39131 : node39128;
														assign node39128 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node39131 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node39134 = (inp[0]) ? node39138 : node39135;
														assign node39135 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node39138 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node39141 = (inp[2]) ? node39157 : node39142;
													assign node39142 = (inp[1]) ? node39152 : node39143;
														assign node39143 = (inp[5]) ? node39145 : 4'b1010;
															assign node39145 = (inp[15]) ? node39149 : node39146;
																assign node39146 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node39149 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node39152 = (inp[0]) ? 4'b1000 : node39153;
															assign node39153 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node39157 = (inp[5]) ? 4'b1000 : node39158;
														assign node39158 = (inp[1]) ? 4'b1000 : node39159;
															assign node39159 = (inp[0]) ? node39163 : node39160;
																assign node39160 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node39163 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node39168 = (inp[6]) ? node39188 : node39169;
											assign node39169 = (inp[13]) ? node39181 : node39170;
												assign node39170 = (inp[1]) ? node39176 : node39171;
													assign node39171 = (inp[2]) ? 4'b0100 : node39172;
														assign node39172 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node39176 = (inp[0]) ? 4'b1000 : node39177;
														assign node39177 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node39181 = (inp[15]) ? node39185 : node39182;
													assign node39182 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node39185 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node39188 = (inp[13]) ? node39200 : node39189;
												assign node39189 = (inp[1]) ? node39191 : 4'b1010;
													assign node39191 = (inp[2]) ? 4'b0010 : node39192;
														assign node39192 = (inp[0]) ? node39196 : node39193;
															assign node39193 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node39196 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node39200 = (inp[1]) ? node39208 : node39201;
													assign node39201 = (inp[0]) ? node39205 : node39202;
														assign node39202 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node39205 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node39208 = (inp[5]) ? node39210 : 4'b0010;
														assign node39210 = (inp[15]) ? node39214 : node39211;
															assign node39211 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node39214 = (inp[0]) ? 4'b0010 : 4'b0000;
								assign node39217 = (inp[12]) ? node39373 : node39218;
									assign node39218 = (inp[6]) ? node39288 : node39219;
										assign node39219 = (inp[11]) ? node39251 : node39220;
											assign node39220 = (inp[13]) ? node39238 : node39221;
												assign node39221 = (inp[1]) ? node39229 : node39222;
													assign node39222 = (inp[15]) ? node39226 : node39223;
														assign node39223 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node39226 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node39229 = (inp[5]) ? node39235 : node39230;
														assign node39230 = (inp[15]) ? node39232 : 4'b0110;
															assign node39232 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node39235 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node39238 = (inp[1]) ? node39246 : node39239;
													assign node39239 = (inp[15]) ? node39243 : node39240;
														assign node39240 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node39243 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node39246 = (inp[5]) ? 4'b0110 : node39247;
														assign node39247 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node39251 = (inp[1]) ? node39267 : node39252;
												assign node39252 = (inp[13]) ? node39260 : node39253;
													assign node39253 = (inp[15]) ? node39257 : node39254;
														assign node39254 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node39257 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node39260 = (inp[5]) ? 4'b1010 : node39261;
														assign node39261 = (inp[15]) ? 4'b1000 : node39262;
															assign node39262 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node39267 = (inp[2]) ? node39281 : node39268;
													assign node39268 = (inp[5]) ? 4'b1000 : node39269;
														assign node39269 = (inp[13]) ? node39275 : node39270;
															assign node39270 = (inp[0]) ? node39272 : 4'b1000;
																assign node39272 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node39275 = (inp[0]) ? 4'b1000 : node39276;
																assign node39276 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node39281 = (inp[0]) ? node39285 : node39282;
														assign node39282 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node39285 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node39288 = (inp[11]) ? node39332 : node39289;
											assign node39289 = (inp[1]) ? node39305 : node39290;
												assign node39290 = (inp[13]) ? node39298 : node39291;
													assign node39291 = (inp[2]) ? 4'b0100 : node39292;
														assign node39292 = (inp[15]) ? 4'b0110 : node39293;
															assign node39293 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node39298 = (inp[15]) ? node39302 : node39299;
														assign node39299 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node39302 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node39305 = (inp[13]) ? node39325 : node39306;
													assign node39306 = (inp[2]) ? node39316 : node39307;
														assign node39307 = (inp[5]) ? node39309 : 4'b1000;
															assign node39309 = (inp[15]) ? node39313 : node39310;
																assign node39310 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node39313 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node39316 = (inp[5]) ? 4'b1010 : node39317;
															assign node39317 = (inp[15]) ? node39321 : node39318;
																assign node39318 = (inp[0]) ? 4'b1000 : 4'b1010;
																assign node39321 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node39325 = (inp[2]) ? 4'b1000 : node39326;
														assign node39326 = (inp[0]) ? node39328 : 4'b1000;
															assign node39328 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node39332 = (inp[13]) ? node39354 : node39333;
												assign node39333 = (inp[1]) ? node39341 : node39334;
													assign node39334 = (inp[15]) ? node39338 : node39335;
														assign node39335 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node39338 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node39341 = (inp[5]) ? node39349 : node39342;
														assign node39342 = (inp[2]) ? 4'b0010 : node39343;
															assign node39343 = (inp[0]) ? node39345 : 4'b0000;
																assign node39345 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node39349 = (inp[15]) ? 4'b0000 : node39350;
															assign node39350 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node39354 = (inp[5]) ? node39364 : node39355;
													assign node39355 = (inp[2]) ? 4'b0000 : node39356;
														assign node39356 = (inp[0]) ? node39360 : node39357;
															assign node39357 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node39360 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node39364 = (inp[2]) ? 4'b0010 : node39365;
														assign node39365 = (inp[15]) ? node39369 : node39366;
															assign node39366 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node39369 = (inp[0]) ? 4'b0010 : 4'b0000;
									assign node39373 = (inp[1]) ? node39463 : node39374;
										assign node39374 = (inp[11]) ? node39422 : node39375;
											assign node39375 = (inp[13]) ? node39405 : node39376;
												assign node39376 = (inp[6]) ? node39392 : node39377;
													assign node39377 = (inp[2]) ? node39385 : node39378;
														assign node39378 = (inp[15]) ? node39382 : node39379;
															assign node39379 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node39382 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node39385 = (inp[0]) ? node39389 : node39386;
															assign node39386 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node39389 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node39392 = (inp[2]) ? node39400 : node39393;
														assign node39393 = (inp[0]) ? node39397 : node39394;
															assign node39394 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node39397 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node39400 = (inp[0]) ? 4'b0010 : node39401;
															assign node39401 = (inp[15]) ? 4'b0000 : 4'b0010;
												assign node39405 = (inp[6]) ? node39415 : node39406;
													assign node39406 = (inp[5]) ? node39408 : 4'b0000;
														assign node39408 = (inp[15]) ? node39412 : node39409;
															assign node39409 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node39412 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node39415 = (inp[0]) ? node39419 : node39416;
														assign node39416 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node39419 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node39422 = (inp[5]) ? node39452 : node39423;
												assign node39423 = (inp[2]) ? node39437 : node39424;
													assign node39424 = (inp[13]) ? node39430 : node39425;
														assign node39425 = (inp[0]) ? node39427 : 4'b1000;
															assign node39427 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node39430 = (inp[0]) ? node39434 : node39431;
															assign node39431 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node39434 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node39437 = (inp[13]) ? node39445 : node39438;
														assign node39438 = (inp[6]) ? node39440 : 4'b0010;
															assign node39440 = (inp[0]) ? node39442 : 4'b1000;
																assign node39442 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node39445 = (inp[6]) ? node39447 : 4'b1000;
															assign node39447 = (inp[15]) ? 4'b0010 : node39448;
																assign node39448 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node39452 = (inp[6]) ? node39456 : node39453;
													assign node39453 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node39456 = (inp[13]) ? node39458 : 4'b1000;
														assign node39458 = (inp[15]) ? 4'b0000 : node39459;
															assign node39459 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node39463 = (inp[0]) ? node39493 : node39464;
											assign node39464 = (inp[15]) ? node39486 : node39465;
												assign node39465 = (inp[2]) ? node39481 : node39466;
													assign node39466 = (inp[5]) ? node39474 : node39467;
														assign node39467 = (inp[13]) ? 4'b0010 : node39468;
															assign node39468 = (inp[6]) ? 4'b0010 : node39469;
																assign node39469 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node39474 = (inp[11]) ? node39478 : node39475;
															assign node39475 = (inp[6]) ? 4'b1010 : 4'b0010;
															assign node39478 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node39481 = (inp[13]) ? 4'b1010 : node39482;
														assign node39482 = (inp[6]) ? 4'b1010 : 4'b0010;
												assign node39486 = (inp[6]) ? node39490 : node39487;
													assign node39487 = (inp[11]) ? 4'b1000 : 4'b0000;
													assign node39490 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node39493 = (inp[15]) ? node39519 : node39494;
												assign node39494 = (inp[2]) ? node39506 : node39495;
													assign node39495 = (inp[13]) ? node39501 : node39496;
														assign node39496 = (inp[11]) ? node39498 : 4'b0000;
															assign node39498 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node39501 = (inp[11]) ? 4'b0000 : node39502;
															assign node39502 = (inp[6]) ? 4'b1000 : 4'b0000;
													assign node39506 = (inp[5]) ? node39514 : node39507;
														assign node39507 = (inp[11]) ? node39511 : node39508;
															assign node39508 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node39511 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node39514 = (inp[6]) ? 4'b0000 : node39515;
															assign node39515 = (inp[11]) ? 4'b1000 : 4'b0000;
												assign node39519 = (inp[5]) ? node39531 : node39520;
													assign node39520 = (inp[2]) ? node39526 : node39521;
														assign node39521 = (inp[11]) ? 4'b1010 : node39522;
															assign node39522 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node39526 = (inp[11]) ? 4'b0010 : node39527;
															assign node39527 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node39531 = (inp[6]) ? node39535 : node39532;
														assign node39532 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node39535 = (inp[11]) ? 4'b0010 : 4'b1010;
							assign node39538 = (inp[12]) ? node39902 : node39539;
								assign node39539 = (inp[10]) ? node39751 : node39540;
									assign node39540 = (inp[2]) ? node39628 : node39541;
										assign node39541 = (inp[11]) ? node39593 : node39542;
											assign node39542 = (inp[6]) ? node39576 : node39543;
												assign node39543 = (inp[1]) ? node39559 : node39544;
													assign node39544 = (inp[13]) ? node39554 : node39545;
														assign node39545 = (inp[5]) ? node39551 : node39546;
															assign node39546 = (inp[15]) ? 4'b1000 : node39547;
																assign node39547 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node39551 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node39554 = (inp[0]) ? node39556 : 4'b0010;
															assign node39556 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node39559 = (inp[5]) ? node39569 : node39560;
														assign node39560 = (inp[13]) ? 4'b0010 : node39561;
															assign node39561 = (inp[0]) ? node39565 : node39562;
																assign node39562 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node39565 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node39569 = (inp[13]) ? 4'b0000 : node39570;
															assign node39570 = (inp[0]) ? node39572 : 4'b0010;
																assign node39572 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node39576 = (inp[1]) ? node39586 : node39577;
													assign node39577 = (inp[13]) ? node39583 : node39578;
														assign node39578 = (inp[0]) ? 4'b0010 : node39579;
															assign node39579 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node39583 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node39586 = (inp[15]) ? node39590 : node39587;
														assign node39587 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node39590 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node39593 = (inp[6]) ? node39607 : node39594;
												assign node39594 = (inp[13]) ? node39600 : node39595;
													assign node39595 = (inp[0]) ? 4'b1000 : node39596;
														assign node39596 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node39600 = (inp[5]) ? 4'b1000 : node39601;
														assign node39601 = (inp[15]) ? node39603 : 4'b1010;
															assign node39603 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node39607 = (inp[13]) ? node39621 : node39608;
													assign node39608 = (inp[1]) ? node39616 : node39609;
														assign node39609 = (inp[15]) ? node39613 : node39610;
															assign node39610 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node39613 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node39616 = (inp[0]) ? 4'b0010 : node39617;
															assign node39617 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node39621 = (inp[15]) ? node39625 : node39622;
														assign node39622 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node39625 = (inp[0]) ? 4'b0010 : 4'b0000;
										assign node39628 = (inp[5]) ? node39694 : node39629;
											assign node39629 = (inp[11]) ? node39655 : node39630;
												assign node39630 = (inp[6]) ? node39640 : node39631;
													assign node39631 = (inp[1]) ? node39635 : node39632;
														assign node39632 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node39635 = (inp[15]) ? node39637 : 4'b0010;
															assign node39637 = (inp[13]) ? 4'b0010 : 4'b0000;
													assign node39640 = (inp[1]) ? node39648 : node39641;
														assign node39641 = (inp[13]) ? 4'b1000 : node39642;
															assign node39642 = (inp[15]) ? 4'b0000 : node39643;
																assign node39643 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node39648 = (inp[13]) ? node39650 : 4'b1000;
															assign node39650 = (inp[15]) ? node39652 : 4'b1000;
																assign node39652 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node39655 = (inp[6]) ? node39679 : node39656;
													assign node39656 = (inp[13]) ? node39668 : node39657;
														assign node39657 = (inp[1]) ? node39663 : node39658;
															assign node39658 = (inp[0]) ? node39660 : 4'b0010;
																assign node39660 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node39663 = (inp[15]) ? 4'b1010 : node39664;
																assign node39664 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node39668 = (inp[1]) ? node39674 : node39669;
															assign node39669 = (inp[15]) ? 4'b1000 : node39670;
																assign node39670 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node39674 = (inp[15]) ? node39676 : 4'b1000;
																assign node39676 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node39679 = (inp[13]) ? node39689 : node39680;
														assign node39680 = (inp[1]) ? node39686 : node39681;
															assign node39681 = (inp[15]) ? node39683 : 4'b1010;
																assign node39683 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node39686 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node39689 = (inp[15]) ? 4'b0000 : node39690;
															assign node39690 = (inp[0]) ? 4'b0000 : 4'b0010;
											assign node39694 = (inp[6]) ? node39720 : node39695;
												assign node39695 = (inp[11]) ? node39711 : node39696;
													assign node39696 = (inp[13]) ? node39706 : node39697;
														assign node39697 = (inp[1]) ? node39699 : 4'b1010;
															assign node39699 = (inp[0]) ? node39703 : node39700;
																assign node39700 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node39703 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node39706 = (inp[0]) ? node39708 : 4'b0000;
															assign node39708 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node39711 = (inp[13]) ? node39715 : node39712;
														assign node39712 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node39715 = (inp[0]) ? 4'b1010 : node39716;
															assign node39716 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node39720 = (inp[11]) ? node39736 : node39721;
													assign node39721 = (inp[1]) ? node39723 : 4'b1010;
														assign node39723 = (inp[13]) ? node39729 : node39724;
															assign node39724 = (inp[0]) ? node39726 : 4'b1010;
																assign node39726 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node39729 = (inp[0]) ? node39733 : node39730;
																assign node39730 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node39733 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node39736 = (inp[13]) ? node39744 : node39737;
														assign node39737 = (inp[1]) ? 4'b0010 : node39738;
															assign node39738 = (inp[0]) ? 4'b1000 : node39739;
																assign node39739 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node39744 = (inp[1]) ? node39746 : 4'b0000;
															assign node39746 = (inp[15]) ? node39748 : 4'b0000;
																assign node39748 = (inp[0]) ? 4'b0010 : 4'b0000;
									assign node39751 = (inp[11]) ? node39827 : node39752;
										assign node39752 = (inp[6]) ? node39786 : node39753;
											assign node39753 = (inp[13]) ? node39779 : node39754;
												assign node39754 = (inp[1]) ? node39762 : node39755;
													assign node39755 = (inp[15]) ? node39759 : node39756;
														assign node39756 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node39759 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node39762 = (inp[2]) ? node39770 : node39763;
														assign node39763 = (inp[5]) ? node39767 : node39764;
															assign node39764 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node39767 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node39770 = (inp[5]) ? node39774 : node39771;
															assign node39771 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node39774 = (inp[15]) ? 4'b0000 : node39775;
																assign node39775 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node39779 = (inp[0]) ? node39783 : node39780;
													assign node39780 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node39783 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node39786 = (inp[13]) ? node39804 : node39787;
												assign node39787 = (inp[1]) ? node39799 : node39788;
													assign node39788 = (inp[5]) ? node39794 : node39789;
														assign node39789 = (inp[15]) ? 4'b0010 : node39790;
															assign node39790 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node39794 = (inp[15]) ? 4'b0000 : node39795;
															assign node39795 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node39799 = (inp[0]) ? 4'b1110 : node39800;
														assign node39800 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node39804 = (inp[1]) ? node39816 : node39805;
													assign node39805 = (inp[15]) ? node39811 : node39806;
														assign node39806 = (inp[2]) ? node39808 : 4'b1110;
															assign node39808 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node39811 = (inp[0]) ? 4'b1100 : node39812;
															assign node39812 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node39816 = (inp[5]) ? 4'b1110 : node39817;
														assign node39817 = (inp[2]) ? 4'b1110 : node39818;
															assign node39818 = (inp[15]) ? node39822 : node39819;
																assign node39819 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node39822 = (inp[0]) ? 4'b1110 : 4'b1100;
										assign node39827 = (inp[6]) ? node39861 : node39828;
											assign node39828 = (inp[1]) ? node39838 : node39829;
												assign node39829 = (inp[13]) ? node39835 : node39830;
													assign node39830 = (inp[0]) ? node39832 : 4'b0000;
														assign node39832 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node39835 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node39838 = (inp[15]) ? node39854 : node39839;
													assign node39839 = (inp[13]) ? node39847 : node39840;
														assign node39840 = (inp[2]) ? node39842 : 4'b1100;
															assign node39842 = (inp[0]) ? node39844 : 4'b1110;
																assign node39844 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node39847 = (inp[2]) ? 4'b1100 : node39848;
															assign node39848 = (inp[5]) ? 4'b1110 : node39849;
																assign node39849 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node39854 = (inp[5]) ? node39858 : node39855;
														assign node39855 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node39858 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node39861 = (inp[1]) ? node39879 : node39862;
												assign node39862 = (inp[13]) ? node39874 : node39863;
													assign node39863 = (inp[0]) ? node39869 : node39864;
														assign node39864 = (inp[15]) ? node39866 : 4'b1110;
															assign node39866 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node39869 = (inp[5]) ? 4'b1100 : node39870;
															assign node39870 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node39874 = (inp[2]) ? node39876 : 4'b0110;
														assign node39876 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node39879 = (inp[13]) ? node39893 : node39880;
													assign node39880 = (inp[15]) ? node39886 : node39881;
														assign node39881 = (inp[0]) ? node39883 : 4'b0100;
															assign node39883 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node39886 = (inp[2]) ? node39888 : 4'b0110;
															assign node39888 = (inp[0]) ? 4'b0100 : node39889;
																assign node39889 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node39893 = (inp[0]) ? 4'b0110 : node39894;
														assign node39894 = (inp[5]) ? node39898 : node39895;
															assign node39895 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node39898 = (inp[15]) ? 4'b0110 : 4'b0100;
								assign node39902 = (inp[10]) ? node40052 : node39903;
									assign node39903 = (inp[11]) ? node39961 : node39904;
										assign node39904 = (inp[6]) ? node39930 : node39905;
											assign node39905 = (inp[13]) ? node39915 : node39906;
												assign node39906 = (inp[1]) ? node39910 : node39907;
													assign node39907 = (inp[2]) ? 4'b1000 : 4'b1010;
													assign node39910 = (inp[15]) ? 4'b0010 : node39911;
														assign node39911 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node39915 = (inp[1]) ? node39923 : node39916;
													assign node39916 = (inp[15]) ? node39920 : node39917;
														assign node39917 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node39920 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node39923 = (inp[15]) ? node39927 : node39924;
														assign node39924 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node39927 = (inp[0]) ? 4'b0010 : 4'b0000;
											assign node39930 = (inp[1]) ? node39952 : node39931;
												assign node39931 = (inp[13]) ? node39945 : node39932;
													assign node39932 = (inp[5]) ? node39940 : node39933;
														assign node39933 = (inp[0]) ? node39937 : node39934;
															assign node39934 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node39937 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node39940 = (inp[0]) ? 4'b0000 : node39941;
															assign node39941 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node39945 = (inp[0]) ? node39947 : 4'b1100;
														assign node39947 = (inp[5]) ? node39949 : 4'b1100;
															assign node39949 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node39952 = (inp[0]) ? node39954 : 4'b1100;
													assign node39954 = (inp[15]) ? node39958 : node39955;
														assign node39955 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node39958 = (inp[5]) ? 4'b1100 : 4'b1110;
										assign node39961 = (inp[6]) ? node40001 : node39962;
											assign node39962 = (inp[13]) ? node39992 : node39963;
												assign node39963 = (inp[1]) ? node39971 : node39964;
													assign node39964 = (inp[5]) ? node39966 : 4'b0010;
														assign node39966 = (inp[0]) ? 4'b0000 : node39967;
															assign node39967 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node39971 = (inp[2]) ? node39985 : node39972;
														assign node39972 = (inp[5]) ? node39980 : node39973;
															assign node39973 = (inp[0]) ? node39977 : node39974;
																assign node39974 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node39977 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node39980 = (inp[15]) ? 4'b1110 : node39981;
																assign node39981 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node39985 = (inp[5]) ? node39987 : 4'b1110;
															assign node39987 = (inp[15]) ? node39989 : 4'b1110;
																assign node39989 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node39992 = (inp[15]) ? 4'b1100 : node39993;
													assign node39993 = (inp[0]) ? node39997 : node39994;
														assign node39994 = (inp[5]) ? 4'b1100 : 4'b1110;
														assign node39997 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node40001 = (inp[1]) ? node40027 : node40002;
												assign node40002 = (inp[13]) ? node40018 : node40003;
													assign node40003 = (inp[2]) ? node40011 : node40004;
														assign node40004 = (inp[5]) ? 4'b1100 : node40005;
															assign node40005 = (inp[15]) ? 4'b1110 : node40006;
																assign node40006 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node40011 = (inp[5]) ? node40013 : 4'b1100;
															assign node40013 = (inp[0]) ? 4'b1100 : node40014;
																assign node40014 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node40018 = (inp[5]) ? node40020 : 4'b0100;
														assign node40020 = (inp[2]) ? node40022 : 4'b0100;
															assign node40022 = (inp[0]) ? 4'b0110 : node40023;
																assign node40023 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node40027 = (inp[13]) ? node40043 : node40028;
													assign node40028 = (inp[2]) ? node40036 : node40029;
														assign node40029 = (inp[15]) ? node40033 : node40030;
															assign node40030 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node40033 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node40036 = (inp[15]) ? node40038 : 4'b0100;
															assign node40038 = (inp[5]) ? 4'b0100 : node40039;
																assign node40039 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node40043 = (inp[0]) ? 4'b0110 : node40044;
														assign node40044 = (inp[5]) ? node40048 : node40045;
															assign node40045 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node40048 = (inp[2]) ? 4'b0110 : 4'b0100;
									assign node40052 = (inp[15]) ? node40142 : node40053;
										assign node40053 = (inp[2]) ? node40097 : node40054;
											assign node40054 = (inp[5]) ? node40072 : node40055;
												assign node40055 = (inp[0]) ? node40067 : node40056;
													assign node40056 = (inp[11]) ? node40058 : 4'b1110;
														assign node40058 = (inp[13]) ? node40064 : node40059;
															assign node40059 = (inp[1]) ? 4'b1110 : node40060;
																assign node40060 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node40064 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node40067 = (inp[11]) ? 4'b1100 : node40068;
														assign node40068 = (inp[6]) ? 4'b1100 : 4'b0100;
												assign node40072 = (inp[0]) ? node40090 : node40073;
													assign node40073 = (inp[13]) ? node40085 : node40074;
														assign node40074 = (inp[6]) ? node40080 : node40075;
															assign node40075 = (inp[1]) ? node40077 : 4'b1100;
																assign node40077 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node40080 = (inp[1]) ? node40082 : 4'b0100;
																assign node40082 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node40085 = (inp[11]) ? 4'b1100 : node40086;
															assign node40086 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node40090 = (inp[1]) ? node40092 : 4'b0110;
														assign node40092 = (inp[11]) ? node40094 : 4'b1110;
															assign node40094 = (inp[6]) ? 4'b0110 : 4'b1110;
											assign node40097 = (inp[5]) ? node40127 : node40098;
												assign node40098 = (inp[0]) ? node40110 : node40099;
													assign node40099 = (inp[1]) ? node40105 : node40100;
														assign node40100 = (inp[6]) ? 4'b0110 : node40101;
															assign node40101 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node40105 = (inp[11]) ? 4'b1110 : node40106;
															assign node40106 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node40110 = (inp[1]) ? node40118 : node40111;
														assign node40111 = (inp[6]) ? node40113 : 4'b1100;
															assign node40113 = (inp[11]) ? node40115 : 4'b1100;
																assign node40115 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node40118 = (inp[13]) ? 4'b1100 : node40119;
															assign node40119 = (inp[11]) ? node40123 : node40120;
																assign node40120 = (inp[6]) ? 4'b1100 : 4'b0100;
																assign node40123 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node40127 = (inp[0]) ? node40131 : node40128;
													assign node40128 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node40131 = (inp[11]) ? node40137 : node40132;
														assign node40132 = (inp[6]) ? 4'b1110 : node40133;
															assign node40133 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node40137 = (inp[6]) ? 4'b0110 : node40138;
															assign node40138 = (inp[1]) ? 4'b1110 : 4'b0110;
										assign node40142 = (inp[0]) ? node40186 : node40143;
											assign node40143 = (inp[5]) ? node40169 : node40144;
												assign node40144 = (inp[13]) ? node40154 : node40145;
													assign node40145 = (inp[11]) ? node40147 : 4'b1100;
														assign node40147 = (inp[1]) ? node40151 : node40148;
															assign node40148 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node40151 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node40154 = (inp[1]) ? node40162 : node40155;
														assign node40155 = (inp[11]) ? node40159 : node40156;
															assign node40156 = (inp[6]) ? 4'b1100 : 4'b0100;
															assign node40159 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node40162 = (inp[6]) ? node40166 : node40163;
															assign node40163 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node40166 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node40169 = (inp[11]) ? node40177 : node40170;
													assign node40170 = (inp[6]) ? 4'b1110 : node40171;
														assign node40171 = (inp[13]) ? 4'b0110 : node40172;
															assign node40172 = (inp[1]) ? 4'b0110 : 4'b1110;
													assign node40177 = (inp[6]) ? node40181 : node40178;
														assign node40178 = (inp[1]) ? 4'b1110 : 4'b0110;
														assign node40181 = (inp[13]) ? 4'b0110 : node40182;
															assign node40182 = (inp[2]) ? 4'b0110 : 4'b1110;
											assign node40186 = (inp[5]) ? node40212 : node40187;
												assign node40187 = (inp[2]) ? node40203 : node40188;
													assign node40188 = (inp[13]) ? node40198 : node40189;
														assign node40189 = (inp[6]) ? node40191 : 4'b1110;
															assign node40191 = (inp[1]) ? node40195 : node40192;
																assign node40192 = (inp[11]) ? 4'b1110 : 4'b0110;
																assign node40195 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node40198 = (inp[6]) ? node40200 : 4'b0110;
															assign node40200 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node40203 = (inp[1]) ? 4'b0110 : node40204;
														assign node40204 = (inp[13]) ? node40206 : 4'b0110;
															assign node40206 = (inp[11]) ? node40208 : 4'b0110;
																assign node40208 = (inp[6]) ? 4'b0110 : 4'b1110;
												assign node40212 = (inp[6]) ? node40218 : node40213;
													assign node40213 = (inp[11]) ? 4'b1100 : node40214;
														assign node40214 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node40218 = (inp[2]) ? node40220 : 4'b0100;
														assign node40220 = (inp[1]) ? 4'b0100 : node40221;
															assign node40221 = (inp[11]) ? node40225 : node40222;
																assign node40222 = (inp[13]) ? 4'b1100 : 4'b0100;
																assign node40225 = (inp[13]) ? 4'b0100 : 4'b1100;
						assign node40229 = (inp[4]) ? node40837 : node40230;
							assign node40230 = (inp[10]) ? node40514 : node40231;
								assign node40231 = (inp[12]) ? node40355 : node40232;
									assign node40232 = (inp[15]) ? node40318 : node40233;
										assign node40233 = (inp[0]) ? node40283 : node40234;
											assign node40234 = (inp[5]) ? node40258 : node40235;
												assign node40235 = (inp[1]) ? node40245 : node40236;
													assign node40236 = (inp[2]) ? node40238 : 4'b0010;
														assign node40238 = (inp[6]) ? 4'b0010 : node40239;
															assign node40239 = (inp[11]) ? node40241 : 4'b0010;
																assign node40241 = (inp[13]) ? 4'b1010 : 4'b0010;
													assign node40245 = (inp[2]) ? node40251 : node40246;
														assign node40246 = (inp[6]) ? 4'b1010 : node40247;
															assign node40247 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node40251 = (inp[11]) ? node40255 : node40252;
															assign node40252 = (inp[13]) ? 4'b1010 : 4'b0010;
															assign node40255 = (inp[6]) ? 4'b0010 : 4'b1010;
												assign node40258 = (inp[6]) ? node40272 : node40259;
													assign node40259 = (inp[1]) ? node40269 : node40260;
														assign node40260 = (inp[2]) ? 4'b1010 : node40261;
															assign node40261 = (inp[11]) ? node40265 : node40262;
																assign node40262 = (inp[13]) ? 4'b0010 : 4'b1010;
																assign node40265 = (inp[13]) ? 4'b1010 : 4'b0010;
														assign node40269 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node40272 = (inp[11]) ? node40278 : node40273;
														assign node40273 = (inp[13]) ? 4'b1010 : node40274;
															assign node40274 = (inp[1]) ? 4'b1010 : 4'b0010;
														assign node40278 = (inp[13]) ? 4'b0010 : node40279;
															assign node40279 = (inp[1]) ? 4'b0010 : 4'b1010;
											assign node40283 = (inp[11]) ? node40293 : node40284;
												assign node40284 = (inp[6]) ? node40290 : node40285;
													assign node40285 = (inp[13]) ? 4'b0000 : node40286;
														assign node40286 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node40290 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node40293 = (inp[2]) ? node40303 : node40294;
													assign node40294 = (inp[13]) ? node40300 : node40295;
														assign node40295 = (inp[5]) ? 4'b1000 : node40296;
															assign node40296 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node40300 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node40303 = (inp[5]) ? node40309 : node40304;
														assign node40304 = (inp[6]) ? 4'b1000 : node40305;
															assign node40305 = (inp[1]) ? 4'b1000 : 4'b0000;
														assign node40309 = (inp[6]) ? node40313 : node40310;
															assign node40310 = (inp[1]) ? 4'b1000 : 4'b0000;
															assign node40313 = (inp[13]) ? 4'b0000 : node40314;
																assign node40314 = (inp[1]) ? 4'b0000 : 4'b1000;
										assign node40318 = (inp[0]) ? node40342 : node40319;
											assign node40319 = (inp[11]) ? node40331 : node40320;
												assign node40320 = (inp[6]) ? node40326 : node40321;
													assign node40321 = (inp[13]) ? 4'b0000 : node40322;
														assign node40322 = (inp[1]) ? 4'b0000 : 4'b1000;
													assign node40326 = (inp[1]) ? 4'b1000 : node40327;
														assign node40327 = (inp[13]) ? 4'b1000 : 4'b0000;
												assign node40331 = (inp[6]) ? node40337 : node40332;
													assign node40332 = (inp[1]) ? 4'b1000 : node40333;
														assign node40333 = (inp[13]) ? 4'b1000 : 4'b0000;
													assign node40337 = (inp[1]) ? 4'b0000 : node40338;
														assign node40338 = (inp[13]) ? 4'b0000 : 4'b1000;
											assign node40342 = (inp[6]) ? node40348 : node40343;
												assign node40343 = (inp[11]) ? node40345 : 4'b0010;
													assign node40345 = (inp[1]) ? 4'b1010 : 4'b0010;
												assign node40348 = (inp[11]) ? node40350 : 4'b1010;
													assign node40350 = (inp[1]) ? 4'b0010 : node40351;
														assign node40351 = (inp[13]) ? 4'b0010 : 4'b1010;
									assign node40355 = (inp[6]) ? node40427 : node40356;
										assign node40356 = (inp[11]) ? node40394 : node40357;
											assign node40357 = (inp[13]) ? node40373 : node40358;
												assign node40358 = (inp[1]) ? node40366 : node40359;
													assign node40359 = (inp[0]) ? node40363 : node40360;
														assign node40360 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node40363 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node40366 = (inp[15]) ? node40370 : node40367;
														assign node40367 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node40370 = (inp[0]) ? 4'b0010 : 4'b0000;
												assign node40373 = (inp[1]) ? node40387 : node40374;
													assign node40374 = (inp[2]) ? node40382 : node40375;
														assign node40375 = (inp[0]) ? node40379 : node40376;
															assign node40376 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node40379 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node40382 = (inp[0]) ? 4'b0010 : node40383;
															assign node40383 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node40387 = (inp[0]) ? node40391 : node40388;
														assign node40388 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node40391 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node40394 = (inp[1]) ? node40410 : node40395;
												assign node40395 = (inp[13]) ? node40407 : node40396;
													assign node40396 = (inp[2]) ? node40398 : 4'b0010;
														assign node40398 = (inp[5]) ? node40400 : 4'b0000;
															assign node40400 = (inp[15]) ? node40404 : node40401;
																assign node40401 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node40404 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node40407 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node40410 = (inp[2]) ? node40418 : node40411;
													assign node40411 = (inp[5]) ? 4'b1110 : node40412;
														assign node40412 = (inp[15]) ? node40414 : 4'b1100;
															assign node40414 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node40418 = (inp[13]) ? 4'b1100 : node40419;
														assign node40419 = (inp[5]) ? node40421 : 4'b1100;
															assign node40421 = (inp[15]) ? 4'b1110 : node40422;
																assign node40422 = (inp[0]) ? 4'b1110 : 4'b1100;
										assign node40427 = (inp[11]) ? node40477 : node40428;
											assign node40428 = (inp[1]) ? node40452 : node40429;
												assign node40429 = (inp[13]) ? node40443 : node40430;
													assign node40430 = (inp[2]) ? node40436 : node40431;
														assign node40431 = (inp[15]) ? node40433 : 4'b0000;
															assign node40433 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node40436 = (inp[15]) ? node40440 : node40437;
															assign node40437 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node40440 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node40443 = (inp[5]) ? 4'b1110 : node40444;
														assign node40444 = (inp[15]) ? node40448 : node40445;
															assign node40445 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node40448 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node40452 = (inp[5]) ? node40468 : node40453;
													assign node40453 = (inp[2]) ? node40461 : node40454;
														assign node40454 = (inp[0]) ? node40458 : node40455;
															assign node40455 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node40458 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node40461 = (inp[0]) ? node40465 : node40462;
															assign node40462 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node40465 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node40468 = (inp[2]) ? 4'b1100 : node40469;
														assign node40469 = (inp[15]) ? node40473 : node40470;
															assign node40470 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node40473 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node40477 = (inp[1]) ? node40493 : node40478;
												assign node40478 = (inp[13]) ? node40486 : node40479;
													assign node40479 = (inp[5]) ? node40481 : 4'b1110;
														assign node40481 = (inp[0]) ? 4'b1100 : node40482;
															assign node40482 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node40486 = (inp[0]) ? 4'b0110 : node40487;
														assign node40487 = (inp[5]) ? node40489 : 4'b0100;
															assign node40489 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node40493 = (inp[15]) ? node40501 : node40494;
													assign node40494 = (inp[0]) ? node40498 : node40495;
														assign node40495 = (inp[5]) ? 4'b0100 : 4'b0110;
														assign node40498 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node40501 = (inp[13]) ? node40507 : node40502;
														assign node40502 = (inp[5]) ? node40504 : 4'b0110;
															assign node40504 = (inp[2]) ? 4'b0100 : 4'b0110;
														assign node40507 = (inp[0]) ? node40511 : node40508;
															assign node40508 = (inp[5]) ? 4'b0110 : 4'b0100;
															assign node40511 = (inp[5]) ? 4'b0100 : 4'b0110;
								assign node40514 = (inp[12]) ? node40660 : node40515;
									assign node40515 = (inp[11]) ? node40587 : node40516;
										assign node40516 = (inp[6]) ? node40552 : node40517;
											assign node40517 = (inp[13]) ? node40529 : node40518;
												assign node40518 = (inp[1]) ? node40526 : node40519;
													assign node40519 = (inp[0]) ? node40523 : node40520;
														assign node40520 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node40523 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node40526 = (inp[2]) ? 4'b0010 : 4'b0000;
												assign node40529 = (inp[2]) ? node40545 : node40530;
													assign node40530 = (inp[5]) ? 4'b0010 : node40531;
														assign node40531 = (inp[1]) ? node40537 : node40532;
															assign node40532 = (inp[15]) ? 4'b0010 : node40533;
																assign node40533 = (inp[0]) ? 4'b0000 : 4'b0010;
															assign node40537 = (inp[0]) ? node40541 : node40538;
																assign node40538 = (inp[15]) ? 4'b0000 : 4'b0010;
																assign node40541 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node40545 = (inp[5]) ? node40547 : 4'b0010;
														assign node40547 = (inp[0]) ? node40549 : 4'b0000;
															assign node40549 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node40552 = (inp[1]) ? node40570 : node40553;
												assign node40553 = (inp[13]) ? node40561 : node40554;
													assign node40554 = (inp[0]) ? node40558 : node40555;
														assign node40555 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node40558 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node40561 = (inp[2]) ? 4'b1110 : node40562;
														assign node40562 = (inp[5]) ? node40564 : 4'b1100;
															assign node40564 = (inp[15]) ? 4'b1110 : node40565;
																assign node40565 = (inp[0]) ? 4'b1110 : 4'b1100;
												assign node40570 = (inp[5]) ? node40580 : node40571;
													assign node40571 = (inp[2]) ? node40573 : 4'b1100;
														assign node40573 = (inp[15]) ? node40577 : node40574;
															assign node40574 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node40577 = (inp[13]) ? 4'b1110 : 4'b1100;
													assign node40580 = (inp[0]) ? node40584 : node40581;
														assign node40581 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node40584 = (inp[15]) ? 4'b1100 : 4'b1110;
										assign node40587 = (inp[6]) ? node40621 : node40588;
											assign node40588 = (inp[13]) ? node40604 : node40589;
												assign node40589 = (inp[1]) ? node40595 : node40590;
													assign node40590 = (inp[0]) ? 4'b0010 : node40591;
														assign node40591 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node40595 = (inp[0]) ? node40597 : 4'b1110;
														assign node40597 = (inp[5]) ? node40601 : node40598;
															assign node40598 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node40601 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node40604 = (inp[2]) ? node40614 : node40605;
													assign node40605 = (inp[15]) ? 4'b1110 : node40606;
														assign node40606 = (inp[5]) ? node40610 : node40607;
															assign node40607 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node40610 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node40614 = (inp[1]) ? 4'b1100 : node40615;
														assign node40615 = (inp[5]) ? 4'b1110 : node40616;
															assign node40616 = (inp[15]) ? 4'b1110 : 4'b1100;
											assign node40621 = (inp[13]) ? node40639 : node40622;
												assign node40622 = (inp[1]) ? node40630 : node40623;
													assign node40623 = (inp[15]) ? node40625 : 4'b1100;
														assign node40625 = (inp[0]) ? node40627 : 4'b1100;
															assign node40627 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node40630 = (inp[5]) ? node40632 : 4'b0110;
														assign node40632 = (inp[15]) ? node40636 : node40633;
															assign node40633 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node40636 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node40639 = (inp[1]) ? node40655 : node40640;
													assign node40640 = (inp[5]) ? node40650 : node40641;
														assign node40641 = (inp[2]) ? 4'b0100 : node40642;
															assign node40642 = (inp[0]) ? node40646 : node40643;
																assign node40643 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node40646 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node40650 = (inp[15]) ? 4'b0110 : node40651;
															assign node40651 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node40655 = (inp[15]) ? node40657 : 4'b0110;
														assign node40657 = (inp[0]) ? 4'b0110 : 4'b0100;
									assign node40660 = (inp[15]) ? node40764 : node40661;
										assign node40661 = (inp[1]) ? node40715 : node40662;
											assign node40662 = (inp[11]) ? node40688 : node40663;
												assign node40663 = (inp[6]) ? node40681 : node40664;
													assign node40664 = (inp[13]) ? 4'b0110 : node40665;
														assign node40665 = (inp[2]) ? node40673 : node40666;
															assign node40666 = (inp[5]) ? node40670 : node40667;
																assign node40667 = (inp[0]) ? 4'b1100 : 4'b1110;
																assign node40670 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node40673 = (inp[0]) ? node40677 : node40674;
																assign node40674 = (inp[5]) ? 4'b1100 : 4'b1110;
																assign node40677 = (inp[5]) ? 4'b1110 : 4'b1100;
													assign node40681 = (inp[13]) ? node40685 : node40682;
														assign node40682 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node40685 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node40688 = (inp[0]) ? node40704 : node40689;
													assign node40689 = (inp[5]) ? node40697 : node40690;
														assign node40690 = (inp[2]) ? node40692 : 4'b1110;
															assign node40692 = (inp[13]) ? node40694 : 4'b1110;
																assign node40694 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node40697 = (inp[6]) ? node40701 : node40698;
															assign node40698 = (inp[2]) ? 4'b1100 : 4'b0100;
															assign node40701 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node40704 = (inp[5]) ? node40708 : node40705;
														assign node40705 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node40708 = (inp[13]) ? node40712 : node40709;
															assign node40709 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node40712 = (inp[6]) ? 4'b0110 : 4'b1110;
											assign node40715 = (inp[5]) ? node40739 : node40716;
												assign node40716 = (inp[0]) ? node40724 : node40717;
													assign node40717 = (inp[11]) ? node40721 : node40718;
														assign node40718 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node40721 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node40724 = (inp[13]) ? 4'b0100 : node40725;
														assign node40725 = (inp[2]) ? node40733 : node40726;
															assign node40726 = (inp[6]) ? node40730 : node40727;
																assign node40727 = (inp[11]) ? 4'b1100 : 4'b0100;
																assign node40730 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node40733 = (inp[6]) ? node40735 : 4'b0100;
																assign node40735 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node40739 = (inp[0]) ? node40747 : node40740;
													assign node40740 = (inp[6]) ? node40744 : node40741;
														assign node40741 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node40744 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node40747 = (inp[13]) ? node40759 : node40748;
														assign node40748 = (inp[2]) ? node40754 : node40749;
															assign node40749 = (inp[11]) ? node40751 : 4'b1110;
																assign node40751 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node40754 = (inp[6]) ? 4'b1110 : node40755;
																assign node40755 = (inp[11]) ? 4'b1110 : 4'b0110;
														assign node40759 = (inp[11]) ? 4'b0110 : node40760;
															assign node40760 = (inp[6]) ? 4'b1110 : 4'b0110;
										assign node40764 = (inp[6]) ? node40792 : node40765;
											assign node40765 = (inp[11]) ? node40777 : node40766;
												assign node40766 = (inp[5]) ? node40774 : node40767;
													assign node40767 = (inp[0]) ? node40769 : 4'b0100;
														assign node40769 = (inp[1]) ? 4'b0110 : node40770;
															assign node40770 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node40774 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node40777 = (inp[13]) ? node40787 : node40778;
													assign node40778 = (inp[1]) ? node40782 : node40779;
														assign node40779 = (inp[2]) ? 4'b0100 : 4'b0110;
														assign node40782 = (inp[2]) ? node40784 : 4'b1100;
															assign node40784 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node40787 = (inp[0]) ? 4'b1110 : node40788;
														assign node40788 = (inp[5]) ? 4'b1110 : 4'b1100;
											assign node40792 = (inp[11]) ? node40812 : node40793;
												assign node40793 = (inp[13]) ? node40805 : node40794;
													assign node40794 = (inp[1]) ? node40800 : node40795;
														assign node40795 = (inp[5]) ? 4'b0100 : node40796;
															assign node40796 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node40800 = (inp[2]) ? 4'b1100 : node40801;
															assign node40801 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node40805 = (inp[0]) ? node40809 : node40806;
														assign node40806 = (inp[5]) ? 4'b1110 : 4'b1100;
														assign node40809 = (inp[5]) ? 4'b1100 : 4'b1110;
												assign node40812 = (inp[2]) ? node40822 : node40813;
													assign node40813 = (inp[5]) ? node40819 : node40814;
														assign node40814 = (inp[13]) ? 4'b0100 : node40815;
															assign node40815 = (inp[1]) ? 4'b0100 : 4'b1100;
														assign node40819 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node40822 = (inp[13]) ? node40828 : node40823;
														assign node40823 = (inp[0]) ? 4'b0100 : node40824;
															assign node40824 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node40828 = (inp[1]) ? 4'b0110 : node40829;
															assign node40829 = (inp[5]) ? node40833 : node40830;
																assign node40830 = (inp[0]) ? 4'b0110 : 4'b0100;
																assign node40833 = (inp[0]) ? 4'b0100 : 4'b0110;
							assign node40837 = (inp[10]) ? node41173 : node40838;
								assign node40838 = (inp[12]) ? node41022 : node40839;
									assign node40839 = (inp[6]) ? node40921 : node40840;
										assign node40840 = (inp[11]) ? node40880 : node40841;
											assign node40841 = (inp[1]) ? node40863 : node40842;
												assign node40842 = (inp[13]) ? node40852 : node40843;
													assign node40843 = (inp[5]) ? 4'b1100 : node40844;
														assign node40844 = (inp[2]) ? node40846 : 4'b1110;
															assign node40846 = (inp[15]) ? node40848 : 4'b1100;
																assign node40848 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node40852 = (inp[2]) ? node40854 : 4'b0110;
														assign node40854 = (inp[15]) ? 4'b0110 : node40855;
															assign node40855 = (inp[0]) ? node40859 : node40856;
																assign node40856 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node40859 = (inp[5]) ? 4'b0110 : 4'b0100;
												assign node40863 = (inp[5]) ? node40873 : node40864;
													assign node40864 = (inp[13]) ? 4'b0110 : node40865;
														assign node40865 = (inp[0]) ? node40869 : node40866;
															assign node40866 = (inp[15]) ? 4'b0100 : 4'b0110;
															assign node40869 = (inp[15]) ? 4'b0110 : 4'b0100;
													assign node40873 = (inp[15]) ? node40877 : node40874;
														assign node40874 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node40877 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node40880 = (inp[1]) ? node40902 : node40881;
												assign node40881 = (inp[13]) ? node40893 : node40882;
													assign node40882 = (inp[15]) ? 4'b0110 : node40883;
														assign node40883 = (inp[2]) ? 4'b0110 : node40884;
															assign node40884 = (inp[0]) ? node40888 : node40885;
																assign node40885 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node40888 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node40893 = (inp[5]) ? node40895 : 4'b1100;
														assign node40895 = (inp[2]) ? 4'b1100 : node40896;
															assign node40896 = (inp[0]) ? node40898 : 4'b1110;
																assign node40898 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node40902 = (inp[2]) ? node40916 : node40903;
													assign node40903 = (inp[5]) ? 4'b1110 : node40904;
														assign node40904 = (inp[13]) ? node40910 : node40905;
															assign node40905 = (inp[0]) ? 4'b1100 : node40906;
																assign node40906 = (inp[15]) ? 4'b1100 : 4'b1110;
															assign node40910 = (inp[15]) ? node40912 : 4'b1110;
																assign node40912 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node40916 = (inp[0]) ? node40918 : 4'b1100;
														assign node40918 = (inp[15]) ? 4'b1110 : 4'b1100;
										assign node40921 = (inp[11]) ? node40973 : node40922;
											assign node40922 = (inp[1]) ? node40946 : node40923;
												assign node40923 = (inp[13]) ? node40941 : node40924;
													assign node40924 = (inp[5]) ? node40934 : node40925;
														assign node40925 = (inp[2]) ? node40929 : node40926;
															assign node40926 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node40929 = (inp[0]) ? 4'b0100 : node40930;
																assign node40930 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node40934 = (inp[2]) ? node40936 : 4'b0110;
															assign node40936 = (inp[15]) ? node40938 : 4'b0110;
																assign node40938 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node40941 = (inp[5]) ? 4'b1110 : node40942;
														assign node40942 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node40946 = (inp[2]) ? node40962 : node40947;
													assign node40947 = (inp[5]) ? node40957 : node40948;
														assign node40948 = (inp[13]) ? node40952 : node40949;
															assign node40949 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node40952 = (inp[15]) ? node40954 : 4'b1110;
																assign node40954 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node40957 = (inp[15]) ? node40959 : 4'b1100;
															assign node40959 = (inp[13]) ? 4'b1110 : 4'b1100;
													assign node40962 = (inp[15]) ? node40964 : 4'b1110;
														assign node40964 = (inp[13]) ? node40970 : node40965;
															assign node40965 = (inp[0]) ? node40967 : 4'b1110;
																assign node40967 = (inp[5]) ? 4'b1100 : 4'b1110;
															assign node40970 = (inp[0]) ? 4'b1110 : 4'b1100;
											assign node40973 = (inp[1]) ? node40995 : node40974;
												assign node40974 = (inp[13]) ? node40986 : node40975;
													assign node40975 = (inp[0]) ? node40977 : 4'b1110;
														assign node40977 = (inp[2]) ? node40979 : 4'b1100;
															assign node40979 = (inp[5]) ? node40983 : node40980;
																assign node40980 = (inp[15]) ? 4'b1110 : 4'b1100;
																assign node40983 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node40986 = (inp[2]) ? 4'b0110 : node40987;
														assign node40987 = (inp[0]) ? 4'b0110 : node40988;
															assign node40988 = (inp[5]) ? node40990 : 4'b0100;
																assign node40990 = (inp[15]) ? 4'b0110 : 4'b0100;
												assign node40995 = (inp[0]) ? node41015 : node40996;
													assign node40996 = (inp[13]) ? node41010 : node40997;
														assign node40997 = (inp[2]) ? node41005 : node40998;
															assign node40998 = (inp[5]) ? node41002 : node40999;
																assign node40999 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node41002 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node41005 = (inp[5]) ? 4'b0110 : node41006;
																assign node41006 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node41010 = (inp[15]) ? 4'b0110 : node41011;
															assign node41011 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node41015 = (inp[13]) ? node41019 : node41016;
														assign node41016 = (inp[5]) ? 4'b0110 : 4'b0100;
														assign node41019 = (inp[5]) ? 4'b0100 : 4'b0110;
									assign node41022 = (inp[6]) ? node41100 : node41023;
										assign node41023 = (inp[11]) ? node41055 : node41024;
											assign node41024 = (inp[13]) ? node41044 : node41025;
												assign node41025 = (inp[1]) ? node41033 : node41026;
													assign node41026 = (inp[0]) ? 4'b1110 : node41027;
														assign node41027 = (inp[15]) ? 4'b1100 : node41028;
															assign node41028 = (inp[5]) ? 4'b1100 : 4'b1110;
													assign node41033 = (inp[15]) ? node41035 : 4'b0110;
														assign node41035 = (inp[2]) ? node41037 : 4'b0110;
															assign node41037 = (inp[0]) ? node41041 : node41038;
																assign node41038 = (inp[5]) ? 4'b0110 : 4'b0100;
																assign node41041 = (inp[5]) ? 4'b0100 : 4'b0110;
												assign node41044 = (inp[5]) ? node41050 : node41045;
													assign node41045 = (inp[15]) ? 4'b0110 : node41046;
														assign node41046 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node41050 = (inp[15]) ? node41052 : 4'b0100;
														assign node41052 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node41055 = (inp[13]) ? node41085 : node41056;
												assign node41056 = (inp[1]) ? node41074 : node41057;
													assign node41057 = (inp[2]) ? node41065 : node41058;
														assign node41058 = (inp[0]) ? node41060 : 4'b0110;
															assign node41060 = (inp[5]) ? node41062 : 4'b0110;
																assign node41062 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node41065 = (inp[0]) ? 4'b0110 : node41066;
															assign node41066 = (inp[15]) ? node41070 : node41067;
																assign node41067 = (inp[5]) ? 4'b0100 : 4'b0110;
																assign node41070 = (inp[5]) ? 4'b0110 : 4'b0100;
													assign node41074 = (inp[0]) ? 4'b1000 : node41075;
														assign node41075 = (inp[2]) ? node41079 : node41076;
															assign node41076 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node41079 = (inp[15]) ? 4'b1000 : node41080;
																assign node41080 = (inp[5]) ? 4'b1000 : 4'b1010;
												assign node41085 = (inp[5]) ? node41093 : node41086;
													assign node41086 = (inp[0]) ? node41090 : node41087;
														assign node41087 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node41090 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node41093 = (inp[0]) ? node41097 : node41094;
														assign node41094 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node41097 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node41100 = (inp[11]) ? node41138 : node41101;
											assign node41101 = (inp[1]) ? node41125 : node41102;
												assign node41102 = (inp[13]) ? node41114 : node41103;
													assign node41103 = (inp[15]) ? node41105 : 4'b0110;
														assign node41105 = (inp[2]) ? node41107 : 4'b0100;
															assign node41107 = (inp[0]) ? node41111 : node41108;
																assign node41108 = (inp[5]) ? 4'b0110 : 4'b0100;
																assign node41111 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node41114 = (inp[15]) ? node41116 : 4'b1000;
														assign node41116 = (inp[2]) ? node41118 : 4'b1000;
															assign node41118 = (inp[5]) ? node41122 : node41119;
																assign node41119 = (inp[0]) ? 4'b1010 : 4'b1000;
																assign node41122 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node41125 = (inp[5]) ? node41133 : node41126;
													assign node41126 = (inp[0]) ? node41130 : node41127;
														assign node41127 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node41130 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node41133 = (inp[2]) ? node41135 : 4'b1000;
														assign node41135 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node41138 = (inp[13]) ? node41152 : node41139;
												assign node41139 = (inp[1]) ? node41145 : node41140;
													assign node41140 = (inp[0]) ? 4'b1000 : node41141;
														assign node41141 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node41145 = (inp[0]) ? node41147 : 4'b0000;
														assign node41147 = (inp[5]) ? 4'b0000 : node41148;
															assign node41148 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node41152 = (inp[0]) ? node41160 : node41153;
													assign node41153 = (inp[5]) ? node41157 : node41154;
														assign node41154 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node41157 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node41160 = (inp[2]) ? node41168 : node41161;
														assign node41161 = (inp[1]) ? node41163 : 4'b0000;
															assign node41163 = (inp[5]) ? node41165 : 4'b0000;
																assign node41165 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node41168 = (inp[5]) ? 4'b0010 : node41169;
															assign node41169 = (inp[15]) ? 4'b0010 : 4'b0000;
								assign node41173 = (inp[12]) ? node41341 : node41174;
									assign node41174 = (inp[6]) ? node41242 : node41175;
										assign node41175 = (inp[11]) ? node41205 : node41176;
											assign node41176 = (inp[1]) ? node41192 : node41177;
												assign node41177 = (inp[13]) ? node41181 : node41178;
													assign node41178 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node41181 = (inp[5]) ? node41187 : node41182;
														assign node41182 = (inp[0]) ? node41184 : 4'b0100;
															assign node41184 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node41187 = (inp[15]) ? node41189 : 4'b0110;
															assign node41189 = (inp[2]) ? 4'b0100 : 4'b0110;
												assign node41192 = (inp[15]) ? node41200 : node41193;
													assign node41193 = (inp[5]) ? node41197 : node41194;
														assign node41194 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node41197 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node41200 = (inp[0]) ? 4'b0100 : node41201;
														assign node41201 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node41205 = (inp[13]) ? node41229 : node41206;
												assign node41206 = (inp[1]) ? node41220 : node41207;
													assign node41207 = (inp[5]) ? node41213 : node41208;
														assign node41208 = (inp[15]) ? node41210 : 4'b0100;
															assign node41210 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node41213 = (inp[0]) ? node41217 : node41214;
															assign node41214 = (inp[2]) ? 4'b0110 : 4'b0100;
															assign node41217 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node41220 = (inp[0]) ? node41222 : 4'b1010;
														assign node41222 = (inp[5]) ? node41226 : node41223;
															assign node41223 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node41226 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node41229 = (inp[15]) ? node41237 : node41230;
													assign node41230 = (inp[0]) ? node41234 : node41231;
														assign node41231 = (inp[5]) ? 4'b1000 : 4'b1010;
														assign node41234 = (inp[5]) ? 4'b1010 : 4'b1000;
													assign node41237 = (inp[5]) ? node41239 : 4'b1010;
														assign node41239 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node41242 = (inp[11]) ? node41302 : node41243;
											assign node41243 = (inp[13]) ? node41269 : node41244;
												assign node41244 = (inp[1]) ? node41260 : node41245;
													assign node41245 = (inp[2]) ? node41255 : node41246;
														assign node41246 = (inp[5]) ? 4'b0100 : node41247;
															assign node41247 = (inp[0]) ? node41251 : node41248;
																assign node41248 = (inp[15]) ? 4'b0100 : 4'b0110;
																assign node41251 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node41255 = (inp[5]) ? 4'b0110 : node41256;
															assign node41256 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node41260 = (inp[5]) ? node41264 : node41261;
														assign node41261 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node41264 = (inp[0]) ? node41266 : 4'b1000;
															assign node41266 = (inp[15]) ? 4'b1000 : 4'b1010;
												assign node41269 = (inp[2]) ? node41283 : node41270;
													assign node41270 = (inp[15]) ? node41272 : 4'b1010;
														assign node41272 = (inp[1]) ? node41278 : node41273;
															assign node41273 = (inp[0]) ? 4'b1000 : node41274;
																assign node41274 = (inp[5]) ? 4'b1010 : 4'b1000;
															assign node41278 = (inp[5]) ? 4'b1010 : node41279;
																assign node41279 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node41283 = (inp[1]) ? node41293 : node41284;
														assign node41284 = (inp[15]) ? 4'b1010 : node41285;
															assign node41285 = (inp[0]) ? node41289 : node41286;
																assign node41286 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node41289 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node41293 = (inp[0]) ? node41295 : 4'b1000;
															assign node41295 = (inp[5]) ? node41299 : node41296;
																assign node41296 = (inp[15]) ? 4'b1010 : 4'b1000;
																assign node41299 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node41302 = (inp[1]) ? node41322 : node41303;
												assign node41303 = (inp[13]) ? node41313 : node41304;
													assign node41304 = (inp[2]) ? node41308 : node41305;
														assign node41305 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node41308 = (inp[5]) ? 4'b1010 : node41309;
															assign node41309 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node41313 = (inp[15]) ? node41317 : node41314;
														assign node41314 = (inp[2]) ? 4'b0000 : 4'b0010;
														assign node41317 = (inp[0]) ? node41319 : 4'b0010;
															assign node41319 = (inp[2]) ? 4'b0010 : 4'b0000;
												assign node41322 = (inp[15]) ? node41334 : node41323;
													assign node41323 = (inp[2]) ? node41329 : node41324;
														assign node41324 = (inp[0]) ? 4'b0010 : node41325;
															assign node41325 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node41329 = (inp[0]) ? node41331 : 4'b0000;
															assign node41331 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node41334 = (inp[0]) ? node41338 : node41335;
														assign node41335 = (inp[5]) ? 4'b0010 : 4'b0000;
														assign node41338 = (inp[5]) ? 4'b0000 : 4'b0010;
									assign node41341 = (inp[6]) ? node41409 : node41342;
										assign node41342 = (inp[11]) ? node41374 : node41343;
											assign node41343 = (inp[13]) ? node41359 : node41344;
												assign node41344 = (inp[1]) ? node41352 : node41345;
													assign node41345 = (inp[2]) ? node41347 : 4'b1000;
														assign node41347 = (inp[15]) ? node41349 : 4'b1010;
															assign node41349 = (inp[5]) ? 4'b1000 : 4'b1010;
													assign node41352 = (inp[0]) ? node41354 : 4'b0010;
														assign node41354 = (inp[15]) ? node41356 : 4'b0000;
															assign node41356 = (inp[5]) ? 4'b0000 : 4'b0010;
												assign node41359 = (inp[5]) ? node41367 : node41360;
													assign node41360 = (inp[15]) ? node41364 : node41361;
														assign node41361 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node41364 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node41367 = (inp[1]) ? 4'b0010 : node41368;
														assign node41368 = (inp[0]) ? 4'b0000 : node41369;
															assign node41369 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node41374 = (inp[13]) ? node41398 : node41375;
												assign node41375 = (inp[1]) ? node41389 : node41376;
													assign node41376 = (inp[5]) ? node41382 : node41377;
														assign node41377 = (inp[15]) ? 4'b0010 : node41378;
															assign node41378 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node41382 = (inp[15]) ? node41386 : node41383;
															assign node41383 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node41386 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node41389 = (inp[5]) ? node41391 : 4'b1000;
														assign node41391 = (inp[15]) ? node41395 : node41392;
															assign node41392 = (inp[0]) ? 4'b1010 : 4'b1000;
															assign node41395 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node41398 = (inp[5]) ? node41404 : node41399;
													assign node41399 = (inp[1]) ? node41401 : 4'b1010;
														assign node41401 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node41404 = (inp[15]) ? node41406 : 4'b1000;
														assign node41406 = (inp[0]) ? 4'b1000 : 4'b1010;
										assign node41409 = (inp[11]) ? node41453 : node41410;
											assign node41410 = (inp[1]) ? node41430 : node41411;
												assign node41411 = (inp[13]) ? node41423 : node41412;
													assign node41412 = (inp[5]) ? node41418 : node41413;
														assign node41413 = (inp[15]) ? node41415 : 4'b0010;
															assign node41415 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node41418 = (inp[0]) ? 4'b0000 : node41419;
															assign node41419 = (inp[15]) ? 4'b0010 : 4'b0000;
													assign node41423 = (inp[2]) ? 4'b1000 : node41424;
														assign node41424 = (inp[0]) ? node41426 : 4'b1010;
															assign node41426 = (inp[5]) ? 4'b1010 : 4'b1000;
												assign node41430 = (inp[5]) ? node41446 : node41431;
													assign node41431 = (inp[13]) ? node41439 : node41432;
														assign node41432 = (inp[15]) ? node41436 : node41433;
															assign node41433 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node41436 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node41439 = (inp[0]) ? node41443 : node41440;
															assign node41440 = (inp[15]) ? 4'b1000 : 4'b1010;
															assign node41443 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node41446 = (inp[0]) ? node41450 : node41447;
														assign node41447 = (inp[15]) ? 4'b1010 : 4'b1000;
														assign node41450 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node41453 = (inp[1]) ? node41469 : node41454;
												assign node41454 = (inp[13]) ? node41462 : node41455;
													assign node41455 = (inp[5]) ? 4'b1000 : node41456;
														assign node41456 = (inp[0]) ? node41458 : 4'b1010;
															assign node41458 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node41462 = (inp[0]) ? node41464 : 4'b0000;
														assign node41464 = (inp[5]) ? 4'b0010 : node41465;
															assign node41465 = (inp[15]) ? 4'b0010 : 4'b0000;
												assign node41469 = (inp[2]) ? node41487 : node41470;
													assign node41470 = (inp[13]) ? node41474 : node41471;
														assign node41471 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node41474 = (inp[15]) ? node41482 : node41475;
															assign node41475 = (inp[5]) ? node41479 : node41476;
																assign node41476 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node41479 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node41482 = (inp[0]) ? 4'b0010 : node41483;
																assign node41483 = (inp[5]) ? 4'b0010 : 4'b0000;
													assign node41487 = (inp[0]) ? node41489 : 4'b0010;
														assign node41489 = (inp[15]) ? node41493 : node41490;
															assign node41490 = (inp[5]) ? 4'b0010 : 4'b0000;
															assign node41493 = (inp[5]) ? 4'b0000 : 4'b0010;
					assign node41496 = (inp[1]) ? node42972 : node41497;
						assign node41497 = (inp[15]) ? node42251 : node41498;
							assign node41498 = (inp[0]) ? node41882 : node41499;
								assign node41499 = (inp[5]) ? node41695 : node41500;
									assign node41500 = (inp[9]) ? node41594 : node41501;
										assign node41501 = (inp[4]) ? node41545 : node41502;
											assign node41502 = (inp[10]) ? node41524 : node41503;
												assign node41503 = (inp[12]) ? node41515 : node41504;
													assign node41504 = (inp[6]) ? node41506 : 4'b1110;
														assign node41506 = (inp[2]) ? 4'b0110 : node41507;
															assign node41507 = (inp[11]) ? node41511 : node41508;
																assign node41508 = (inp[13]) ? 4'b1110 : 4'b0110;
																assign node41511 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node41515 = (inp[6]) ? node41519 : node41516;
														assign node41516 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node41519 = (inp[11]) ? node41521 : 4'b1010;
															assign node41521 = (inp[13]) ? 4'b0010 : 4'b1010;
												assign node41524 = (inp[11]) ? node41538 : node41525;
													assign node41525 = (inp[12]) ? node41533 : node41526;
														assign node41526 = (inp[2]) ? node41528 : 4'b0110;
															assign node41528 = (inp[13]) ? 4'b1010 : node41529;
																assign node41529 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node41533 = (inp[13]) ? node41535 : 4'b0010;
															assign node41535 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node41538 = (inp[13]) ? node41542 : node41539;
														assign node41539 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node41542 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node41545 = (inp[12]) ? node41573 : node41546;
												assign node41546 = (inp[10]) ? node41558 : node41547;
													assign node41547 = (inp[2]) ? node41549 : 4'b1010;
														assign node41549 = (inp[13]) ? 4'b1010 : node41550;
															assign node41550 = (inp[6]) ? node41554 : node41551;
																assign node41551 = (inp[11]) ? 4'b0010 : 4'b1010;
																assign node41554 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node41558 = (inp[6]) ? node41566 : node41559;
														assign node41559 = (inp[11]) ? node41563 : node41560;
															assign node41560 = (inp[13]) ? 4'b0010 : 4'b1010;
															assign node41563 = (inp[13]) ? 4'b1100 : 4'b0010;
														assign node41566 = (inp[11]) ? node41570 : node41567;
															assign node41567 = (inp[13]) ? 4'b1100 : 4'b0010;
															assign node41570 = (inp[13]) ? 4'b0100 : 4'b1100;
												assign node41573 = (inp[10]) ? node41583 : node41574;
													assign node41574 = (inp[6]) ? node41576 : 4'b0010;
														assign node41576 = (inp[2]) ? 4'b0100 : node41577;
															assign node41577 = (inp[11]) ? 4'b1100 : node41578;
																assign node41578 = (inp[13]) ? 4'b1100 : 4'b0010;
													assign node41583 = (inp[6]) ? node41589 : node41584;
														assign node41584 = (inp[13]) ? node41586 : 4'b1100;
															assign node41586 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node41589 = (inp[13]) ? 4'b0100 : node41590;
															assign node41590 = (inp[11]) ? 4'b1100 : 4'b0100;
										assign node41594 = (inp[4]) ? node41644 : node41595;
											assign node41595 = (inp[12]) ? node41623 : node41596;
												assign node41596 = (inp[10]) ? node41610 : node41597;
													assign node41597 = (inp[2]) ? node41605 : node41598;
														assign node41598 = (inp[6]) ? 4'b0010 : node41599;
															assign node41599 = (inp[13]) ? node41601 : 4'b1010;
																assign node41601 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node41605 = (inp[6]) ? 4'b1010 : node41606;
															assign node41606 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node41610 = (inp[11]) ? node41618 : node41611;
														assign node41611 = (inp[6]) ? node41615 : node41612;
															assign node41612 = (inp[13]) ? 4'b0010 : 4'b1010;
															assign node41615 = (inp[13]) ? 4'b1100 : 4'b0010;
														assign node41618 = (inp[13]) ? 4'b1100 : node41619;
															assign node41619 = (inp[6]) ? 4'b1100 : 4'b0010;
												assign node41623 = (inp[10]) ? node41633 : node41624;
													assign node41624 = (inp[13]) ? node41630 : node41625;
														assign node41625 = (inp[6]) ? node41627 : 4'b0010;
															assign node41627 = (inp[11]) ? 4'b1100 : 4'b0010;
														assign node41630 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node41633 = (inp[2]) ? 4'b1100 : node41634;
														assign node41634 = (inp[6]) ? 4'b1100 : node41635;
															assign node41635 = (inp[11]) ? node41639 : node41636;
																assign node41636 = (inp[13]) ? 4'b0100 : 4'b1100;
																assign node41639 = (inp[13]) ? 4'b1100 : 4'b0100;
											assign node41644 = (inp[12]) ? node41674 : node41645;
												assign node41645 = (inp[10]) ? node41661 : node41646;
													assign node41646 = (inp[2]) ? node41656 : node41647;
														assign node41647 = (inp[6]) ? 4'b1100 : node41648;
															assign node41648 = (inp[13]) ? node41652 : node41649;
																assign node41649 = (inp[11]) ? 4'b0100 : 4'b1100;
																assign node41652 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node41656 = (inp[6]) ? 4'b0100 : node41657;
															assign node41657 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node41661 = (inp[11]) ? node41667 : node41662;
														assign node41662 = (inp[2]) ? node41664 : 4'b0100;
															assign node41664 = (inp[13]) ? 4'b1000 : 4'b0100;
														assign node41667 = (inp[13]) ? node41671 : node41668;
															assign node41668 = (inp[6]) ? 4'b1000 : 4'b0100;
															assign node41671 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node41674 = (inp[10]) ? node41686 : node41675;
													assign node41675 = (inp[13]) ? node41681 : node41676;
														assign node41676 = (inp[2]) ? node41678 : 4'b0100;
															assign node41678 = (inp[11]) ? 4'b1000 : 4'b0100;
														assign node41681 = (inp[6]) ? node41683 : 4'b1000;
															assign node41683 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node41686 = (inp[11]) ? node41688 : 4'b0000;
														assign node41688 = (inp[6]) ? node41692 : node41689;
															assign node41689 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node41692 = (inp[13]) ? 4'b0000 : 4'b1000;
									assign node41695 = (inp[13]) ? node41793 : node41696;
										assign node41696 = (inp[12]) ? node41754 : node41697;
											assign node41697 = (inp[2]) ? node41721 : node41698;
												assign node41698 = (inp[6]) ? node41712 : node41699;
													assign node41699 = (inp[11]) ? node41705 : node41700;
														assign node41700 = (inp[9]) ? node41702 : 4'b1000;
															assign node41702 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node41705 = (inp[4]) ? node41709 : node41706;
															assign node41706 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node41709 = (inp[9]) ? 4'b0100 : 4'b0000;
													assign node41712 = (inp[11]) ? 4'b1100 : node41713;
														assign node41713 = (inp[4]) ? node41717 : node41714;
															assign node41714 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node41717 = (inp[9]) ? 4'b0100 : 4'b0000;
												assign node41721 = (inp[9]) ? node41737 : node41722;
													assign node41722 = (inp[4]) ? node41730 : node41723;
														assign node41723 = (inp[6]) ? node41727 : node41724;
															assign node41724 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node41727 = (inp[10]) ? 4'b1000 : 4'b1100;
														assign node41730 = (inp[11]) ? node41734 : node41731;
															assign node41731 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node41734 = (inp[10]) ? 4'b1100 : 4'b1000;
													assign node41737 = (inp[4]) ? node41749 : node41738;
														assign node41738 = (inp[10]) ? node41744 : node41739;
															assign node41739 = (inp[6]) ? 4'b1000 : node41740;
																assign node41740 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node41744 = (inp[6]) ? node41746 : 4'b0000;
																assign node41746 = (inp[11]) ? 4'b1100 : 4'b0000;
														assign node41749 = (inp[11]) ? 4'b0100 : node41750;
															assign node41750 = (inp[6]) ? 4'b0100 : 4'b1100;
											assign node41754 = (inp[9]) ? node41770 : node41755;
												assign node41755 = (inp[4]) ? node41763 : node41756;
													assign node41756 = (inp[10]) ? 4'b1000 : node41757;
														assign node41757 = (inp[11]) ? 4'b1000 : node41758;
															assign node41758 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node41763 = (inp[2]) ? node41765 : 4'b1100;
														assign node41765 = (inp[10]) ? 4'b0100 : node41766;
															assign node41766 = (inp[11]) ? 4'b0000 : 4'b1000;
												assign node41770 = (inp[6]) ? node41784 : node41771;
													assign node41771 = (inp[11]) ? node41779 : node41772;
														assign node41772 = (inp[10]) ? node41776 : node41773;
															assign node41773 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node41776 = (inp[4]) ? 4'b1000 : 4'b1100;
														assign node41779 = (inp[10]) ? node41781 : 4'b0000;
															assign node41781 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node41784 = (inp[11]) ? node41790 : node41785;
														assign node41785 = (inp[4]) ? node41787 : 4'b0000;
															assign node41787 = (inp[2]) ? 4'b0000 : 4'b0100;
														assign node41790 = (inp[4]) ? 4'b1000 : 4'b1100;
										assign node41793 = (inp[9]) ? node41839 : node41794;
											assign node41794 = (inp[12]) ? node41822 : node41795;
												assign node41795 = (inp[10]) ? node41805 : node41796;
													assign node41796 = (inp[4]) ? 4'b1000 : node41797;
														assign node41797 = (inp[6]) ? node41801 : node41798;
															assign node41798 = (inp[11]) ? 4'b1100 : 4'b0100;
															assign node41801 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node41805 = (inp[4]) ? node41817 : node41806;
														assign node41806 = (inp[2]) ? node41812 : node41807;
															assign node41807 = (inp[11]) ? 4'b1000 : node41808;
																assign node41808 = (inp[6]) ? 4'b1000 : 4'b0100;
															assign node41812 = (inp[6]) ? node41814 : 4'b1000;
																assign node41814 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node41817 = (inp[2]) ? 4'b1100 : node41818;
															assign node41818 = (inp[6]) ? 4'b1100 : 4'b0000;
												assign node41822 = (inp[4]) ? node41832 : node41823;
													assign node41823 = (inp[11]) ? node41829 : node41824;
														assign node41824 = (inp[6]) ? 4'b1000 : node41825;
															assign node41825 = (inp[10]) ? 4'b0000 : 4'b0100;
														assign node41829 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node41832 = (inp[11]) ? node41836 : node41833;
														assign node41833 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node41836 = (inp[2]) ? 4'b1100 : 4'b0100;
											assign node41839 = (inp[2]) ? node41865 : node41840;
												assign node41840 = (inp[10]) ? node41852 : node41841;
													assign node41841 = (inp[6]) ? node41847 : node41842;
														assign node41842 = (inp[11]) ? node41844 : 4'b0100;
															assign node41844 = (inp[4]) ? 4'b1100 : 4'b1000;
														assign node41847 = (inp[4]) ? node41849 : 4'b1100;
															assign node41849 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node41852 = (inp[4]) ? 4'b0000 : node41853;
														assign node41853 = (inp[12]) ? node41859 : node41854;
															assign node41854 = (inp[6]) ? node41856 : 4'b0000;
																assign node41856 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node41859 = (inp[6]) ? node41861 : 4'b1100;
																assign node41861 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node41865 = (inp[4]) ? node41875 : node41866;
													assign node41866 = (inp[12]) ? 4'b0100 : node41867;
														assign node41867 = (inp[10]) ? node41869 : 4'b1000;
															assign node41869 = (inp[6]) ? node41871 : 4'b0000;
																assign node41871 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node41875 = (inp[11]) ? 4'b0000 : node41876;
														assign node41876 = (inp[10]) ? node41878 : 4'b0100;
															assign node41878 = (inp[12]) ? 4'b0000 : 4'b0100;
								assign node41882 = (inp[5]) ? node42070 : node41883;
									assign node41883 = (inp[9]) ? node41989 : node41884;
										assign node41884 = (inp[4]) ? node41938 : node41885;
											assign node41885 = (inp[12]) ? node41911 : node41886;
												assign node41886 = (inp[10]) ? node41896 : node41887;
													assign node41887 = (inp[13]) ? 4'b0100 : node41888;
														assign node41888 = (inp[11]) ? node41892 : node41889;
															assign node41889 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node41892 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node41896 = (inp[11]) ? node41906 : node41897;
														assign node41897 = (inp[2]) ? node41901 : node41898;
															assign node41898 = (inp[13]) ? 4'b1000 : 4'b0100;
															assign node41901 = (inp[13]) ? 4'b0100 : node41902;
																assign node41902 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node41906 = (inp[13]) ? 4'b1000 : node41907;
															assign node41907 = (inp[6]) ? 4'b1000 : 4'b0100;
												assign node41911 = (inp[10]) ? node41929 : node41912;
													assign node41912 = (inp[11]) ? node41922 : node41913;
														assign node41913 = (inp[2]) ? node41917 : node41914;
															assign node41914 = (inp[13]) ? 4'b1000 : 4'b0100;
															assign node41917 = (inp[6]) ? 4'b0100 : node41918;
																assign node41918 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node41922 = (inp[6]) ? node41926 : node41923;
															assign node41923 = (inp[13]) ? 4'b1000 : 4'b0100;
															assign node41926 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node41929 = (inp[13]) ? node41931 : 4'b0000;
														assign node41931 = (inp[11]) ? node41935 : node41932;
															assign node41932 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node41935 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node41938 = (inp[10]) ? node41968 : node41939;
												assign node41939 = (inp[12]) ? node41957 : node41940;
													assign node41940 = (inp[6]) ? node41948 : node41941;
														assign node41941 = (inp[13]) ? node41945 : node41942;
															assign node41942 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node41945 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node41948 = (inp[2]) ? node41952 : node41949;
															assign node41949 = (inp[11]) ? 4'b1000 : 4'b0000;
															assign node41952 = (inp[13]) ? node41954 : 4'b1000;
																assign node41954 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node41957 = (inp[6]) ? node41965 : node41958;
														assign node41958 = (inp[11]) ? node41962 : node41959;
															assign node41959 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node41962 = (inp[13]) ? 4'b1110 : 4'b0000;
														assign node41965 = (inp[2]) ? 4'b1110 : 4'b0110;
												assign node41968 = (inp[12]) ? node41978 : node41969;
													assign node41969 = (inp[13]) ? node41971 : 4'b0000;
														assign node41971 = (inp[6]) ? node41975 : node41972;
															assign node41972 = (inp[11]) ? 4'b1110 : 4'b0000;
															assign node41975 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node41978 = (inp[11]) ? node41984 : node41979;
														assign node41979 = (inp[6]) ? 4'b0110 : node41980;
															assign node41980 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node41984 = (inp[6]) ? 4'b1110 : node41985;
															assign node41985 = (inp[13]) ? 4'b1110 : 4'b0110;
										assign node41989 = (inp[4]) ? node42027 : node41990;
											assign node41990 = (inp[10]) ? node42006 : node41991;
												assign node41991 = (inp[2]) ? node42003 : node41992;
													assign node41992 = (inp[11]) ? node41994 : 4'b0000;
														assign node41994 = (inp[12]) ? node42000 : node41995;
															assign node41995 = (inp[6]) ? node41997 : 4'b0000;
																assign node41997 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node42000 = (inp[13]) ? 4'b1110 : 4'b0000;
													assign node42003 = (inp[12]) ? 4'b1110 : 4'b1000;
												assign node42006 = (inp[12]) ? node42018 : node42007;
													assign node42007 = (inp[6]) ? node42013 : node42008;
														assign node42008 = (inp[2]) ? node42010 : 4'b0000;
															assign node42010 = (inp[11]) ? 4'b1110 : 4'b1000;
														assign node42013 = (inp[2]) ? node42015 : 4'b1110;
															assign node42015 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node42018 = (inp[11]) ? node42020 : 4'b0110;
														assign node42020 = (inp[2]) ? node42022 : 4'b1110;
															assign node42022 = (inp[6]) ? 4'b0110 : node42023;
																assign node42023 = (inp[13]) ? 4'b1110 : 4'b0110;
											assign node42027 = (inp[12]) ? node42047 : node42028;
												assign node42028 = (inp[13]) ? node42036 : node42029;
													assign node42029 = (inp[2]) ? node42031 : 4'b1110;
														assign node42031 = (inp[6]) ? 4'b0110 : node42032;
															assign node42032 = (inp[11]) ? 4'b0110 : 4'b1110;
													assign node42036 = (inp[10]) ? node42040 : node42037;
														assign node42037 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node42040 = (inp[2]) ? node42042 : 4'b1010;
															assign node42042 = (inp[6]) ? node42044 : 4'b0110;
																assign node42044 = (inp[11]) ? 4'b0010 : 4'b1010;
												assign node42047 = (inp[10]) ? node42057 : node42048;
													assign node42048 = (inp[13]) ? node42054 : node42049;
														assign node42049 = (inp[11]) ? 4'b1010 : node42050;
															assign node42050 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node42054 = (inp[2]) ? 4'b0010 : 4'b1010;
													assign node42057 = (inp[13]) ? node42065 : node42058;
														assign node42058 = (inp[2]) ? node42060 : 4'b1010;
															assign node42060 = (inp[6]) ? node42062 : 4'b0010;
																assign node42062 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node42065 = (inp[11]) ? node42067 : 4'b1010;
															assign node42067 = (inp[6]) ? 4'b0010 : 4'b1010;
									assign node42070 = (inp[6]) ? node42152 : node42071;
										assign node42071 = (inp[12]) ? node42103 : node42072;
											assign node42072 = (inp[13]) ? node42090 : node42073;
												assign node42073 = (inp[11]) ? node42079 : node42074;
													assign node42074 = (inp[2]) ? node42076 : 4'b1110;
														assign node42076 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node42079 = (inp[10]) ? node42085 : node42080;
														assign node42080 = (inp[4]) ? node42082 : 4'b0010;
															assign node42082 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node42085 = (inp[4]) ? 4'b0010 : node42086;
															assign node42086 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node42090 = (inp[11]) ? node42098 : node42091;
													assign node42091 = (inp[4]) ? node42095 : node42092;
														assign node42092 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node42095 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node42098 = (inp[2]) ? 4'b1110 : node42099;
														assign node42099 = (inp[9]) ? 4'b1010 : 4'b1110;
											assign node42103 = (inp[11]) ? node42127 : node42104;
												assign node42104 = (inp[13]) ? node42120 : node42105;
													assign node42105 = (inp[4]) ? node42113 : node42106;
														assign node42106 = (inp[9]) ? node42110 : node42107;
															assign node42107 = (inp[10]) ? 4'b1010 : 4'b1110;
															assign node42110 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node42113 = (inp[9]) ? node42117 : node42114;
															assign node42114 = (inp[10]) ? 4'b1110 : 4'b1010;
															assign node42117 = (inp[10]) ? 4'b1010 : 4'b1110;
													assign node42120 = (inp[2]) ? node42122 : 4'b0010;
														assign node42122 = (inp[10]) ? node42124 : 4'b0110;
															assign node42124 = (inp[4]) ? 4'b0010 : 4'b0110;
												assign node42127 = (inp[13]) ? node42141 : node42128;
													assign node42128 = (inp[4]) ? node42136 : node42129;
														assign node42129 = (inp[10]) ? node42133 : node42130;
															assign node42130 = (inp[2]) ? 4'b0010 : 4'b0110;
															assign node42133 = (inp[9]) ? 4'b0110 : 4'b0010;
														assign node42136 = (inp[10]) ? 4'b0110 : node42137;
															assign node42137 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node42141 = (inp[10]) ? node42147 : node42142;
														assign node42142 = (inp[2]) ? 4'b1010 : node42143;
															assign node42143 = (inp[4]) ? 4'b1110 : 4'b1010;
														assign node42147 = (inp[9]) ? 4'b1110 : node42148;
															assign node42148 = (inp[2]) ? 4'b1110 : 4'b1010;
										assign node42152 = (inp[13]) ? node42204 : node42153;
											assign node42153 = (inp[11]) ? node42181 : node42154;
												assign node42154 = (inp[12]) ? node42174 : node42155;
													assign node42155 = (inp[2]) ? node42161 : node42156;
														assign node42156 = (inp[10]) ? 4'b0110 : node42157;
															assign node42157 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node42161 = (inp[10]) ? node42169 : node42162;
															assign node42162 = (inp[9]) ? node42166 : node42163;
																assign node42163 = (inp[4]) ? 4'b0010 : 4'b0110;
																assign node42166 = (inp[4]) ? 4'b0110 : 4'b0010;
															assign node42169 = (inp[9]) ? node42171 : 4'b0010;
																assign node42171 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node42174 = (inp[4]) ? 4'b0010 : node42175;
														assign node42175 = (inp[10]) ? node42177 : 4'b0010;
															assign node42177 = (inp[2]) ? 4'b0110 : 4'b0010;
												assign node42181 = (inp[9]) ? node42195 : node42182;
													assign node42182 = (inp[2]) ? node42188 : node42183;
														assign node42183 = (inp[4]) ? node42185 : 4'b1010;
															assign node42185 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node42188 = (inp[10]) ? 4'b1110 : node42189;
															assign node42189 = (inp[4]) ? node42191 : 4'b1110;
																assign node42191 = (inp[12]) ? 4'b1110 : 4'b1010;
													assign node42195 = (inp[4]) ? node42199 : node42196;
														assign node42196 = (inp[10]) ? 4'b1110 : 4'b1010;
														assign node42199 = (inp[10]) ? 4'b1010 : node42200;
															assign node42200 = (inp[12]) ? 4'b1010 : 4'b1110;
											assign node42204 = (inp[11]) ? node42234 : node42205;
												assign node42205 = (inp[12]) ? node42221 : node42206;
													assign node42206 = (inp[2]) ? 4'b1010 : node42207;
														assign node42207 = (inp[9]) ? node42215 : node42208;
															assign node42208 = (inp[10]) ? node42212 : node42209;
																assign node42209 = (inp[4]) ? 4'b1010 : 4'b1110;
																assign node42212 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node42215 = (inp[10]) ? node42217 : 4'b1010;
																assign node42217 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node42221 = (inp[2]) ? node42229 : node42222;
														assign node42222 = (inp[9]) ? node42226 : node42223;
															assign node42223 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node42226 = (inp[4]) ? 4'b1010 : 4'b1110;
														assign node42229 = (inp[9]) ? 4'b1110 : node42230;
															assign node42230 = (inp[4]) ? 4'b1110 : 4'b1010;
												assign node42234 = (inp[2]) ? node42244 : node42235;
													assign node42235 = (inp[12]) ? 4'b0010 : node42236;
														assign node42236 = (inp[4]) ? 4'b0010 : node42237;
															assign node42237 = (inp[9]) ? 4'b0010 : node42238;
																assign node42238 = (inp[10]) ? 4'b0010 : 4'b0110;
													assign node42244 = (inp[12]) ? node42246 : 4'b0110;
														assign node42246 = (inp[4]) ? 4'b0010 : node42247;
															assign node42247 = (inp[9]) ? 4'b0110 : 4'b0010;
							assign node42251 = (inp[0]) ? node42573 : node42252;
								assign node42252 = (inp[5]) ? node42408 : node42253;
									assign node42253 = (inp[4]) ? node42325 : node42254;
										assign node42254 = (inp[9]) ? node42290 : node42255;
											assign node42255 = (inp[12]) ? node42277 : node42256;
												assign node42256 = (inp[6]) ? node42266 : node42257;
													assign node42257 = (inp[2]) ? node42259 : 4'b0100;
														assign node42259 = (inp[11]) ? node42263 : node42260;
															assign node42260 = (inp[13]) ? 4'b0100 : 4'b1100;
															assign node42263 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node42266 = (inp[10]) ? node42272 : node42267;
														assign node42267 = (inp[11]) ? 4'b0100 : node42268;
															assign node42268 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node42272 = (inp[13]) ? 4'b1000 : node42273;
															assign node42273 = (inp[11]) ? 4'b1000 : 4'b0100;
												assign node42277 = (inp[10]) ? node42285 : node42278;
													assign node42278 = (inp[6]) ? 4'b1000 : node42279;
														assign node42279 = (inp[13]) ? 4'b1000 : node42280;
															assign node42280 = (inp[2]) ? 4'b1100 : 4'b0100;
													assign node42285 = (inp[6]) ? node42287 : 4'b0000;
														assign node42287 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node42290 = (inp[10]) ? node42304 : node42291;
												assign node42291 = (inp[12]) ? node42301 : node42292;
													assign node42292 = (inp[13]) ? 4'b1000 : node42293;
														assign node42293 = (inp[2]) ? node42295 : 4'b0000;
															assign node42295 = (inp[11]) ? 4'b1000 : node42296;
																assign node42296 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node42301 = (inp[6]) ? 4'b1110 : 4'b0000;
												assign node42304 = (inp[11]) ? node42318 : node42305;
													assign node42305 = (inp[12]) ? node42313 : node42306;
														assign node42306 = (inp[13]) ? node42310 : node42307;
															assign node42307 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node42310 = (inp[6]) ? 4'b1110 : 4'b0000;
														assign node42313 = (inp[6]) ? 4'b0110 : node42314;
															assign node42314 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node42318 = (inp[6]) ? node42322 : node42319;
														assign node42319 = (inp[13]) ? 4'b1110 : 4'b0110;
														assign node42322 = (inp[13]) ? 4'b0110 : 4'b1110;
										assign node42325 = (inp[9]) ? node42369 : node42326;
											assign node42326 = (inp[12]) ? node42350 : node42327;
												assign node42327 = (inp[10]) ? node42341 : node42328;
													assign node42328 = (inp[11]) ? node42336 : node42329;
														assign node42329 = (inp[13]) ? node42333 : node42330;
															assign node42330 = (inp[6]) ? 4'b0000 : 4'b1000;
															assign node42333 = (inp[6]) ? 4'b1000 : 4'b0000;
														assign node42336 = (inp[6]) ? node42338 : 4'b0000;
															assign node42338 = (inp[13]) ? 4'b0000 : 4'b1000;
													assign node42341 = (inp[11]) ? 4'b1110 : node42342;
														assign node42342 = (inp[6]) ? node42346 : node42343;
															assign node42343 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node42346 = (inp[13]) ? 4'b1110 : 4'b0000;
												assign node42350 = (inp[13]) ? node42362 : node42351;
													assign node42351 = (inp[10]) ? node42357 : node42352;
														assign node42352 = (inp[6]) ? node42354 : 4'b0000;
															assign node42354 = (inp[11]) ? 4'b1110 : 4'b0000;
														assign node42357 = (inp[6]) ? node42359 : 4'b0110;
															assign node42359 = (inp[11]) ? 4'b1110 : 4'b0110;
													assign node42362 = (inp[11]) ? node42366 : node42363;
														assign node42363 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node42366 = (inp[6]) ? 4'b0110 : 4'b1110;
											assign node42369 = (inp[12]) ? node42385 : node42370;
												assign node42370 = (inp[6]) ? node42376 : node42371;
													assign node42371 = (inp[11]) ? 4'b0110 : node42372;
														assign node42372 = (inp[10]) ? 4'b0110 : 4'b1110;
													assign node42376 = (inp[11]) ? node42380 : node42377;
														assign node42377 = (inp[13]) ? 4'b1110 : 4'b0110;
														assign node42380 = (inp[10]) ? 4'b1010 : node42381;
															assign node42381 = (inp[13]) ? 4'b0110 : 4'b1110;
												assign node42385 = (inp[10]) ? node42397 : node42386;
													assign node42386 = (inp[11]) ? node42390 : node42387;
														assign node42387 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node42390 = (inp[2]) ? 4'b1010 : node42391;
															assign node42391 = (inp[13]) ? node42393 : 4'b0110;
																assign node42393 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node42397 = (inp[6]) ? node42403 : node42398;
														assign node42398 = (inp[13]) ? node42400 : 4'b0010;
															assign node42400 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node42403 = (inp[11]) ? node42405 : 4'b1010;
															assign node42405 = (inp[13]) ? 4'b0010 : 4'b1010;
									assign node42408 = (inp[4]) ? node42498 : node42409;
										assign node42409 = (inp[2]) ? node42457 : node42410;
											assign node42410 = (inp[10]) ? node42440 : node42411;
												assign node42411 = (inp[9]) ? node42425 : node42412;
													assign node42412 = (inp[11]) ? node42418 : node42413;
														assign node42413 = (inp[13]) ? node42415 : 4'b1110;
															assign node42415 = (inp[6]) ? 4'b1110 : 4'b0110;
														assign node42418 = (inp[12]) ? node42420 : 4'b1110;
															assign node42420 = (inp[13]) ? node42422 : 4'b0110;
																assign node42422 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node42425 = (inp[12]) ? node42435 : node42426;
														assign node42426 = (inp[13]) ? node42428 : 4'b0010;
															assign node42428 = (inp[6]) ? node42432 : node42429;
																assign node42429 = (inp[11]) ? 4'b1010 : 4'b0010;
																assign node42432 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node42435 = (inp[11]) ? node42437 : 4'b0010;
															assign node42437 = (inp[13]) ? 4'b0110 : 4'b1110;
												assign node42440 = (inp[9]) ? node42454 : node42441;
													assign node42441 = (inp[12]) ? node42443 : 4'b0010;
														assign node42443 = (inp[11]) ? node42449 : node42444;
															assign node42444 = (inp[13]) ? 4'b0010 : node42445;
																assign node42445 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node42449 = (inp[6]) ? 4'b1010 : node42450;
																assign node42450 = (inp[13]) ? 4'b1010 : 4'b0010;
													assign node42454 = (inp[12]) ? 4'b0110 : 4'b0010;
											assign node42457 = (inp[6]) ? node42481 : node42458;
												assign node42458 = (inp[9]) ? node42472 : node42459;
													assign node42459 = (inp[10]) ? node42465 : node42460;
														assign node42460 = (inp[11]) ? 4'b0110 : node42461;
															assign node42461 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node42465 = (inp[12]) ? node42469 : node42466;
															assign node42466 = (inp[11]) ? 4'b1010 : 4'b0110;
															assign node42469 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node42472 = (inp[12]) ? node42478 : node42473;
														assign node42473 = (inp[13]) ? 4'b0010 : node42474;
															assign node42474 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node42478 = (inp[10]) ? 4'b0110 : 4'b0010;
												assign node42481 = (inp[9]) ? node42495 : node42482;
													assign node42482 = (inp[12]) ? node42488 : node42483;
														assign node42483 = (inp[11]) ? node42485 : 4'b0110;
															assign node42485 = (inp[13]) ? 4'b0110 : 4'b1110;
														assign node42488 = (inp[10]) ? node42490 : 4'b1010;
															assign node42490 = (inp[13]) ? 4'b0010 : node42491;
																assign node42491 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node42495 = (inp[10]) ? 4'b1110 : 4'b0110;
										assign node42498 = (inp[12]) ? node42528 : node42499;
											assign node42499 = (inp[9]) ? node42515 : node42500;
												assign node42500 = (inp[10]) ? node42510 : node42501;
													assign node42501 = (inp[11]) ? 4'b1010 : node42502;
														assign node42502 = (inp[13]) ? node42506 : node42503;
															assign node42503 = (inp[6]) ? 4'b0010 : 4'b1010;
															assign node42506 = (inp[6]) ? 4'b1010 : 4'b0010;
													assign node42510 = (inp[13]) ? node42512 : 4'b0010;
														assign node42512 = (inp[6]) ? 4'b1110 : 4'b0010;
												assign node42515 = (inp[11]) ? node42521 : node42516;
													assign node42516 = (inp[13]) ? 4'b0110 : node42517;
														assign node42517 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node42521 = (inp[2]) ? node42523 : 4'b1010;
														assign node42523 = (inp[6]) ? node42525 : 4'b0110;
															assign node42525 = (inp[13]) ? 4'b0110 : 4'b1010;
											assign node42528 = (inp[9]) ? node42548 : node42529;
												assign node42529 = (inp[10]) ? node42543 : node42530;
													assign node42530 = (inp[13]) ? node42538 : node42531;
														assign node42531 = (inp[2]) ? 4'b0010 : node42532;
															assign node42532 = (inp[11]) ? 4'b0010 : node42533;
																assign node42533 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node42538 = (inp[11]) ? node42540 : 4'b0010;
															assign node42540 = (inp[2]) ? 4'b0110 : 4'b1110;
													assign node42543 = (inp[13]) ? 4'b0110 : node42544;
														assign node42544 = (inp[6]) ? 4'b1110 : 4'b0110;
												assign node42548 = (inp[10]) ? node42560 : node42549;
													assign node42549 = (inp[6]) ? node42555 : node42550;
														assign node42550 = (inp[13]) ? 4'b0110 : node42551;
															assign node42551 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node42555 = (inp[2]) ? 4'b1010 : node42556;
															assign node42556 = (inp[13]) ? 4'b0010 : 4'b0110;
													assign node42560 = (inp[11]) ? node42566 : node42561;
														assign node42561 = (inp[13]) ? node42563 : 4'b0010;
															assign node42563 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node42566 = (inp[2]) ? 4'b1010 : node42567;
															assign node42567 = (inp[13]) ? 4'b0010 : node42568;
																assign node42568 = (inp[6]) ? 4'b1010 : 4'b0010;
								assign node42573 = (inp[5]) ? node42761 : node42574;
									assign node42574 = (inp[4]) ? node42666 : node42575;
										assign node42575 = (inp[9]) ? node42617 : node42576;
											assign node42576 = (inp[12]) ? node42596 : node42577;
												assign node42577 = (inp[10]) ? node42587 : node42578;
													assign node42578 = (inp[11]) ? node42580 : 4'b1110;
														assign node42580 = (inp[6]) ? node42584 : node42581;
															assign node42581 = (inp[13]) ? 4'b1110 : 4'b0110;
															assign node42584 = (inp[13]) ? 4'b0110 : 4'b1110;
													assign node42587 = (inp[13]) ? 4'b1010 : node42588;
														assign node42588 = (inp[6]) ? node42592 : node42589;
															assign node42589 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node42592 = (inp[11]) ? 4'b1010 : 4'b0110;
												assign node42596 = (inp[11]) ? node42606 : node42597;
													assign node42597 = (inp[13]) ? node42603 : node42598;
														assign node42598 = (inp[6]) ? node42600 : 4'b1110;
															assign node42600 = (inp[10]) ? 4'b0010 : 4'b0110;
														assign node42603 = (inp[6]) ? 4'b1010 : 4'b0110;
													assign node42606 = (inp[2]) ? node42612 : node42607;
														assign node42607 = (inp[10]) ? node42609 : 4'b1010;
															assign node42609 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node42612 = (inp[13]) ? 4'b0010 : node42613;
															assign node42613 = (inp[6]) ? 4'b1010 : 4'b0010;
											assign node42617 = (inp[12]) ? node42645 : node42618;
												assign node42618 = (inp[6]) ? node42632 : node42619;
													assign node42619 = (inp[2]) ? node42625 : node42620;
														assign node42620 = (inp[10]) ? 4'b0010 : node42621;
															assign node42621 = (inp[13]) ? 4'b0010 : 4'b1010;
														assign node42625 = (inp[13]) ? node42629 : node42626;
															assign node42626 = (inp[11]) ? 4'b0010 : 4'b1010;
															assign node42629 = (inp[11]) ? 4'b1010 : 4'b0010;
													assign node42632 = (inp[10]) ? node42636 : node42633;
														assign node42633 = (inp[13]) ? 4'b0010 : 4'b1010;
														assign node42636 = (inp[2]) ? node42640 : node42637;
															assign node42637 = (inp[11]) ? 4'b1100 : 4'b0010;
															assign node42640 = (inp[11]) ? node42642 : 4'b1100;
																assign node42642 = (inp[13]) ? 4'b0100 : 4'b1100;
												assign node42645 = (inp[10]) ? node42651 : node42646;
													assign node42646 = (inp[11]) ? 4'b1100 : node42647;
														assign node42647 = (inp[13]) ? 4'b1100 : 4'b1010;
													assign node42651 = (inp[11]) ? node42661 : node42652;
														assign node42652 = (inp[2]) ? 4'b0100 : node42653;
															assign node42653 = (inp[13]) ? node42657 : node42654;
																assign node42654 = (inp[6]) ? 4'b0100 : 4'b1100;
																assign node42657 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node42661 = (inp[13]) ? 4'b1100 : node42662;
															assign node42662 = (inp[6]) ? 4'b1100 : 4'b0100;
										assign node42666 = (inp[9]) ? node42712 : node42667;
											assign node42667 = (inp[12]) ? node42683 : node42668;
												assign node42668 = (inp[10]) ? node42676 : node42669;
													assign node42669 = (inp[2]) ? 4'b0010 : node42670;
														assign node42670 = (inp[13]) ? 4'b0010 : node42671;
															assign node42671 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node42676 = (inp[13]) ? node42680 : node42677;
														assign node42677 = (inp[6]) ? 4'b0010 : 4'b1010;
														assign node42680 = (inp[6]) ? 4'b1100 : 4'b0010;
												assign node42683 = (inp[10]) ? node42693 : node42684;
													assign node42684 = (inp[6]) ? node42690 : node42685;
														assign node42685 = (inp[11]) ? 4'b0010 : node42686;
															assign node42686 = (inp[13]) ? 4'b0010 : 4'b1010;
														assign node42690 = (inp[13]) ? 4'b0100 : 4'b1100;
													assign node42693 = (inp[6]) ? node42705 : node42694;
														assign node42694 = (inp[2]) ? node42700 : node42695;
															assign node42695 = (inp[11]) ? node42697 : 4'b0100;
																assign node42697 = (inp[13]) ? 4'b1100 : 4'b0100;
															assign node42700 = (inp[11]) ? 4'b0100 : node42701;
																assign node42701 = (inp[13]) ? 4'b0100 : 4'b1100;
														assign node42705 = (inp[11]) ? node42709 : node42706;
															assign node42706 = (inp[2]) ? 4'b0100 : 4'b1100;
															assign node42709 = (inp[2]) ? 4'b1100 : 4'b0100;
											assign node42712 = (inp[10]) ? node42736 : node42713;
												assign node42713 = (inp[12]) ? node42725 : node42714;
													assign node42714 = (inp[13]) ? node42720 : node42715;
														assign node42715 = (inp[2]) ? 4'b1100 : node42716;
															assign node42716 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node42720 = (inp[11]) ? 4'b0100 : node42721;
															assign node42721 = (inp[6]) ? 4'b1100 : 4'b0100;
													assign node42725 = (inp[13]) ? node42731 : node42726;
														assign node42726 = (inp[2]) ? 4'b0100 : node42727;
															assign node42727 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node42731 = (inp[11]) ? node42733 : 4'b0100;
															assign node42733 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node42736 = (inp[12]) ? node42746 : node42737;
													assign node42737 = (inp[13]) ? node42741 : node42738;
														assign node42738 = (inp[2]) ? 4'b1100 : 4'b0100;
														assign node42741 = (inp[6]) ? node42743 : 4'b1000;
															assign node42743 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node42746 = (inp[11]) ? node42756 : node42747;
														assign node42747 = (inp[2]) ? node42753 : node42748;
															assign node42748 = (inp[6]) ? node42750 : 4'b0000;
																assign node42750 = (inp[13]) ? 4'b1000 : 4'b0000;
															assign node42753 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node42756 = (inp[13]) ? node42758 : 4'b1000;
															assign node42758 = (inp[6]) ? 4'b0000 : 4'b1000;
									assign node42761 = (inp[4]) ? node42867 : node42762;
										assign node42762 = (inp[2]) ? node42818 : node42763;
											assign node42763 = (inp[6]) ? node42799 : node42764;
												assign node42764 = (inp[12]) ? node42778 : node42765;
													assign node42765 = (inp[13]) ? node42773 : node42766;
														assign node42766 = (inp[11]) ? node42770 : node42767;
															assign node42767 = (inp[9]) ? 4'b1000 : 4'b1100;
															assign node42770 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node42773 = (inp[10]) ? node42775 : 4'b1000;
															assign node42775 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node42778 = (inp[11]) ? node42790 : node42779;
														assign node42779 = (inp[13]) ? node42783 : node42780;
															assign node42780 = (inp[10]) ? 4'b1100 : 4'b1000;
															assign node42783 = (inp[9]) ? node42787 : node42784;
																assign node42784 = (inp[10]) ? 4'b0000 : 4'b0100;
																assign node42787 = (inp[10]) ? 4'b0100 : 4'b0000;
														assign node42790 = (inp[13]) ? node42796 : node42791;
															assign node42791 = (inp[9]) ? 4'b0000 : node42792;
																assign node42792 = (inp[10]) ? 4'b0000 : 4'b0100;
															assign node42796 = (inp[9]) ? 4'b1100 : 4'b1000;
												assign node42799 = (inp[12]) ? node42807 : node42800;
													assign node42800 = (inp[13]) ? node42804 : node42801;
														assign node42801 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node42804 = (inp[11]) ? 4'b0100 : 4'b1000;
													assign node42807 = (inp[9]) ? node42813 : node42808;
														assign node42808 = (inp[11]) ? 4'b1000 : node42809;
															assign node42809 = (inp[13]) ? 4'b1000 : 4'b0100;
														assign node42813 = (inp[13]) ? node42815 : 4'b1100;
															assign node42815 = (inp[11]) ? 4'b0100 : 4'b1100;
											assign node42818 = (inp[11]) ? node42848 : node42819;
												assign node42819 = (inp[12]) ? node42835 : node42820;
													assign node42820 = (inp[9]) ? node42828 : node42821;
														assign node42821 = (inp[10]) ? 4'b0100 : node42822;
															assign node42822 = (inp[6]) ? node42824 : 4'b0100;
																assign node42824 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node42828 = (inp[6]) ? node42832 : node42829;
															assign node42829 = (inp[13]) ? 4'b0000 : 4'b1000;
															assign node42832 = (inp[13]) ? 4'b1100 : 4'b0000;
													assign node42835 = (inp[10]) ? node42843 : node42836;
														assign node42836 = (inp[9]) ? node42838 : 4'b1000;
															assign node42838 = (inp[13]) ? 4'b0000 : node42839;
																assign node42839 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node42843 = (inp[9]) ? 4'b1100 : node42844;
															assign node42844 = (inp[13]) ? 4'b0000 : 4'b1000;
												assign node42848 = (inp[12]) ? node42862 : node42849;
													assign node42849 = (inp[6]) ? node42855 : node42850;
														assign node42850 = (inp[13]) ? 4'b1000 : node42851;
															assign node42851 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node42855 = (inp[13]) ? 4'b0000 : node42856;
															assign node42856 = (inp[10]) ? node42858 : 4'b1000;
																assign node42858 = (inp[9]) ? 4'b1100 : 4'b1000;
													assign node42862 = (inp[9]) ? 4'b0100 : node42863;
														assign node42863 = (inp[6]) ? 4'b0000 : 4'b0100;
										assign node42867 = (inp[12]) ? node42915 : node42868;
											assign node42868 = (inp[9]) ? node42888 : node42869;
												assign node42869 = (inp[10]) ? node42875 : node42870;
													assign node42870 = (inp[13]) ? 4'b0000 : node42871;
														assign node42871 = (inp[2]) ? 4'b1000 : 4'b0000;
													assign node42875 = (inp[13]) ? node42881 : node42876;
														assign node42876 = (inp[2]) ? node42878 : 4'b0000;
															assign node42878 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node42881 = (inp[11]) ? node42885 : node42882;
															assign node42882 = (inp[6]) ? 4'b1100 : 4'b0000;
															assign node42885 = (inp[6]) ? 4'b0100 : 4'b1100;
												assign node42888 = (inp[10]) ? node42900 : node42889;
													assign node42889 = (inp[13]) ? node42895 : node42890;
														assign node42890 = (inp[11]) ? node42892 : 4'b1100;
															assign node42892 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node42895 = (inp[6]) ? 4'b0100 : node42896;
															assign node42896 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node42900 = (inp[13]) ? node42908 : node42901;
														assign node42901 = (inp[2]) ? 4'b0100 : node42902;
															assign node42902 = (inp[11]) ? 4'b0100 : node42903;
																assign node42903 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node42908 = (inp[6]) ? node42912 : node42909;
															assign node42909 = (inp[11]) ? 4'b1000 : 4'b0100;
															assign node42912 = (inp[11]) ? 4'b0000 : 4'b1000;
											assign node42915 = (inp[9]) ? node42945 : node42916;
												assign node42916 = (inp[10]) ? node42932 : node42917;
													assign node42917 = (inp[6]) ? node42921 : node42918;
														assign node42918 = (inp[13]) ? 4'b0000 : 4'b1000;
														assign node42921 = (inp[2]) ? node42927 : node42922;
															assign node42922 = (inp[13]) ? node42924 : 4'b1100;
																assign node42924 = (inp[11]) ? 4'b0100 : 4'b1100;
															assign node42927 = (inp[13]) ? node42929 : 4'b0000;
																assign node42929 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node42932 = (inp[6]) ? node42940 : node42933;
														assign node42933 = (inp[11]) ? node42937 : node42934;
															assign node42934 = (inp[13]) ? 4'b0100 : 4'b1100;
															assign node42937 = (inp[13]) ? 4'b1100 : 4'b0100;
														assign node42940 = (inp[11]) ? node42942 : 4'b0100;
															assign node42942 = (inp[13]) ? 4'b0100 : 4'b1100;
												assign node42945 = (inp[10]) ? node42957 : node42946;
													assign node42946 = (inp[13]) ? node42950 : node42947;
														assign node42947 = (inp[6]) ? 4'b0100 : 4'b1100;
														assign node42950 = (inp[11]) ? node42954 : node42951;
															assign node42951 = (inp[6]) ? 4'b1000 : 4'b0100;
															assign node42954 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node42957 = (inp[2]) ? node42965 : node42958;
														assign node42958 = (inp[11]) ? 4'b1000 : node42959;
															assign node42959 = (inp[6]) ? node42961 : 4'b1000;
																assign node42961 = (inp[13]) ? 4'b1000 : 4'b0000;
														assign node42965 = (inp[11]) ? 4'b0000 : node42966;
															assign node42966 = (inp[13]) ? node42968 : 4'b1000;
																assign node42968 = (inp[6]) ? 4'b1000 : 4'b0000;
						assign node42972 = (inp[2]) ? node43656 : node42973;
							assign node42973 = (inp[9]) ? node43343 : node42974;
								assign node42974 = (inp[4]) ? node43156 : node42975;
									assign node42975 = (inp[10]) ? node43067 : node42976;
										assign node42976 = (inp[12]) ? node43030 : node42977;
											assign node42977 = (inp[11]) ? node43009 : node42978;
												assign node42978 = (inp[6]) ? node42988 : node42979;
													assign node42979 = (inp[5]) ? node42985 : node42980;
														assign node42980 = (inp[0]) ? 4'b0100 : node42981;
															assign node42981 = (inp[15]) ? 4'b0100 : 4'b0110;
														assign node42985 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node42988 = (inp[13]) ? node43002 : node42989;
														assign node42989 = (inp[0]) ? node42997 : node42990;
															assign node42990 = (inp[5]) ? node42994 : node42991;
																assign node42991 = (inp[15]) ? 4'b1100 : 4'b1110;
																assign node42994 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node42997 = (inp[5]) ? node42999 : 4'b1110;
																assign node42999 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node43002 = (inp[0]) ? 4'b1100 : node43003;
															assign node43003 = (inp[15]) ? node43005 : 4'b1100;
																assign node43005 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node43009 = (inp[6]) ? node43013 : node43010;
													assign node43010 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node43013 = (inp[15]) ? node43025 : node43014;
														assign node43014 = (inp[13]) ? node43020 : node43015;
															assign node43015 = (inp[5]) ? node43017 : 4'b0110;
																assign node43017 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node43020 = (inp[5]) ? 4'b0110 : node43021;
																assign node43021 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node43025 = (inp[0]) ? 4'b0100 : node43026;
															assign node43026 = (inp[5]) ? 4'b0110 : 4'b0100;
											assign node43030 = (inp[6]) ? node43050 : node43031;
												assign node43031 = (inp[11]) ? node43045 : node43032;
													assign node43032 = (inp[5]) ? node43040 : node43033;
														assign node43033 = (inp[0]) ? node43037 : node43034;
															assign node43034 = (inp[13]) ? 4'b0100 : 4'b0110;
															assign node43037 = (inp[13]) ? 4'b0110 : 4'b0100;
														assign node43040 = (inp[0]) ? 4'b0110 : node43041;
															assign node43041 = (inp[13]) ? 4'b0100 : 4'b0110;
													assign node43045 = (inp[13]) ? 4'b1010 : node43046;
														assign node43046 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node43050 = (inp[11]) ? node43054 : node43051;
													assign node43051 = (inp[13]) ? 4'b1000 : 4'b1010;
													assign node43054 = (inp[15]) ? node43060 : node43055;
														assign node43055 = (inp[5]) ? node43057 : 4'b0000;
															assign node43057 = (inp[13]) ? 4'b0010 : 4'b0000;
														assign node43060 = (inp[5]) ? node43064 : node43061;
															assign node43061 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node43064 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node43067 = (inp[11]) ? node43113 : node43068;
											assign node43068 = (inp[6]) ? node43096 : node43069;
												assign node43069 = (inp[12]) ? node43083 : node43070;
													assign node43070 = (inp[13]) ? node43078 : node43071;
														assign node43071 = (inp[0]) ? 4'b0110 : node43072;
															assign node43072 = (inp[5]) ? node43074 : 4'b0100;
																assign node43074 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node43078 = (inp[0]) ? 4'b0100 : node43079;
															assign node43079 = (inp[5]) ? 4'b0100 : 4'b0110;
													assign node43083 = (inp[5]) ? node43091 : node43084;
														assign node43084 = (inp[0]) ? node43088 : node43085;
															assign node43085 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node43088 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node43091 = (inp[15]) ? node43093 : 4'b0010;
															assign node43093 = (inp[0]) ? 4'b0000 : 4'b0010;
												assign node43096 = (inp[5]) ? node43108 : node43097;
													assign node43097 = (inp[12]) ? node43099 : 4'b1010;
														assign node43099 = (inp[13]) ? node43101 : 4'b1010;
															assign node43101 = (inp[0]) ? node43105 : node43102;
																assign node43102 = (inp[15]) ? 4'b1000 : 4'b1010;
																assign node43105 = (inp[15]) ? 4'b1010 : 4'b1000;
													assign node43108 = (inp[15]) ? 4'b1000 : node43109;
														assign node43109 = (inp[0]) ? 4'b1010 : 4'b1000;
											assign node43113 = (inp[6]) ? node43139 : node43114;
												assign node43114 = (inp[13]) ? node43130 : node43115;
													assign node43115 = (inp[12]) ? node43125 : node43116;
														assign node43116 = (inp[0]) ? 4'b1010 : node43117;
															assign node43117 = (inp[15]) ? node43121 : node43118;
																assign node43118 = (inp[5]) ? 4'b1000 : 4'b1010;
																assign node43121 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node43125 = (inp[5]) ? node43127 : 4'b1010;
															assign node43127 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node43130 = (inp[5]) ? 4'b1000 : node43131;
														assign node43131 = (inp[15]) ? node43135 : node43132;
															assign node43132 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node43135 = (inp[0]) ? 4'b1010 : 4'b1000;
												assign node43139 = (inp[12]) ? node43151 : node43140;
													assign node43140 = (inp[15]) ? 4'b0010 : node43141;
														assign node43141 = (inp[13]) ? 4'b0000 : node43142;
															assign node43142 = (inp[5]) ? node43146 : node43143;
																assign node43143 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node43146 = (inp[0]) ? 4'b0010 : 4'b0000;
													assign node43151 = (inp[5]) ? node43153 : 4'b0000;
														assign node43153 = (inp[13]) ? 4'b0010 : 4'b0000;
									assign node43156 = (inp[10]) ? node43272 : node43157;
										assign node43157 = (inp[12]) ? node43227 : node43158;
											assign node43158 = (inp[13]) ? node43194 : node43159;
												assign node43159 = (inp[15]) ? node43175 : node43160;
													assign node43160 = (inp[6]) ? node43168 : node43161;
														assign node43161 = (inp[5]) ? node43165 : node43162;
															assign node43162 = (inp[0]) ? 4'b1000 : 4'b1010;
															assign node43165 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node43168 = (inp[11]) ? 4'b0010 : node43169;
															assign node43169 = (inp[5]) ? node43171 : 4'b1010;
																assign node43171 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node43175 = (inp[0]) ? node43187 : node43176;
														assign node43176 = (inp[5]) ? node43182 : node43177;
															assign node43177 = (inp[6]) ? node43179 : 4'b1000;
																assign node43179 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node43182 = (inp[11]) ? 4'b1010 : node43183;
																assign node43183 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node43187 = (inp[11]) ? node43191 : node43188;
															assign node43188 = (inp[6]) ? 4'b1000 : 4'b0000;
															assign node43191 = (inp[6]) ? 4'b0000 : 4'b1000;
												assign node43194 = (inp[5]) ? node43208 : node43195;
													assign node43195 = (inp[0]) ? node43203 : node43196;
														assign node43196 = (inp[15]) ? node43198 : 4'b0010;
															assign node43198 = (inp[6]) ? 4'b0000 : node43199;
																assign node43199 = (inp[11]) ? 4'b1000 : 4'b0000;
														assign node43203 = (inp[6]) ? node43205 : 4'b0000;
															assign node43205 = (inp[11]) ? 4'b0000 : 4'b1000;
													assign node43208 = (inp[0]) ? node43220 : node43209;
														assign node43209 = (inp[15]) ? node43215 : node43210;
															assign node43210 = (inp[6]) ? node43212 : 4'b1000;
																assign node43212 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node43215 = (inp[6]) ? 4'b0010 : node43216;
																assign node43216 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node43220 = (inp[15]) ? 4'b0000 : node43221;
															assign node43221 = (inp[6]) ? node43223 : 4'b0010;
																assign node43223 = (inp[11]) ? 4'b0010 : 4'b1010;
											assign node43227 = (inp[6]) ? node43245 : node43228;
												assign node43228 = (inp[11]) ? node43240 : node43229;
													assign node43229 = (inp[5]) ? node43235 : node43230;
														assign node43230 = (inp[0]) ? 4'b0010 : node43231;
															assign node43231 = (inp[15]) ? 4'b0000 : 4'b0010;
														assign node43235 = (inp[15]) ? node43237 : 4'b0000;
															assign node43237 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node43240 = (inp[5]) ? 4'b1100 : node43241;
														assign node43241 = (inp[13]) ? 4'b1110 : 4'b1100;
												assign node43245 = (inp[11]) ? node43259 : node43246;
													assign node43246 = (inp[5]) ? node43254 : node43247;
														assign node43247 = (inp[13]) ? 4'b1100 : node43248;
															assign node43248 = (inp[15]) ? node43250 : 4'b1100;
																assign node43250 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node43254 = (inp[0]) ? node43256 : 4'b1110;
															assign node43256 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node43259 = (inp[5]) ? node43265 : node43260;
														assign node43260 = (inp[15]) ? node43262 : 4'b0110;
															assign node43262 = (inp[13]) ? 4'b0100 : 4'b0110;
														assign node43265 = (inp[13]) ? 4'b0110 : node43266;
															assign node43266 = (inp[0]) ? node43268 : 4'b0100;
																assign node43268 = (inp[15]) ? 4'b0100 : 4'b0110;
										assign node43272 = (inp[6]) ? node43294 : node43273;
											assign node43273 = (inp[11]) ? node43287 : node43274;
												assign node43274 = (inp[12]) ? node43280 : node43275;
													assign node43275 = (inp[5]) ? node43277 : 4'b0000;
														assign node43277 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node43280 = (inp[15]) ? node43284 : node43281;
														assign node43281 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node43284 = (inp[0]) ? 4'b0100 : 4'b0110;
												assign node43287 = (inp[15]) ? node43291 : node43288;
													assign node43288 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node43291 = (inp[0]) ? 4'b1100 : 4'b1110;
											assign node43294 = (inp[11]) ? node43322 : node43295;
												assign node43295 = (inp[5]) ? node43315 : node43296;
													assign node43296 = (inp[12]) ? node43310 : node43297;
														assign node43297 = (inp[13]) ? node43305 : node43298;
															assign node43298 = (inp[15]) ? node43302 : node43299;
																assign node43299 = (inp[0]) ? 4'b1110 : 4'b1100;
																assign node43302 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node43305 = (inp[0]) ? node43307 : 4'b1100;
																assign node43307 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node43310 = (inp[15]) ? node43312 : 4'b1100;
															assign node43312 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node43315 = (inp[13]) ? node43317 : 4'b1100;
														assign node43317 = (inp[0]) ? node43319 : 4'b1110;
															assign node43319 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node43322 = (inp[12]) ? node43330 : node43323;
													assign node43323 = (inp[15]) ? node43327 : node43324;
														assign node43324 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node43327 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node43330 = (inp[13]) ? node43336 : node43331;
														assign node43331 = (inp[5]) ? node43333 : 4'b0110;
															assign node43333 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node43336 = (inp[0]) ? node43340 : node43337;
															assign node43337 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node43340 = (inp[15]) ? 4'b0100 : 4'b0110;
								assign node43343 = (inp[4]) ? node43511 : node43344;
									assign node43344 = (inp[12]) ? node43438 : node43345;
										assign node43345 = (inp[10]) ? node43393 : node43346;
											assign node43346 = (inp[11]) ? node43370 : node43347;
												assign node43347 = (inp[6]) ? node43359 : node43348;
													assign node43348 = (inp[5]) ? 4'b0010 : node43349;
														assign node43349 = (inp[13]) ? node43353 : node43350;
															assign node43350 = (inp[15]) ? 4'b0010 : 4'b0000;
															assign node43353 = (inp[0]) ? 4'b0010 : node43354;
																assign node43354 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node43359 = (inp[0]) ? node43365 : node43360;
														assign node43360 = (inp[13]) ? node43362 : 4'b1000;
															assign node43362 = (inp[5]) ? 4'b1010 : 4'b1000;
														assign node43365 = (inp[5]) ? node43367 : 4'b1010;
															assign node43367 = (inp[13]) ? 4'b1010 : 4'b1000;
												assign node43370 = (inp[6]) ? node43380 : node43371;
													assign node43371 = (inp[15]) ? 4'b1000 : node43372;
														assign node43372 = (inp[13]) ? 4'b1000 : node43373;
															assign node43373 = (inp[5]) ? 4'b1010 : node43374;
																assign node43374 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node43380 = (inp[0]) ? node43386 : node43381;
														assign node43381 = (inp[5]) ? node43383 : 4'b0000;
															assign node43383 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node43386 = (inp[13]) ? node43390 : node43387;
															assign node43387 = (inp[15]) ? 4'b0000 : 4'b0010;
															assign node43390 = (inp[15]) ? 4'b0010 : 4'b0000;
											assign node43393 = (inp[11]) ? node43413 : node43394;
												assign node43394 = (inp[6]) ? node43410 : node43395;
													assign node43395 = (inp[5]) ? node43405 : node43396;
														assign node43396 = (inp[13]) ? node43398 : 4'b0010;
															assign node43398 = (inp[15]) ? node43402 : node43399;
																assign node43399 = (inp[0]) ? 4'b0000 : 4'b0010;
																assign node43402 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node43405 = (inp[13]) ? node43407 : 4'b0000;
															assign node43407 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node43410 = (inp[5]) ? 4'b1110 : 4'b1100;
												assign node43413 = (inp[6]) ? node43431 : node43414;
													assign node43414 = (inp[13]) ? node43424 : node43415;
														assign node43415 = (inp[5]) ? node43421 : node43416;
															assign node43416 = (inp[15]) ? node43418 : 4'b1110;
																assign node43418 = (inp[0]) ? 4'b1100 : 4'b1110;
															assign node43421 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node43424 = (inp[15]) ? node43428 : node43425;
															assign node43425 = (inp[0]) ? 4'b1110 : 4'b1100;
															assign node43428 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node43431 = (inp[5]) ? node43433 : 4'b0110;
														assign node43433 = (inp[0]) ? 4'b0100 : node43434;
															assign node43434 = (inp[15]) ? 4'b0110 : 4'b0100;
										assign node43438 = (inp[6]) ? node43484 : node43439;
											assign node43439 = (inp[11]) ? node43463 : node43440;
												assign node43440 = (inp[10]) ? node43450 : node43441;
													assign node43441 = (inp[15]) ? node43447 : node43442;
														assign node43442 = (inp[0]) ? 4'b0010 : node43443;
															assign node43443 = (inp[5]) ? 4'b0000 : 4'b0010;
														assign node43447 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node43450 = (inp[13]) ? node43458 : node43451;
														assign node43451 = (inp[5]) ? 4'b0100 : node43452;
															assign node43452 = (inp[15]) ? 4'b0110 : node43453;
																assign node43453 = (inp[0]) ? 4'b0110 : 4'b0100;
														assign node43458 = (inp[15]) ? 4'b0110 : node43459;
															assign node43459 = (inp[0]) ? 4'b0110 : 4'b0100;
												assign node43463 = (inp[13]) ? node43471 : node43464;
													assign node43464 = (inp[0]) ? node43468 : node43465;
														assign node43465 = (inp[15]) ? 4'b1110 : 4'b1100;
														assign node43468 = (inp[15]) ? 4'b1100 : 4'b1110;
													assign node43471 = (inp[10]) ? node43477 : node43472;
														assign node43472 = (inp[0]) ? node43474 : 4'b1110;
															assign node43474 = (inp[15]) ? 4'b1100 : 4'b1110;
														assign node43477 = (inp[0]) ? node43481 : node43478;
															assign node43478 = (inp[15]) ? 4'b1110 : 4'b1100;
															assign node43481 = (inp[15]) ? 4'b1100 : 4'b1110;
											assign node43484 = (inp[11]) ? node43492 : node43485;
												assign node43485 = (inp[15]) ? node43489 : node43486;
													assign node43486 = (inp[0]) ? 4'b1110 : 4'b1100;
													assign node43489 = (inp[0]) ? 4'b1100 : 4'b1110;
												assign node43492 = (inp[10]) ? node43498 : node43493;
													assign node43493 = (inp[15]) ? 4'b0110 : node43494;
														assign node43494 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node43498 = (inp[13]) ? node43504 : node43499;
														assign node43499 = (inp[15]) ? node43501 : 4'b0100;
															assign node43501 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node43504 = (inp[0]) ? node43508 : node43505;
															assign node43505 = (inp[15]) ? 4'b0110 : 4'b0100;
															assign node43508 = (inp[15]) ? 4'b0100 : 4'b0110;
									assign node43511 = (inp[12]) ? node43605 : node43512;
										assign node43512 = (inp[10]) ? node43558 : node43513;
											assign node43513 = (inp[15]) ? node43539 : node43514;
												assign node43514 = (inp[0]) ? node43522 : node43515;
													assign node43515 = (inp[6]) ? node43519 : node43516;
														assign node43516 = (inp[11]) ? 4'b1100 : 4'b0100;
														assign node43519 = (inp[11]) ? 4'b0100 : 4'b1100;
													assign node43522 = (inp[13]) ? node43532 : node43523;
														assign node43523 = (inp[5]) ? node43527 : node43524;
															assign node43524 = (inp[11]) ? 4'b0110 : 4'b1110;
															assign node43527 = (inp[11]) ? node43529 : 4'b0110;
																assign node43529 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node43532 = (inp[6]) ? node43536 : node43533;
															assign node43533 = (inp[11]) ? 4'b1110 : 4'b0110;
															assign node43536 = (inp[11]) ? 4'b0110 : 4'b1110;
												assign node43539 = (inp[0]) ? node43551 : node43540;
													assign node43540 = (inp[13]) ? node43544 : node43541;
														assign node43541 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node43544 = (inp[5]) ? 4'b1110 : node43545;
															assign node43545 = (inp[11]) ? 4'b1110 : node43546;
																assign node43546 = (inp[6]) ? 4'b1110 : 4'b0110;
													assign node43551 = (inp[11]) ? node43555 : node43552;
														assign node43552 = (inp[6]) ? 4'b1100 : 4'b0100;
														assign node43555 = (inp[6]) ? 4'b0100 : 4'b1100;
											assign node43558 = (inp[6]) ? node43582 : node43559;
												assign node43559 = (inp[11]) ? node43567 : node43560;
													assign node43560 = (inp[13]) ? 4'b0100 : node43561;
														assign node43561 = (inp[15]) ? 4'b0100 : node43562;
															assign node43562 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node43567 = (inp[13]) ? node43575 : node43568;
														assign node43568 = (inp[15]) ? node43572 : node43569;
															assign node43569 = (inp[5]) ? 4'b1000 : 4'b1010;
															assign node43572 = (inp[0]) ? 4'b1000 : 4'b1010;
														assign node43575 = (inp[5]) ? 4'b1000 : node43576;
															assign node43576 = (inp[0]) ? 4'b1000 : node43577;
																assign node43577 = (inp[15]) ? 4'b1010 : 4'b1000;
												assign node43582 = (inp[11]) ? node43596 : node43583;
													assign node43583 = (inp[5]) ? node43585 : 4'b1010;
														assign node43585 = (inp[13]) ? node43591 : node43586;
															assign node43586 = (inp[0]) ? 4'b1000 : node43587;
																assign node43587 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node43591 = (inp[15]) ? 4'b1010 : node43592;
																assign node43592 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node43596 = (inp[5]) ? 4'b0010 : node43597;
														assign node43597 = (inp[15]) ? node43601 : node43598;
															assign node43598 = (inp[13]) ? 4'b0010 : 4'b0000;
															assign node43601 = (inp[0]) ? 4'b0000 : 4'b0010;
										assign node43605 = (inp[6]) ? node43633 : node43606;
											assign node43606 = (inp[11]) ? node43622 : node43607;
												assign node43607 = (inp[10]) ? node43617 : node43608;
													assign node43608 = (inp[5]) ? node43610 : 4'b0110;
														assign node43610 = (inp[13]) ? 4'b0100 : node43611;
															assign node43611 = (inp[15]) ? 4'b0110 : node43612;
																assign node43612 = (inp[0]) ? 4'b0110 : 4'b0100;
													assign node43617 = (inp[13]) ? node43619 : 4'b0000;
														assign node43619 = (inp[5]) ? 4'b0010 : 4'b0000;
												assign node43622 = (inp[13]) ? node43628 : node43623;
													assign node43623 = (inp[15]) ? node43625 : 4'b1000;
														assign node43625 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node43628 = (inp[0]) ? 4'b1010 : node43629;
														assign node43629 = (inp[15]) ? 4'b1010 : 4'b1000;
											assign node43633 = (inp[11]) ? node43641 : node43634;
												assign node43634 = (inp[15]) ? node43638 : node43635;
													assign node43635 = (inp[0]) ? 4'b1010 : 4'b1000;
													assign node43638 = (inp[0]) ? 4'b1000 : 4'b1010;
												assign node43641 = (inp[10]) ? node43649 : node43642;
													assign node43642 = (inp[15]) ? node43646 : node43643;
														assign node43643 = (inp[0]) ? 4'b0010 : 4'b0000;
														assign node43646 = (inp[0]) ? 4'b0000 : 4'b0010;
													assign node43649 = (inp[13]) ? node43651 : 4'b0010;
														assign node43651 = (inp[15]) ? 4'b0000 : node43652;
															assign node43652 = (inp[0]) ? 4'b0010 : 4'b0000;
							assign node43656 = (inp[10]) ? node44018 : node43657;
								assign node43657 = (inp[15]) ? node43839 : node43658;
									assign node43658 = (inp[0]) ? node43752 : node43659;
										assign node43659 = (inp[5]) ? node43705 : node43660;
											assign node43660 = (inp[9]) ? node43686 : node43661;
												assign node43661 = (inp[4]) ? node43675 : node43662;
													assign node43662 = (inp[12]) ? node43668 : node43663;
														assign node43663 = (inp[6]) ? node43665 : 4'b0110;
															assign node43665 = (inp[11]) ? 4'b0110 : 4'b1110;
														assign node43668 = (inp[11]) ? node43672 : node43669;
															assign node43669 = (inp[6]) ? 4'b1010 : 4'b0110;
															assign node43672 = (inp[6]) ? 4'b0010 : 4'b1010;
													assign node43675 = (inp[12]) ? node43681 : node43676;
														assign node43676 = (inp[6]) ? node43678 : 4'b1010;
															assign node43678 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node43681 = (inp[6]) ? node43683 : 4'b0010;
															assign node43683 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node43686 = (inp[4]) ? node43696 : node43687;
													assign node43687 = (inp[11]) ? node43691 : node43688;
														assign node43688 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node43691 = (inp[12]) ? node43693 : 4'b0010;
															assign node43693 = (inp[6]) ? 4'b0100 : 4'b1100;
													assign node43696 = (inp[12]) ? node43698 : 4'b0100;
														assign node43698 = (inp[11]) ? node43702 : node43699;
															assign node43699 = (inp[6]) ? 4'b1000 : 4'b0100;
															assign node43702 = (inp[6]) ? 4'b0000 : 4'b1000;
											assign node43705 = (inp[6]) ? node43723 : node43706;
												assign node43706 = (inp[11]) ? node43714 : node43707;
													assign node43707 = (inp[9]) ? node43711 : node43708;
														assign node43708 = (inp[4]) ? 4'b0000 : 4'b0100;
														assign node43711 = (inp[4]) ? 4'b0100 : 4'b0000;
													assign node43714 = (inp[12]) ? node43716 : 4'b1000;
														assign node43716 = (inp[9]) ? node43720 : node43717;
															assign node43717 = (inp[4]) ? 4'b1100 : 4'b1000;
															assign node43720 = (inp[4]) ? 4'b1000 : 4'b1100;
												assign node43723 = (inp[11]) ? node43733 : node43724;
													assign node43724 = (inp[4]) ? node43726 : 4'b1100;
														assign node43726 = (inp[9]) ? node43730 : node43727;
															assign node43727 = (inp[12]) ? 4'b1100 : 4'b1000;
															assign node43730 = (inp[12]) ? 4'b1000 : 4'b1100;
													assign node43733 = (inp[9]) ? node43739 : node43734;
														assign node43734 = (inp[12]) ? node43736 : 4'b0100;
															assign node43736 = (inp[4]) ? 4'b0100 : 4'b0000;
														assign node43739 = (inp[13]) ? node43747 : node43740;
															assign node43740 = (inp[12]) ? node43744 : node43741;
																assign node43741 = (inp[4]) ? 4'b0100 : 4'b0000;
																assign node43744 = (inp[4]) ? 4'b0000 : 4'b0100;
															assign node43747 = (inp[4]) ? 4'b0100 : node43748;
																assign node43748 = (inp[12]) ? 4'b0100 : 4'b0000;
										assign node43752 = (inp[5]) ? node43796 : node43753;
											assign node43753 = (inp[9]) ? node43781 : node43754;
												assign node43754 = (inp[13]) ? node43766 : node43755;
													assign node43755 = (inp[4]) ? node43759 : node43756;
														assign node43756 = (inp[12]) ? 4'b1000 : 4'b0100;
														assign node43759 = (inp[12]) ? 4'b0000 : node43760;
															assign node43760 = (inp[11]) ? node43762 : 4'b1000;
																assign node43762 = (inp[6]) ? 4'b0000 : 4'b1000;
													assign node43766 = (inp[12]) ? node43776 : node43767;
														assign node43767 = (inp[4]) ? node43773 : node43768;
															assign node43768 = (inp[11]) ? node43770 : 4'b0100;
																assign node43770 = (inp[6]) ? 4'b0100 : 4'b1100;
															assign node43773 = (inp[6]) ? 4'b0000 : 4'b1000;
														assign node43776 = (inp[4]) ? node43778 : 4'b0100;
															assign node43778 = (inp[11]) ? 4'b0110 : 4'b1110;
												assign node43781 = (inp[11]) ? node43783 : 4'b0110;
													assign node43783 = (inp[6]) ? node43791 : node43784;
														assign node43784 = (inp[13]) ? node43786 : 4'b1110;
															assign node43786 = (inp[4]) ? node43788 : 4'b1000;
																assign node43788 = (inp[12]) ? 4'b1010 : 4'b1110;
														assign node43791 = (inp[12]) ? node43793 : 4'b0000;
															assign node43793 = (inp[4]) ? 4'b0010 : 4'b0110;
											assign node43796 = (inp[4]) ? node43816 : node43797;
												assign node43797 = (inp[9]) ? node43805 : node43798;
													assign node43798 = (inp[11]) ? node43800 : 4'b0110;
														assign node43800 = (inp[12]) ? node43802 : 4'b0110;
															assign node43802 = (inp[13]) ? 4'b1010 : 4'b0010;
													assign node43805 = (inp[12]) ? node43813 : node43806;
														assign node43806 = (inp[13]) ? node43808 : 4'b0010;
															assign node43808 = (inp[6]) ? 4'b1010 : node43809;
																assign node43809 = (inp[11]) ? 4'b1010 : 4'b0010;
														assign node43813 = (inp[11]) ? 4'b0110 : 4'b0010;
												assign node43816 = (inp[13]) ? node43828 : node43817;
													assign node43817 = (inp[6]) ? node43825 : node43818;
														assign node43818 = (inp[11]) ? node43820 : 4'b0010;
															assign node43820 = (inp[12]) ? node43822 : 4'b1010;
																assign node43822 = (inp[9]) ? 4'b1010 : 4'b1110;
														assign node43825 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node43828 = (inp[9]) ? node43834 : node43829;
														assign node43829 = (inp[11]) ? 4'b0010 : node43830;
															assign node43830 = (inp[6]) ? 4'b1010 : 4'b0010;
														assign node43834 = (inp[6]) ? node43836 : 4'b0110;
															assign node43836 = (inp[11]) ? 4'b0110 : 4'b1110;
									assign node43839 = (inp[0]) ? node43935 : node43840;
										assign node43840 = (inp[5]) ? node43888 : node43841;
											assign node43841 = (inp[9]) ? node43861 : node43842;
												assign node43842 = (inp[13]) ? node43850 : node43843;
													assign node43843 = (inp[4]) ? node43847 : node43844;
														assign node43844 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node43847 = (inp[6]) ? 4'b0110 : 4'b1110;
													assign node43850 = (inp[4]) ? node43852 : 4'b0100;
														assign node43852 = (inp[12]) ? node43858 : node43853;
															assign node43853 = (inp[6]) ? node43855 : 4'b1000;
																assign node43855 = (inp[11]) ? 4'b0000 : 4'b1000;
															assign node43858 = (inp[11]) ? 4'b0110 : 4'b0000;
												assign node43861 = (inp[4]) ? node43877 : node43862;
													assign node43862 = (inp[12]) ? node43868 : node43863;
														assign node43863 = (inp[6]) ? node43865 : 4'b0000;
															assign node43865 = (inp[11]) ? 4'b0000 : 4'b1000;
														assign node43868 = (inp[13]) ? node43874 : node43869;
															assign node43869 = (inp[11]) ? node43871 : 4'b1110;
																assign node43871 = (inp[6]) ? 4'b0110 : 4'b1110;
															assign node43874 = (inp[6]) ? 4'b0110 : 4'b0000;
													assign node43877 = (inp[12]) ? node43881 : node43878;
														assign node43878 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node43881 = (inp[11]) ? node43885 : node43882;
															assign node43882 = (inp[6]) ? 4'b1010 : 4'b0110;
															assign node43885 = (inp[6]) ? 4'b0010 : 4'b1010;
											assign node43888 = (inp[11]) ? node43908 : node43889;
												assign node43889 = (inp[6]) ? node43897 : node43890;
													assign node43890 = (inp[4]) ? node43894 : node43891;
														assign node43891 = (inp[9]) ? 4'b0010 : 4'b0110;
														assign node43894 = (inp[9]) ? 4'b0110 : 4'b0010;
													assign node43897 = (inp[12]) ? node43903 : node43898;
														assign node43898 = (inp[4]) ? node43900 : 4'b1010;
															assign node43900 = (inp[9]) ? 4'b1110 : 4'b1010;
														assign node43903 = (inp[9]) ? node43905 : 4'b1110;
															assign node43905 = (inp[4]) ? 4'b1010 : 4'b1110;
												assign node43908 = (inp[6]) ? node43918 : node43909;
													assign node43909 = (inp[12]) ? 4'b1110 : node43910;
														assign node43910 = (inp[4]) ? node43914 : node43911;
															assign node43911 = (inp[9]) ? 4'b1010 : 4'b1110;
															assign node43914 = (inp[9]) ? 4'b1110 : 4'b1010;
													assign node43918 = (inp[9]) ? node43926 : node43919;
														assign node43919 = (inp[12]) ? node43923 : node43920;
															assign node43920 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node43923 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node43926 = (inp[13]) ? node43928 : 4'b0110;
															assign node43928 = (inp[12]) ? node43932 : node43929;
																assign node43929 = (inp[4]) ? 4'b0110 : 4'b0010;
																assign node43932 = (inp[4]) ? 4'b0010 : 4'b0110;
										assign node43935 = (inp[5]) ? node43985 : node43936;
											assign node43936 = (inp[4]) ? node43966 : node43937;
												assign node43937 = (inp[9]) ? node43953 : node43938;
													assign node43938 = (inp[12]) ? node43946 : node43939;
														assign node43939 = (inp[11]) ? node43943 : node43940;
															assign node43940 = (inp[6]) ? 4'b1110 : 4'b0110;
															assign node43943 = (inp[6]) ? 4'b0110 : 4'b1110;
														assign node43946 = (inp[6]) ? node43950 : node43947;
															assign node43947 = (inp[11]) ? 4'b1010 : 4'b0110;
															assign node43950 = (inp[11]) ? 4'b0010 : 4'b1010;
													assign node43953 = (inp[12]) ? node43961 : node43954;
														assign node43954 = (inp[13]) ? node43956 : 4'b1010;
															assign node43956 = (inp[6]) ? node43958 : 4'b0010;
																assign node43958 = (inp[11]) ? 4'b0010 : 4'b1010;
														assign node43961 = (inp[6]) ? node43963 : 4'b0010;
															assign node43963 = (inp[11]) ? 4'b0100 : 4'b1100;
												assign node43966 = (inp[9]) ? node43974 : node43967;
													assign node43967 = (inp[12]) ? node43969 : 4'b1010;
														assign node43969 = (inp[6]) ? node43971 : 4'b1100;
															assign node43971 = (inp[13]) ? 4'b1100 : 4'b0100;
													assign node43974 = (inp[12]) ? node43980 : node43975;
														assign node43975 = (inp[6]) ? node43977 : 4'b0100;
															assign node43977 = (inp[11]) ? 4'b0100 : 4'b1100;
														assign node43980 = (inp[13]) ? node43982 : 4'b1000;
															assign node43982 = (inp[11]) ? 4'b0000 : 4'b0100;
											assign node43985 = (inp[13]) ? node43993 : node43986;
												assign node43986 = (inp[9]) ? node43990 : node43987;
													assign node43987 = (inp[11]) ? 4'b1100 : 4'b0100;
													assign node43990 = (inp[4]) ? 4'b0100 : 4'b1100;
												assign node43993 = (inp[11]) ? node44005 : node43994;
													assign node43994 = (inp[6]) ? node44000 : node43995;
														assign node43995 = (inp[4]) ? 4'b0100 : node43996;
															assign node43996 = (inp[9]) ? 4'b0000 : 4'b0100;
														assign node44000 = (inp[4]) ? node44002 : 4'b1100;
															assign node44002 = (inp[9]) ? 4'b1000 : 4'b1100;
													assign node44005 = (inp[6]) ? node44013 : node44006;
														assign node44006 = (inp[9]) ? 4'b1100 : node44007;
															assign node44007 = (inp[4]) ? 4'b1000 : node44008;
																assign node44008 = (inp[12]) ? 4'b1000 : 4'b1100;
														assign node44013 = (inp[12]) ? node44015 : 4'b0000;
															assign node44015 = (inp[4]) ? 4'b0100 : 4'b0000;
								assign node44018 = (inp[5]) ? node44164 : node44019;
									assign node44019 = (inp[11]) ? node44105 : node44020;
										assign node44020 = (inp[6]) ? node44078 : node44021;
											assign node44021 = (inp[15]) ? node44049 : node44022;
												assign node44022 = (inp[4]) ? node44038 : node44023;
													assign node44023 = (inp[0]) ? node44031 : node44024;
														assign node44024 = (inp[9]) ? node44028 : node44025;
															assign node44025 = (inp[12]) ? 4'b0010 : 4'b0110;
															assign node44028 = (inp[12]) ? 4'b0100 : 4'b0010;
														assign node44031 = (inp[12]) ? node44035 : node44032;
															assign node44032 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node44035 = (inp[9]) ? 4'b0110 : 4'b0000;
													assign node44038 = (inp[0]) ? node44044 : node44039;
														assign node44039 = (inp[12]) ? 4'b0100 : node44040;
															assign node44040 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node44044 = (inp[12]) ? node44046 : 4'b0110;
															assign node44046 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node44049 = (inp[13]) ? node44065 : node44050;
													assign node44050 = (inp[4]) ? node44058 : node44051;
														assign node44051 = (inp[9]) ? node44055 : node44052;
															assign node44052 = (inp[0]) ? 4'b0110 : 4'b0100;
															assign node44055 = (inp[0]) ? 4'b0100 : 4'b0110;
														assign node44058 = (inp[12]) ? node44062 : node44059;
															assign node44059 = (inp[9]) ? 4'b0100 : 4'b0000;
															assign node44062 = (inp[0]) ? 4'b0100 : 4'b0110;
													assign node44065 = (inp[12]) ? 4'b0000 : node44066;
														assign node44066 = (inp[4]) ? node44070 : node44067;
															assign node44067 = (inp[9]) ? 4'b0000 : 4'b0100;
															assign node44070 = (inp[9]) ? node44074 : node44071;
																assign node44071 = (inp[0]) ? 4'b0010 : 4'b0000;
																assign node44074 = (inp[0]) ? 4'b0100 : 4'b0110;
											assign node44078 = (inp[4]) ? node44094 : node44079;
												assign node44079 = (inp[9]) ? node44089 : node44080;
													assign node44080 = (inp[12]) ? node44086 : node44081;
														assign node44081 = (inp[15]) ? node44083 : 4'b1010;
															assign node44083 = (inp[13]) ? 4'b1010 : 4'b1000;
														assign node44086 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node44089 = (inp[0]) ? 4'b1110 : node44090;
														assign node44090 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node44094 = (inp[9]) ? node44102 : node44095;
													assign node44095 = (inp[15]) ? node44099 : node44096;
														assign node44096 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node44099 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node44102 = (inp[15]) ? 4'b1000 : 4'b1010;
										assign node44105 = (inp[6]) ? node44135 : node44106;
											assign node44106 = (inp[4]) ? node44118 : node44107;
												assign node44107 = (inp[9]) ? node44113 : node44108;
													assign node44108 = (inp[0]) ? 4'b1000 : node44109;
														assign node44109 = (inp[15]) ? 4'b1000 : 4'b1010;
													assign node44113 = (inp[12]) ? 4'b1100 : node44114;
														assign node44114 = (inp[15]) ? 4'b1110 : 4'b1100;
												assign node44118 = (inp[9]) ? node44126 : node44119;
													assign node44119 = (inp[15]) ? node44123 : node44120;
														assign node44120 = (inp[0]) ? 4'b1110 : 4'b1100;
														assign node44123 = (inp[0]) ? 4'b1100 : 4'b1110;
													assign node44126 = (inp[12]) ? 4'b1010 : node44127;
														assign node44127 = (inp[0]) ? node44131 : node44128;
															assign node44128 = (inp[15]) ? 4'b1010 : 4'b1000;
															assign node44131 = (inp[15]) ? 4'b1000 : 4'b1010;
											assign node44135 = (inp[15]) ? node44149 : node44136;
												assign node44136 = (inp[0]) ? node44144 : node44137;
													assign node44137 = (inp[4]) ? node44141 : node44138;
														assign node44138 = (inp[9]) ? 4'b0100 : 4'b0010;
														assign node44141 = (inp[9]) ? 4'b0000 : 4'b0100;
													assign node44144 = (inp[4]) ? node44146 : 4'b0000;
														assign node44146 = (inp[13]) ? 4'b0010 : 4'b0110;
												assign node44149 = (inp[0]) ? node44157 : node44150;
													assign node44150 = (inp[9]) ? node44154 : node44151;
														assign node44151 = (inp[4]) ? 4'b0110 : 4'b0000;
														assign node44154 = (inp[4]) ? 4'b0010 : 4'b0110;
													assign node44157 = (inp[12]) ? 4'b0010 : node44158;
														assign node44158 = (inp[13]) ? node44160 : 4'b0100;
															assign node44160 = (inp[4]) ? 4'b0000 : 4'b0100;
									assign node44164 = (inp[11]) ? node44262 : node44165;
										assign node44165 = (inp[6]) ? node44223 : node44166;
											assign node44166 = (inp[0]) ? node44188 : node44167;
												assign node44167 = (inp[15]) ? node44173 : node44168;
													assign node44168 = (inp[9]) ? node44170 : 4'b0100;
														assign node44170 = (inp[4]) ? 4'b0000 : 4'b0100;
													assign node44173 = (inp[12]) ? node44181 : node44174;
														assign node44174 = (inp[9]) ? node44178 : node44175;
															assign node44175 = (inp[4]) ? 4'b0010 : 4'b0110;
															assign node44178 = (inp[4]) ? 4'b0110 : 4'b0010;
														assign node44181 = (inp[4]) ? node44185 : node44182;
															assign node44182 = (inp[9]) ? 4'b0110 : 4'b0010;
															assign node44185 = (inp[9]) ? 4'b0010 : 4'b0110;
												assign node44188 = (inp[15]) ? node44202 : node44189;
													assign node44189 = (inp[13]) ? node44195 : node44190;
														assign node44190 = (inp[9]) ? 4'b0010 : node44191;
															assign node44191 = (inp[12]) ? 4'b0010 : 4'b0110;
														assign node44195 = (inp[12]) ? node44197 : 4'b0010;
															assign node44197 = (inp[9]) ? 4'b0110 : node44198;
																assign node44198 = (inp[4]) ? 4'b0110 : 4'b0010;
													assign node44202 = (inp[9]) ? node44216 : node44203;
														assign node44203 = (inp[13]) ? node44209 : node44204;
															assign node44204 = (inp[4]) ? node44206 : 4'b0000;
																assign node44206 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node44209 = (inp[4]) ? node44213 : node44210;
																assign node44210 = (inp[12]) ? 4'b0000 : 4'b0100;
																assign node44213 = (inp[12]) ? 4'b0100 : 4'b0000;
														assign node44216 = (inp[4]) ? node44220 : node44217;
															assign node44217 = (inp[12]) ? 4'b0100 : 4'b0000;
															assign node44220 = (inp[12]) ? 4'b0000 : 4'b0100;
											assign node44223 = (inp[4]) ? node44235 : node44224;
												assign node44224 = (inp[9]) ? node44232 : node44225;
													assign node44225 = (inp[15]) ? node44229 : node44226;
														assign node44226 = (inp[0]) ? 4'b1010 : 4'b1000;
														assign node44229 = (inp[0]) ? 4'b1000 : 4'b1010;
													assign node44232 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node44235 = (inp[9]) ? node44249 : node44236;
													assign node44236 = (inp[13]) ? node44242 : node44237;
														assign node44237 = (inp[15]) ? node44239 : 4'b1100;
															assign node44239 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node44242 = (inp[12]) ? 4'b1110 : node44243;
															assign node44243 = (inp[0]) ? 4'b1100 : node44244;
																assign node44244 = (inp[15]) ? 4'b1110 : 4'b1100;
													assign node44249 = (inp[13]) ? node44257 : node44250;
														assign node44250 = (inp[12]) ? node44252 : 4'b1010;
															assign node44252 = (inp[0]) ? node44254 : 4'b1000;
																assign node44254 = (inp[15]) ? 4'b1000 : 4'b1010;
														assign node44257 = (inp[0]) ? 4'b1000 : node44258;
															assign node44258 = (inp[15]) ? 4'b1010 : 4'b1000;
										assign node44262 = (inp[6]) ? node44304 : node44263;
											assign node44263 = (inp[13]) ? node44285 : node44264;
												assign node44264 = (inp[12]) ? node44276 : node44265;
													assign node44265 = (inp[4]) ? node44273 : node44266;
														assign node44266 = (inp[9]) ? node44268 : 4'b1010;
															assign node44268 = (inp[15]) ? node44270 : 4'b1110;
																assign node44270 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node44273 = (inp[9]) ? 4'b1010 : 4'b1100;
													assign node44276 = (inp[9]) ? node44282 : node44277;
														assign node44277 = (inp[4]) ? node44279 : 4'b1000;
															assign node44279 = (inp[0]) ? 4'b1100 : 4'b1110;
														assign node44282 = (inp[15]) ? 4'b1100 : 4'b1110;
												assign node44285 = (inp[15]) ? node44299 : node44286;
													assign node44286 = (inp[0]) ? node44292 : node44287;
														assign node44287 = (inp[9]) ? node44289 : 4'b1100;
															assign node44289 = (inp[12]) ? 4'b1100 : 4'b1000;
														assign node44292 = (inp[9]) ? node44296 : node44293;
															assign node44293 = (inp[4]) ? 4'b1110 : 4'b1010;
															assign node44296 = (inp[4]) ? 4'b1010 : 4'b1110;
													assign node44299 = (inp[4]) ? 4'b1010 : node44300;
														assign node44300 = (inp[9]) ? 4'b1110 : 4'b1010;
											assign node44304 = (inp[9]) ? node44326 : node44305;
												assign node44305 = (inp[4]) ? node44319 : node44306;
													assign node44306 = (inp[13]) ? node44314 : node44307;
														assign node44307 = (inp[15]) ? node44311 : node44308;
															assign node44308 = (inp[0]) ? 4'b0010 : 4'b0000;
															assign node44311 = (inp[0]) ? 4'b0000 : 4'b0010;
														assign node44314 = (inp[0]) ? node44316 : 4'b0000;
															assign node44316 = (inp[15]) ? 4'b0000 : 4'b0010;
													assign node44319 = (inp[0]) ? node44323 : node44320;
														assign node44320 = (inp[12]) ? 4'b0110 : 4'b0100;
														assign node44323 = (inp[12]) ? 4'b0100 : 4'b0110;
												assign node44326 = (inp[4]) ? node44334 : node44327;
													assign node44327 = (inp[0]) ? node44331 : node44328;
														assign node44328 = (inp[15]) ? 4'b0110 : 4'b0100;
														assign node44331 = (inp[15]) ? 4'b0100 : 4'b0110;
													assign node44334 = (inp[0]) ? node44338 : node44335;
														assign node44335 = (inp[15]) ? 4'b0010 : 4'b0000;
														assign node44338 = (inp[15]) ? 4'b0000 : 4'b0010;

endmodule