module dtc_split5_bm27 (
	input  wire [16-1:0] inp,
	output wire [16-1:0] outp
);

	wire [16-1:0] node1;
	wire [16-1:0] node2;
	wire [16-1:0] node3;
	wire [16-1:0] node4;
	wire [16-1:0] node5;
	wire [16-1:0] node6;
	wire [16-1:0] node7;
	wire [16-1:0] node8;
	wire [16-1:0] node9;
	wire [16-1:0] node10;
	wire [16-1:0] node11;
	wire [16-1:0] node12;
	wire [16-1:0] node13;
	wire [16-1:0] node16;
	wire [16-1:0] node19;
	wire [16-1:0] node20;
	wire [16-1:0] node23;
	wire [16-1:0] node26;
	wire [16-1:0] node27;
	wire [16-1:0] node28;
	wire [16-1:0] node31;
	wire [16-1:0] node34;
	wire [16-1:0] node35;
	wire [16-1:0] node38;
	wire [16-1:0] node41;
	wire [16-1:0] node42;
	wire [16-1:0] node43;
	wire [16-1:0] node44;
	wire [16-1:0] node47;
	wire [16-1:0] node50;
	wire [16-1:0] node51;
	wire [16-1:0] node54;
	wire [16-1:0] node57;
	wire [16-1:0] node58;
	wire [16-1:0] node59;
	wire [16-1:0] node62;
	wire [16-1:0] node65;
	wire [16-1:0] node66;
	wire [16-1:0] node69;
	wire [16-1:0] node72;
	wire [16-1:0] node73;
	wire [16-1:0] node74;
	wire [16-1:0] node75;
	wire [16-1:0] node76;
	wire [16-1:0] node80;
	wire [16-1:0] node81;
	wire [16-1:0] node84;
	wire [16-1:0] node87;
	wire [16-1:0] node88;
	wire [16-1:0] node89;
	wire [16-1:0] node92;
	wire [16-1:0] node95;
	wire [16-1:0] node96;
	wire [16-1:0] node99;
	wire [16-1:0] node102;
	wire [16-1:0] node103;
	wire [16-1:0] node104;
	wire [16-1:0] node105;
	wire [16-1:0] node108;
	wire [16-1:0] node111;
	wire [16-1:0] node112;
	wire [16-1:0] node115;
	wire [16-1:0] node118;
	wire [16-1:0] node119;
	wire [16-1:0] node120;
	wire [16-1:0] node123;
	wire [16-1:0] node126;
	wire [16-1:0] node127;
	wire [16-1:0] node130;
	wire [16-1:0] node133;
	wire [16-1:0] node134;
	wire [16-1:0] node135;
	wire [16-1:0] node136;
	wire [16-1:0] node137;
	wire [16-1:0] node138;
	wire [16-1:0] node141;
	wire [16-1:0] node144;
	wire [16-1:0] node145;
	wire [16-1:0] node148;
	wire [16-1:0] node151;
	wire [16-1:0] node152;
	wire [16-1:0] node153;
	wire [16-1:0] node156;
	wire [16-1:0] node159;
	wire [16-1:0] node160;
	wire [16-1:0] node163;
	wire [16-1:0] node166;
	wire [16-1:0] node167;
	wire [16-1:0] node168;
	wire [16-1:0] node169;
	wire [16-1:0] node172;
	wire [16-1:0] node175;
	wire [16-1:0] node176;
	wire [16-1:0] node179;
	wire [16-1:0] node182;
	wire [16-1:0] node183;
	wire [16-1:0] node185;
	wire [16-1:0] node188;
	wire [16-1:0] node189;
	wire [16-1:0] node192;
	wire [16-1:0] node195;
	wire [16-1:0] node196;
	wire [16-1:0] node197;
	wire [16-1:0] node198;
	wire [16-1:0] node199;
	wire [16-1:0] node202;
	wire [16-1:0] node205;
	wire [16-1:0] node206;
	wire [16-1:0] node209;
	wire [16-1:0] node212;
	wire [16-1:0] node213;
	wire [16-1:0] node214;
	wire [16-1:0] node217;
	wire [16-1:0] node220;
	wire [16-1:0] node221;
	wire [16-1:0] node224;
	wire [16-1:0] node227;
	wire [16-1:0] node228;
	wire [16-1:0] node229;
	wire [16-1:0] node230;
	wire [16-1:0] node233;
	wire [16-1:0] node236;
	wire [16-1:0] node237;
	wire [16-1:0] node240;
	wire [16-1:0] node243;
	wire [16-1:0] node244;
	wire [16-1:0] node246;
	wire [16-1:0] node249;
	wire [16-1:0] node250;
	wire [16-1:0] node253;
	wire [16-1:0] node256;
	wire [16-1:0] node257;
	wire [16-1:0] node258;
	wire [16-1:0] node259;
	wire [16-1:0] node260;
	wire [16-1:0] node261;
	wire [16-1:0] node262;
	wire [16-1:0] node265;
	wire [16-1:0] node268;
	wire [16-1:0] node269;
	wire [16-1:0] node272;
	wire [16-1:0] node275;
	wire [16-1:0] node276;
	wire [16-1:0] node277;
	wire [16-1:0] node280;
	wire [16-1:0] node283;
	wire [16-1:0] node285;
	wire [16-1:0] node288;
	wire [16-1:0] node289;
	wire [16-1:0] node290;
	wire [16-1:0] node291;
	wire [16-1:0] node294;
	wire [16-1:0] node297;
	wire [16-1:0] node298;
	wire [16-1:0] node302;
	wire [16-1:0] node303;
	wire [16-1:0] node305;
	wire [16-1:0] node308;
	wire [16-1:0] node309;
	wire [16-1:0] node313;
	wire [16-1:0] node314;
	wire [16-1:0] node315;
	wire [16-1:0] node316;
	wire [16-1:0] node317;
	wire [16-1:0] node320;
	wire [16-1:0] node323;
	wire [16-1:0] node324;
	wire [16-1:0] node327;
	wire [16-1:0] node330;
	wire [16-1:0] node331;
	wire [16-1:0] node333;
	wire [16-1:0] node336;
	wire [16-1:0] node338;
	wire [16-1:0] node341;
	wire [16-1:0] node342;
	wire [16-1:0] node343;
	wire [16-1:0] node344;
	wire [16-1:0] node347;
	wire [16-1:0] node350;
	wire [16-1:0] node351;
	wire [16-1:0] node354;
	wire [16-1:0] node357;
	wire [16-1:0] node358;
	wire [16-1:0] node359;
	wire [16-1:0] node362;
	wire [16-1:0] node365;
	wire [16-1:0] node366;
	wire [16-1:0] node369;
	wire [16-1:0] node372;
	wire [16-1:0] node373;
	wire [16-1:0] node374;
	wire [16-1:0] node375;
	wire [16-1:0] node376;
	wire [16-1:0] node377;
	wire [16-1:0] node381;
	wire [16-1:0] node382;
	wire [16-1:0] node385;
	wire [16-1:0] node388;
	wire [16-1:0] node389;
	wire [16-1:0] node390;
	wire [16-1:0] node393;
	wire [16-1:0] node396;
	wire [16-1:0] node397;
	wire [16-1:0] node401;
	wire [16-1:0] node402;
	wire [16-1:0] node403;
	wire [16-1:0] node406;
	wire [16-1:0] node407;
	wire [16-1:0] node411;
	wire [16-1:0] node412;
	wire [16-1:0] node413;
	wire [16-1:0] node416;
	wire [16-1:0] node419;
	wire [16-1:0] node420;
	wire [16-1:0] node423;
	wire [16-1:0] node426;
	wire [16-1:0] node427;
	wire [16-1:0] node428;
	wire [16-1:0] node429;
	wire [16-1:0] node430;
	wire [16-1:0] node433;
	wire [16-1:0] node436;
	wire [16-1:0] node437;
	wire [16-1:0] node440;
	wire [16-1:0] node443;
	wire [16-1:0] node444;
	wire [16-1:0] node445;
	wire [16-1:0] node448;
	wire [16-1:0] node451;
	wire [16-1:0] node452;
	wire [16-1:0] node455;
	wire [16-1:0] node458;
	wire [16-1:0] node459;
	wire [16-1:0] node461;
	wire [16-1:0] node462;
	wire [16-1:0] node465;
	wire [16-1:0] node468;
	wire [16-1:0] node469;
	wire [16-1:0] node471;
	wire [16-1:0] node474;
	wire [16-1:0] node475;
	wire [16-1:0] node478;
	wire [16-1:0] node481;
	wire [16-1:0] node482;
	wire [16-1:0] node483;
	wire [16-1:0] node484;
	wire [16-1:0] node485;
	wire [16-1:0] node486;
	wire [16-1:0] node487;
	wire [16-1:0] node488;
	wire [16-1:0] node491;
	wire [16-1:0] node494;
	wire [16-1:0] node495;
	wire [16-1:0] node499;
	wire [16-1:0] node500;
	wire [16-1:0] node501;
	wire [16-1:0] node504;
	wire [16-1:0] node507;
	wire [16-1:0] node508;
	wire [16-1:0] node511;
	wire [16-1:0] node514;
	wire [16-1:0] node515;
	wire [16-1:0] node516;
	wire [16-1:0] node517;
	wire [16-1:0] node521;
	wire [16-1:0] node522;
	wire [16-1:0] node526;
	wire [16-1:0] node527;
	wire [16-1:0] node528;
	wire [16-1:0] node531;
	wire [16-1:0] node534;
	wire [16-1:0] node535;
	wire [16-1:0] node539;
	wire [16-1:0] node540;
	wire [16-1:0] node541;
	wire [16-1:0] node542;
	wire [16-1:0] node543;
	wire [16-1:0] node546;
	wire [16-1:0] node549;
	wire [16-1:0] node550;
	wire [16-1:0] node553;
	wire [16-1:0] node556;
	wire [16-1:0] node557;
	wire [16-1:0] node558;
	wire [16-1:0] node561;
	wire [16-1:0] node564;
	wire [16-1:0] node565;
	wire [16-1:0] node568;
	wire [16-1:0] node571;
	wire [16-1:0] node572;
	wire [16-1:0] node573;
	wire [16-1:0] node574;
	wire [16-1:0] node577;
	wire [16-1:0] node580;
	wire [16-1:0] node581;
	wire [16-1:0] node585;
	wire [16-1:0] node586;
	wire [16-1:0] node587;
	wire [16-1:0] node590;
	wire [16-1:0] node593;
	wire [16-1:0] node594;
	wire [16-1:0] node597;
	wire [16-1:0] node600;
	wire [16-1:0] node601;
	wire [16-1:0] node602;
	wire [16-1:0] node603;
	wire [16-1:0] node604;
	wire [16-1:0] node605;
	wire [16-1:0] node608;
	wire [16-1:0] node611;
	wire [16-1:0] node612;
	wire [16-1:0] node615;
	wire [16-1:0] node618;
	wire [16-1:0] node619;
	wire [16-1:0] node620;
	wire [16-1:0] node623;
	wire [16-1:0] node626;
	wire [16-1:0] node627;
	wire [16-1:0] node630;
	wire [16-1:0] node633;
	wire [16-1:0] node634;
	wire [16-1:0] node635;
	wire [16-1:0] node636;
	wire [16-1:0] node639;
	wire [16-1:0] node642;
	wire [16-1:0] node643;
	wire [16-1:0] node646;
	wire [16-1:0] node649;
	wire [16-1:0] node650;
	wire [16-1:0] node651;
	wire [16-1:0] node654;
	wire [16-1:0] node657;
	wire [16-1:0] node658;
	wire [16-1:0] node661;
	wire [16-1:0] node664;
	wire [16-1:0] node665;
	wire [16-1:0] node666;
	wire [16-1:0] node667;
	wire [16-1:0] node668;
	wire [16-1:0] node671;
	wire [16-1:0] node674;
	wire [16-1:0] node675;
	wire [16-1:0] node678;
	wire [16-1:0] node681;
	wire [16-1:0] node682;
	wire [16-1:0] node683;
	wire [16-1:0] node686;
	wire [16-1:0] node689;
	wire [16-1:0] node690;
	wire [16-1:0] node693;
	wire [16-1:0] node696;
	wire [16-1:0] node697;
	wire [16-1:0] node698;
	wire [16-1:0] node699;
	wire [16-1:0] node702;
	wire [16-1:0] node705;
	wire [16-1:0] node706;
	wire [16-1:0] node709;
	wire [16-1:0] node712;
	wire [16-1:0] node713;
	wire [16-1:0] node714;
	wire [16-1:0] node717;
	wire [16-1:0] node720;
	wire [16-1:0] node721;
	wire [16-1:0] node724;
	wire [16-1:0] node727;
	wire [16-1:0] node728;
	wire [16-1:0] node729;
	wire [16-1:0] node730;
	wire [16-1:0] node731;
	wire [16-1:0] node732;
	wire [16-1:0] node733;
	wire [16-1:0] node736;
	wire [16-1:0] node739;
	wire [16-1:0] node740;
	wire [16-1:0] node743;
	wire [16-1:0] node746;
	wire [16-1:0] node747;
	wire [16-1:0] node748;
	wire [16-1:0] node751;
	wire [16-1:0] node754;
	wire [16-1:0] node755;
	wire [16-1:0] node758;
	wire [16-1:0] node761;
	wire [16-1:0] node762;
	wire [16-1:0] node763;
	wire [16-1:0] node764;
	wire [16-1:0] node767;
	wire [16-1:0] node770;
	wire [16-1:0] node771;
	wire [16-1:0] node774;
	wire [16-1:0] node777;
	wire [16-1:0] node778;
	wire [16-1:0] node779;
	wire [16-1:0] node782;
	wire [16-1:0] node785;
	wire [16-1:0] node787;
	wire [16-1:0] node790;
	wire [16-1:0] node791;
	wire [16-1:0] node792;
	wire [16-1:0] node793;
	wire [16-1:0] node794;
	wire [16-1:0] node797;
	wire [16-1:0] node800;
	wire [16-1:0] node801;
	wire [16-1:0] node805;
	wire [16-1:0] node806;
	wire [16-1:0] node807;
	wire [16-1:0] node810;
	wire [16-1:0] node813;
	wire [16-1:0] node814;
	wire [16-1:0] node817;
	wire [16-1:0] node820;
	wire [16-1:0] node821;
	wire [16-1:0] node822;
	wire [16-1:0] node823;
	wire [16-1:0] node827;
	wire [16-1:0] node828;
	wire [16-1:0] node831;
	wire [16-1:0] node834;
	wire [16-1:0] node835;
	wire [16-1:0] node836;
	wire [16-1:0] node839;
	wire [16-1:0] node842;
	wire [16-1:0] node843;
	wire [16-1:0] node846;
	wire [16-1:0] node849;
	wire [16-1:0] node850;
	wire [16-1:0] node851;
	wire [16-1:0] node852;
	wire [16-1:0] node853;
	wire [16-1:0] node854;
	wire [16-1:0] node857;
	wire [16-1:0] node860;
	wire [16-1:0] node861;
	wire [16-1:0] node864;
	wire [16-1:0] node867;
	wire [16-1:0] node868;
	wire [16-1:0] node869;
	wire [16-1:0] node872;
	wire [16-1:0] node875;
	wire [16-1:0] node876;
	wire [16-1:0] node879;
	wire [16-1:0] node882;
	wire [16-1:0] node883;
	wire [16-1:0] node884;
	wire [16-1:0] node885;
	wire [16-1:0] node888;
	wire [16-1:0] node891;
	wire [16-1:0] node892;
	wire [16-1:0] node896;
	wire [16-1:0] node897;
	wire [16-1:0] node898;
	wire [16-1:0] node901;
	wire [16-1:0] node904;
	wire [16-1:0] node905;
	wire [16-1:0] node908;
	wire [16-1:0] node911;
	wire [16-1:0] node912;
	wire [16-1:0] node913;
	wire [16-1:0] node914;
	wire [16-1:0] node915;
	wire [16-1:0] node918;
	wire [16-1:0] node921;
	wire [16-1:0] node922;
	wire [16-1:0] node925;
	wire [16-1:0] node928;
	wire [16-1:0] node929;
	wire [16-1:0] node930;
	wire [16-1:0] node933;
	wire [16-1:0] node936;
	wire [16-1:0] node938;
	wire [16-1:0] node941;
	wire [16-1:0] node942;
	wire [16-1:0] node943;
	wire [16-1:0] node944;
	wire [16-1:0] node947;
	wire [16-1:0] node950;
	wire [16-1:0] node951;
	wire [16-1:0] node954;
	wire [16-1:0] node957;
	wire [16-1:0] node958;
	wire [16-1:0] node959;
	wire [16-1:0] node962;
	wire [16-1:0] node965;
	wire [16-1:0] node966;
	wire [16-1:0] node969;
	wire [16-1:0] node972;
	wire [16-1:0] node973;
	wire [16-1:0] node974;
	wire [16-1:0] node975;
	wire [16-1:0] node976;
	wire [16-1:0] node977;
	wire [16-1:0] node978;
	wire [16-1:0] node979;
	wire [16-1:0] node980;
	wire [16-1:0] node983;
	wire [16-1:0] node986;
	wire [16-1:0] node987;
	wire [16-1:0] node990;
	wire [16-1:0] node993;
	wire [16-1:0] node994;
	wire [16-1:0] node995;
	wire [16-1:0] node998;
	wire [16-1:0] node1001;
	wire [16-1:0] node1002;
	wire [16-1:0] node1005;
	wire [16-1:0] node1008;
	wire [16-1:0] node1009;
	wire [16-1:0] node1010;
	wire [16-1:0] node1011;
	wire [16-1:0] node1014;
	wire [16-1:0] node1017;
	wire [16-1:0] node1018;
	wire [16-1:0] node1021;
	wire [16-1:0] node1024;
	wire [16-1:0] node1025;
	wire [16-1:0] node1026;
	wire [16-1:0] node1029;
	wire [16-1:0] node1032;
	wire [16-1:0] node1033;
	wire [16-1:0] node1036;
	wire [16-1:0] node1039;
	wire [16-1:0] node1040;
	wire [16-1:0] node1041;
	wire [16-1:0] node1042;
	wire [16-1:0] node1043;
	wire [16-1:0] node1046;
	wire [16-1:0] node1049;
	wire [16-1:0] node1050;
	wire [16-1:0] node1053;
	wire [16-1:0] node1056;
	wire [16-1:0] node1057;
	wire [16-1:0] node1058;
	wire [16-1:0] node1061;
	wire [16-1:0] node1064;
	wire [16-1:0] node1065;
	wire [16-1:0] node1068;
	wire [16-1:0] node1071;
	wire [16-1:0] node1072;
	wire [16-1:0] node1073;
	wire [16-1:0] node1074;
	wire [16-1:0] node1077;
	wire [16-1:0] node1080;
	wire [16-1:0] node1081;
	wire [16-1:0] node1084;
	wire [16-1:0] node1087;
	wire [16-1:0] node1088;
	wire [16-1:0] node1089;
	wire [16-1:0] node1092;
	wire [16-1:0] node1095;
	wire [16-1:0] node1096;
	wire [16-1:0] node1099;
	wire [16-1:0] node1102;
	wire [16-1:0] node1103;
	wire [16-1:0] node1104;
	wire [16-1:0] node1105;
	wire [16-1:0] node1106;
	wire [16-1:0] node1107;
	wire [16-1:0] node1110;
	wire [16-1:0] node1113;
	wire [16-1:0] node1114;
	wire [16-1:0] node1118;
	wire [16-1:0] node1119;
	wire [16-1:0] node1120;
	wire [16-1:0] node1123;
	wire [16-1:0] node1126;
	wire [16-1:0] node1127;
	wire [16-1:0] node1130;
	wire [16-1:0] node1133;
	wire [16-1:0] node1134;
	wire [16-1:0] node1135;
	wire [16-1:0] node1136;
	wire [16-1:0] node1139;
	wire [16-1:0] node1142;
	wire [16-1:0] node1143;
	wire [16-1:0] node1146;
	wire [16-1:0] node1149;
	wire [16-1:0] node1150;
	wire [16-1:0] node1151;
	wire [16-1:0] node1154;
	wire [16-1:0] node1157;
	wire [16-1:0] node1158;
	wire [16-1:0] node1161;
	wire [16-1:0] node1164;
	wire [16-1:0] node1165;
	wire [16-1:0] node1166;
	wire [16-1:0] node1167;
	wire [16-1:0] node1168;
	wire [16-1:0] node1171;
	wire [16-1:0] node1174;
	wire [16-1:0] node1175;
	wire [16-1:0] node1178;
	wire [16-1:0] node1181;
	wire [16-1:0] node1182;
	wire [16-1:0] node1184;
	wire [16-1:0] node1187;
	wire [16-1:0] node1188;
	wire [16-1:0] node1192;
	wire [16-1:0] node1193;
	wire [16-1:0] node1194;
	wire [16-1:0] node1195;
	wire [16-1:0] node1198;
	wire [16-1:0] node1201;
	wire [16-1:0] node1202;
	wire [16-1:0] node1205;
	wire [16-1:0] node1208;
	wire [16-1:0] node1209;
	wire [16-1:0] node1210;
	wire [16-1:0] node1213;
	wire [16-1:0] node1216;
	wire [16-1:0] node1217;
	wire [16-1:0] node1220;
	wire [16-1:0] node1223;
	wire [16-1:0] node1224;
	wire [16-1:0] node1225;
	wire [16-1:0] node1226;
	wire [16-1:0] node1227;
	wire [16-1:0] node1228;
	wire [16-1:0] node1229;
	wire [16-1:0] node1232;
	wire [16-1:0] node1235;
	wire [16-1:0] node1236;
	wire [16-1:0] node1239;
	wire [16-1:0] node1242;
	wire [16-1:0] node1243;
	wire [16-1:0] node1244;
	wire [16-1:0] node1247;
	wire [16-1:0] node1250;
	wire [16-1:0] node1251;
	wire [16-1:0] node1254;
	wire [16-1:0] node1257;
	wire [16-1:0] node1258;
	wire [16-1:0] node1259;
	wire [16-1:0] node1260;
	wire [16-1:0] node1263;
	wire [16-1:0] node1266;
	wire [16-1:0] node1267;
	wire [16-1:0] node1270;
	wire [16-1:0] node1273;
	wire [16-1:0] node1274;
	wire [16-1:0] node1275;
	wire [16-1:0] node1278;
	wire [16-1:0] node1281;
	wire [16-1:0] node1282;
	wire [16-1:0] node1285;
	wire [16-1:0] node1288;
	wire [16-1:0] node1289;
	wire [16-1:0] node1290;
	wire [16-1:0] node1291;
	wire [16-1:0] node1292;
	wire [16-1:0] node1295;
	wire [16-1:0] node1298;
	wire [16-1:0] node1299;
	wire [16-1:0] node1302;
	wire [16-1:0] node1305;
	wire [16-1:0] node1306;
	wire [16-1:0] node1307;
	wire [16-1:0] node1310;
	wire [16-1:0] node1313;
	wire [16-1:0] node1314;
	wire [16-1:0] node1317;
	wire [16-1:0] node1320;
	wire [16-1:0] node1321;
	wire [16-1:0] node1322;
	wire [16-1:0] node1323;
	wire [16-1:0] node1326;
	wire [16-1:0] node1329;
	wire [16-1:0] node1330;
	wire [16-1:0] node1333;
	wire [16-1:0] node1336;
	wire [16-1:0] node1337;
	wire [16-1:0] node1338;
	wire [16-1:0] node1341;
	wire [16-1:0] node1344;
	wire [16-1:0] node1345;
	wire [16-1:0] node1348;
	wire [16-1:0] node1351;
	wire [16-1:0] node1352;
	wire [16-1:0] node1353;
	wire [16-1:0] node1354;
	wire [16-1:0] node1355;
	wire [16-1:0] node1357;
	wire [16-1:0] node1360;
	wire [16-1:0] node1361;
	wire [16-1:0] node1364;
	wire [16-1:0] node1367;
	wire [16-1:0] node1368;
	wire [16-1:0] node1369;
	wire [16-1:0] node1372;
	wire [16-1:0] node1375;
	wire [16-1:0] node1376;
	wire [16-1:0] node1379;
	wire [16-1:0] node1382;
	wire [16-1:0] node1383;
	wire [16-1:0] node1384;
	wire [16-1:0] node1386;
	wire [16-1:0] node1389;
	wire [16-1:0] node1390;
	wire [16-1:0] node1393;
	wire [16-1:0] node1396;
	wire [16-1:0] node1397;
	wire [16-1:0] node1398;
	wire [16-1:0] node1401;
	wire [16-1:0] node1404;
	wire [16-1:0] node1405;
	wire [16-1:0] node1408;
	wire [16-1:0] node1411;
	wire [16-1:0] node1412;
	wire [16-1:0] node1413;
	wire [16-1:0] node1414;
	wire [16-1:0] node1415;
	wire [16-1:0] node1418;
	wire [16-1:0] node1421;
	wire [16-1:0] node1422;
	wire [16-1:0] node1425;
	wire [16-1:0] node1428;
	wire [16-1:0] node1429;
	wire [16-1:0] node1431;
	wire [16-1:0] node1434;
	wire [16-1:0] node1435;
	wire [16-1:0] node1438;
	wire [16-1:0] node1441;
	wire [16-1:0] node1442;
	wire [16-1:0] node1443;
	wire [16-1:0] node1444;
	wire [16-1:0] node1447;
	wire [16-1:0] node1450;
	wire [16-1:0] node1451;
	wire [16-1:0] node1454;
	wire [16-1:0] node1457;
	wire [16-1:0] node1458;
	wire [16-1:0] node1460;
	wire [16-1:0] node1463;
	wire [16-1:0] node1464;
	wire [16-1:0] node1467;
	wire [16-1:0] node1470;
	wire [16-1:0] node1471;
	wire [16-1:0] node1472;
	wire [16-1:0] node1473;
	wire [16-1:0] node1474;
	wire [16-1:0] node1475;
	wire [16-1:0] node1476;
	wire [16-1:0] node1477;
	wire [16-1:0] node1480;
	wire [16-1:0] node1483;
	wire [16-1:0] node1484;
	wire [16-1:0] node1487;
	wire [16-1:0] node1490;
	wire [16-1:0] node1491;
	wire [16-1:0] node1492;
	wire [16-1:0] node1495;
	wire [16-1:0] node1498;
	wire [16-1:0] node1499;
	wire [16-1:0] node1503;
	wire [16-1:0] node1504;
	wire [16-1:0] node1505;
	wire [16-1:0] node1506;
	wire [16-1:0] node1510;
	wire [16-1:0] node1511;
	wire [16-1:0] node1514;
	wire [16-1:0] node1517;
	wire [16-1:0] node1518;
	wire [16-1:0] node1519;
	wire [16-1:0] node1523;
	wire [16-1:0] node1524;
	wire [16-1:0] node1527;
	wire [16-1:0] node1530;
	wire [16-1:0] node1531;
	wire [16-1:0] node1532;
	wire [16-1:0] node1533;
	wire [16-1:0] node1534;
	wire [16-1:0] node1537;
	wire [16-1:0] node1540;
	wire [16-1:0] node1541;
	wire [16-1:0] node1544;
	wire [16-1:0] node1547;
	wire [16-1:0] node1548;
	wire [16-1:0] node1549;
	wire [16-1:0] node1552;
	wire [16-1:0] node1555;
	wire [16-1:0] node1556;
	wire [16-1:0] node1559;
	wire [16-1:0] node1562;
	wire [16-1:0] node1563;
	wire [16-1:0] node1564;
	wire [16-1:0] node1565;
	wire [16-1:0] node1568;
	wire [16-1:0] node1571;
	wire [16-1:0] node1572;
	wire [16-1:0] node1575;
	wire [16-1:0] node1578;
	wire [16-1:0] node1579;
	wire [16-1:0] node1580;
	wire [16-1:0] node1583;
	wire [16-1:0] node1586;
	wire [16-1:0] node1587;
	wire [16-1:0] node1590;
	wire [16-1:0] node1593;
	wire [16-1:0] node1594;
	wire [16-1:0] node1595;
	wire [16-1:0] node1596;
	wire [16-1:0] node1597;
	wire [16-1:0] node1598;
	wire [16-1:0] node1601;
	wire [16-1:0] node1604;
	wire [16-1:0] node1605;
	wire [16-1:0] node1608;
	wire [16-1:0] node1611;
	wire [16-1:0] node1612;
	wire [16-1:0] node1613;
	wire [16-1:0] node1616;
	wire [16-1:0] node1619;
	wire [16-1:0] node1620;
	wire [16-1:0] node1623;
	wire [16-1:0] node1626;
	wire [16-1:0] node1627;
	wire [16-1:0] node1628;
	wire [16-1:0] node1629;
	wire [16-1:0] node1632;
	wire [16-1:0] node1635;
	wire [16-1:0] node1636;
	wire [16-1:0] node1639;
	wire [16-1:0] node1642;
	wire [16-1:0] node1643;
	wire [16-1:0] node1645;
	wire [16-1:0] node1648;
	wire [16-1:0] node1651;
	wire [16-1:0] node1652;
	wire [16-1:0] node1653;
	wire [16-1:0] node1654;
	wire [16-1:0] node1655;
	wire [16-1:0] node1658;
	wire [16-1:0] node1661;
	wire [16-1:0] node1662;
	wire [16-1:0] node1665;
	wire [16-1:0] node1668;
	wire [16-1:0] node1669;
	wire [16-1:0] node1670;
	wire [16-1:0] node1673;
	wire [16-1:0] node1676;
	wire [16-1:0] node1677;
	wire [16-1:0] node1681;
	wire [16-1:0] node1682;
	wire [16-1:0] node1683;
	wire [16-1:0] node1685;
	wire [16-1:0] node1688;
	wire [16-1:0] node1689;
	wire [16-1:0] node1692;
	wire [16-1:0] node1695;
	wire [16-1:0] node1696;
	wire [16-1:0] node1697;
	wire [16-1:0] node1700;
	wire [16-1:0] node1703;
	wire [16-1:0] node1704;
	wire [16-1:0] node1707;
	wire [16-1:0] node1710;
	wire [16-1:0] node1711;
	wire [16-1:0] node1712;
	wire [16-1:0] node1713;
	wire [16-1:0] node1714;
	wire [16-1:0] node1715;
	wire [16-1:0] node1717;
	wire [16-1:0] node1720;
	wire [16-1:0] node1721;
	wire [16-1:0] node1725;
	wire [16-1:0] node1727;
	wire [16-1:0] node1728;
	wire [16-1:0] node1732;
	wire [16-1:0] node1733;
	wire [16-1:0] node1734;
	wire [16-1:0] node1736;
	wire [16-1:0] node1739;
	wire [16-1:0] node1740;
	wire [16-1:0] node1743;
	wire [16-1:0] node1746;
	wire [16-1:0] node1747;
	wire [16-1:0] node1748;
	wire [16-1:0] node1751;
	wire [16-1:0] node1754;
	wire [16-1:0] node1755;
	wire [16-1:0] node1758;
	wire [16-1:0] node1761;
	wire [16-1:0] node1762;
	wire [16-1:0] node1763;
	wire [16-1:0] node1764;
	wire [16-1:0] node1765;
	wire [16-1:0] node1768;
	wire [16-1:0] node1771;
	wire [16-1:0] node1772;
	wire [16-1:0] node1775;
	wire [16-1:0] node1778;
	wire [16-1:0] node1779;
	wire [16-1:0] node1780;
	wire [16-1:0] node1783;
	wire [16-1:0] node1786;
	wire [16-1:0] node1787;
	wire [16-1:0] node1790;
	wire [16-1:0] node1793;
	wire [16-1:0] node1794;
	wire [16-1:0] node1795;
	wire [16-1:0] node1796;
	wire [16-1:0] node1799;
	wire [16-1:0] node1802;
	wire [16-1:0] node1803;
	wire [16-1:0] node1806;
	wire [16-1:0] node1809;
	wire [16-1:0] node1810;
	wire [16-1:0] node1811;
	wire [16-1:0] node1814;
	wire [16-1:0] node1817;
	wire [16-1:0] node1818;
	wire [16-1:0] node1821;
	wire [16-1:0] node1824;
	wire [16-1:0] node1825;
	wire [16-1:0] node1826;
	wire [16-1:0] node1827;
	wire [16-1:0] node1828;
	wire [16-1:0] node1829;
	wire [16-1:0] node1832;
	wire [16-1:0] node1835;
	wire [16-1:0] node1836;
	wire [16-1:0] node1839;
	wire [16-1:0] node1842;
	wire [16-1:0] node1843;
	wire [16-1:0] node1844;
	wire [16-1:0] node1847;
	wire [16-1:0] node1850;
	wire [16-1:0] node1852;
	wire [16-1:0] node1855;
	wire [16-1:0] node1856;
	wire [16-1:0] node1857;
	wire [16-1:0] node1858;
	wire [16-1:0] node1861;
	wire [16-1:0] node1864;
	wire [16-1:0] node1865;
	wire [16-1:0] node1868;
	wire [16-1:0] node1871;
	wire [16-1:0] node1872;
	wire [16-1:0] node1874;
	wire [16-1:0] node1877;
	wire [16-1:0] node1878;
	wire [16-1:0] node1881;
	wire [16-1:0] node1884;
	wire [16-1:0] node1885;
	wire [16-1:0] node1886;
	wire [16-1:0] node1887;
	wire [16-1:0] node1889;
	wire [16-1:0] node1892;
	wire [16-1:0] node1893;
	wire [16-1:0] node1896;
	wire [16-1:0] node1899;
	wire [16-1:0] node1900;
	wire [16-1:0] node1901;
	wire [16-1:0] node1904;
	wire [16-1:0] node1907;
	wire [16-1:0] node1908;
	wire [16-1:0] node1911;
	wire [16-1:0] node1914;
	wire [16-1:0] node1915;
	wire [16-1:0] node1916;
	wire [16-1:0] node1917;
	wire [16-1:0] node1920;
	wire [16-1:0] node1923;
	wire [16-1:0] node1924;
	wire [16-1:0] node1927;
	wire [16-1:0] node1930;
	wire [16-1:0] node1931;
	wire [16-1:0] node1932;
	wire [16-1:0] node1935;
	wire [16-1:0] node1938;
	wire [16-1:0] node1939;
	wire [16-1:0] node1942;
	wire [16-1:0] node1945;
	wire [16-1:0] node1946;
	wire [16-1:0] node1947;
	wire [16-1:0] node1948;
	wire [16-1:0] node1949;
	wire [16-1:0] node1950;
	wire [16-1:0] node1951;
	wire [16-1:0] node1952;
	wire [16-1:0] node1953;
	wire [16-1:0] node1954;
	wire [16-1:0] node1957;
	wire [16-1:0] node1960;
	wire [16-1:0] node1961;
	wire [16-1:0] node1964;
	wire [16-1:0] node1967;
	wire [16-1:0] node1968;
	wire [16-1:0] node1969;
	wire [16-1:0] node1972;
	wire [16-1:0] node1975;
	wire [16-1:0] node1976;
	wire [16-1:0] node1979;
	wire [16-1:0] node1982;
	wire [16-1:0] node1983;
	wire [16-1:0] node1984;
	wire [16-1:0] node1985;
	wire [16-1:0] node1988;
	wire [16-1:0] node1991;
	wire [16-1:0] node1992;
	wire [16-1:0] node1995;
	wire [16-1:0] node1998;
	wire [16-1:0] node1999;
	wire [16-1:0] node2000;
	wire [16-1:0] node2003;
	wire [16-1:0] node2006;
	wire [16-1:0] node2007;
	wire [16-1:0] node2010;
	wire [16-1:0] node2013;
	wire [16-1:0] node2014;
	wire [16-1:0] node2015;
	wire [16-1:0] node2016;
	wire [16-1:0] node2017;
	wire [16-1:0] node2020;
	wire [16-1:0] node2023;
	wire [16-1:0] node2024;
	wire [16-1:0] node2028;
	wire [16-1:0] node2029;
	wire [16-1:0] node2031;
	wire [16-1:0] node2034;
	wire [16-1:0] node2035;
	wire [16-1:0] node2038;
	wire [16-1:0] node2041;
	wire [16-1:0] node2042;
	wire [16-1:0] node2043;
	wire [16-1:0] node2044;
	wire [16-1:0] node2047;
	wire [16-1:0] node2050;
	wire [16-1:0] node2051;
	wire [16-1:0] node2054;
	wire [16-1:0] node2057;
	wire [16-1:0] node2058;
	wire [16-1:0] node2059;
	wire [16-1:0] node2063;
	wire [16-1:0] node2064;
	wire [16-1:0] node2067;
	wire [16-1:0] node2070;
	wire [16-1:0] node2071;
	wire [16-1:0] node2072;
	wire [16-1:0] node2073;
	wire [16-1:0] node2074;
	wire [16-1:0] node2075;
	wire [16-1:0] node2078;
	wire [16-1:0] node2081;
	wire [16-1:0] node2082;
	wire [16-1:0] node2085;
	wire [16-1:0] node2088;
	wire [16-1:0] node2089;
	wire [16-1:0] node2090;
	wire [16-1:0] node2093;
	wire [16-1:0] node2096;
	wire [16-1:0] node2097;
	wire [16-1:0] node2100;
	wire [16-1:0] node2103;
	wire [16-1:0] node2104;
	wire [16-1:0] node2105;
	wire [16-1:0] node2106;
	wire [16-1:0] node2109;
	wire [16-1:0] node2112;
	wire [16-1:0] node2113;
	wire [16-1:0] node2116;
	wire [16-1:0] node2119;
	wire [16-1:0] node2120;
	wire [16-1:0] node2121;
	wire [16-1:0] node2124;
	wire [16-1:0] node2127;
	wire [16-1:0] node2128;
	wire [16-1:0] node2131;
	wire [16-1:0] node2134;
	wire [16-1:0] node2135;
	wire [16-1:0] node2136;
	wire [16-1:0] node2137;
	wire [16-1:0] node2138;
	wire [16-1:0] node2141;
	wire [16-1:0] node2144;
	wire [16-1:0] node2145;
	wire [16-1:0] node2148;
	wire [16-1:0] node2151;
	wire [16-1:0] node2152;
	wire [16-1:0] node2153;
	wire [16-1:0] node2157;
	wire [16-1:0] node2158;
	wire [16-1:0] node2161;
	wire [16-1:0] node2164;
	wire [16-1:0] node2165;
	wire [16-1:0] node2166;
	wire [16-1:0] node2167;
	wire [16-1:0] node2170;
	wire [16-1:0] node2173;
	wire [16-1:0] node2174;
	wire [16-1:0] node2177;
	wire [16-1:0] node2180;
	wire [16-1:0] node2181;
	wire [16-1:0] node2182;
	wire [16-1:0] node2185;
	wire [16-1:0] node2188;
	wire [16-1:0] node2189;
	wire [16-1:0] node2192;
	wire [16-1:0] node2195;
	wire [16-1:0] node2196;
	wire [16-1:0] node2197;
	wire [16-1:0] node2198;
	wire [16-1:0] node2199;
	wire [16-1:0] node2200;
	wire [16-1:0] node2201;
	wire [16-1:0] node2204;
	wire [16-1:0] node2207;
	wire [16-1:0] node2208;
	wire [16-1:0] node2211;
	wire [16-1:0] node2214;
	wire [16-1:0] node2215;
	wire [16-1:0] node2216;
	wire [16-1:0] node2219;
	wire [16-1:0] node2222;
	wire [16-1:0] node2223;
	wire [16-1:0] node2226;
	wire [16-1:0] node2229;
	wire [16-1:0] node2230;
	wire [16-1:0] node2231;
	wire [16-1:0] node2232;
	wire [16-1:0] node2235;
	wire [16-1:0] node2238;
	wire [16-1:0] node2239;
	wire [16-1:0] node2242;
	wire [16-1:0] node2245;
	wire [16-1:0] node2246;
	wire [16-1:0] node2247;
	wire [16-1:0] node2251;
	wire [16-1:0] node2252;
	wire [16-1:0] node2256;
	wire [16-1:0] node2257;
	wire [16-1:0] node2258;
	wire [16-1:0] node2259;
	wire [16-1:0] node2260;
	wire [16-1:0] node2263;
	wire [16-1:0] node2266;
	wire [16-1:0] node2267;
	wire [16-1:0] node2270;
	wire [16-1:0] node2273;
	wire [16-1:0] node2274;
	wire [16-1:0] node2275;
	wire [16-1:0] node2278;
	wire [16-1:0] node2281;
	wire [16-1:0] node2282;
	wire [16-1:0] node2285;
	wire [16-1:0] node2288;
	wire [16-1:0] node2289;
	wire [16-1:0] node2290;
	wire [16-1:0] node2291;
	wire [16-1:0] node2294;
	wire [16-1:0] node2297;
	wire [16-1:0] node2298;
	wire [16-1:0] node2301;
	wire [16-1:0] node2304;
	wire [16-1:0] node2305;
	wire [16-1:0] node2306;
	wire [16-1:0] node2309;
	wire [16-1:0] node2312;
	wire [16-1:0] node2313;
	wire [16-1:0] node2316;
	wire [16-1:0] node2319;
	wire [16-1:0] node2320;
	wire [16-1:0] node2321;
	wire [16-1:0] node2322;
	wire [16-1:0] node2323;
	wire [16-1:0] node2324;
	wire [16-1:0] node2327;
	wire [16-1:0] node2330;
	wire [16-1:0] node2331;
	wire [16-1:0] node2334;
	wire [16-1:0] node2337;
	wire [16-1:0] node2338;
	wire [16-1:0] node2339;
	wire [16-1:0] node2342;
	wire [16-1:0] node2345;
	wire [16-1:0] node2346;
	wire [16-1:0] node2349;
	wire [16-1:0] node2352;
	wire [16-1:0] node2353;
	wire [16-1:0] node2354;
	wire [16-1:0] node2355;
	wire [16-1:0] node2358;
	wire [16-1:0] node2361;
	wire [16-1:0] node2362;
	wire [16-1:0] node2366;
	wire [16-1:0] node2367;
	wire [16-1:0] node2368;
	wire [16-1:0] node2372;
	wire [16-1:0] node2373;
	wire [16-1:0] node2376;
	wire [16-1:0] node2379;
	wire [16-1:0] node2380;
	wire [16-1:0] node2381;
	wire [16-1:0] node2382;
	wire [16-1:0] node2383;
	wire [16-1:0] node2386;
	wire [16-1:0] node2389;
	wire [16-1:0] node2390;
	wire [16-1:0] node2393;
	wire [16-1:0] node2396;
	wire [16-1:0] node2397;
	wire [16-1:0] node2398;
	wire [16-1:0] node2401;
	wire [16-1:0] node2404;
	wire [16-1:0] node2405;
	wire [16-1:0] node2408;
	wire [16-1:0] node2411;
	wire [16-1:0] node2412;
	wire [16-1:0] node2413;
	wire [16-1:0] node2414;
	wire [16-1:0] node2417;
	wire [16-1:0] node2420;
	wire [16-1:0] node2421;
	wire [16-1:0] node2424;
	wire [16-1:0] node2427;
	wire [16-1:0] node2428;
	wire [16-1:0] node2430;
	wire [16-1:0] node2433;
	wire [16-1:0] node2434;
	wire [16-1:0] node2437;
	wire [16-1:0] node2440;
	wire [16-1:0] node2441;
	wire [16-1:0] node2442;
	wire [16-1:0] node2443;
	wire [16-1:0] node2444;
	wire [16-1:0] node2445;
	wire [16-1:0] node2446;
	wire [16-1:0] node2447;
	wire [16-1:0] node2451;
	wire [16-1:0] node2452;
	wire [16-1:0] node2455;
	wire [16-1:0] node2458;
	wire [16-1:0] node2459;
	wire [16-1:0] node2460;
	wire [16-1:0] node2463;
	wire [16-1:0] node2466;
	wire [16-1:0] node2467;
	wire [16-1:0] node2471;
	wire [16-1:0] node2472;
	wire [16-1:0] node2473;
	wire [16-1:0] node2474;
	wire [16-1:0] node2477;
	wire [16-1:0] node2480;
	wire [16-1:0] node2481;
	wire [16-1:0] node2484;
	wire [16-1:0] node2487;
	wire [16-1:0] node2488;
	wire [16-1:0] node2489;
	wire [16-1:0] node2492;
	wire [16-1:0] node2495;
	wire [16-1:0] node2496;
	wire [16-1:0] node2500;
	wire [16-1:0] node2501;
	wire [16-1:0] node2502;
	wire [16-1:0] node2503;
	wire [16-1:0] node2504;
	wire [16-1:0] node2507;
	wire [16-1:0] node2510;
	wire [16-1:0] node2511;
	wire [16-1:0] node2515;
	wire [16-1:0] node2516;
	wire [16-1:0] node2517;
	wire [16-1:0] node2520;
	wire [16-1:0] node2523;
	wire [16-1:0] node2524;
	wire [16-1:0] node2527;
	wire [16-1:0] node2530;
	wire [16-1:0] node2531;
	wire [16-1:0] node2532;
	wire [16-1:0] node2533;
	wire [16-1:0] node2537;
	wire [16-1:0] node2538;
	wire [16-1:0] node2542;
	wire [16-1:0] node2543;
	wire [16-1:0] node2544;
	wire [16-1:0] node2547;
	wire [16-1:0] node2550;
	wire [16-1:0] node2552;
	wire [16-1:0] node2555;
	wire [16-1:0] node2556;
	wire [16-1:0] node2557;
	wire [16-1:0] node2558;
	wire [16-1:0] node2559;
	wire [16-1:0] node2560;
	wire [16-1:0] node2563;
	wire [16-1:0] node2566;
	wire [16-1:0] node2567;
	wire [16-1:0] node2570;
	wire [16-1:0] node2573;
	wire [16-1:0] node2574;
	wire [16-1:0] node2575;
	wire [16-1:0] node2578;
	wire [16-1:0] node2581;
	wire [16-1:0] node2582;
	wire [16-1:0] node2585;
	wire [16-1:0] node2588;
	wire [16-1:0] node2589;
	wire [16-1:0] node2590;
	wire [16-1:0] node2591;
	wire [16-1:0] node2594;
	wire [16-1:0] node2597;
	wire [16-1:0] node2598;
	wire [16-1:0] node2601;
	wire [16-1:0] node2604;
	wire [16-1:0] node2605;
	wire [16-1:0] node2606;
	wire [16-1:0] node2609;
	wire [16-1:0] node2613;
	wire [16-1:0] node2614;
	wire [16-1:0] node2615;
	wire [16-1:0] node2616;
	wire [16-1:0] node2617;
	wire [16-1:0] node2620;
	wire [16-1:0] node2623;
	wire [16-1:0] node2624;
	wire [16-1:0] node2628;
	wire [16-1:0] node2629;
	wire [16-1:0] node2630;
	wire [16-1:0] node2633;
	wire [16-1:0] node2636;
	wire [16-1:0] node2637;
	wire [16-1:0] node2640;
	wire [16-1:0] node2643;
	wire [16-1:0] node2644;
	wire [16-1:0] node2645;
	wire [16-1:0] node2646;
	wire [16-1:0] node2649;
	wire [16-1:0] node2652;
	wire [16-1:0] node2653;
	wire [16-1:0] node2656;
	wire [16-1:0] node2659;
	wire [16-1:0] node2660;
	wire [16-1:0] node2661;
	wire [16-1:0] node2664;
	wire [16-1:0] node2667;
	wire [16-1:0] node2669;
	wire [16-1:0] node2672;
	wire [16-1:0] node2673;
	wire [16-1:0] node2674;
	wire [16-1:0] node2675;
	wire [16-1:0] node2676;
	wire [16-1:0] node2677;
	wire [16-1:0] node2678;
	wire [16-1:0] node2681;
	wire [16-1:0] node2684;
	wire [16-1:0] node2685;
	wire [16-1:0] node2688;
	wire [16-1:0] node2691;
	wire [16-1:0] node2692;
	wire [16-1:0] node2693;
	wire [16-1:0] node2696;
	wire [16-1:0] node2699;
	wire [16-1:0] node2700;
	wire [16-1:0] node2703;
	wire [16-1:0] node2706;
	wire [16-1:0] node2707;
	wire [16-1:0] node2708;
	wire [16-1:0] node2709;
	wire [16-1:0] node2712;
	wire [16-1:0] node2715;
	wire [16-1:0] node2716;
	wire [16-1:0] node2719;
	wire [16-1:0] node2722;
	wire [16-1:0] node2723;
	wire [16-1:0] node2724;
	wire [16-1:0] node2727;
	wire [16-1:0] node2730;
	wire [16-1:0] node2731;
	wire [16-1:0] node2734;
	wire [16-1:0] node2737;
	wire [16-1:0] node2738;
	wire [16-1:0] node2739;
	wire [16-1:0] node2740;
	wire [16-1:0] node2741;
	wire [16-1:0] node2744;
	wire [16-1:0] node2747;
	wire [16-1:0] node2748;
	wire [16-1:0] node2752;
	wire [16-1:0] node2753;
	wire [16-1:0] node2754;
	wire [16-1:0] node2757;
	wire [16-1:0] node2760;
	wire [16-1:0] node2761;
	wire [16-1:0] node2764;
	wire [16-1:0] node2767;
	wire [16-1:0] node2768;
	wire [16-1:0] node2769;
	wire [16-1:0] node2770;
	wire [16-1:0] node2773;
	wire [16-1:0] node2776;
	wire [16-1:0] node2777;
	wire [16-1:0] node2781;
	wire [16-1:0] node2782;
	wire [16-1:0] node2783;
	wire [16-1:0] node2786;
	wire [16-1:0] node2789;
	wire [16-1:0] node2790;
	wire [16-1:0] node2793;
	wire [16-1:0] node2796;
	wire [16-1:0] node2797;
	wire [16-1:0] node2798;
	wire [16-1:0] node2799;
	wire [16-1:0] node2800;
	wire [16-1:0] node2801;
	wire [16-1:0] node2804;
	wire [16-1:0] node2807;
	wire [16-1:0] node2810;
	wire [16-1:0] node2811;
	wire [16-1:0] node2812;
	wire [16-1:0] node2815;
	wire [16-1:0] node2818;
	wire [16-1:0] node2819;
	wire [16-1:0] node2822;
	wire [16-1:0] node2825;
	wire [16-1:0] node2826;
	wire [16-1:0] node2827;
	wire [16-1:0] node2828;
	wire [16-1:0] node2831;
	wire [16-1:0] node2834;
	wire [16-1:0] node2835;
	wire [16-1:0] node2838;
	wire [16-1:0] node2841;
	wire [16-1:0] node2842;
	wire [16-1:0] node2843;
	wire [16-1:0] node2846;
	wire [16-1:0] node2849;
	wire [16-1:0] node2850;
	wire [16-1:0] node2853;
	wire [16-1:0] node2856;
	wire [16-1:0] node2857;
	wire [16-1:0] node2858;
	wire [16-1:0] node2859;
	wire [16-1:0] node2860;
	wire [16-1:0] node2863;
	wire [16-1:0] node2866;
	wire [16-1:0] node2867;
	wire [16-1:0] node2870;
	wire [16-1:0] node2873;
	wire [16-1:0] node2874;
	wire [16-1:0] node2875;
	wire [16-1:0] node2878;
	wire [16-1:0] node2882;
	wire [16-1:0] node2883;
	wire [16-1:0] node2884;
	wire [16-1:0] node2885;
	wire [16-1:0] node2888;
	wire [16-1:0] node2891;
	wire [16-1:0] node2892;
	wire [16-1:0] node2895;
	wire [16-1:0] node2898;
	wire [16-1:0] node2899;
	wire [16-1:0] node2901;
	wire [16-1:0] node2904;
	wire [16-1:0] node2905;
	wire [16-1:0] node2908;
	wire [16-1:0] node2911;
	wire [16-1:0] node2912;
	wire [16-1:0] node2913;
	wire [16-1:0] node2914;
	wire [16-1:0] node2915;
	wire [16-1:0] node2916;
	wire [16-1:0] node2917;
	wire [16-1:0] node2918;
	wire [16-1:0] node2919;
	wire [16-1:0] node2922;
	wire [16-1:0] node2925;
	wire [16-1:0] node2927;
	wire [16-1:0] node2930;
	wire [16-1:0] node2931;
	wire [16-1:0] node2932;
	wire [16-1:0] node2936;
	wire [16-1:0] node2937;
	wire [16-1:0] node2941;
	wire [16-1:0] node2942;
	wire [16-1:0] node2943;
	wire [16-1:0] node2944;
	wire [16-1:0] node2947;
	wire [16-1:0] node2950;
	wire [16-1:0] node2951;
	wire [16-1:0] node2954;
	wire [16-1:0] node2957;
	wire [16-1:0] node2958;
	wire [16-1:0] node2960;
	wire [16-1:0] node2963;
	wire [16-1:0] node2964;
	wire [16-1:0] node2967;
	wire [16-1:0] node2970;
	wire [16-1:0] node2971;
	wire [16-1:0] node2972;
	wire [16-1:0] node2973;
	wire [16-1:0] node2974;
	wire [16-1:0] node2977;
	wire [16-1:0] node2980;
	wire [16-1:0] node2981;
	wire [16-1:0] node2984;
	wire [16-1:0] node2987;
	wire [16-1:0] node2988;
	wire [16-1:0] node2989;
	wire [16-1:0] node2992;
	wire [16-1:0] node2995;
	wire [16-1:0] node2996;
	wire [16-1:0] node2999;
	wire [16-1:0] node3002;
	wire [16-1:0] node3003;
	wire [16-1:0] node3004;
	wire [16-1:0] node3005;
	wire [16-1:0] node3008;
	wire [16-1:0] node3011;
	wire [16-1:0] node3012;
	wire [16-1:0] node3015;
	wire [16-1:0] node3018;
	wire [16-1:0] node3019;
	wire [16-1:0] node3020;
	wire [16-1:0] node3023;
	wire [16-1:0] node3026;
	wire [16-1:0] node3027;
	wire [16-1:0] node3030;
	wire [16-1:0] node3033;
	wire [16-1:0] node3034;
	wire [16-1:0] node3035;
	wire [16-1:0] node3036;
	wire [16-1:0] node3037;
	wire [16-1:0] node3038;
	wire [16-1:0] node3041;
	wire [16-1:0] node3044;
	wire [16-1:0] node3045;
	wire [16-1:0] node3048;
	wire [16-1:0] node3051;
	wire [16-1:0] node3052;
	wire [16-1:0] node3053;
	wire [16-1:0] node3056;
	wire [16-1:0] node3059;
	wire [16-1:0] node3060;
	wire [16-1:0] node3063;
	wire [16-1:0] node3066;
	wire [16-1:0] node3067;
	wire [16-1:0] node3068;
	wire [16-1:0] node3069;
	wire [16-1:0] node3072;
	wire [16-1:0] node3075;
	wire [16-1:0] node3076;
	wire [16-1:0] node3079;
	wire [16-1:0] node3082;
	wire [16-1:0] node3083;
	wire [16-1:0] node3084;
	wire [16-1:0] node3087;
	wire [16-1:0] node3090;
	wire [16-1:0] node3091;
	wire [16-1:0] node3095;
	wire [16-1:0] node3096;
	wire [16-1:0] node3097;
	wire [16-1:0] node3098;
	wire [16-1:0] node3099;
	wire [16-1:0] node3102;
	wire [16-1:0] node3105;
	wire [16-1:0] node3106;
	wire [16-1:0] node3109;
	wire [16-1:0] node3112;
	wire [16-1:0] node3113;
	wire [16-1:0] node3114;
	wire [16-1:0] node3117;
	wire [16-1:0] node3120;
	wire [16-1:0] node3121;
	wire [16-1:0] node3124;
	wire [16-1:0] node3127;
	wire [16-1:0] node3128;
	wire [16-1:0] node3129;
	wire [16-1:0] node3131;
	wire [16-1:0] node3134;
	wire [16-1:0] node3136;
	wire [16-1:0] node3139;
	wire [16-1:0] node3140;
	wire [16-1:0] node3141;
	wire [16-1:0] node3144;
	wire [16-1:0] node3147;
	wire [16-1:0] node3148;
	wire [16-1:0] node3151;
	wire [16-1:0] node3154;
	wire [16-1:0] node3155;
	wire [16-1:0] node3156;
	wire [16-1:0] node3157;
	wire [16-1:0] node3158;
	wire [16-1:0] node3159;
	wire [16-1:0] node3160;
	wire [16-1:0] node3163;
	wire [16-1:0] node3166;
	wire [16-1:0] node3167;
	wire [16-1:0] node3170;
	wire [16-1:0] node3173;
	wire [16-1:0] node3174;
	wire [16-1:0] node3175;
	wire [16-1:0] node3178;
	wire [16-1:0] node3181;
	wire [16-1:0] node3182;
	wire [16-1:0] node3185;
	wire [16-1:0] node3188;
	wire [16-1:0] node3189;
	wire [16-1:0] node3190;
	wire [16-1:0] node3191;
	wire [16-1:0] node3194;
	wire [16-1:0] node3197;
	wire [16-1:0] node3198;
	wire [16-1:0] node3201;
	wire [16-1:0] node3204;
	wire [16-1:0] node3205;
	wire [16-1:0] node3206;
	wire [16-1:0] node3209;
	wire [16-1:0] node3212;
	wire [16-1:0] node3214;
	wire [16-1:0] node3217;
	wire [16-1:0] node3218;
	wire [16-1:0] node3219;
	wire [16-1:0] node3220;
	wire [16-1:0] node3221;
	wire [16-1:0] node3224;
	wire [16-1:0] node3227;
	wire [16-1:0] node3228;
	wire [16-1:0] node3231;
	wire [16-1:0] node3234;
	wire [16-1:0] node3235;
	wire [16-1:0] node3236;
	wire [16-1:0] node3239;
	wire [16-1:0] node3242;
	wire [16-1:0] node3243;
	wire [16-1:0] node3246;
	wire [16-1:0] node3249;
	wire [16-1:0] node3250;
	wire [16-1:0] node3251;
	wire [16-1:0] node3252;
	wire [16-1:0] node3255;
	wire [16-1:0] node3258;
	wire [16-1:0] node3259;
	wire [16-1:0] node3262;
	wire [16-1:0] node3265;
	wire [16-1:0] node3266;
	wire [16-1:0] node3267;
	wire [16-1:0] node3270;
	wire [16-1:0] node3273;
	wire [16-1:0] node3274;
	wire [16-1:0] node3277;
	wire [16-1:0] node3280;
	wire [16-1:0] node3281;
	wire [16-1:0] node3282;
	wire [16-1:0] node3283;
	wire [16-1:0] node3284;
	wire [16-1:0] node3285;
	wire [16-1:0] node3288;
	wire [16-1:0] node3291;
	wire [16-1:0] node3292;
	wire [16-1:0] node3295;
	wire [16-1:0] node3298;
	wire [16-1:0] node3299;
	wire [16-1:0] node3300;
	wire [16-1:0] node3303;
	wire [16-1:0] node3306;
	wire [16-1:0] node3307;
	wire [16-1:0] node3310;
	wire [16-1:0] node3313;
	wire [16-1:0] node3314;
	wire [16-1:0] node3315;
	wire [16-1:0] node3316;
	wire [16-1:0] node3319;
	wire [16-1:0] node3322;
	wire [16-1:0] node3323;
	wire [16-1:0] node3326;
	wire [16-1:0] node3329;
	wire [16-1:0] node3330;
	wire [16-1:0] node3331;
	wire [16-1:0] node3334;
	wire [16-1:0] node3337;
	wire [16-1:0] node3338;
	wire [16-1:0] node3341;
	wire [16-1:0] node3344;
	wire [16-1:0] node3345;
	wire [16-1:0] node3346;
	wire [16-1:0] node3347;
	wire [16-1:0] node3348;
	wire [16-1:0] node3351;
	wire [16-1:0] node3354;
	wire [16-1:0] node3355;
	wire [16-1:0] node3358;
	wire [16-1:0] node3361;
	wire [16-1:0] node3362;
	wire [16-1:0] node3364;
	wire [16-1:0] node3367;
	wire [16-1:0] node3368;
	wire [16-1:0] node3372;
	wire [16-1:0] node3373;
	wire [16-1:0] node3374;
	wire [16-1:0] node3375;
	wire [16-1:0] node3378;
	wire [16-1:0] node3381;
	wire [16-1:0] node3382;
	wire [16-1:0] node3385;
	wire [16-1:0] node3388;
	wire [16-1:0] node3389;
	wire [16-1:0] node3390;
	wire [16-1:0] node3393;
	wire [16-1:0] node3396;
	wire [16-1:0] node3397;
	wire [16-1:0] node3400;
	wire [16-1:0] node3403;
	wire [16-1:0] node3404;
	wire [16-1:0] node3405;
	wire [16-1:0] node3406;
	wire [16-1:0] node3407;
	wire [16-1:0] node3408;
	wire [16-1:0] node3409;
	wire [16-1:0] node3410;
	wire [16-1:0] node3413;
	wire [16-1:0] node3416;
	wire [16-1:0] node3417;
	wire [16-1:0] node3420;
	wire [16-1:0] node3423;
	wire [16-1:0] node3424;
	wire [16-1:0] node3425;
	wire [16-1:0] node3428;
	wire [16-1:0] node3431;
	wire [16-1:0] node3432;
	wire [16-1:0] node3436;
	wire [16-1:0] node3437;
	wire [16-1:0] node3438;
	wire [16-1:0] node3439;
	wire [16-1:0] node3442;
	wire [16-1:0] node3445;
	wire [16-1:0] node3446;
	wire [16-1:0] node3450;
	wire [16-1:0] node3451;
	wire [16-1:0] node3452;
	wire [16-1:0] node3455;
	wire [16-1:0] node3458;
	wire [16-1:0] node3459;
	wire [16-1:0] node3462;
	wire [16-1:0] node3465;
	wire [16-1:0] node3466;
	wire [16-1:0] node3467;
	wire [16-1:0] node3468;
	wire [16-1:0] node3469;
	wire [16-1:0] node3472;
	wire [16-1:0] node3475;
	wire [16-1:0] node3476;
	wire [16-1:0] node3479;
	wire [16-1:0] node3482;
	wire [16-1:0] node3483;
	wire [16-1:0] node3484;
	wire [16-1:0] node3487;
	wire [16-1:0] node3490;
	wire [16-1:0] node3491;
	wire [16-1:0] node3494;
	wire [16-1:0] node3497;
	wire [16-1:0] node3498;
	wire [16-1:0] node3499;
	wire [16-1:0] node3500;
	wire [16-1:0] node3503;
	wire [16-1:0] node3506;
	wire [16-1:0] node3507;
	wire [16-1:0] node3510;
	wire [16-1:0] node3513;
	wire [16-1:0] node3514;
	wire [16-1:0] node3515;
	wire [16-1:0] node3519;
	wire [16-1:0] node3520;
	wire [16-1:0] node3523;
	wire [16-1:0] node3526;
	wire [16-1:0] node3527;
	wire [16-1:0] node3528;
	wire [16-1:0] node3529;
	wire [16-1:0] node3530;
	wire [16-1:0] node3531;
	wire [16-1:0] node3534;
	wire [16-1:0] node3537;
	wire [16-1:0] node3538;
	wire [16-1:0] node3541;
	wire [16-1:0] node3544;
	wire [16-1:0] node3545;
	wire [16-1:0] node3546;
	wire [16-1:0] node3549;
	wire [16-1:0] node3552;
	wire [16-1:0] node3553;
	wire [16-1:0] node3556;
	wire [16-1:0] node3559;
	wire [16-1:0] node3560;
	wire [16-1:0] node3561;
	wire [16-1:0] node3562;
	wire [16-1:0] node3565;
	wire [16-1:0] node3568;
	wire [16-1:0] node3569;
	wire [16-1:0] node3572;
	wire [16-1:0] node3575;
	wire [16-1:0] node3576;
	wire [16-1:0] node3578;
	wire [16-1:0] node3581;
	wire [16-1:0] node3582;
	wire [16-1:0] node3585;
	wire [16-1:0] node3588;
	wire [16-1:0] node3589;
	wire [16-1:0] node3590;
	wire [16-1:0] node3591;
	wire [16-1:0] node3592;
	wire [16-1:0] node3595;
	wire [16-1:0] node3598;
	wire [16-1:0] node3599;
	wire [16-1:0] node3602;
	wire [16-1:0] node3605;
	wire [16-1:0] node3606;
	wire [16-1:0] node3607;
	wire [16-1:0] node3610;
	wire [16-1:0] node3613;
	wire [16-1:0] node3616;
	wire [16-1:0] node3617;
	wire [16-1:0] node3618;
	wire [16-1:0] node3619;
	wire [16-1:0] node3622;
	wire [16-1:0] node3625;
	wire [16-1:0] node3626;
	wire [16-1:0] node3629;
	wire [16-1:0] node3632;
	wire [16-1:0] node3633;
	wire [16-1:0] node3635;
	wire [16-1:0] node3638;
	wire [16-1:0] node3639;
	wire [16-1:0] node3642;
	wire [16-1:0] node3645;
	wire [16-1:0] node3646;
	wire [16-1:0] node3647;
	wire [16-1:0] node3648;
	wire [16-1:0] node3649;
	wire [16-1:0] node3650;
	wire [16-1:0] node3651;
	wire [16-1:0] node3654;
	wire [16-1:0] node3657;
	wire [16-1:0] node3658;
	wire [16-1:0] node3662;
	wire [16-1:0] node3663;
	wire [16-1:0] node3664;
	wire [16-1:0] node3667;
	wire [16-1:0] node3670;
	wire [16-1:0] node3671;
	wire [16-1:0] node3674;
	wire [16-1:0] node3677;
	wire [16-1:0] node3678;
	wire [16-1:0] node3679;
	wire [16-1:0] node3680;
	wire [16-1:0] node3683;
	wire [16-1:0] node3686;
	wire [16-1:0] node3687;
	wire [16-1:0] node3690;
	wire [16-1:0] node3693;
	wire [16-1:0] node3694;
	wire [16-1:0] node3695;
	wire [16-1:0] node3698;
	wire [16-1:0] node3701;
	wire [16-1:0] node3702;
	wire [16-1:0] node3705;
	wire [16-1:0] node3708;
	wire [16-1:0] node3709;
	wire [16-1:0] node3710;
	wire [16-1:0] node3711;
	wire [16-1:0] node3712;
	wire [16-1:0] node3715;
	wire [16-1:0] node3718;
	wire [16-1:0] node3719;
	wire [16-1:0] node3722;
	wire [16-1:0] node3725;
	wire [16-1:0] node3726;
	wire [16-1:0] node3727;
	wire [16-1:0] node3730;
	wire [16-1:0] node3733;
	wire [16-1:0] node3734;
	wire [16-1:0] node3737;
	wire [16-1:0] node3740;
	wire [16-1:0] node3741;
	wire [16-1:0] node3742;
	wire [16-1:0] node3743;
	wire [16-1:0] node3746;
	wire [16-1:0] node3749;
	wire [16-1:0] node3750;
	wire [16-1:0] node3753;
	wire [16-1:0] node3756;
	wire [16-1:0] node3757;
	wire [16-1:0] node3758;
	wire [16-1:0] node3761;
	wire [16-1:0] node3764;
	wire [16-1:0] node3765;
	wire [16-1:0] node3768;
	wire [16-1:0] node3771;
	wire [16-1:0] node3772;
	wire [16-1:0] node3773;
	wire [16-1:0] node3774;
	wire [16-1:0] node3775;
	wire [16-1:0] node3776;
	wire [16-1:0] node3780;
	wire [16-1:0] node3781;
	wire [16-1:0] node3784;
	wire [16-1:0] node3787;
	wire [16-1:0] node3788;
	wire [16-1:0] node3789;
	wire [16-1:0] node3792;
	wire [16-1:0] node3795;
	wire [16-1:0] node3796;
	wire [16-1:0] node3800;
	wire [16-1:0] node3801;
	wire [16-1:0] node3802;
	wire [16-1:0] node3803;
	wire [16-1:0] node3806;
	wire [16-1:0] node3809;
	wire [16-1:0] node3810;
	wire [16-1:0] node3813;
	wire [16-1:0] node3816;
	wire [16-1:0] node3817;
	wire [16-1:0] node3818;
	wire [16-1:0] node3821;
	wire [16-1:0] node3824;
	wire [16-1:0] node3825;
	wire [16-1:0] node3828;
	wire [16-1:0] node3831;
	wire [16-1:0] node3832;
	wire [16-1:0] node3833;
	wire [16-1:0] node3834;
	wire [16-1:0] node3836;
	wire [16-1:0] node3839;
	wire [16-1:0] node3841;
	wire [16-1:0] node3844;
	wire [16-1:0] node3845;
	wire [16-1:0] node3846;
	wire [16-1:0] node3849;
	wire [16-1:0] node3852;
	wire [16-1:0] node3853;
	wire [16-1:0] node3856;
	wire [16-1:0] node3859;
	wire [16-1:0] node3860;
	wire [16-1:0] node3861;
	wire [16-1:0] node3863;
	wire [16-1:0] node3866;
	wire [16-1:0] node3867;
	wire [16-1:0] node3870;
	wire [16-1:0] node3873;
	wire [16-1:0] node3874;
	wire [16-1:0] node3875;
	wire [16-1:0] node3878;
	wire [16-1:0] node3881;
	wire [16-1:0] node3882;
	wire [16-1:0] node3885;
	wire [16-1:0] node3888;
	wire [16-1:0] node3889;
	wire [16-1:0] node3890;
	wire [16-1:0] node3891;
	wire [16-1:0] node3892;
	wire [16-1:0] node3893;
	wire [16-1:0] node3894;
	wire [16-1:0] node3895;
	wire [16-1:0] node3896;
	wire [16-1:0] node3897;
	wire [16-1:0] node3898;
	wire [16-1:0] node3901;
	wire [16-1:0] node3904;
	wire [16-1:0] node3905;
	wire [16-1:0] node3908;
	wire [16-1:0] node3911;
	wire [16-1:0] node3912;
	wire [16-1:0] node3913;
	wire [16-1:0] node3916;
	wire [16-1:0] node3919;
	wire [16-1:0] node3920;
	wire [16-1:0] node3923;
	wire [16-1:0] node3926;
	wire [16-1:0] node3927;
	wire [16-1:0] node3928;
	wire [16-1:0] node3929;
	wire [16-1:0] node3932;
	wire [16-1:0] node3935;
	wire [16-1:0] node3936;
	wire [16-1:0] node3940;
	wire [16-1:0] node3941;
	wire [16-1:0] node3943;
	wire [16-1:0] node3946;
	wire [16-1:0] node3947;
	wire [16-1:0] node3950;
	wire [16-1:0] node3953;
	wire [16-1:0] node3954;
	wire [16-1:0] node3955;
	wire [16-1:0] node3956;
	wire [16-1:0] node3957;
	wire [16-1:0] node3960;
	wire [16-1:0] node3963;
	wire [16-1:0] node3964;
	wire [16-1:0] node3967;
	wire [16-1:0] node3970;
	wire [16-1:0] node3971;
	wire [16-1:0] node3972;
	wire [16-1:0] node3975;
	wire [16-1:0] node3978;
	wire [16-1:0] node3979;
	wire [16-1:0] node3982;
	wire [16-1:0] node3985;
	wire [16-1:0] node3986;
	wire [16-1:0] node3987;
	wire [16-1:0] node3988;
	wire [16-1:0] node3991;
	wire [16-1:0] node3994;
	wire [16-1:0] node3995;
	wire [16-1:0] node3998;
	wire [16-1:0] node4001;
	wire [16-1:0] node4002;
	wire [16-1:0] node4003;
	wire [16-1:0] node4006;
	wire [16-1:0] node4009;
	wire [16-1:0] node4010;
	wire [16-1:0] node4014;
	wire [16-1:0] node4015;
	wire [16-1:0] node4016;
	wire [16-1:0] node4017;
	wire [16-1:0] node4018;
	wire [16-1:0] node4019;
	wire [16-1:0] node4022;
	wire [16-1:0] node4025;
	wire [16-1:0] node4026;
	wire [16-1:0] node4029;
	wire [16-1:0] node4032;
	wire [16-1:0] node4033;
	wire [16-1:0] node4034;
	wire [16-1:0] node4037;
	wire [16-1:0] node4040;
	wire [16-1:0] node4041;
	wire [16-1:0] node4044;
	wire [16-1:0] node4047;
	wire [16-1:0] node4048;
	wire [16-1:0] node4049;
	wire [16-1:0] node4050;
	wire [16-1:0] node4054;
	wire [16-1:0] node4055;
	wire [16-1:0] node4058;
	wire [16-1:0] node4061;
	wire [16-1:0] node4062;
	wire [16-1:0] node4063;
	wire [16-1:0] node4066;
	wire [16-1:0] node4069;
	wire [16-1:0] node4070;
	wire [16-1:0] node4073;
	wire [16-1:0] node4076;
	wire [16-1:0] node4077;
	wire [16-1:0] node4078;
	wire [16-1:0] node4079;
	wire [16-1:0] node4080;
	wire [16-1:0] node4083;
	wire [16-1:0] node4086;
	wire [16-1:0] node4087;
	wire [16-1:0] node4090;
	wire [16-1:0] node4093;
	wire [16-1:0] node4094;
	wire [16-1:0] node4095;
	wire [16-1:0] node4098;
	wire [16-1:0] node4101;
	wire [16-1:0] node4102;
	wire [16-1:0] node4105;
	wire [16-1:0] node4108;
	wire [16-1:0] node4109;
	wire [16-1:0] node4110;
	wire [16-1:0] node4111;
	wire [16-1:0] node4115;
	wire [16-1:0] node4116;
	wire [16-1:0] node4119;
	wire [16-1:0] node4122;
	wire [16-1:0] node4123;
	wire [16-1:0] node4124;
	wire [16-1:0] node4127;
	wire [16-1:0] node4130;
	wire [16-1:0] node4131;
	wire [16-1:0] node4134;
	wire [16-1:0] node4137;
	wire [16-1:0] node4138;
	wire [16-1:0] node4139;
	wire [16-1:0] node4140;
	wire [16-1:0] node4141;
	wire [16-1:0] node4142;
	wire [16-1:0] node4143;
	wire [16-1:0] node4146;
	wire [16-1:0] node4149;
	wire [16-1:0] node4150;
	wire [16-1:0] node4153;
	wire [16-1:0] node4156;
	wire [16-1:0] node4157;
	wire [16-1:0] node4158;
	wire [16-1:0] node4161;
	wire [16-1:0] node4164;
	wire [16-1:0] node4165;
	wire [16-1:0] node4168;
	wire [16-1:0] node4171;
	wire [16-1:0] node4172;
	wire [16-1:0] node4173;
	wire [16-1:0] node4174;
	wire [16-1:0] node4177;
	wire [16-1:0] node4180;
	wire [16-1:0] node4181;
	wire [16-1:0] node4184;
	wire [16-1:0] node4187;
	wire [16-1:0] node4188;
	wire [16-1:0] node4189;
	wire [16-1:0] node4192;
	wire [16-1:0] node4195;
	wire [16-1:0] node4196;
	wire [16-1:0] node4199;
	wire [16-1:0] node4202;
	wire [16-1:0] node4203;
	wire [16-1:0] node4204;
	wire [16-1:0] node4205;
	wire [16-1:0] node4206;
	wire [16-1:0] node4209;
	wire [16-1:0] node4212;
	wire [16-1:0] node4213;
	wire [16-1:0] node4217;
	wire [16-1:0] node4218;
	wire [16-1:0] node4219;
	wire [16-1:0] node4222;
	wire [16-1:0] node4225;
	wire [16-1:0] node4226;
	wire [16-1:0] node4229;
	wire [16-1:0] node4232;
	wire [16-1:0] node4233;
	wire [16-1:0] node4234;
	wire [16-1:0] node4235;
	wire [16-1:0] node4238;
	wire [16-1:0] node4241;
	wire [16-1:0] node4242;
	wire [16-1:0] node4245;
	wire [16-1:0] node4248;
	wire [16-1:0] node4249;
	wire [16-1:0] node4250;
	wire [16-1:0] node4253;
	wire [16-1:0] node4256;
	wire [16-1:0] node4257;
	wire [16-1:0] node4260;
	wire [16-1:0] node4263;
	wire [16-1:0] node4264;
	wire [16-1:0] node4265;
	wire [16-1:0] node4266;
	wire [16-1:0] node4267;
	wire [16-1:0] node4268;
	wire [16-1:0] node4271;
	wire [16-1:0] node4274;
	wire [16-1:0] node4275;
	wire [16-1:0] node4278;
	wire [16-1:0] node4281;
	wire [16-1:0] node4282;
	wire [16-1:0] node4283;
	wire [16-1:0] node4286;
	wire [16-1:0] node4289;
	wire [16-1:0] node4290;
	wire [16-1:0] node4293;
	wire [16-1:0] node4296;
	wire [16-1:0] node4297;
	wire [16-1:0] node4298;
	wire [16-1:0] node4299;
	wire [16-1:0] node4302;
	wire [16-1:0] node4305;
	wire [16-1:0] node4306;
	wire [16-1:0] node4309;
	wire [16-1:0] node4312;
	wire [16-1:0] node4313;
	wire [16-1:0] node4315;
	wire [16-1:0] node4318;
	wire [16-1:0] node4319;
	wire [16-1:0] node4322;
	wire [16-1:0] node4325;
	wire [16-1:0] node4326;
	wire [16-1:0] node4327;
	wire [16-1:0] node4328;
	wire [16-1:0] node4330;
	wire [16-1:0] node4333;
	wire [16-1:0] node4334;
	wire [16-1:0] node4337;
	wire [16-1:0] node4340;
	wire [16-1:0] node4341;
	wire [16-1:0] node4342;
	wire [16-1:0] node4345;
	wire [16-1:0] node4348;
	wire [16-1:0] node4349;
	wire [16-1:0] node4352;
	wire [16-1:0] node4355;
	wire [16-1:0] node4356;
	wire [16-1:0] node4357;
	wire [16-1:0] node4358;
	wire [16-1:0] node4361;
	wire [16-1:0] node4364;
	wire [16-1:0] node4365;
	wire [16-1:0] node4368;
	wire [16-1:0] node4371;
	wire [16-1:0] node4372;
	wire [16-1:0] node4373;
	wire [16-1:0] node4376;
	wire [16-1:0] node4379;
	wire [16-1:0] node4380;
	wire [16-1:0] node4383;
	wire [16-1:0] node4386;
	wire [16-1:0] node4387;
	wire [16-1:0] node4388;
	wire [16-1:0] node4389;
	wire [16-1:0] node4390;
	wire [16-1:0] node4391;
	wire [16-1:0] node4392;
	wire [16-1:0] node4393;
	wire [16-1:0] node4396;
	wire [16-1:0] node4399;
	wire [16-1:0] node4400;
	wire [16-1:0] node4403;
	wire [16-1:0] node4406;
	wire [16-1:0] node4407;
	wire [16-1:0] node4408;
	wire [16-1:0] node4411;
	wire [16-1:0] node4414;
	wire [16-1:0] node4415;
	wire [16-1:0] node4418;
	wire [16-1:0] node4421;
	wire [16-1:0] node4422;
	wire [16-1:0] node4423;
	wire [16-1:0] node4424;
	wire [16-1:0] node4427;
	wire [16-1:0] node4430;
	wire [16-1:0] node4431;
	wire [16-1:0] node4434;
	wire [16-1:0] node4437;
	wire [16-1:0] node4438;
	wire [16-1:0] node4440;
	wire [16-1:0] node4443;
	wire [16-1:0] node4444;
	wire [16-1:0] node4447;
	wire [16-1:0] node4450;
	wire [16-1:0] node4451;
	wire [16-1:0] node4452;
	wire [16-1:0] node4453;
	wire [16-1:0] node4454;
	wire [16-1:0] node4458;
	wire [16-1:0] node4459;
	wire [16-1:0] node4463;
	wire [16-1:0] node4464;
	wire [16-1:0] node4465;
	wire [16-1:0] node4468;
	wire [16-1:0] node4471;
	wire [16-1:0] node4472;
	wire [16-1:0] node4475;
	wire [16-1:0] node4478;
	wire [16-1:0] node4479;
	wire [16-1:0] node4480;
	wire [16-1:0] node4481;
	wire [16-1:0] node4484;
	wire [16-1:0] node4487;
	wire [16-1:0] node4488;
	wire [16-1:0] node4491;
	wire [16-1:0] node4494;
	wire [16-1:0] node4495;
	wire [16-1:0] node4496;
	wire [16-1:0] node4499;
	wire [16-1:0] node4502;
	wire [16-1:0] node4503;
	wire [16-1:0] node4506;
	wire [16-1:0] node4509;
	wire [16-1:0] node4510;
	wire [16-1:0] node4511;
	wire [16-1:0] node4512;
	wire [16-1:0] node4513;
	wire [16-1:0] node4514;
	wire [16-1:0] node4517;
	wire [16-1:0] node4520;
	wire [16-1:0] node4521;
	wire [16-1:0] node4524;
	wire [16-1:0] node4527;
	wire [16-1:0] node4528;
	wire [16-1:0] node4529;
	wire [16-1:0] node4532;
	wire [16-1:0] node4535;
	wire [16-1:0] node4536;
	wire [16-1:0] node4539;
	wire [16-1:0] node4542;
	wire [16-1:0] node4543;
	wire [16-1:0] node4544;
	wire [16-1:0] node4545;
	wire [16-1:0] node4548;
	wire [16-1:0] node4551;
	wire [16-1:0] node4552;
	wire [16-1:0] node4555;
	wire [16-1:0] node4558;
	wire [16-1:0] node4559;
	wire [16-1:0] node4560;
	wire [16-1:0] node4563;
	wire [16-1:0] node4566;
	wire [16-1:0] node4567;
	wire [16-1:0] node4570;
	wire [16-1:0] node4573;
	wire [16-1:0] node4574;
	wire [16-1:0] node4575;
	wire [16-1:0] node4576;
	wire [16-1:0] node4577;
	wire [16-1:0] node4580;
	wire [16-1:0] node4583;
	wire [16-1:0] node4584;
	wire [16-1:0] node4588;
	wire [16-1:0] node4589;
	wire [16-1:0] node4590;
	wire [16-1:0] node4593;
	wire [16-1:0] node4596;
	wire [16-1:0] node4597;
	wire [16-1:0] node4600;
	wire [16-1:0] node4603;
	wire [16-1:0] node4604;
	wire [16-1:0] node4605;
	wire [16-1:0] node4606;
	wire [16-1:0] node4609;
	wire [16-1:0] node4612;
	wire [16-1:0] node4613;
	wire [16-1:0] node4616;
	wire [16-1:0] node4619;
	wire [16-1:0] node4620;
	wire [16-1:0] node4621;
	wire [16-1:0] node4624;
	wire [16-1:0] node4627;
	wire [16-1:0] node4628;
	wire [16-1:0] node4631;
	wire [16-1:0] node4634;
	wire [16-1:0] node4635;
	wire [16-1:0] node4636;
	wire [16-1:0] node4637;
	wire [16-1:0] node4638;
	wire [16-1:0] node4639;
	wire [16-1:0] node4641;
	wire [16-1:0] node4644;
	wire [16-1:0] node4645;
	wire [16-1:0] node4649;
	wire [16-1:0] node4650;
	wire [16-1:0] node4651;
	wire [16-1:0] node4654;
	wire [16-1:0] node4657;
	wire [16-1:0] node4658;
	wire [16-1:0] node4661;
	wire [16-1:0] node4664;
	wire [16-1:0] node4665;
	wire [16-1:0] node4666;
	wire [16-1:0] node4667;
	wire [16-1:0] node4670;
	wire [16-1:0] node4673;
	wire [16-1:0] node4674;
	wire [16-1:0] node4677;
	wire [16-1:0] node4680;
	wire [16-1:0] node4681;
	wire [16-1:0] node4682;
	wire [16-1:0] node4685;
	wire [16-1:0] node4688;
	wire [16-1:0] node4689;
	wire [16-1:0] node4692;
	wire [16-1:0] node4695;
	wire [16-1:0] node4696;
	wire [16-1:0] node4697;
	wire [16-1:0] node4698;
	wire [16-1:0] node4699;
	wire [16-1:0] node4702;
	wire [16-1:0] node4705;
	wire [16-1:0] node4706;
	wire [16-1:0] node4710;
	wire [16-1:0] node4711;
	wire [16-1:0] node4713;
	wire [16-1:0] node4716;
	wire [16-1:0] node4717;
	wire [16-1:0] node4720;
	wire [16-1:0] node4723;
	wire [16-1:0] node4724;
	wire [16-1:0] node4725;
	wire [16-1:0] node4726;
	wire [16-1:0] node4729;
	wire [16-1:0] node4732;
	wire [16-1:0] node4733;
	wire [16-1:0] node4736;
	wire [16-1:0] node4739;
	wire [16-1:0] node4740;
	wire [16-1:0] node4741;
	wire [16-1:0] node4744;
	wire [16-1:0] node4747;
	wire [16-1:0] node4748;
	wire [16-1:0] node4751;
	wire [16-1:0] node4754;
	wire [16-1:0] node4755;
	wire [16-1:0] node4756;
	wire [16-1:0] node4757;
	wire [16-1:0] node4758;
	wire [16-1:0] node4759;
	wire [16-1:0] node4762;
	wire [16-1:0] node4765;
	wire [16-1:0] node4766;
	wire [16-1:0] node4769;
	wire [16-1:0] node4772;
	wire [16-1:0] node4773;
	wire [16-1:0] node4774;
	wire [16-1:0] node4777;
	wire [16-1:0] node4780;
	wire [16-1:0] node4781;
	wire [16-1:0] node4784;
	wire [16-1:0] node4787;
	wire [16-1:0] node4788;
	wire [16-1:0] node4789;
	wire [16-1:0] node4790;
	wire [16-1:0] node4793;
	wire [16-1:0] node4796;
	wire [16-1:0] node4797;
	wire [16-1:0] node4800;
	wire [16-1:0] node4803;
	wire [16-1:0] node4804;
	wire [16-1:0] node4805;
	wire [16-1:0] node4808;
	wire [16-1:0] node4811;
	wire [16-1:0] node4812;
	wire [16-1:0] node4815;
	wire [16-1:0] node4818;
	wire [16-1:0] node4819;
	wire [16-1:0] node4820;
	wire [16-1:0] node4821;
	wire [16-1:0] node4822;
	wire [16-1:0] node4826;
	wire [16-1:0] node4827;
	wire [16-1:0] node4830;
	wire [16-1:0] node4833;
	wire [16-1:0] node4834;
	wire [16-1:0] node4835;
	wire [16-1:0] node4838;
	wire [16-1:0] node4841;
	wire [16-1:0] node4843;
	wire [16-1:0] node4846;
	wire [16-1:0] node4847;
	wire [16-1:0] node4848;
	wire [16-1:0] node4849;
	wire [16-1:0] node4852;
	wire [16-1:0] node4855;
	wire [16-1:0] node4856;
	wire [16-1:0] node4859;
	wire [16-1:0] node4862;
	wire [16-1:0] node4863;
	wire [16-1:0] node4864;
	wire [16-1:0] node4867;
	wire [16-1:0] node4870;
	wire [16-1:0] node4871;
	wire [16-1:0] node4874;
	wire [16-1:0] node4877;
	wire [16-1:0] node4878;
	wire [16-1:0] node4879;
	wire [16-1:0] node4880;
	wire [16-1:0] node4881;
	wire [16-1:0] node4882;
	wire [16-1:0] node4883;
	wire [16-1:0] node4884;
	wire [16-1:0] node4885;
	wire [16-1:0] node4888;
	wire [16-1:0] node4891;
	wire [16-1:0] node4892;
	wire [16-1:0] node4895;
	wire [16-1:0] node4898;
	wire [16-1:0] node4899;
	wire [16-1:0] node4901;
	wire [16-1:0] node4904;
	wire [16-1:0] node4905;
	wire [16-1:0] node4908;
	wire [16-1:0] node4911;
	wire [16-1:0] node4912;
	wire [16-1:0] node4913;
	wire [16-1:0] node4915;
	wire [16-1:0] node4918;
	wire [16-1:0] node4919;
	wire [16-1:0] node4922;
	wire [16-1:0] node4925;
	wire [16-1:0] node4926;
	wire [16-1:0] node4927;
	wire [16-1:0] node4930;
	wire [16-1:0] node4933;
	wire [16-1:0] node4934;
	wire [16-1:0] node4937;
	wire [16-1:0] node4940;
	wire [16-1:0] node4941;
	wire [16-1:0] node4942;
	wire [16-1:0] node4943;
	wire [16-1:0] node4944;
	wire [16-1:0] node4947;
	wire [16-1:0] node4950;
	wire [16-1:0] node4952;
	wire [16-1:0] node4955;
	wire [16-1:0] node4956;
	wire [16-1:0] node4957;
	wire [16-1:0] node4960;
	wire [16-1:0] node4963;
	wire [16-1:0] node4964;
	wire [16-1:0] node4967;
	wire [16-1:0] node4970;
	wire [16-1:0] node4971;
	wire [16-1:0] node4972;
	wire [16-1:0] node4973;
	wire [16-1:0] node4976;
	wire [16-1:0] node4979;
	wire [16-1:0] node4980;
	wire [16-1:0] node4983;
	wire [16-1:0] node4986;
	wire [16-1:0] node4987;
	wire [16-1:0] node4988;
	wire [16-1:0] node4991;
	wire [16-1:0] node4994;
	wire [16-1:0] node4995;
	wire [16-1:0] node4998;
	wire [16-1:0] node5001;
	wire [16-1:0] node5002;
	wire [16-1:0] node5003;
	wire [16-1:0] node5004;
	wire [16-1:0] node5005;
	wire [16-1:0] node5006;
	wire [16-1:0] node5009;
	wire [16-1:0] node5012;
	wire [16-1:0] node5013;
	wire [16-1:0] node5016;
	wire [16-1:0] node5019;
	wire [16-1:0] node5020;
	wire [16-1:0] node5021;
	wire [16-1:0] node5024;
	wire [16-1:0] node5027;
	wire [16-1:0] node5028;
	wire [16-1:0] node5031;
	wire [16-1:0] node5034;
	wire [16-1:0] node5035;
	wire [16-1:0] node5036;
	wire [16-1:0] node5037;
	wire [16-1:0] node5040;
	wire [16-1:0] node5043;
	wire [16-1:0] node5044;
	wire [16-1:0] node5047;
	wire [16-1:0] node5050;
	wire [16-1:0] node5051;
	wire [16-1:0] node5053;
	wire [16-1:0] node5056;
	wire [16-1:0] node5057;
	wire [16-1:0] node5060;
	wire [16-1:0] node5063;
	wire [16-1:0] node5064;
	wire [16-1:0] node5065;
	wire [16-1:0] node5066;
	wire [16-1:0] node5067;
	wire [16-1:0] node5070;
	wire [16-1:0] node5073;
	wire [16-1:0] node5074;
	wire [16-1:0] node5077;
	wire [16-1:0] node5080;
	wire [16-1:0] node5081;
	wire [16-1:0] node5082;
	wire [16-1:0] node5085;
	wire [16-1:0] node5088;
	wire [16-1:0] node5089;
	wire [16-1:0] node5092;
	wire [16-1:0] node5095;
	wire [16-1:0] node5096;
	wire [16-1:0] node5097;
	wire [16-1:0] node5099;
	wire [16-1:0] node5102;
	wire [16-1:0] node5103;
	wire [16-1:0] node5106;
	wire [16-1:0] node5109;
	wire [16-1:0] node5110;
	wire [16-1:0] node5111;
	wire [16-1:0] node5114;
	wire [16-1:0] node5117;
	wire [16-1:0] node5118;
	wire [16-1:0] node5121;
	wire [16-1:0] node5124;
	wire [16-1:0] node5125;
	wire [16-1:0] node5126;
	wire [16-1:0] node5127;
	wire [16-1:0] node5128;
	wire [16-1:0] node5129;
	wire [16-1:0] node5130;
	wire [16-1:0] node5133;
	wire [16-1:0] node5136;
	wire [16-1:0] node5137;
	wire [16-1:0] node5140;
	wire [16-1:0] node5143;
	wire [16-1:0] node5144;
	wire [16-1:0] node5145;
	wire [16-1:0] node5148;
	wire [16-1:0] node5151;
	wire [16-1:0] node5152;
	wire [16-1:0] node5156;
	wire [16-1:0] node5157;
	wire [16-1:0] node5158;
	wire [16-1:0] node5159;
	wire [16-1:0] node5162;
	wire [16-1:0] node5165;
	wire [16-1:0] node5166;
	wire [16-1:0] node5169;
	wire [16-1:0] node5172;
	wire [16-1:0] node5173;
	wire [16-1:0] node5174;
	wire [16-1:0] node5177;
	wire [16-1:0] node5180;
	wire [16-1:0] node5181;
	wire [16-1:0] node5184;
	wire [16-1:0] node5187;
	wire [16-1:0] node5188;
	wire [16-1:0] node5189;
	wire [16-1:0] node5190;
	wire [16-1:0] node5191;
	wire [16-1:0] node5194;
	wire [16-1:0] node5197;
	wire [16-1:0] node5198;
	wire [16-1:0] node5201;
	wire [16-1:0] node5204;
	wire [16-1:0] node5205;
	wire [16-1:0] node5206;
	wire [16-1:0] node5209;
	wire [16-1:0] node5212;
	wire [16-1:0] node5213;
	wire [16-1:0] node5216;
	wire [16-1:0] node5219;
	wire [16-1:0] node5220;
	wire [16-1:0] node5221;
	wire [16-1:0] node5223;
	wire [16-1:0] node5226;
	wire [16-1:0] node5227;
	wire [16-1:0] node5230;
	wire [16-1:0] node5233;
	wire [16-1:0] node5234;
	wire [16-1:0] node5235;
	wire [16-1:0] node5238;
	wire [16-1:0] node5241;
	wire [16-1:0] node5242;
	wire [16-1:0] node5246;
	wire [16-1:0] node5247;
	wire [16-1:0] node5248;
	wire [16-1:0] node5249;
	wire [16-1:0] node5250;
	wire [16-1:0] node5251;
	wire [16-1:0] node5255;
	wire [16-1:0] node5256;
	wire [16-1:0] node5259;
	wire [16-1:0] node5262;
	wire [16-1:0] node5263;
	wire [16-1:0] node5264;
	wire [16-1:0] node5267;
	wire [16-1:0] node5270;
	wire [16-1:0] node5271;
	wire [16-1:0] node5275;
	wire [16-1:0] node5276;
	wire [16-1:0] node5277;
	wire [16-1:0] node5278;
	wire [16-1:0] node5281;
	wire [16-1:0] node5284;
	wire [16-1:0] node5285;
	wire [16-1:0] node5288;
	wire [16-1:0] node5291;
	wire [16-1:0] node5292;
	wire [16-1:0] node5293;
	wire [16-1:0] node5296;
	wire [16-1:0] node5299;
	wire [16-1:0] node5300;
	wire [16-1:0] node5303;
	wire [16-1:0] node5306;
	wire [16-1:0] node5307;
	wire [16-1:0] node5308;
	wire [16-1:0] node5309;
	wire [16-1:0] node5311;
	wire [16-1:0] node5314;
	wire [16-1:0] node5315;
	wire [16-1:0] node5318;
	wire [16-1:0] node5321;
	wire [16-1:0] node5322;
	wire [16-1:0] node5323;
	wire [16-1:0] node5326;
	wire [16-1:0] node5329;
	wire [16-1:0] node5330;
	wire [16-1:0] node5333;
	wire [16-1:0] node5336;
	wire [16-1:0] node5337;
	wire [16-1:0] node5339;
	wire [16-1:0] node5341;
	wire [16-1:0] node5344;
	wire [16-1:0] node5345;
	wire [16-1:0] node5346;
	wire [16-1:0] node5349;
	wire [16-1:0] node5352;
	wire [16-1:0] node5353;
	wire [16-1:0] node5356;
	wire [16-1:0] node5359;
	wire [16-1:0] node5360;
	wire [16-1:0] node5361;
	wire [16-1:0] node5362;
	wire [16-1:0] node5363;
	wire [16-1:0] node5364;
	wire [16-1:0] node5365;
	wire [16-1:0] node5366;
	wire [16-1:0] node5369;
	wire [16-1:0] node5372;
	wire [16-1:0] node5373;
	wire [16-1:0] node5376;
	wire [16-1:0] node5379;
	wire [16-1:0] node5380;
	wire [16-1:0] node5381;
	wire [16-1:0] node5384;
	wire [16-1:0] node5387;
	wire [16-1:0] node5390;
	wire [16-1:0] node5391;
	wire [16-1:0] node5392;
	wire [16-1:0] node5393;
	wire [16-1:0] node5396;
	wire [16-1:0] node5399;
	wire [16-1:0] node5402;
	wire [16-1:0] node5403;
	wire [16-1:0] node5404;
	wire [16-1:0] node5407;
	wire [16-1:0] node5410;
	wire [16-1:0] node5412;
	wire [16-1:0] node5415;
	wire [16-1:0] node5416;
	wire [16-1:0] node5417;
	wire [16-1:0] node5418;
	wire [16-1:0] node5419;
	wire [16-1:0] node5422;
	wire [16-1:0] node5425;
	wire [16-1:0] node5426;
	wire [16-1:0] node5429;
	wire [16-1:0] node5432;
	wire [16-1:0] node5433;
	wire [16-1:0] node5434;
	wire [16-1:0] node5437;
	wire [16-1:0] node5440;
	wire [16-1:0] node5441;
	wire [16-1:0] node5444;
	wire [16-1:0] node5447;
	wire [16-1:0] node5448;
	wire [16-1:0] node5449;
	wire [16-1:0] node5450;
	wire [16-1:0] node5453;
	wire [16-1:0] node5456;
	wire [16-1:0] node5457;
	wire [16-1:0] node5460;
	wire [16-1:0] node5463;
	wire [16-1:0] node5464;
	wire [16-1:0] node5465;
	wire [16-1:0] node5468;
	wire [16-1:0] node5471;
	wire [16-1:0] node5472;
	wire [16-1:0] node5475;
	wire [16-1:0] node5478;
	wire [16-1:0] node5479;
	wire [16-1:0] node5480;
	wire [16-1:0] node5481;
	wire [16-1:0] node5482;
	wire [16-1:0] node5483;
	wire [16-1:0] node5486;
	wire [16-1:0] node5489;
	wire [16-1:0] node5490;
	wire [16-1:0] node5493;
	wire [16-1:0] node5496;
	wire [16-1:0] node5497;
	wire [16-1:0] node5498;
	wire [16-1:0] node5501;
	wire [16-1:0] node5504;
	wire [16-1:0] node5505;
	wire [16-1:0] node5508;
	wire [16-1:0] node5511;
	wire [16-1:0] node5512;
	wire [16-1:0] node5513;
	wire [16-1:0] node5514;
	wire [16-1:0] node5517;
	wire [16-1:0] node5520;
	wire [16-1:0] node5521;
	wire [16-1:0] node5524;
	wire [16-1:0] node5527;
	wire [16-1:0] node5528;
	wire [16-1:0] node5530;
	wire [16-1:0] node5533;
	wire [16-1:0] node5534;
	wire [16-1:0] node5537;
	wire [16-1:0] node5540;
	wire [16-1:0] node5541;
	wire [16-1:0] node5542;
	wire [16-1:0] node5543;
	wire [16-1:0] node5544;
	wire [16-1:0] node5547;
	wire [16-1:0] node5550;
	wire [16-1:0] node5551;
	wire [16-1:0] node5554;
	wire [16-1:0] node5557;
	wire [16-1:0] node5558;
	wire [16-1:0] node5559;
	wire [16-1:0] node5562;
	wire [16-1:0] node5565;
	wire [16-1:0] node5566;
	wire [16-1:0] node5569;
	wire [16-1:0] node5572;
	wire [16-1:0] node5573;
	wire [16-1:0] node5574;
	wire [16-1:0] node5576;
	wire [16-1:0] node5579;
	wire [16-1:0] node5580;
	wire [16-1:0] node5583;
	wire [16-1:0] node5586;
	wire [16-1:0] node5587;
	wire [16-1:0] node5588;
	wire [16-1:0] node5591;
	wire [16-1:0] node5594;
	wire [16-1:0] node5595;
	wire [16-1:0] node5598;
	wire [16-1:0] node5601;
	wire [16-1:0] node5602;
	wire [16-1:0] node5603;
	wire [16-1:0] node5604;
	wire [16-1:0] node5605;
	wire [16-1:0] node5606;
	wire [16-1:0] node5608;
	wire [16-1:0] node5611;
	wire [16-1:0] node5612;
	wire [16-1:0] node5615;
	wire [16-1:0] node5618;
	wire [16-1:0] node5619;
	wire [16-1:0] node5620;
	wire [16-1:0] node5623;
	wire [16-1:0] node5626;
	wire [16-1:0] node5628;
	wire [16-1:0] node5631;
	wire [16-1:0] node5632;
	wire [16-1:0] node5633;
	wire [16-1:0] node5634;
	wire [16-1:0] node5637;
	wire [16-1:0] node5640;
	wire [16-1:0] node5641;
	wire [16-1:0] node5644;
	wire [16-1:0] node5647;
	wire [16-1:0] node5648;
	wire [16-1:0] node5649;
	wire [16-1:0] node5652;
	wire [16-1:0] node5655;
	wire [16-1:0] node5656;
	wire [16-1:0] node5659;
	wire [16-1:0] node5662;
	wire [16-1:0] node5663;
	wire [16-1:0] node5664;
	wire [16-1:0] node5665;
	wire [16-1:0] node5666;
	wire [16-1:0] node5669;
	wire [16-1:0] node5672;
	wire [16-1:0] node5673;
	wire [16-1:0] node5676;
	wire [16-1:0] node5679;
	wire [16-1:0] node5680;
	wire [16-1:0] node5682;
	wire [16-1:0] node5685;
	wire [16-1:0] node5686;
	wire [16-1:0] node5689;
	wire [16-1:0] node5692;
	wire [16-1:0] node5693;
	wire [16-1:0] node5694;
	wire [16-1:0] node5695;
	wire [16-1:0] node5698;
	wire [16-1:0] node5701;
	wire [16-1:0] node5702;
	wire [16-1:0] node5705;
	wire [16-1:0] node5708;
	wire [16-1:0] node5709;
	wire [16-1:0] node5710;
	wire [16-1:0] node5713;
	wire [16-1:0] node5716;
	wire [16-1:0] node5717;
	wire [16-1:0] node5720;
	wire [16-1:0] node5723;
	wire [16-1:0] node5724;
	wire [16-1:0] node5725;
	wire [16-1:0] node5726;
	wire [16-1:0] node5727;
	wire [16-1:0] node5729;
	wire [16-1:0] node5732;
	wire [16-1:0] node5733;
	wire [16-1:0] node5736;
	wire [16-1:0] node5739;
	wire [16-1:0] node5740;
	wire [16-1:0] node5741;
	wire [16-1:0] node5744;
	wire [16-1:0] node5747;
	wire [16-1:0] node5748;
	wire [16-1:0] node5751;
	wire [16-1:0] node5754;
	wire [16-1:0] node5755;
	wire [16-1:0] node5756;
	wire [16-1:0] node5757;
	wire [16-1:0] node5761;
	wire [16-1:0] node5762;
	wire [16-1:0] node5765;
	wire [16-1:0] node5768;
	wire [16-1:0] node5769;
	wire [16-1:0] node5770;
	wire [16-1:0] node5773;
	wire [16-1:0] node5776;
	wire [16-1:0] node5777;
	wire [16-1:0] node5780;
	wire [16-1:0] node5783;
	wire [16-1:0] node5784;
	wire [16-1:0] node5785;
	wire [16-1:0] node5786;
	wire [16-1:0] node5787;
	wire [16-1:0] node5790;
	wire [16-1:0] node5793;
	wire [16-1:0] node5794;
	wire [16-1:0] node5797;
	wire [16-1:0] node5800;
	wire [16-1:0] node5801;
	wire [16-1:0] node5802;
	wire [16-1:0] node5805;
	wire [16-1:0] node5808;
	wire [16-1:0] node5809;
	wire [16-1:0] node5812;
	wire [16-1:0] node5815;
	wire [16-1:0] node5816;
	wire [16-1:0] node5817;
	wire [16-1:0] node5818;
	wire [16-1:0] node5821;
	wire [16-1:0] node5824;
	wire [16-1:0] node5825;
	wire [16-1:0] node5828;
	wire [16-1:0] node5831;
	wire [16-1:0] node5832;
	wire [16-1:0] node5833;
	wire [16-1:0] node5836;
	wire [16-1:0] node5839;
	wire [16-1:0] node5840;
	wire [16-1:0] node5843;
	wire [16-1:0] node5846;
	wire [16-1:0] node5847;
	wire [16-1:0] node5848;
	wire [16-1:0] node5849;
	wire [16-1:0] node5850;
	wire [16-1:0] node5851;
	wire [16-1:0] node5852;
	wire [16-1:0] node5853;
	wire [16-1:0] node5854;
	wire [16-1:0] node5855;
	wire [16-1:0] node5858;
	wire [16-1:0] node5861;
	wire [16-1:0] node5862;
	wire [16-1:0] node5865;
	wire [16-1:0] node5868;
	wire [16-1:0] node5869;
	wire [16-1:0] node5870;
	wire [16-1:0] node5873;
	wire [16-1:0] node5876;
	wire [16-1:0] node5877;
	wire [16-1:0] node5880;
	wire [16-1:0] node5883;
	wire [16-1:0] node5884;
	wire [16-1:0] node5885;
	wire [16-1:0] node5886;
	wire [16-1:0] node5889;
	wire [16-1:0] node5892;
	wire [16-1:0] node5893;
	wire [16-1:0] node5897;
	wire [16-1:0] node5898;
	wire [16-1:0] node5899;
	wire [16-1:0] node5902;
	wire [16-1:0] node5905;
	wire [16-1:0] node5906;
	wire [16-1:0] node5910;
	wire [16-1:0] node5911;
	wire [16-1:0] node5912;
	wire [16-1:0] node5913;
	wire [16-1:0] node5914;
	wire [16-1:0] node5918;
	wire [16-1:0] node5919;
	wire [16-1:0] node5922;
	wire [16-1:0] node5925;
	wire [16-1:0] node5926;
	wire [16-1:0] node5927;
	wire [16-1:0] node5930;
	wire [16-1:0] node5933;
	wire [16-1:0] node5934;
	wire [16-1:0] node5937;
	wire [16-1:0] node5940;
	wire [16-1:0] node5941;
	wire [16-1:0] node5942;
	wire [16-1:0] node5943;
	wire [16-1:0] node5947;
	wire [16-1:0] node5948;
	wire [16-1:0] node5951;
	wire [16-1:0] node5954;
	wire [16-1:0] node5955;
	wire [16-1:0] node5956;
	wire [16-1:0] node5959;
	wire [16-1:0] node5962;
	wire [16-1:0] node5963;
	wire [16-1:0] node5966;
	wire [16-1:0] node5969;
	wire [16-1:0] node5970;
	wire [16-1:0] node5971;
	wire [16-1:0] node5972;
	wire [16-1:0] node5973;
	wire [16-1:0] node5974;
	wire [16-1:0] node5977;
	wire [16-1:0] node5980;
	wire [16-1:0] node5981;
	wire [16-1:0] node5985;
	wire [16-1:0] node5986;
	wire [16-1:0] node5987;
	wire [16-1:0] node5990;
	wire [16-1:0] node5993;
	wire [16-1:0] node5994;
	wire [16-1:0] node5997;
	wire [16-1:0] node6000;
	wire [16-1:0] node6001;
	wire [16-1:0] node6002;
	wire [16-1:0] node6003;
	wire [16-1:0] node6006;
	wire [16-1:0] node6009;
	wire [16-1:0] node6011;
	wire [16-1:0] node6014;
	wire [16-1:0] node6015;
	wire [16-1:0] node6016;
	wire [16-1:0] node6020;
	wire [16-1:0] node6021;
	wire [16-1:0] node6024;
	wire [16-1:0] node6027;
	wire [16-1:0] node6028;
	wire [16-1:0] node6029;
	wire [16-1:0] node6030;
	wire [16-1:0] node6031;
	wire [16-1:0] node6034;
	wire [16-1:0] node6037;
	wire [16-1:0] node6038;
	wire [16-1:0] node6041;
	wire [16-1:0] node6044;
	wire [16-1:0] node6045;
	wire [16-1:0] node6046;
	wire [16-1:0] node6049;
	wire [16-1:0] node6052;
	wire [16-1:0] node6053;
	wire [16-1:0] node6057;
	wire [16-1:0] node6058;
	wire [16-1:0] node6059;
	wire [16-1:0] node6060;
	wire [16-1:0] node6063;
	wire [16-1:0] node6066;
	wire [16-1:0] node6067;
	wire [16-1:0] node6070;
	wire [16-1:0] node6073;
	wire [16-1:0] node6074;
	wire [16-1:0] node6075;
	wire [16-1:0] node6078;
	wire [16-1:0] node6081;
	wire [16-1:0] node6082;
	wire [16-1:0] node6086;
	wire [16-1:0] node6087;
	wire [16-1:0] node6088;
	wire [16-1:0] node6089;
	wire [16-1:0] node6090;
	wire [16-1:0] node6091;
	wire [16-1:0] node6092;
	wire [16-1:0] node6095;
	wire [16-1:0] node6098;
	wire [16-1:0] node6099;
	wire [16-1:0] node6103;
	wire [16-1:0] node6104;
	wire [16-1:0] node6105;
	wire [16-1:0] node6108;
	wire [16-1:0] node6111;
	wire [16-1:0] node6112;
	wire [16-1:0] node6115;
	wire [16-1:0] node6118;
	wire [16-1:0] node6119;
	wire [16-1:0] node6120;
	wire [16-1:0] node6121;
	wire [16-1:0] node6125;
	wire [16-1:0] node6126;
	wire [16-1:0] node6129;
	wire [16-1:0] node6132;
	wire [16-1:0] node6133;
	wire [16-1:0] node6134;
	wire [16-1:0] node6137;
	wire [16-1:0] node6140;
	wire [16-1:0] node6141;
	wire [16-1:0] node6144;
	wire [16-1:0] node6147;
	wire [16-1:0] node6148;
	wire [16-1:0] node6149;
	wire [16-1:0] node6150;
	wire [16-1:0] node6151;
	wire [16-1:0] node6154;
	wire [16-1:0] node6157;
	wire [16-1:0] node6158;
	wire [16-1:0] node6162;
	wire [16-1:0] node6163;
	wire [16-1:0] node6164;
	wire [16-1:0] node6167;
	wire [16-1:0] node6170;
	wire [16-1:0] node6171;
	wire [16-1:0] node6174;
	wire [16-1:0] node6177;
	wire [16-1:0] node6178;
	wire [16-1:0] node6179;
	wire [16-1:0] node6180;
	wire [16-1:0] node6183;
	wire [16-1:0] node6186;
	wire [16-1:0] node6187;
	wire [16-1:0] node6190;
	wire [16-1:0] node6193;
	wire [16-1:0] node6194;
	wire [16-1:0] node6195;
	wire [16-1:0] node6198;
	wire [16-1:0] node6201;
	wire [16-1:0] node6202;
	wire [16-1:0] node6205;
	wire [16-1:0] node6208;
	wire [16-1:0] node6209;
	wire [16-1:0] node6210;
	wire [16-1:0] node6211;
	wire [16-1:0] node6212;
	wire [16-1:0] node6213;
	wire [16-1:0] node6216;
	wire [16-1:0] node6219;
	wire [16-1:0] node6220;
	wire [16-1:0] node6223;
	wire [16-1:0] node6226;
	wire [16-1:0] node6227;
	wire [16-1:0] node6229;
	wire [16-1:0] node6232;
	wire [16-1:0] node6233;
	wire [16-1:0] node6236;
	wire [16-1:0] node6239;
	wire [16-1:0] node6240;
	wire [16-1:0] node6241;
	wire [16-1:0] node6242;
	wire [16-1:0] node6245;
	wire [16-1:0] node6248;
	wire [16-1:0] node6249;
	wire [16-1:0] node6252;
	wire [16-1:0] node6255;
	wire [16-1:0] node6256;
	wire [16-1:0] node6257;
	wire [16-1:0] node6260;
	wire [16-1:0] node6263;
	wire [16-1:0] node6264;
	wire [16-1:0] node6267;
	wire [16-1:0] node6270;
	wire [16-1:0] node6271;
	wire [16-1:0] node6272;
	wire [16-1:0] node6273;
	wire [16-1:0] node6274;
	wire [16-1:0] node6277;
	wire [16-1:0] node6280;
	wire [16-1:0] node6281;
	wire [16-1:0] node6284;
	wire [16-1:0] node6287;
	wire [16-1:0] node6288;
	wire [16-1:0] node6290;
	wire [16-1:0] node6293;
	wire [16-1:0] node6294;
	wire [16-1:0] node6297;
	wire [16-1:0] node6300;
	wire [16-1:0] node6301;
	wire [16-1:0] node6302;
	wire [16-1:0] node6303;
	wire [16-1:0] node6306;
	wire [16-1:0] node6309;
	wire [16-1:0] node6311;
	wire [16-1:0] node6314;
	wire [16-1:0] node6315;
	wire [16-1:0] node6316;
	wire [16-1:0] node6319;
	wire [16-1:0] node6322;
	wire [16-1:0] node6323;
	wire [16-1:0] node6326;
	wire [16-1:0] node6329;
	wire [16-1:0] node6330;
	wire [16-1:0] node6331;
	wire [16-1:0] node6332;
	wire [16-1:0] node6333;
	wire [16-1:0] node6334;
	wire [16-1:0] node6335;
	wire [16-1:0] node6336;
	wire [16-1:0] node6339;
	wire [16-1:0] node6342;
	wire [16-1:0] node6343;
	wire [16-1:0] node6346;
	wire [16-1:0] node6349;
	wire [16-1:0] node6350;
	wire [16-1:0] node6351;
	wire [16-1:0] node6354;
	wire [16-1:0] node6357;
	wire [16-1:0] node6358;
	wire [16-1:0] node6361;
	wire [16-1:0] node6364;
	wire [16-1:0] node6365;
	wire [16-1:0] node6366;
	wire [16-1:0] node6367;
	wire [16-1:0] node6370;
	wire [16-1:0] node6373;
	wire [16-1:0] node6374;
	wire [16-1:0] node6377;
	wire [16-1:0] node6380;
	wire [16-1:0] node6381;
	wire [16-1:0] node6382;
	wire [16-1:0] node6385;
	wire [16-1:0] node6388;
	wire [16-1:0] node6389;
	wire [16-1:0] node6393;
	wire [16-1:0] node6394;
	wire [16-1:0] node6395;
	wire [16-1:0] node6396;
	wire [16-1:0] node6397;
	wire [16-1:0] node6400;
	wire [16-1:0] node6403;
	wire [16-1:0] node6404;
	wire [16-1:0] node6407;
	wire [16-1:0] node6410;
	wire [16-1:0] node6411;
	wire [16-1:0] node6412;
	wire [16-1:0] node6415;
	wire [16-1:0] node6418;
	wire [16-1:0] node6419;
	wire [16-1:0] node6422;
	wire [16-1:0] node6425;
	wire [16-1:0] node6426;
	wire [16-1:0] node6427;
	wire [16-1:0] node6428;
	wire [16-1:0] node6432;
	wire [16-1:0] node6433;
	wire [16-1:0] node6436;
	wire [16-1:0] node6439;
	wire [16-1:0] node6440;
	wire [16-1:0] node6441;
	wire [16-1:0] node6444;
	wire [16-1:0] node6447;
	wire [16-1:0] node6448;
	wire [16-1:0] node6451;
	wire [16-1:0] node6454;
	wire [16-1:0] node6455;
	wire [16-1:0] node6456;
	wire [16-1:0] node6457;
	wire [16-1:0] node6458;
	wire [16-1:0] node6459;
	wire [16-1:0] node6462;
	wire [16-1:0] node6465;
	wire [16-1:0] node6466;
	wire [16-1:0] node6469;
	wire [16-1:0] node6472;
	wire [16-1:0] node6473;
	wire [16-1:0] node6474;
	wire [16-1:0] node6477;
	wire [16-1:0] node6480;
	wire [16-1:0] node6481;
	wire [16-1:0] node6484;
	wire [16-1:0] node6487;
	wire [16-1:0] node6488;
	wire [16-1:0] node6489;
	wire [16-1:0] node6490;
	wire [16-1:0] node6493;
	wire [16-1:0] node6496;
	wire [16-1:0] node6497;
	wire [16-1:0] node6500;
	wire [16-1:0] node6503;
	wire [16-1:0] node6504;
	wire [16-1:0] node6505;
	wire [16-1:0] node6508;
	wire [16-1:0] node6511;
	wire [16-1:0] node6512;
	wire [16-1:0] node6515;
	wire [16-1:0] node6518;
	wire [16-1:0] node6519;
	wire [16-1:0] node6520;
	wire [16-1:0] node6521;
	wire [16-1:0] node6522;
	wire [16-1:0] node6525;
	wire [16-1:0] node6528;
	wire [16-1:0] node6529;
	wire [16-1:0] node6532;
	wire [16-1:0] node6535;
	wire [16-1:0] node6536;
	wire [16-1:0] node6538;
	wire [16-1:0] node6541;
	wire [16-1:0] node6542;
	wire [16-1:0] node6545;
	wire [16-1:0] node6548;
	wire [16-1:0] node6549;
	wire [16-1:0] node6550;
	wire [16-1:0] node6551;
	wire [16-1:0] node6554;
	wire [16-1:0] node6557;
	wire [16-1:0] node6558;
	wire [16-1:0] node6561;
	wire [16-1:0] node6564;
	wire [16-1:0] node6565;
	wire [16-1:0] node6566;
	wire [16-1:0] node6569;
	wire [16-1:0] node6572;
	wire [16-1:0] node6573;
	wire [16-1:0] node6576;
	wire [16-1:0] node6579;
	wire [16-1:0] node6580;
	wire [16-1:0] node6581;
	wire [16-1:0] node6582;
	wire [16-1:0] node6583;
	wire [16-1:0] node6584;
	wire [16-1:0] node6585;
	wire [16-1:0] node6588;
	wire [16-1:0] node6591;
	wire [16-1:0] node6592;
	wire [16-1:0] node6595;
	wire [16-1:0] node6598;
	wire [16-1:0] node6599;
	wire [16-1:0] node6600;
	wire [16-1:0] node6603;
	wire [16-1:0] node6606;
	wire [16-1:0] node6607;
	wire [16-1:0] node6610;
	wire [16-1:0] node6613;
	wire [16-1:0] node6614;
	wire [16-1:0] node6615;
	wire [16-1:0] node6616;
	wire [16-1:0] node6619;
	wire [16-1:0] node6622;
	wire [16-1:0] node6623;
	wire [16-1:0] node6627;
	wire [16-1:0] node6628;
	wire [16-1:0] node6629;
	wire [16-1:0] node6632;
	wire [16-1:0] node6635;
	wire [16-1:0] node6636;
	wire [16-1:0] node6640;
	wire [16-1:0] node6641;
	wire [16-1:0] node6642;
	wire [16-1:0] node6643;
	wire [16-1:0] node6644;
	wire [16-1:0] node6647;
	wire [16-1:0] node6650;
	wire [16-1:0] node6651;
	wire [16-1:0] node6654;
	wire [16-1:0] node6657;
	wire [16-1:0] node6658;
	wire [16-1:0] node6659;
	wire [16-1:0] node6662;
	wire [16-1:0] node6665;
	wire [16-1:0] node6666;
	wire [16-1:0] node6669;
	wire [16-1:0] node6672;
	wire [16-1:0] node6673;
	wire [16-1:0] node6674;
	wire [16-1:0] node6675;
	wire [16-1:0] node6679;
	wire [16-1:0] node6680;
	wire [16-1:0] node6683;
	wire [16-1:0] node6686;
	wire [16-1:0] node6687;
	wire [16-1:0] node6688;
	wire [16-1:0] node6691;
	wire [16-1:0] node6694;
	wire [16-1:0] node6695;
	wire [16-1:0] node6698;
	wire [16-1:0] node6701;
	wire [16-1:0] node6702;
	wire [16-1:0] node6703;
	wire [16-1:0] node6704;
	wire [16-1:0] node6705;
	wire [16-1:0] node6706;
	wire [16-1:0] node6709;
	wire [16-1:0] node6712;
	wire [16-1:0] node6713;
	wire [16-1:0] node6716;
	wire [16-1:0] node6719;
	wire [16-1:0] node6720;
	wire [16-1:0] node6722;
	wire [16-1:0] node6725;
	wire [16-1:0] node6726;
	wire [16-1:0] node6729;
	wire [16-1:0] node6732;
	wire [16-1:0] node6733;
	wire [16-1:0] node6734;
	wire [16-1:0] node6735;
	wire [16-1:0] node6738;
	wire [16-1:0] node6741;
	wire [16-1:0] node6742;
	wire [16-1:0] node6745;
	wire [16-1:0] node6748;
	wire [16-1:0] node6749;
	wire [16-1:0] node6750;
	wire [16-1:0] node6753;
	wire [16-1:0] node6756;
	wire [16-1:0] node6757;
	wire [16-1:0] node6760;
	wire [16-1:0] node6763;
	wire [16-1:0] node6764;
	wire [16-1:0] node6765;
	wire [16-1:0] node6766;
	wire [16-1:0] node6767;
	wire [16-1:0] node6770;
	wire [16-1:0] node6773;
	wire [16-1:0] node6774;
	wire [16-1:0] node6777;
	wire [16-1:0] node6780;
	wire [16-1:0] node6781;
	wire [16-1:0] node6782;
	wire [16-1:0] node6785;
	wire [16-1:0] node6788;
	wire [16-1:0] node6789;
	wire [16-1:0] node6792;
	wire [16-1:0] node6795;
	wire [16-1:0] node6796;
	wire [16-1:0] node6797;
	wire [16-1:0] node6798;
	wire [16-1:0] node6801;
	wire [16-1:0] node6804;
	wire [16-1:0] node6805;
	wire [16-1:0] node6809;
	wire [16-1:0] node6810;
	wire [16-1:0] node6811;
	wire [16-1:0] node6814;
	wire [16-1:0] node6817;
	wire [16-1:0] node6818;
	wire [16-1:0] node6821;
	wire [16-1:0] node6824;
	wire [16-1:0] node6825;
	wire [16-1:0] node6826;
	wire [16-1:0] node6827;
	wire [16-1:0] node6828;
	wire [16-1:0] node6829;
	wire [16-1:0] node6830;
	wire [16-1:0] node6831;
	wire [16-1:0] node6832;
	wire [16-1:0] node6835;
	wire [16-1:0] node6838;
	wire [16-1:0] node6839;
	wire [16-1:0] node6842;
	wire [16-1:0] node6845;
	wire [16-1:0] node6846;
	wire [16-1:0] node6848;
	wire [16-1:0] node6851;
	wire [16-1:0] node6852;
	wire [16-1:0] node6856;
	wire [16-1:0] node6857;
	wire [16-1:0] node6858;
	wire [16-1:0] node6859;
	wire [16-1:0] node6863;
	wire [16-1:0] node6864;
	wire [16-1:0] node6867;
	wire [16-1:0] node6870;
	wire [16-1:0] node6871;
	wire [16-1:0] node6872;
	wire [16-1:0] node6875;
	wire [16-1:0] node6878;
	wire [16-1:0] node6879;
	wire [16-1:0] node6882;
	wire [16-1:0] node6885;
	wire [16-1:0] node6886;
	wire [16-1:0] node6887;
	wire [16-1:0] node6888;
	wire [16-1:0] node6889;
	wire [16-1:0] node6893;
	wire [16-1:0] node6894;
	wire [16-1:0] node6897;
	wire [16-1:0] node6900;
	wire [16-1:0] node6901;
	wire [16-1:0] node6902;
	wire [16-1:0] node6905;
	wire [16-1:0] node6908;
	wire [16-1:0] node6909;
	wire [16-1:0] node6913;
	wire [16-1:0] node6914;
	wire [16-1:0] node6915;
	wire [16-1:0] node6916;
	wire [16-1:0] node6919;
	wire [16-1:0] node6922;
	wire [16-1:0] node6923;
	wire [16-1:0] node6926;
	wire [16-1:0] node6929;
	wire [16-1:0] node6930;
	wire [16-1:0] node6931;
	wire [16-1:0] node6934;
	wire [16-1:0] node6937;
	wire [16-1:0] node6938;
	wire [16-1:0] node6941;
	wire [16-1:0] node6944;
	wire [16-1:0] node6945;
	wire [16-1:0] node6946;
	wire [16-1:0] node6947;
	wire [16-1:0] node6948;
	wire [16-1:0] node6949;
	wire [16-1:0] node6952;
	wire [16-1:0] node6955;
	wire [16-1:0] node6957;
	wire [16-1:0] node6960;
	wire [16-1:0] node6961;
	wire [16-1:0] node6963;
	wire [16-1:0] node6966;
	wire [16-1:0] node6967;
	wire [16-1:0] node6970;
	wire [16-1:0] node6973;
	wire [16-1:0] node6974;
	wire [16-1:0] node6975;
	wire [16-1:0] node6976;
	wire [16-1:0] node6979;
	wire [16-1:0] node6982;
	wire [16-1:0] node6983;
	wire [16-1:0] node6986;
	wire [16-1:0] node6989;
	wire [16-1:0] node6990;
	wire [16-1:0] node6991;
	wire [16-1:0] node6994;
	wire [16-1:0] node6997;
	wire [16-1:0] node6998;
	wire [16-1:0] node7001;
	wire [16-1:0] node7004;
	wire [16-1:0] node7005;
	wire [16-1:0] node7006;
	wire [16-1:0] node7007;
	wire [16-1:0] node7008;
	wire [16-1:0] node7011;
	wire [16-1:0] node7014;
	wire [16-1:0] node7015;
	wire [16-1:0] node7018;
	wire [16-1:0] node7021;
	wire [16-1:0] node7022;
	wire [16-1:0] node7023;
	wire [16-1:0] node7026;
	wire [16-1:0] node7029;
	wire [16-1:0] node7031;
	wire [16-1:0] node7034;
	wire [16-1:0] node7035;
	wire [16-1:0] node7036;
	wire [16-1:0] node7037;
	wire [16-1:0] node7040;
	wire [16-1:0] node7043;
	wire [16-1:0] node7044;
	wire [16-1:0] node7047;
	wire [16-1:0] node7050;
	wire [16-1:0] node7051;
	wire [16-1:0] node7052;
	wire [16-1:0] node7055;
	wire [16-1:0] node7058;
	wire [16-1:0] node7059;
	wire [16-1:0] node7062;
	wire [16-1:0] node7065;
	wire [16-1:0] node7066;
	wire [16-1:0] node7067;
	wire [16-1:0] node7068;
	wire [16-1:0] node7069;
	wire [16-1:0] node7070;
	wire [16-1:0] node7071;
	wire [16-1:0] node7074;
	wire [16-1:0] node7077;
	wire [16-1:0] node7078;
	wire [16-1:0] node7081;
	wire [16-1:0] node7084;
	wire [16-1:0] node7085;
	wire [16-1:0] node7086;
	wire [16-1:0] node7090;
	wire [16-1:0] node7091;
	wire [16-1:0] node7095;
	wire [16-1:0] node7096;
	wire [16-1:0] node7097;
	wire [16-1:0] node7098;
	wire [16-1:0] node7101;
	wire [16-1:0] node7104;
	wire [16-1:0] node7105;
	wire [16-1:0] node7108;
	wire [16-1:0] node7111;
	wire [16-1:0] node7112;
	wire [16-1:0] node7113;
	wire [16-1:0] node7116;
	wire [16-1:0] node7119;
	wire [16-1:0] node7121;
	wire [16-1:0] node7124;
	wire [16-1:0] node7125;
	wire [16-1:0] node7126;
	wire [16-1:0] node7127;
	wire [16-1:0] node7128;
	wire [16-1:0] node7131;
	wire [16-1:0] node7134;
	wire [16-1:0] node7135;
	wire [16-1:0] node7138;
	wire [16-1:0] node7141;
	wire [16-1:0] node7142;
	wire [16-1:0] node7143;
	wire [16-1:0] node7146;
	wire [16-1:0] node7149;
	wire [16-1:0] node7150;
	wire [16-1:0] node7153;
	wire [16-1:0] node7156;
	wire [16-1:0] node7157;
	wire [16-1:0] node7158;
	wire [16-1:0] node7159;
	wire [16-1:0] node7162;
	wire [16-1:0] node7165;
	wire [16-1:0] node7166;
	wire [16-1:0] node7169;
	wire [16-1:0] node7172;
	wire [16-1:0] node7173;
	wire [16-1:0] node7174;
	wire [16-1:0] node7177;
	wire [16-1:0] node7180;
	wire [16-1:0] node7181;
	wire [16-1:0] node7184;
	wire [16-1:0] node7187;
	wire [16-1:0] node7188;
	wire [16-1:0] node7189;
	wire [16-1:0] node7190;
	wire [16-1:0] node7191;
	wire [16-1:0] node7192;
	wire [16-1:0] node7196;
	wire [16-1:0] node7197;
	wire [16-1:0] node7200;
	wire [16-1:0] node7203;
	wire [16-1:0] node7204;
	wire [16-1:0] node7205;
	wire [16-1:0] node7208;
	wire [16-1:0] node7211;
	wire [16-1:0] node7213;
	wire [16-1:0] node7216;
	wire [16-1:0] node7217;
	wire [16-1:0] node7218;
	wire [16-1:0] node7219;
	wire [16-1:0] node7222;
	wire [16-1:0] node7225;
	wire [16-1:0] node7226;
	wire [16-1:0] node7229;
	wire [16-1:0] node7232;
	wire [16-1:0] node7233;
	wire [16-1:0] node7234;
	wire [16-1:0] node7237;
	wire [16-1:0] node7240;
	wire [16-1:0] node7241;
	wire [16-1:0] node7244;
	wire [16-1:0] node7247;
	wire [16-1:0] node7248;
	wire [16-1:0] node7249;
	wire [16-1:0] node7250;
	wire [16-1:0] node7251;
	wire [16-1:0] node7255;
	wire [16-1:0] node7256;
	wire [16-1:0] node7259;
	wire [16-1:0] node7262;
	wire [16-1:0] node7263;
	wire [16-1:0] node7264;
	wire [16-1:0] node7267;
	wire [16-1:0] node7270;
	wire [16-1:0] node7271;
	wire [16-1:0] node7274;
	wire [16-1:0] node7277;
	wire [16-1:0] node7278;
	wire [16-1:0] node7279;
	wire [16-1:0] node7280;
	wire [16-1:0] node7283;
	wire [16-1:0] node7286;
	wire [16-1:0] node7287;
	wire [16-1:0] node7290;
	wire [16-1:0] node7293;
	wire [16-1:0] node7294;
	wire [16-1:0] node7295;
	wire [16-1:0] node7298;
	wire [16-1:0] node7301;
	wire [16-1:0] node7302;
	wire [16-1:0] node7305;
	wire [16-1:0] node7308;
	wire [16-1:0] node7309;
	wire [16-1:0] node7310;
	wire [16-1:0] node7311;
	wire [16-1:0] node7312;
	wire [16-1:0] node7313;
	wire [16-1:0] node7314;
	wire [16-1:0] node7315;
	wire [16-1:0] node7318;
	wire [16-1:0] node7321;
	wire [16-1:0] node7322;
	wire [16-1:0] node7325;
	wire [16-1:0] node7328;
	wire [16-1:0] node7329;
	wire [16-1:0] node7330;
	wire [16-1:0] node7333;
	wire [16-1:0] node7336;
	wire [16-1:0] node7337;
	wire [16-1:0] node7341;
	wire [16-1:0] node7342;
	wire [16-1:0] node7343;
	wire [16-1:0] node7345;
	wire [16-1:0] node7348;
	wire [16-1:0] node7349;
	wire [16-1:0] node7352;
	wire [16-1:0] node7355;
	wire [16-1:0] node7356;
	wire [16-1:0] node7357;
	wire [16-1:0] node7361;
	wire [16-1:0] node7362;
	wire [16-1:0] node7365;
	wire [16-1:0] node7368;
	wire [16-1:0] node7369;
	wire [16-1:0] node7370;
	wire [16-1:0] node7371;
	wire [16-1:0] node7372;
	wire [16-1:0] node7375;
	wire [16-1:0] node7378;
	wire [16-1:0] node7379;
	wire [16-1:0] node7382;
	wire [16-1:0] node7385;
	wire [16-1:0] node7386;
	wire [16-1:0] node7387;
	wire [16-1:0] node7390;
	wire [16-1:0] node7393;
	wire [16-1:0] node7394;
	wire [16-1:0] node7397;
	wire [16-1:0] node7400;
	wire [16-1:0] node7401;
	wire [16-1:0] node7402;
	wire [16-1:0] node7403;
	wire [16-1:0] node7407;
	wire [16-1:0] node7408;
	wire [16-1:0] node7411;
	wire [16-1:0] node7414;
	wire [16-1:0] node7415;
	wire [16-1:0] node7416;
	wire [16-1:0] node7419;
	wire [16-1:0] node7422;
	wire [16-1:0] node7423;
	wire [16-1:0] node7426;
	wire [16-1:0] node7429;
	wire [16-1:0] node7430;
	wire [16-1:0] node7431;
	wire [16-1:0] node7432;
	wire [16-1:0] node7433;
	wire [16-1:0] node7435;
	wire [16-1:0] node7438;
	wire [16-1:0] node7439;
	wire [16-1:0] node7442;
	wire [16-1:0] node7445;
	wire [16-1:0] node7446;
	wire [16-1:0] node7447;
	wire [16-1:0] node7450;
	wire [16-1:0] node7453;
	wire [16-1:0] node7455;
	wire [16-1:0] node7458;
	wire [16-1:0] node7459;
	wire [16-1:0] node7460;
	wire [16-1:0] node7461;
	wire [16-1:0] node7464;
	wire [16-1:0] node7467;
	wire [16-1:0] node7468;
	wire [16-1:0] node7471;
	wire [16-1:0] node7474;
	wire [16-1:0] node7475;
	wire [16-1:0] node7476;
	wire [16-1:0] node7479;
	wire [16-1:0] node7482;
	wire [16-1:0] node7484;
	wire [16-1:0] node7487;
	wire [16-1:0] node7488;
	wire [16-1:0] node7489;
	wire [16-1:0] node7490;
	wire [16-1:0] node7491;
	wire [16-1:0] node7494;
	wire [16-1:0] node7497;
	wire [16-1:0] node7498;
	wire [16-1:0] node7501;
	wire [16-1:0] node7504;
	wire [16-1:0] node7505;
	wire [16-1:0] node7506;
	wire [16-1:0] node7509;
	wire [16-1:0] node7512;
	wire [16-1:0] node7513;
	wire [16-1:0] node7516;
	wire [16-1:0] node7519;
	wire [16-1:0] node7520;
	wire [16-1:0] node7521;
	wire [16-1:0] node7522;
	wire [16-1:0] node7525;
	wire [16-1:0] node7528;
	wire [16-1:0] node7529;
	wire [16-1:0] node7532;
	wire [16-1:0] node7535;
	wire [16-1:0] node7536;
	wire [16-1:0] node7537;
	wire [16-1:0] node7540;
	wire [16-1:0] node7543;
	wire [16-1:0] node7545;
	wire [16-1:0] node7548;
	wire [16-1:0] node7549;
	wire [16-1:0] node7550;
	wire [16-1:0] node7551;
	wire [16-1:0] node7552;
	wire [16-1:0] node7553;
	wire [16-1:0] node7554;
	wire [16-1:0] node7557;
	wire [16-1:0] node7560;
	wire [16-1:0] node7561;
	wire [16-1:0] node7564;
	wire [16-1:0] node7567;
	wire [16-1:0] node7568;
	wire [16-1:0] node7569;
	wire [16-1:0] node7572;
	wire [16-1:0] node7575;
	wire [16-1:0] node7576;
	wire [16-1:0] node7579;
	wire [16-1:0] node7582;
	wire [16-1:0] node7583;
	wire [16-1:0] node7584;
	wire [16-1:0] node7585;
	wire [16-1:0] node7588;
	wire [16-1:0] node7591;
	wire [16-1:0] node7592;
	wire [16-1:0] node7595;
	wire [16-1:0] node7598;
	wire [16-1:0] node7599;
	wire [16-1:0] node7600;
	wire [16-1:0] node7603;
	wire [16-1:0] node7606;
	wire [16-1:0] node7607;
	wire [16-1:0] node7610;
	wire [16-1:0] node7613;
	wire [16-1:0] node7614;
	wire [16-1:0] node7615;
	wire [16-1:0] node7616;
	wire [16-1:0] node7617;
	wire [16-1:0] node7620;
	wire [16-1:0] node7623;
	wire [16-1:0] node7624;
	wire [16-1:0] node7627;
	wire [16-1:0] node7630;
	wire [16-1:0] node7631;
	wire [16-1:0] node7632;
	wire [16-1:0] node7635;
	wire [16-1:0] node7638;
	wire [16-1:0] node7639;
	wire [16-1:0] node7642;
	wire [16-1:0] node7645;
	wire [16-1:0] node7646;
	wire [16-1:0] node7647;
	wire [16-1:0] node7649;
	wire [16-1:0] node7652;
	wire [16-1:0] node7653;
	wire [16-1:0] node7656;
	wire [16-1:0] node7659;
	wire [16-1:0] node7660;
	wire [16-1:0] node7662;
	wire [16-1:0] node7665;
	wire [16-1:0] node7668;
	wire [16-1:0] node7669;
	wire [16-1:0] node7670;
	wire [16-1:0] node7671;
	wire [16-1:0] node7672;
	wire [16-1:0] node7675;
	wire [16-1:0] node7676;
	wire [16-1:0] node7679;
	wire [16-1:0] node7682;
	wire [16-1:0] node7683;
	wire [16-1:0] node7684;
	wire [16-1:0] node7687;
	wire [16-1:0] node7690;
	wire [16-1:0] node7691;
	wire [16-1:0] node7694;
	wire [16-1:0] node7697;
	wire [16-1:0] node7698;
	wire [16-1:0] node7699;
	wire [16-1:0] node7700;
	wire [16-1:0] node7703;
	wire [16-1:0] node7706;
	wire [16-1:0] node7707;
	wire [16-1:0] node7710;
	wire [16-1:0] node7713;
	wire [16-1:0] node7714;
	wire [16-1:0] node7716;
	wire [16-1:0] node7719;
	wire [16-1:0] node7720;
	wire [16-1:0] node7723;
	wire [16-1:0] node7726;
	wire [16-1:0] node7727;
	wire [16-1:0] node7728;
	wire [16-1:0] node7729;
	wire [16-1:0] node7730;
	wire [16-1:0] node7733;
	wire [16-1:0] node7736;
	wire [16-1:0] node7737;
	wire [16-1:0] node7740;
	wire [16-1:0] node7743;
	wire [16-1:0] node7744;
	wire [16-1:0] node7745;
	wire [16-1:0] node7748;
	wire [16-1:0] node7751;
	wire [16-1:0] node7753;
	wire [16-1:0] node7756;
	wire [16-1:0] node7757;
	wire [16-1:0] node7758;
	wire [16-1:0] node7759;
	wire [16-1:0] node7762;
	wire [16-1:0] node7765;
	wire [16-1:0] node7766;
	wire [16-1:0] node7769;
	wire [16-1:0] node7772;
	wire [16-1:0] node7773;
	wire [16-1:0] node7775;
	wire [16-1:0] node7778;
	wire [16-1:0] node7779;
	wire [16-1:0] node7782;
	wire [16-1:0] node7785;
	wire [16-1:0] node7786;
	wire [16-1:0] node7787;
	wire [16-1:0] node7788;
	wire [16-1:0] node7789;
	wire [16-1:0] node7790;
	wire [16-1:0] node7791;
	wire [16-1:0] node7792;
	wire [16-1:0] node7793;
	wire [16-1:0] node7794;
	wire [16-1:0] node7795;
	wire [16-1:0] node7796;
	wire [16-1:0] node7799;
	wire [16-1:0] node7802;
	wire [16-1:0] node7803;
	wire [16-1:0] node7806;
	wire [16-1:0] node7809;
	wire [16-1:0] node7810;
	wire [16-1:0] node7811;
	wire [16-1:0] node7814;
	wire [16-1:0] node7817;
	wire [16-1:0] node7818;
	wire [16-1:0] node7821;
	wire [16-1:0] node7824;
	wire [16-1:0] node7825;
	wire [16-1:0] node7826;
	wire [16-1:0] node7827;
	wire [16-1:0] node7830;
	wire [16-1:0] node7833;
	wire [16-1:0] node7834;
	wire [16-1:0] node7837;
	wire [16-1:0] node7840;
	wire [16-1:0] node7841;
	wire [16-1:0] node7842;
	wire [16-1:0] node7845;
	wire [16-1:0] node7848;
	wire [16-1:0] node7849;
	wire [16-1:0] node7852;
	wire [16-1:0] node7855;
	wire [16-1:0] node7856;
	wire [16-1:0] node7857;
	wire [16-1:0] node7858;
	wire [16-1:0] node7859;
	wire [16-1:0] node7862;
	wire [16-1:0] node7865;
	wire [16-1:0] node7866;
	wire [16-1:0] node7869;
	wire [16-1:0] node7872;
	wire [16-1:0] node7873;
	wire [16-1:0] node7874;
	wire [16-1:0] node7877;
	wire [16-1:0] node7880;
	wire [16-1:0] node7881;
	wire [16-1:0] node7884;
	wire [16-1:0] node7887;
	wire [16-1:0] node7888;
	wire [16-1:0] node7889;
	wire [16-1:0] node7890;
	wire [16-1:0] node7893;
	wire [16-1:0] node7896;
	wire [16-1:0] node7897;
	wire [16-1:0] node7900;
	wire [16-1:0] node7903;
	wire [16-1:0] node7904;
	wire [16-1:0] node7905;
	wire [16-1:0] node7908;
	wire [16-1:0] node7911;
	wire [16-1:0] node7912;
	wire [16-1:0] node7915;
	wire [16-1:0] node7918;
	wire [16-1:0] node7919;
	wire [16-1:0] node7920;
	wire [16-1:0] node7921;
	wire [16-1:0] node7922;
	wire [16-1:0] node7923;
	wire [16-1:0] node7926;
	wire [16-1:0] node7929;
	wire [16-1:0] node7930;
	wire [16-1:0] node7933;
	wire [16-1:0] node7936;
	wire [16-1:0] node7937;
	wire [16-1:0] node7938;
	wire [16-1:0] node7942;
	wire [16-1:0] node7943;
	wire [16-1:0] node7946;
	wire [16-1:0] node7949;
	wire [16-1:0] node7950;
	wire [16-1:0] node7951;
	wire [16-1:0] node7953;
	wire [16-1:0] node7956;
	wire [16-1:0] node7957;
	wire [16-1:0] node7960;
	wire [16-1:0] node7963;
	wire [16-1:0] node7964;
	wire [16-1:0] node7965;
	wire [16-1:0] node7968;
	wire [16-1:0] node7971;
	wire [16-1:0] node7972;
	wire [16-1:0] node7976;
	wire [16-1:0] node7977;
	wire [16-1:0] node7978;
	wire [16-1:0] node7979;
	wire [16-1:0] node7980;
	wire [16-1:0] node7983;
	wire [16-1:0] node7986;
	wire [16-1:0] node7987;
	wire [16-1:0] node7991;
	wire [16-1:0] node7992;
	wire [16-1:0] node7993;
	wire [16-1:0] node7996;
	wire [16-1:0] node7999;
	wire [16-1:0] node8000;
	wire [16-1:0] node8003;
	wire [16-1:0] node8006;
	wire [16-1:0] node8007;
	wire [16-1:0] node8008;
	wire [16-1:0] node8009;
	wire [16-1:0] node8012;
	wire [16-1:0] node8015;
	wire [16-1:0] node8017;
	wire [16-1:0] node8020;
	wire [16-1:0] node8021;
	wire [16-1:0] node8023;
	wire [16-1:0] node8026;
	wire [16-1:0] node8027;
	wire [16-1:0] node8030;
	wire [16-1:0] node8033;
	wire [16-1:0] node8034;
	wire [16-1:0] node8035;
	wire [16-1:0] node8036;
	wire [16-1:0] node8037;
	wire [16-1:0] node8038;
	wire [16-1:0] node8039;
	wire [16-1:0] node8042;
	wire [16-1:0] node8045;
	wire [16-1:0] node8046;
	wire [16-1:0] node8049;
	wire [16-1:0] node8052;
	wire [16-1:0] node8053;
	wire [16-1:0] node8054;
	wire [16-1:0] node8057;
	wire [16-1:0] node8060;
	wire [16-1:0] node8061;
	wire [16-1:0] node8064;
	wire [16-1:0] node8067;
	wire [16-1:0] node8068;
	wire [16-1:0] node8069;
	wire [16-1:0] node8070;
	wire [16-1:0] node8073;
	wire [16-1:0] node8076;
	wire [16-1:0] node8077;
	wire [16-1:0] node8081;
	wire [16-1:0] node8082;
	wire [16-1:0] node8083;
	wire [16-1:0] node8086;
	wire [16-1:0] node8089;
	wire [16-1:0] node8090;
	wire [16-1:0] node8093;
	wire [16-1:0] node8096;
	wire [16-1:0] node8097;
	wire [16-1:0] node8098;
	wire [16-1:0] node8099;
	wire [16-1:0] node8100;
	wire [16-1:0] node8103;
	wire [16-1:0] node8106;
	wire [16-1:0] node8107;
	wire [16-1:0] node8110;
	wire [16-1:0] node8113;
	wire [16-1:0] node8114;
	wire [16-1:0] node8115;
	wire [16-1:0] node8118;
	wire [16-1:0] node8121;
	wire [16-1:0] node8123;
	wire [16-1:0] node8126;
	wire [16-1:0] node8127;
	wire [16-1:0] node8128;
	wire [16-1:0] node8129;
	wire [16-1:0] node8133;
	wire [16-1:0] node8134;
	wire [16-1:0] node8137;
	wire [16-1:0] node8140;
	wire [16-1:0] node8141;
	wire [16-1:0] node8142;
	wire [16-1:0] node8146;
	wire [16-1:0] node8147;
	wire [16-1:0] node8150;
	wire [16-1:0] node8153;
	wire [16-1:0] node8154;
	wire [16-1:0] node8155;
	wire [16-1:0] node8156;
	wire [16-1:0] node8157;
	wire [16-1:0] node8159;
	wire [16-1:0] node8162;
	wire [16-1:0] node8163;
	wire [16-1:0] node8166;
	wire [16-1:0] node8169;
	wire [16-1:0] node8170;
	wire [16-1:0] node8171;
	wire [16-1:0] node8174;
	wire [16-1:0] node8177;
	wire [16-1:0] node8178;
	wire [16-1:0] node8181;
	wire [16-1:0] node8184;
	wire [16-1:0] node8185;
	wire [16-1:0] node8186;
	wire [16-1:0] node8187;
	wire [16-1:0] node8190;
	wire [16-1:0] node8193;
	wire [16-1:0] node8194;
	wire [16-1:0] node8197;
	wire [16-1:0] node8200;
	wire [16-1:0] node8201;
	wire [16-1:0] node8204;
	wire [16-1:0] node8206;
	wire [16-1:0] node8209;
	wire [16-1:0] node8210;
	wire [16-1:0] node8211;
	wire [16-1:0] node8212;
	wire [16-1:0] node8213;
	wire [16-1:0] node8216;
	wire [16-1:0] node8219;
	wire [16-1:0] node8220;
	wire [16-1:0] node8223;
	wire [16-1:0] node8226;
	wire [16-1:0] node8227;
	wire [16-1:0] node8228;
	wire [16-1:0] node8231;
	wire [16-1:0] node8234;
	wire [16-1:0] node8235;
	wire [16-1:0] node8238;
	wire [16-1:0] node8241;
	wire [16-1:0] node8242;
	wire [16-1:0] node8243;
	wire [16-1:0] node8244;
	wire [16-1:0] node8247;
	wire [16-1:0] node8250;
	wire [16-1:0] node8251;
	wire [16-1:0] node8254;
	wire [16-1:0] node8257;
	wire [16-1:0] node8258;
	wire [16-1:0] node8259;
	wire [16-1:0] node8262;
	wire [16-1:0] node8265;
	wire [16-1:0] node8266;
	wire [16-1:0] node8269;
	wire [16-1:0] node8272;
	wire [16-1:0] node8273;
	wire [16-1:0] node8274;
	wire [16-1:0] node8275;
	wire [16-1:0] node8276;
	wire [16-1:0] node8277;
	wire [16-1:0] node8278;
	wire [16-1:0] node8279;
	wire [16-1:0] node8282;
	wire [16-1:0] node8285;
	wire [16-1:0] node8286;
	wire [16-1:0] node8289;
	wire [16-1:0] node8292;
	wire [16-1:0] node8293;
	wire [16-1:0] node8295;
	wire [16-1:0] node8298;
	wire [16-1:0] node8299;
	wire [16-1:0] node8302;
	wire [16-1:0] node8305;
	wire [16-1:0] node8306;
	wire [16-1:0] node8307;
	wire [16-1:0] node8308;
	wire [16-1:0] node8311;
	wire [16-1:0] node8314;
	wire [16-1:0] node8315;
	wire [16-1:0] node8318;
	wire [16-1:0] node8321;
	wire [16-1:0] node8322;
	wire [16-1:0] node8323;
	wire [16-1:0] node8326;
	wire [16-1:0] node8329;
	wire [16-1:0] node8330;
	wire [16-1:0] node8333;
	wire [16-1:0] node8336;
	wire [16-1:0] node8337;
	wire [16-1:0] node8338;
	wire [16-1:0] node8339;
	wire [16-1:0] node8340;
	wire [16-1:0] node8343;
	wire [16-1:0] node8346;
	wire [16-1:0] node8347;
	wire [16-1:0] node8350;
	wire [16-1:0] node8353;
	wire [16-1:0] node8354;
	wire [16-1:0] node8355;
	wire [16-1:0] node8358;
	wire [16-1:0] node8361;
	wire [16-1:0] node8362;
	wire [16-1:0] node8365;
	wire [16-1:0] node8368;
	wire [16-1:0] node8369;
	wire [16-1:0] node8370;
	wire [16-1:0] node8371;
	wire [16-1:0] node8374;
	wire [16-1:0] node8377;
	wire [16-1:0] node8378;
	wire [16-1:0] node8381;
	wire [16-1:0] node8384;
	wire [16-1:0] node8385;
	wire [16-1:0] node8386;
	wire [16-1:0] node8389;
	wire [16-1:0] node8392;
	wire [16-1:0] node8393;
	wire [16-1:0] node8396;
	wire [16-1:0] node8399;
	wire [16-1:0] node8400;
	wire [16-1:0] node8401;
	wire [16-1:0] node8402;
	wire [16-1:0] node8403;
	wire [16-1:0] node8405;
	wire [16-1:0] node8408;
	wire [16-1:0] node8409;
	wire [16-1:0] node8412;
	wire [16-1:0] node8415;
	wire [16-1:0] node8416;
	wire [16-1:0] node8417;
	wire [16-1:0] node8420;
	wire [16-1:0] node8423;
	wire [16-1:0] node8424;
	wire [16-1:0] node8428;
	wire [16-1:0] node8429;
	wire [16-1:0] node8430;
	wire [16-1:0] node8431;
	wire [16-1:0] node8434;
	wire [16-1:0] node8437;
	wire [16-1:0] node8439;
	wire [16-1:0] node8442;
	wire [16-1:0] node8443;
	wire [16-1:0] node8444;
	wire [16-1:0] node8447;
	wire [16-1:0] node8450;
	wire [16-1:0] node8451;
	wire [16-1:0] node8454;
	wire [16-1:0] node8457;
	wire [16-1:0] node8458;
	wire [16-1:0] node8459;
	wire [16-1:0] node8460;
	wire [16-1:0] node8461;
	wire [16-1:0] node8464;
	wire [16-1:0] node8467;
	wire [16-1:0] node8468;
	wire [16-1:0] node8471;
	wire [16-1:0] node8474;
	wire [16-1:0] node8475;
	wire [16-1:0] node8476;
	wire [16-1:0] node8479;
	wire [16-1:0] node8482;
	wire [16-1:0] node8483;
	wire [16-1:0] node8486;
	wire [16-1:0] node8489;
	wire [16-1:0] node8490;
	wire [16-1:0] node8491;
	wire [16-1:0] node8492;
	wire [16-1:0] node8495;
	wire [16-1:0] node8498;
	wire [16-1:0] node8499;
	wire [16-1:0] node8502;
	wire [16-1:0] node8505;
	wire [16-1:0] node8506;
	wire [16-1:0] node8508;
	wire [16-1:0] node8511;
	wire [16-1:0] node8512;
	wire [16-1:0] node8515;
	wire [16-1:0] node8518;
	wire [16-1:0] node8519;
	wire [16-1:0] node8520;
	wire [16-1:0] node8521;
	wire [16-1:0] node8522;
	wire [16-1:0] node8523;
	wire [16-1:0] node8524;
	wire [16-1:0] node8527;
	wire [16-1:0] node8530;
	wire [16-1:0] node8531;
	wire [16-1:0] node8534;
	wire [16-1:0] node8537;
	wire [16-1:0] node8538;
	wire [16-1:0] node8539;
	wire [16-1:0] node8542;
	wire [16-1:0] node8545;
	wire [16-1:0] node8546;
	wire [16-1:0] node8549;
	wire [16-1:0] node8552;
	wire [16-1:0] node8553;
	wire [16-1:0] node8554;
	wire [16-1:0] node8555;
	wire [16-1:0] node8558;
	wire [16-1:0] node8561;
	wire [16-1:0] node8562;
	wire [16-1:0] node8565;
	wire [16-1:0] node8568;
	wire [16-1:0] node8569;
	wire [16-1:0] node8570;
	wire [16-1:0] node8573;
	wire [16-1:0] node8576;
	wire [16-1:0] node8577;
	wire [16-1:0] node8580;
	wire [16-1:0] node8583;
	wire [16-1:0] node8584;
	wire [16-1:0] node8585;
	wire [16-1:0] node8586;
	wire [16-1:0] node8588;
	wire [16-1:0] node8591;
	wire [16-1:0] node8592;
	wire [16-1:0] node8595;
	wire [16-1:0] node8598;
	wire [16-1:0] node8599;
	wire [16-1:0] node8600;
	wire [16-1:0] node8603;
	wire [16-1:0] node8606;
	wire [16-1:0] node8607;
	wire [16-1:0] node8611;
	wire [16-1:0] node8612;
	wire [16-1:0] node8613;
	wire [16-1:0] node8614;
	wire [16-1:0] node8617;
	wire [16-1:0] node8620;
	wire [16-1:0] node8621;
	wire [16-1:0] node8624;
	wire [16-1:0] node8627;
	wire [16-1:0] node8628;
	wire [16-1:0] node8629;
	wire [16-1:0] node8632;
	wire [16-1:0] node8635;
	wire [16-1:0] node8636;
	wire [16-1:0] node8639;
	wire [16-1:0] node8642;
	wire [16-1:0] node8643;
	wire [16-1:0] node8644;
	wire [16-1:0] node8645;
	wire [16-1:0] node8646;
	wire [16-1:0] node8647;
	wire [16-1:0] node8650;
	wire [16-1:0] node8653;
	wire [16-1:0] node8654;
	wire [16-1:0] node8657;
	wire [16-1:0] node8660;
	wire [16-1:0] node8661;
	wire [16-1:0] node8662;
	wire [16-1:0] node8666;
	wire [16-1:0] node8667;
	wire [16-1:0] node8670;
	wire [16-1:0] node8673;
	wire [16-1:0] node8674;
	wire [16-1:0] node8675;
	wire [16-1:0] node8676;
	wire [16-1:0] node8679;
	wire [16-1:0] node8682;
	wire [16-1:0] node8683;
	wire [16-1:0] node8686;
	wire [16-1:0] node8689;
	wire [16-1:0] node8690;
	wire [16-1:0] node8691;
	wire [16-1:0] node8694;
	wire [16-1:0] node8697;
	wire [16-1:0] node8698;
	wire [16-1:0] node8701;
	wire [16-1:0] node8704;
	wire [16-1:0] node8705;
	wire [16-1:0] node8706;
	wire [16-1:0] node8707;
	wire [16-1:0] node8709;
	wire [16-1:0] node8712;
	wire [16-1:0] node8713;
	wire [16-1:0] node8716;
	wire [16-1:0] node8719;
	wire [16-1:0] node8720;
	wire [16-1:0] node8722;
	wire [16-1:0] node8726;
	wire [16-1:0] node8727;
	wire [16-1:0] node8728;
	wire [16-1:0] node8729;
	wire [16-1:0] node8732;
	wire [16-1:0] node8735;
	wire [16-1:0] node8736;
	wire [16-1:0] node8739;
	wire [16-1:0] node8742;
	wire [16-1:0] node8743;
	wire [16-1:0] node8744;
	wire [16-1:0] node8747;
	wire [16-1:0] node8750;
	wire [16-1:0] node8751;
	wire [16-1:0] node8754;
	wire [16-1:0] node8757;
	wire [16-1:0] node8758;
	wire [16-1:0] node8759;
	wire [16-1:0] node8760;
	wire [16-1:0] node8761;
	wire [16-1:0] node8762;
	wire [16-1:0] node8763;
	wire [16-1:0] node8764;
	wire [16-1:0] node8765;
	wire [16-1:0] node8768;
	wire [16-1:0] node8771;
	wire [16-1:0] node8772;
	wire [16-1:0] node8776;
	wire [16-1:0] node8777;
	wire [16-1:0] node8778;
	wire [16-1:0] node8782;
	wire [16-1:0] node8783;
	wire [16-1:0] node8786;
	wire [16-1:0] node8789;
	wire [16-1:0] node8790;
	wire [16-1:0] node8791;
	wire [16-1:0] node8792;
	wire [16-1:0] node8795;
	wire [16-1:0] node8798;
	wire [16-1:0] node8799;
	wire [16-1:0] node8802;
	wire [16-1:0] node8805;
	wire [16-1:0] node8806;
	wire [16-1:0] node8807;
	wire [16-1:0] node8810;
	wire [16-1:0] node8813;
	wire [16-1:0] node8814;
	wire [16-1:0] node8817;
	wire [16-1:0] node8820;
	wire [16-1:0] node8821;
	wire [16-1:0] node8822;
	wire [16-1:0] node8823;
	wire [16-1:0] node8824;
	wire [16-1:0] node8827;
	wire [16-1:0] node8830;
	wire [16-1:0] node8831;
	wire [16-1:0] node8835;
	wire [16-1:0] node8836;
	wire [16-1:0] node8837;
	wire [16-1:0] node8840;
	wire [16-1:0] node8843;
	wire [16-1:0] node8844;
	wire [16-1:0] node8848;
	wire [16-1:0] node8849;
	wire [16-1:0] node8850;
	wire [16-1:0] node8851;
	wire [16-1:0] node8854;
	wire [16-1:0] node8857;
	wire [16-1:0] node8858;
	wire [16-1:0] node8861;
	wire [16-1:0] node8864;
	wire [16-1:0] node8865;
	wire [16-1:0] node8867;
	wire [16-1:0] node8870;
	wire [16-1:0] node8871;
	wire [16-1:0] node8874;
	wire [16-1:0] node8877;
	wire [16-1:0] node8878;
	wire [16-1:0] node8879;
	wire [16-1:0] node8880;
	wire [16-1:0] node8881;
	wire [16-1:0] node8882;
	wire [16-1:0] node8885;
	wire [16-1:0] node8888;
	wire [16-1:0] node8889;
	wire [16-1:0] node8892;
	wire [16-1:0] node8895;
	wire [16-1:0] node8896;
	wire [16-1:0] node8897;
	wire [16-1:0] node8900;
	wire [16-1:0] node8903;
	wire [16-1:0] node8904;
	wire [16-1:0] node8907;
	wire [16-1:0] node8910;
	wire [16-1:0] node8911;
	wire [16-1:0] node8912;
	wire [16-1:0] node8913;
	wire [16-1:0] node8916;
	wire [16-1:0] node8919;
	wire [16-1:0] node8920;
	wire [16-1:0] node8923;
	wire [16-1:0] node8926;
	wire [16-1:0] node8927;
	wire [16-1:0] node8929;
	wire [16-1:0] node8932;
	wire [16-1:0] node8933;
	wire [16-1:0] node8936;
	wire [16-1:0] node8939;
	wire [16-1:0] node8940;
	wire [16-1:0] node8941;
	wire [16-1:0] node8942;
	wire [16-1:0] node8943;
	wire [16-1:0] node8946;
	wire [16-1:0] node8949;
	wire [16-1:0] node8950;
	wire [16-1:0] node8953;
	wire [16-1:0] node8956;
	wire [16-1:0] node8957;
	wire [16-1:0] node8958;
	wire [16-1:0] node8961;
	wire [16-1:0] node8964;
	wire [16-1:0] node8965;
	wire [16-1:0] node8968;
	wire [16-1:0] node8971;
	wire [16-1:0] node8972;
	wire [16-1:0] node8973;
	wire [16-1:0] node8974;
	wire [16-1:0] node8977;
	wire [16-1:0] node8980;
	wire [16-1:0] node8981;
	wire [16-1:0] node8985;
	wire [16-1:0] node8986;
	wire [16-1:0] node8988;
	wire [16-1:0] node8991;
	wire [16-1:0] node8992;
	wire [16-1:0] node8995;
	wire [16-1:0] node8998;
	wire [16-1:0] node8999;
	wire [16-1:0] node9000;
	wire [16-1:0] node9001;
	wire [16-1:0] node9002;
	wire [16-1:0] node9003;
	wire [16-1:0] node9004;
	wire [16-1:0] node9007;
	wire [16-1:0] node9010;
	wire [16-1:0] node9011;
	wire [16-1:0] node9014;
	wire [16-1:0] node9017;
	wire [16-1:0] node9018;
	wire [16-1:0] node9019;
	wire [16-1:0] node9023;
	wire [16-1:0] node9024;
	wire [16-1:0] node9027;
	wire [16-1:0] node9030;
	wire [16-1:0] node9031;
	wire [16-1:0] node9032;
	wire [16-1:0] node9033;
	wire [16-1:0] node9036;
	wire [16-1:0] node9039;
	wire [16-1:0] node9041;
	wire [16-1:0] node9044;
	wire [16-1:0] node9045;
	wire [16-1:0] node9046;
	wire [16-1:0] node9049;
	wire [16-1:0] node9052;
	wire [16-1:0] node9053;
	wire [16-1:0] node9056;
	wire [16-1:0] node9059;
	wire [16-1:0] node9060;
	wire [16-1:0] node9061;
	wire [16-1:0] node9062;
	wire [16-1:0] node9063;
	wire [16-1:0] node9066;
	wire [16-1:0] node9069;
	wire [16-1:0] node9070;
	wire [16-1:0] node9073;
	wire [16-1:0] node9076;
	wire [16-1:0] node9077;
	wire [16-1:0] node9078;
	wire [16-1:0] node9081;
	wire [16-1:0] node9084;
	wire [16-1:0] node9085;
	wire [16-1:0] node9088;
	wire [16-1:0] node9091;
	wire [16-1:0] node9092;
	wire [16-1:0] node9093;
	wire [16-1:0] node9094;
	wire [16-1:0] node9098;
	wire [16-1:0] node9099;
	wire [16-1:0] node9102;
	wire [16-1:0] node9105;
	wire [16-1:0] node9106;
	wire [16-1:0] node9107;
	wire [16-1:0] node9110;
	wire [16-1:0] node9113;
	wire [16-1:0] node9114;
	wire [16-1:0] node9117;
	wire [16-1:0] node9120;
	wire [16-1:0] node9121;
	wire [16-1:0] node9122;
	wire [16-1:0] node9123;
	wire [16-1:0] node9124;
	wire [16-1:0] node9125;
	wire [16-1:0] node9128;
	wire [16-1:0] node9131;
	wire [16-1:0] node9132;
	wire [16-1:0] node9135;
	wire [16-1:0] node9138;
	wire [16-1:0] node9139;
	wire [16-1:0] node9140;
	wire [16-1:0] node9143;
	wire [16-1:0] node9146;
	wire [16-1:0] node9147;
	wire [16-1:0] node9150;
	wire [16-1:0] node9153;
	wire [16-1:0] node9154;
	wire [16-1:0] node9155;
	wire [16-1:0] node9157;
	wire [16-1:0] node9160;
	wire [16-1:0] node9161;
	wire [16-1:0] node9164;
	wire [16-1:0] node9167;
	wire [16-1:0] node9168;
	wire [16-1:0] node9169;
	wire [16-1:0] node9172;
	wire [16-1:0] node9175;
	wire [16-1:0] node9176;
	wire [16-1:0] node9179;
	wire [16-1:0] node9182;
	wire [16-1:0] node9183;
	wire [16-1:0] node9184;
	wire [16-1:0] node9185;
	wire [16-1:0] node9187;
	wire [16-1:0] node9190;
	wire [16-1:0] node9191;
	wire [16-1:0] node9194;
	wire [16-1:0] node9197;
	wire [16-1:0] node9198;
	wire [16-1:0] node9199;
	wire [16-1:0] node9202;
	wire [16-1:0] node9205;
	wire [16-1:0] node9206;
	wire [16-1:0] node9209;
	wire [16-1:0] node9212;
	wire [16-1:0] node9213;
	wire [16-1:0] node9214;
	wire [16-1:0] node9215;
	wire [16-1:0] node9218;
	wire [16-1:0] node9221;
	wire [16-1:0] node9223;
	wire [16-1:0] node9226;
	wire [16-1:0] node9227;
	wire [16-1:0] node9228;
	wire [16-1:0] node9231;
	wire [16-1:0] node9234;
	wire [16-1:0] node9235;
	wire [16-1:0] node9238;
	wire [16-1:0] node9241;
	wire [16-1:0] node9242;
	wire [16-1:0] node9243;
	wire [16-1:0] node9244;
	wire [16-1:0] node9245;
	wire [16-1:0] node9246;
	wire [16-1:0] node9247;
	wire [16-1:0] node9248;
	wire [16-1:0] node9251;
	wire [16-1:0] node9254;
	wire [16-1:0] node9255;
	wire [16-1:0] node9258;
	wire [16-1:0] node9261;
	wire [16-1:0] node9262;
	wire [16-1:0] node9263;
	wire [16-1:0] node9266;
	wire [16-1:0] node9270;
	wire [16-1:0] node9271;
	wire [16-1:0] node9272;
	wire [16-1:0] node9273;
	wire [16-1:0] node9276;
	wire [16-1:0] node9279;
	wire [16-1:0] node9280;
	wire [16-1:0] node9283;
	wire [16-1:0] node9286;
	wire [16-1:0] node9287;
	wire [16-1:0] node9288;
	wire [16-1:0] node9291;
	wire [16-1:0] node9294;
	wire [16-1:0] node9295;
	wire [16-1:0] node9298;
	wire [16-1:0] node9301;
	wire [16-1:0] node9302;
	wire [16-1:0] node9303;
	wire [16-1:0] node9304;
	wire [16-1:0] node9305;
	wire [16-1:0] node9308;
	wire [16-1:0] node9311;
	wire [16-1:0] node9312;
	wire [16-1:0] node9315;
	wire [16-1:0] node9318;
	wire [16-1:0] node9319;
	wire [16-1:0] node9320;
	wire [16-1:0] node9323;
	wire [16-1:0] node9326;
	wire [16-1:0] node9327;
	wire [16-1:0] node9331;
	wire [16-1:0] node9332;
	wire [16-1:0] node9333;
	wire [16-1:0] node9334;
	wire [16-1:0] node9337;
	wire [16-1:0] node9340;
	wire [16-1:0] node9341;
	wire [16-1:0] node9344;
	wire [16-1:0] node9347;
	wire [16-1:0] node9348;
	wire [16-1:0] node9349;
	wire [16-1:0] node9352;
	wire [16-1:0] node9355;
	wire [16-1:0] node9356;
	wire [16-1:0] node9359;
	wire [16-1:0] node9362;
	wire [16-1:0] node9363;
	wire [16-1:0] node9364;
	wire [16-1:0] node9365;
	wire [16-1:0] node9366;
	wire [16-1:0] node9367;
	wire [16-1:0] node9371;
	wire [16-1:0] node9373;
	wire [16-1:0] node9376;
	wire [16-1:0] node9377;
	wire [16-1:0] node9378;
	wire [16-1:0] node9381;
	wire [16-1:0] node9384;
	wire [16-1:0] node9385;
	wire [16-1:0] node9389;
	wire [16-1:0] node9390;
	wire [16-1:0] node9391;
	wire [16-1:0] node9392;
	wire [16-1:0] node9395;
	wire [16-1:0] node9398;
	wire [16-1:0] node9399;
	wire [16-1:0] node9402;
	wire [16-1:0] node9405;
	wire [16-1:0] node9406;
	wire [16-1:0] node9407;
	wire [16-1:0] node9410;
	wire [16-1:0] node9413;
	wire [16-1:0] node9414;
	wire [16-1:0] node9417;
	wire [16-1:0] node9420;
	wire [16-1:0] node9421;
	wire [16-1:0] node9422;
	wire [16-1:0] node9423;
	wire [16-1:0] node9424;
	wire [16-1:0] node9427;
	wire [16-1:0] node9430;
	wire [16-1:0] node9431;
	wire [16-1:0] node9434;
	wire [16-1:0] node9437;
	wire [16-1:0] node9438;
	wire [16-1:0] node9439;
	wire [16-1:0] node9442;
	wire [16-1:0] node9445;
	wire [16-1:0] node9446;
	wire [16-1:0] node9449;
	wire [16-1:0] node9452;
	wire [16-1:0] node9453;
	wire [16-1:0] node9454;
	wire [16-1:0] node9455;
	wire [16-1:0] node9458;
	wire [16-1:0] node9461;
	wire [16-1:0] node9462;
	wire [16-1:0] node9465;
	wire [16-1:0] node9468;
	wire [16-1:0] node9469;
	wire [16-1:0] node9470;
	wire [16-1:0] node9473;
	wire [16-1:0] node9476;
	wire [16-1:0] node9477;
	wire [16-1:0] node9480;
	wire [16-1:0] node9483;
	wire [16-1:0] node9484;
	wire [16-1:0] node9485;
	wire [16-1:0] node9486;
	wire [16-1:0] node9487;
	wire [16-1:0] node9488;
	wire [16-1:0] node9489;
	wire [16-1:0] node9492;
	wire [16-1:0] node9495;
	wire [16-1:0] node9497;
	wire [16-1:0] node9500;
	wire [16-1:0] node9501;
	wire [16-1:0] node9502;
	wire [16-1:0] node9505;
	wire [16-1:0] node9508;
	wire [16-1:0] node9509;
	wire [16-1:0] node9512;
	wire [16-1:0] node9515;
	wire [16-1:0] node9516;
	wire [16-1:0] node9517;
	wire [16-1:0] node9518;
	wire [16-1:0] node9521;
	wire [16-1:0] node9524;
	wire [16-1:0] node9525;
	wire [16-1:0] node9528;
	wire [16-1:0] node9531;
	wire [16-1:0] node9532;
	wire [16-1:0] node9533;
	wire [16-1:0] node9536;
	wire [16-1:0] node9539;
	wire [16-1:0] node9540;
	wire [16-1:0] node9543;
	wire [16-1:0] node9546;
	wire [16-1:0] node9547;
	wire [16-1:0] node9548;
	wire [16-1:0] node9549;
	wire [16-1:0] node9551;
	wire [16-1:0] node9554;
	wire [16-1:0] node9555;
	wire [16-1:0] node9558;
	wire [16-1:0] node9561;
	wire [16-1:0] node9562;
	wire [16-1:0] node9563;
	wire [16-1:0] node9566;
	wire [16-1:0] node9569;
	wire [16-1:0] node9570;
	wire [16-1:0] node9573;
	wire [16-1:0] node9576;
	wire [16-1:0] node9577;
	wire [16-1:0] node9578;
	wire [16-1:0] node9579;
	wire [16-1:0] node9582;
	wire [16-1:0] node9585;
	wire [16-1:0] node9586;
	wire [16-1:0] node9589;
	wire [16-1:0] node9592;
	wire [16-1:0] node9593;
	wire [16-1:0] node9595;
	wire [16-1:0] node9598;
	wire [16-1:0] node9599;
	wire [16-1:0] node9602;
	wire [16-1:0] node9605;
	wire [16-1:0] node9606;
	wire [16-1:0] node9607;
	wire [16-1:0] node9608;
	wire [16-1:0] node9609;
	wire [16-1:0] node9610;
	wire [16-1:0] node9613;
	wire [16-1:0] node9616;
	wire [16-1:0] node9617;
	wire [16-1:0] node9621;
	wire [16-1:0] node9622;
	wire [16-1:0] node9623;
	wire [16-1:0] node9626;
	wire [16-1:0] node9629;
	wire [16-1:0] node9630;
	wire [16-1:0] node9633;
	wire [16-1:0] node9636;
	wire [16-1:0] node9637;
	wire [16-1:0] node9638;
	wire [16-1:0] node9639;
	wire [16-1:0] node9642;
	wire [16-1:0] node9645;
	wire [16-1:0] node9647;
	wire [16-1:0] node9650;
	wire [16-1:0] node9651;
	wire [16-1:0] node9652;
	wire [16-1:0] node9655;
	wire [16-1:0] node9658;
	wire [16-1:0] node9659;
	wire [16-1:0] node9662;
	wire [16-1:0] node9665;
	wire [16-1:0] node9666;
	wire [16-1:0] node9667;
	wire [16-1:0] node9668;
	wire [16-1:0] node9669;
	wire [16-1:0] node9672;
	wire [16-1:0] node9675;
	wire [16-1:0] node9676;
	wire [16-1:0] node9679;
	wire [16-1:0] node9682;
	wire [16-1:0] node9683;
	wire [16-1:0] node9684;
	wire [16-1:0] node9687;
	wire [16-1:0] node9690;
	wire [16-1:0] node9691;
	wire [16-1:0] node9695;
	wire [16-1:0] node9696;
	wire [16-1:0] node9697;
	wire [16-1:0] node9698;
	wire [16-1:0] node9701;
	wire [16-1:0] node9704;
	wire [16-1:0] node9705;
	wire [16-1:0] node9708;
	wire [16-1:0] node9711;
	wire [16-1:0] node9712;
	wire [16-1:0] node9713;
	wire [16-1:0] node9716;
	wire [16-1:0] node9719;
	wire [16-1:0] node9721;
	wire [16-1:0] node9724;
	wire [16-1:0] node9725;
	wire [16-1:0] node9726;
	wire [16-1:0] node9727;
	wire [16-1:0] node9728;
	wire [16-1:0] node9729;
	wire [16-1:0] node9730;
	wire [16-1:0] node9731;
	wire [16-1:0] node9732;
	wire [16-1:0] node9733;
	wire [16-1:0] node9736;
	wire [16-1:0] node9739;
	wire [16-1:0] node9740;
	wire [16-1:0] node9743;
	wire [16-1:0] node9746;
	wire [16-1:0] node9747;
	wire [16-1:0] node9748;
	wire [16-1:0] node9751;
	wire [16-1:0] node9754;
	wire [16-1:0] node9755;
	wire [16-1:0] node9758;
	wire [16-1:0] node9761;
	wire [16-1:0] node9762;
	wire [16-1:0] node9763;
	wire [16-1:0] node9764;
	wire [16-1:0] node9767;
	wire [16-1:0] node9770;
	wire [16-1:0] node9771;
	wire [16-1:0] node9774;
	wire [16-1:0] node9777;
	wire [16-1:0] node9778;
	wire [16-1:0] node9779;
	wire [16-1:0] node9783;
	wire [16-1:0] node9784;
	wire [16-1:0] node9788;
	wire [16-1:0] node9789;
	wire [16-1:0] node9790;
	wire [16-1:0] node9791;
	wire [16-1:0] node9792;
	wire [16-1:0] node9796;
	wire [16-1:0] node9797;
	wire [16-1:0] node9800;
	wire [16-1:0] node9803;
	wire [16-1:0] node9804;
	wire [16-1:0] node9805;
	wire [16-1:0] node9808;
	wire [16-1:0] node9811;
	wire [16-1:0] node9812;
	wire [16-1:0] node9815;
	wire [16-1:0] node9818;
	wire [16-1:0] node9819;
	wire [16-1:0] node9820;
	wire [16-1:0] node9821;
	wire [16-1:0] node9824;
	wire [16-1:0] node9827;
	wire [16-1:0] node9828;
	wire [16-1:0] node9831;
	wire [16-1:0] node9834;
	wire [16-1:0] node9835;
	wire [16-1:0] node9836;
	wire [16-1:0] node9839;
	wire [16-1:0] node9842;
	wire [16-1:0] node9843;
	wire [16-1:0] node9846;
	wire [16-1:0] node9849;
	wire [16-1:0] node9850;
	wire [16-1:0] node9851;
	wire [16-1:0] node9852;
	wire [16-1:0] node9853;
	wire [16-1:0] node9854;
	wire [16-1:0] node9857;
	wire [16-1:0] node9860;
	wire [16-1:0] node9861;
	wire [16-1:0] node9864;
	wire [16-1:0] node9867;
	wire [16-1:0] node9868;
	wire [16-1:0] node9869;
	wire [16-1:0] node9873;
	wire [16-1:0] node9874;
	wire [16-1:0] node9877;
	wire [16-1:0] node9880;
	wire [16-1:0] node9881;
	wire [16-1:0] node9882;
	wire [16-1:0] node9883;
	wire [16-1:0] node9887;
	wire [16-1:0] node9888;
	wire [16-1:0] node9891;
	wire [16-1:0] node9894;
	wire [16-1:0] node9895;
	wire [16-1:0] node9896;
	wire [16-1:0] node9899;
	wire [16-1:0] node9902;
	wire [16-1:0] node9904;
	wire [16-1:0] node9907;
	wire [16-1:0] node9908;
	wire [16-1:0] node9909;
	wire [16-1:0] node9910;
	wire [16-1:0] node9911;
	wire [16-1:0] node9914;
	wire [16-1:0] node9917;
	wire [16-1:0] node9918;
	wire [16-1:0] node9921;
	wire [16-1:0] node9924;
	wire [16-1:0] node9925;
	wire [16-1:0] node9926;
	wire [16-1:0] node9929;
	wire [16-1:0] node9932;
	wire [16-1:0] node9933;
	wire [16-1:0] node9936;
	wire [16-1:0] node9939;
	wire [16-1:0] node9940;
	wire [16-1:0] node9941;
	wire [16-1:0] node9942;
	wire [16-1:0] node9945;
	wire [16-1:0] node9948;
	wire [16-1:0] node9949;
	wire [16-1:0] node9952;
	wire [16-1:0] node9955;
	wire [16-1:0] node9956;
	wire [16-1:0] node9957;
	wire [16-1:0] node9960;
	wire [16-1:0] node9963;
	wire [16-1:0] node9964;
	wire [16-1:0] node9968;
	wire [16-1:0] node9969;
	wire [16-1:0] node9970;
	wire [16-1:0] node9971;
	wire [16-1:0] node9972;
	wire [16-1:0] node9973;
	wire [16-1:0] node9974;
	wire [16-1:0] node9977;
	wire [16-1:0] node9980;
	wire [16-1:0] node9981;
	wire [16-1:0] node9984;
	wire [16-1:0] node9987;
	wire [16-1:0] node9988;
	wire [16-1:0] node9989;
	wire [16-1:0] node9992;
	wire [16-1:0] node9995;
	wire [16-1:0] node9996;
	wire [16-1:0] node9999;
	wire [16-1:0] node10002;
	wire [16-1:0] node10003;
	wire [16-1:0] node10004;
	wire [16-1:0] node10005;
	wire [16-1:0] node10008;
	wire [16-1:0] node10011;
	wire [16-1:0] node10012;
	wire [16-1:0] node10015;
	wire [16-1:0] node10018;
	wire [16-1:0] node10019;
	wire [16-1:0] node10020;
	wire [16-1:0] node10023;
	wire [16-1:0] node10026;
	wire [16-1:0] node10028;
	wire [16-1:0] node10031;
	wire [16-1:0] node10032;
	wire [16-1:0] node10033;
	wire [16-1:0] node10034;
	wire [16-1:0] node10035;
	wire [16-1:0] node10039;
	wire [16-1:0] node10040;
	wire [16-1:0] node10043;
	wire [16-1:0] node10046;
	wire [16-1:0] node10047;
	wire [16-1:0] node10048;
	wire [16-1:0] node10051;
	wire [16-1:0] node10054;
	wire [16-1:0] node10055;
	wire [16-1:0] node10058;
	wire [16-1:0] node10061;
	wire [16-1:0] node10062;
	wire [16-1:0] node10063;
	wire [16-1:0] node10064;
	wire [16-1:0] node10067;
	wire [16-1:0] node10070;
	wire [16-1:0] node10071;
	wire [16-1:0] node10074;
	wire [16-1:0] node10077;
	wire [16-1:0] node10078;
	wire [16-1:0] node10080;
	wire [16-1:0] node10083;
	wire [16-1:0] node10084;
	wire [16-1:0] node10087;
	wire [16-1:0] node10090;
	wire [16-1:0] node10091;
	wire [16-1:0] node10092;
	wire [16-1:0] node10093;
	wire [16-1:0] node10094;
	wire [16-1:0] node10095;
	wire [16-1:0] node10098;
	wire [16-1:0] node10101;
	wire [16-1:0] node10102;
	wire [16-1:0] node10105;
	wire [16-1:0] node10108;
	wire [16-1:0] node10109;
	wire [16-1:0] node10110;
	wire [16-1:0] node10113;
	wire [16-1:0] node10116;
	wire [16-1:0] node10117;
	wire [16-1:0] node10120;
	wire [16-1:0] node10123;
	wire [16-1:0] node10124;
	wire [16-1:0] node10125;
	wire [16-1:0] node10126;
	wire [16-1:0] node10129;
	wire [16-1:0] node10132;
	wire [16-1:0] node10133;
	wire [16-1:0] node10136;
	wire [16-1:0] node10139;
	wire [16-1:0] node10140;
	wire [16-1:0] node10141;
	wire [16-1:0] node10144;
	wire [16-1:0] node10147;
	wire [16-1:0] node10148;
	wire [16-1:0] node10151;
	wire [16-1:0] node10154;
	wire [16-1:0] node10155;
	wire [16-1:0] node10156;
	wire [16-1:0] node10157;
	wire [16-1:0] node10159;
	wire [16-1:0] node10162;
	wire [16-1:0] node10163;
	wire [16-1:0] node10166;
	wire [16-1:0] node10169;
	wire [16-1:0] node10170;
	wire [16-1:0] node10171;
	wire [16-1:0] node10174;
	wire [16-1:0] node10177;
	wire [16-1:0] node10178;
	wire [16-1:0] node10181;
	wire [16-1:0] node10184;
	wire [16-1:0] node10185;
	wire [16-1:0] node10186;
	wire [16-1:0] node10187;
	wire [16-1:0] node10190;
	wire [16-1:0] node10193;
	wire [16-1:0] node10194;
	wire [16-1:0] node10197;
	wire [16-1:0] node10200;
	wire [16-1:0] node10201;
	wire [16-1:0] node10202;
	wire [16-1:0] node10205;
	wire [16-1:0] node10208;
	wire [16-1:0] node10209;
	wire [16-1:0] node10212;
	wire [16-1:0] node10215;
	wire [16-1:0] node10216;
	wire [16-1:0] node10217;
	wire [16-1:0] node10218;
	wire [16-1:0] node10219;
	wire [16-1:0] node10220;
	wire [16-1:0] node10221;
	wire [16-1:0] node10222;
	wire [16-1:0] node10225;
	wire [16-1:0] node10228;
	wire [16-1:0] node10229;
	wire [16-1:0] node10232;
	wire [16-1:0] node10235;
	wire [16-1:0] node10236;
	wire [16-1:0] node10237;
	wire [16-1:0] node10240;
	wire [16-1:0] node10243;
	wire [16-1:0] node10244;
	wire [16-1:0] node10247;
	wire [16-1:0] node10250;
	wire [16-1:0] node10251;
	wire [16-1:0] node10252;
	wire [16-1:0] node10253;
	wire [16-1:0] node10256;
	wire [16-1:0] node10259;
	wire [16-1:0] node10260;
	wire [16-1:0] node10263;
	wire [16-1:0] node10266;
	wire [16-1:0] node10267;
	wire [16-1:0] node10268;
	wire [16-1:0] node10271;
	wire [16-1:0] node10274;
	wire [16-1:0] node10275;
	wire [16-1:0] node10278;
	wire [16-1:0] node10281;
	wire [16-1:0] node10282;
	wire [16-1:0] node10283;
	wire [16-1:0] node10284;
	wire [16-1:0] node10285;
	wire [16-1:0] node10288;
	wire [16-1:0] node10291;
	wire [16-1:0] node10294;
	wire [16-1:0] node10295;
	wire [16-1:0] node10296;
	wire [16-1:0] node10299;
	wire [16-1:0] node10302;
	wire [16-1:0] node10303;
	wire [16-1:0] node10306;
	wire [16-1:0] node10309;
	wire [16-1:0] node10310;
	wire [16-1:0] node10311;
	wire [16-1:0] node10313;
	wire [16-1:0] node10316;
	wire [16-1:0] node10317;
	wire [16-1:0] node10320;
	wire [16-1:0] node10323;
	wire [16-1:0] node10324;
	wire [16-1:0] node10325;
	wire [16-1:0] node10328;
	wire [16-1:0] node10332;
	wire [16-1:0] node10333;
	wire [16-1:0] node10334;
	wire [16-1:0] node10335;
	wire [16-1:0] node10336;
	wire [16-1:0] node10337;
	wire [16-1:0] node10340;
	wire [16-1:0] node10343;
	wire [16-1:0] node10344;
	wire [16-1:0] node10347;
	wire [16-1:0] node10350;
	wire [16-1:0] node10351;
	wire [16-1:0] node10353;
	wire [16-1:0] node10356;
	wire [16-1:0] node10357;
	wire [16-1:0] node10360;
	wire [16-1:0] node10363;
	wire [16-1:0] node10364;
	wire [16-1:0] node10365;
	wire [16-1:0] node10366;
	wire [16-1:0] node10369;
	wire [16-1:0] node10372;
	wire [16-1:0] node10373;
	wire [16-1:0] node10377;
	wire [16-1:0] node10378;
	wire [16-1:0] node10379;
	wire [16-1:0] node10382;
	wire [16-1:0] node10385;
	wire [16-1:0] node10386;
	wire [16-1:0] node10389;
	wire [16-1:0] node10392;
	wire [16-1:0] node10393;
	wire [16-1:0] node10394;
	wire [16-1:0] node10395;
	wire [16-1:0] node10397;
	wire [16-1:0] node10400;
	wire [16-1:0] node10401;
	wire [16-1:0] node10404;
	wire [16-1:0] node10407;
	wire [16-1:0] node10408;
	wire [16-1:0] node10409;
	wire [16-1:0] node10412;
	wire [16-1:0] node10415;
	wire [16-1:0] node10416;
	wire [16-1:0] node10419;
	wire [16-1:0] node10422;
	wire [16-1:0] node10423;
	wire [16-1:0] node10424;
	wire [16-1:0] node10425;
	wire [16-1:0] node10429;
	wire [16-1:0] node10430;
	wire [16-1:0] node10433;
	wire [16-1:0] node10436;
	wire [16-1:0] node10437;
	wire [16-1:0] node10438;
	wire [16-1:0] node10441;
	wire [16-1:0] node10444;
	wire [16-1:0] node10445;
	wire [16-1:0] node10448;
	wire [16-1:0] node10451;
	wire [16-1:0] node10452;
	wire [16-1:0] node10453;
	wire [16-1:0] node10454;
	wire [16-1:0] node10455;
	wire [16-1:0] node10456;
	wire [16-1:0] node10457;
	wire [16-1:0] node10460;
	wire [16-1:0] node10463;
	wire [16-1:0] node10464;
	wire [16-1:0] node10467;
	wire [16-1:0] node10470;
	wire [16-1:0] node10471;
	wire [16-1:0] node10472;
	wire [16-1:0] node10475;
	wire [16-1:0] node10478;
	wire [16-1:0] node10479;
	wire [16-1:0] node10482;
	wire [16-1:0] node10485;
	wire [16-1:0] node10486;
	wire [16-1:0] node10487;
	wire [16-1:0] node10488;
	wire [16-1:0] node10491;
	wire [16-1:0] node10494;
	wire [16-1:0] node10495;
	wire [16-1:0] node10498;
	wire [16-1:0] node10501;
	wire [16-1:0] node10502;
	wire [16-1:0] node10503;
	wire [16-1:0] node10506;
	wire [16-1:0] node10509;
	wire [16-1:0] node10510;
	wire [16-1:0] node10513;
	wire [16-1:0] node10516;
	wire [16-1:0] node10517;
	wire [16-1:0] node10518;
	wire [16-1:0] node10519;
	wire [16-1:0] node10520;
	wire [16-1:0] node10524;
	wire [16-1:0] node10525;
	wire [16-1:0] node10528;
	wire [16-1:0] node10531;
	wire [16-1:0] node10532;
	wire [16-1:0] node10534;
	wire [16-1:0] node10537;
	wire [16-1:0] node10538;
	wire [16-1:0] node10541;
	wire [16-1:0] node10544;
	wire [16-1:0] node10545;
	wire [16-1:0] node10546;
	wire [16-1:0] node10547;
	wire [16-1:0] node10550;
	wire [16-1:0] node10553;
	wire [16-1:0] node10554;
	wire [16-1:0] node10557;
	wire [16-1:0] node10560;
	wire [16-1:0] node10561;
	wire [16-1:0] node10562;
	wire [16-1:0] node10565;
	wire [16-1:0] node10568;
	wire [16-1:0] node10569;
	wire [16-1:0] node10572;
	wire [16-1:0] node10575;
	wire [16-1:0] node10576;
	wire [16-1:0] node10577;
	wire [16-1:0] node10578;
	wire [16-1:0] node10579;
	wire [16-1:0] node10580;
	wire [16-1:0] node10583;
	wire [16-1:0] node10586;
	wire [16-1:0] node10587;
	wire [16-1:0] node10590;
	wire [16-1:0] node10593;
	wire [16-1:0] node10594;
	wire [16-1:0] node10595;
	wire [16-1:0] node10598;
	wire [16-1:0] node10601;
	wire [16-1:0] node10602;
	wire [16-1:0] node10605;
	wire [16-1:0] node10608;
	wire [16-1:0] node10609;
	wire [16-1:0] node10610;
	wire [16-1:0] node10611;
	wire [16-1:0] node10614;
	wire [16-1:0] node10617;
	wire [16-1:0] node10618;
	wire [16-1:0] node10621;
	wire [16-1:0] node10624;
	wire [16-1:0] node10625;
	wire [16-1:0] node10626;
	wire [16-1:0] node10629;
	wire [16-1:0] node10632;
	wire [16-1:0] node10633;
	wire [16-1:0] node10636;
	wire [16-1:0] node10639;
	wire [16-1:0] node10640;
	wire [16-1:0] node10641;
	wire [16-1:0] node10642;
	wire [16-1:0] node10643;
	wire [16-1:0] node10646;
	wire [16-1:0] node10649;
	wire [16-1:0] node10650;
	wire [16-1:0] node10653;
	wire [16-1:0] node10656;
	wire [16-1:0] node10657;
	wire [16-1:0] node10658;
	wire [16-1:0] node10661;
	wire [16-1:0] node10664;
	wire [16-1:0] node10666;
	wire [16-1:0] node10669;
	wire [16-1:0] node10670;
	wire [16-1:0] node10671;
	wire [16-1:0] node10673;
	wire [16-1:0] node10676;
	wire [16-1:0] node10677;
	wire [16-1:0] node10680;
	wire [16-1:0] node10683;
	wire [16-1:0] node10684;
	wire [16-1:0] node10685;
	wire [16-1:0] node10688;
	wire [16-1:0] node10691;
	wire [16-1:0] node10692;
	wire [16-1:0] node10695;
	wire [16-1:0] node10698;
	wire [16-1:0] node10699;
	wire [16-1:0] node10700;
	wire [16-1:0] node10701;
	wire [16-1:0] node10702;
	wire [16-1:0] node10703;
	wire [16-1:0] node10704;
	wire [16-1:0] node10705;
	wire [16-1:0] node10706;
	wire [16-1:0] node10709;
	wire [16-1:0] node10712;
	wire [16-1:0] node10713;
	wire [16-1:0] node10716;
	wire [16-1:0] node10719;
	wire [16-1:0] node10720;
	wire [16-1:0] node10721;
	wire [16-1:0] node10724;
	wire [16-1:0] node10727;
	wire [16-1:0] node10728;
	wire [16-1:0] node10731;
	wire [16-1:0] node10734;
	wire [16-1:0] node10735;
	wire [16-1:0] node10736;
	wire [16-1:0] node10737;
	wire [16-1:0] node10740;
	wire [16-1:0] node10743;
	wire [16-1:0] node10744;
	wire [16-1:0] node10747;
	wire [16-1:0] node10750;
	wire [16-1:0] node10751;
	wire [16-1:0] node10752;
	wire [16-1:0] node10755;
	wire [16-1:0] node10758;
	wire [16-1:0] node10759;
	wire [16-1:0] node10763;
	wire [16-1:0] node10764;
	wire [16-1:0] node10765;
	wire [16-1:0] node10766;
	wire [16-1:0] node10767;
	wire [16-1:0] node10770;
	wire [16-1:0] node10773;
	wire [16-1:0] node10774;
	wire [16-1:0] node10778;
	wire [16-1:0] node10779;
	wire [16-1:0] node10780;
	wire [16-1:0] node10783;
	wire [16-1:0] node10786;
	wire [16-1:0] node10787;
	wire [16-1:0] node10790;
	wire [16-1:0] node10793;
	wire [16-1:0] node10794;
	wire [16-1:0] node10795;
	wire [16-1:0] node10796;
	wire [16-1:0] node10799;
	wire [16-1:0] node10802;
	wire [16-1:0] node10803;
	wire [16-1:0] node10806;
	wire [16-1:0] node10809;
	wire [16-1:0] node10810;
	wire [16-1:0] node10812;
	wire [16-1:0] node10815;
	wire [16-1:0] node10816;
	wire [16-1:0] node10819;
	wire [16-1:0] node10822;
	wire [16-1:0] node10823;
	wire [16-1:0] node10824;
	wire [16-1:0] node10825;
	wire [16-1:0] node10826;
	wire [16-1:0] node10827;
	wire [16-1:0] node10831;
	wire [16-1:0] node10832;
	wire [16-1:0] node10835;
	wire [16-1:0] node10838;
	wire [16-1:0] node10839;
	wire [16-1:0] node10840;
	wire [16-1:0] node10843;
	wire [16-1:0] node10846;
	wire [16-1:0] node10847;
	wire [16-1:0] node10850;
	wire [16-1:0] node10853;
	wire [16-1:0] node10854;
	wire [16-1:0] node10855;
	wire [16-1:0] node10856;
	wire [16-1:0] node10859;
	wire [16-1:0] node10862;
	wire [16-1:0] node10863;
	wire [16-1:0] node10866;
	wire [16-1:0] node10869;
	wire [16-1:0] node10870;
	wire [16-1:0] node10871;
	wire [16-1:0] node10874;
	wire [16-1:0] node10877;
	wire [16-1:0] node10878;
	wire [16-1:0] node10881;
	wire [16-1:0] node10884;
	wire [16-1:0] node10885;
	wire [16-1:0] node10886;
	wire [16-1:0] node10887;
	wire [16-1:0] node10888;
	wire [16-1:0] node10891;
	wire [16-1:0] node10894;
	wire [16-1:0] node10895;
	wire [16-1:0] node10899;
	wire [16-1:0] node10900;
	wire [16-1:0] node10901;
	wire [16-1:0] node10904;
	wire [16-1:0] node10907;
	wire [16-1:0] node10908;
	wire [16-1:0] node10911;
	wire [16-1:0] node10914;
	wire [16-1:0] node10915;
	wire [16-1:0] node10916;
	wire [16-1:0] node10917;
	wire [16-1:0] node10920;
	wire [16-1:0] node10923;
	wire [16-1:0] node10924;
	wire [16-1:0] node10927;
	wire [16-1:0] node10930;
	wire [16-1:0] node10931;
	wire [16-1:0] node10932;
	wire [16-1:0] node10935;
	wire [16-1:0] node10938;
	wire [16-1:0] node10939;
	wire [16-1:0] node10942;
	wire [16-1:0] node10945;
	wire [16-1:0] node10946;
	wire [16-1:0] node10947;
	wire [16-1:0] node10948;
	wire [16-1:0] node10949;
	wire [16-1:0] node10950;
	wire [16-1:0] node10951;
	wire [16-1:0] node10954;
	wire [16-1:0] node10957;
	wire [16-1:0] node10958;
	wire [16-1:0] node10961;
	wire [16-1:0] node10964;
	wire [16-1:0] node10965;
	wire [16-1:0] node10966;
	wire [16-1:0] node10969;
	wire [16-1:0] node10972;
	wire [16-1:0] node10973;
	wire [16-1:0] node10976;
	wire [16-1:0] node10979;
	wire [16-1:0] node10980;
	wire [16-1:0] node10981;
	wire [16-1:0] node10982;
	wire [16-1:0] node10985;
	wire [16-1:0] node10988;
	wire [16-1:0] node10989;
	wire [16-1:0] node10992;
	wire [16-1:0] node10995;
	wire [16-1:0] node10996;
	wire [16-1:0] node10997;
	wire [16-1:0] node11001;
	wire [16-1:0] node11002;
	wire [16-1:0] node11005;
	wire [16-1:0] node11008;
	wire [16-1:0] node11009;
	wire [16-1:0] node11010;
	wire [16-1:0] node11011;
	wire [16-1:0] node11012;
	wire [16-1:0] node11015;
	wire [16-1:0] node11018;
	wire [16-1:0] node11019;
	wire [16-1:0] node11022;
	wire [16-1:0] node11025;
	wire [16-1:0] node11026;
	wire [16-1:0] node11027;
	wire [16-1:0] node11030;
	wire [16-1:0] node11033;
	wire [16-1:0] node11034;
	wire [16-1:0] node11037;
	wire [16-1:0] node11040;
	wire [16-1:0] node11041;
	wire [16-1:0] node11042;
	wire [16-1:0] node11043;
	wire [16-1:0] node11046;
	wire [16-1:0] node11049;
	wire [16-1:0] node11050;
	wire [16-1:0] node11053;
	wire [16-1:0] node11056;
	wire [16-1:0] node11057;
	wire [16-1:0] node11058;
	wire [16-1:0] node11061;
	wire [16-1:0] node11064;
	wire [16-1:0] node11065;
	wire [16-1:0] node11068;
	wire [16-1:0] node11071;
	wire [16-1:0] node11072;
	wire [16-1:0] node11073;
	wire [16-1:0] node11074;
	wire [16-1:0] node11075;
	wire [16-1:0] node11076;
	wire [16-1:0] node11079;
	wire [16-1:0] node11082;
	wire [16-1:0] node11083;
	wire [16-1:0] node11087;
	wire [16-1:0] node11088;
	wire [16-1:0] node11089;
	wire [16-1:0] node11092;
	wire [16-1:0] node11095;
	wire [16-1:0] node11096;
	wire [16-1:0] node11099;
	wire [16-1:0] node11102;
	wire [16-1:0] node11103;
	wire [16-1:0] node11104;
	wire [16-1:0] node11105;
	wire [16-1:0] node11108;
	wire [16-1:0] node11111;
	wire [16-1:0] node11112;
	wire [16-1:0] node11115;
	wire [16-1:0] node11118;
	wire [16-1:0] node11119;
	wire [16-1:0] node11120;
	wire [16-1:0] node11123;
	wire [16-1:0] node11126;
	wire [16-1:0] node11129;
	wire [16-1:0] node11130;
	wire [16-1:0] node11131;
	wire [16-1:0] node11132;
	wire [16-1:0] node11135;
	wire [16-1:0] node11136;
	wire [16-1:0] node11139;
	wire [16-1:0] node11142;
	wire [16-1:0] node11143;
	wire [16-1:0] node11144;
	wire [16-1:0] node11147;
	wire [16-1:0] node11150;
	wire [16-1:0] node11152;
	wire [16-1:0] node11155;
	wire [16-1:0] node11156;
	wire [16-1:0] node11157;
	wire [16-1:0] node11158;
	wire [16-1:0] node11161;
	wire [16-1:0] node11164;
	wire [16-1:0] node11165;
	wire [16-1:0] node11168;
	wire [16-1:0] node11171;
	wire [16-1:0] node11172;
	wire [16-1:0] node11173;
	wire [16-1:0] node11176;
	wire [16-1:0] node11179;
	wire [16-1:0] node11181;
	wire [16-1:0] node11184;
	wire [16-1:0] node11185;
	wire [16-1:0] node11186;
	wire [16-1:0] node11187;
	wire [16-1:0] node11188;
	wire [16-1:0] node11189;
	wire [16-1:0] node11190;
	wire [16-1:0] node11191;
	wire [16-1:0] node11194;
	wire [16-1:0] node11197;
	wire [16-1:0] node11198;
	wire [16-1:0] node11202;
	wire [16-1:0] node11203;
	wire [16-1:0] node11204;
	wire [16-1:0] node11207;
	wire [16-1:0] node11210;
	wire [16-1:0] node11211;
	wire [16-1:0] node11214;
	wire [16-1:0] node11217;
	wire [16-1:0] node11218;
	wire [16-1:0] node11219;
	wire [16-1:0] node11220;
	wire [16-1:0] node11223;
	wire [16-1:0] node11226;
	wire [16-1:0] node11227;
	wire [16-1:0] node11230;
	wire [16-1:0] node11233;
	wire [16-1:0] node11234;
	wire [16-1:0] node11235;
	wire [16-1:0] node11238;
	wire [16-1:0] node11241;
	wire [16-1:0] node11242;
	wire [16-1:0] node11245;
	wire [16-1:0] node11248;
	wire [16-1:0] node11249;
	wire [16-1:0] node11250;
	wire [16-1:0] node11251;
	wire [16-1:0] node11252;
	wire [16-1:0] node11255;
	wire [16-1:0] node11258;
	wire [16-1:0] node11259;
	wire [16-1:0] node11262;
	wire [16-1:0] node11265;
	wire [16-1:0] node11266;
	wire [16-1:0] node11267;
	wire [16-1:0] node11270;
	wire [16-1:0] node11273;
	wire [16-1:0] node11275;
	wire [16-1:0] node11278;
	wire [16-1:0] node11279;
	wire [16-1:0] node11280;
	wire [16-1:0] node11282;
	wire [16-1:0] node11285;
	wire [16-1:0] node11286;
	wire [16-1:0] node11289;
	wire [16-1:0] node11292;
	wire [16-1:0] node11293;
	wire [16-1:0] node11295;
	wire [16-1:0] node11298;
	wire [16-1:0] node11299;
	wire [16-1:0] node11302;
	wire [16-1:0] node11305;
	wire [16-1:0] node11306;
	wire [16-1:0] node11307;
	wire [16-1:0] node11308;
	wire [16-1:0] node11309;
	wire [16-1:0] node11310;
	wire [16-1:0] node11313;
	wire [16-1:0] node11316;
	wire [16-1:0] node11317;
	wire [16-1:0] node11320;
	wire [16-1:0] node11323;
	wire [16-1:0] node11324;
	wire [16-1:0] node11327;
	wire [16-1:0] node11328;
	wire [16-1:0] node11331;
	wire [16-1:0] node11334;
	wire [16-1:0] node11335;
	wire [16-1:0] node11336;
	wire [16-1:0] node11337;
	wire [16-1:0] node11340;
	wire [16-1:0] node11343;
	wire [16-1:0] node11344;
	wire [16-1:0] node11347;
	wire [16-1:0] node11350;
	wire [16-1:0] node11351;
	wire [16-1:0] node11352;
	wire [16-1:0] node11355;
	wire [16-1:0] node11358;
	wire [16-1:0] node11359;
	wire [16-1:0] node11363;
	wire [16-1:0] node11364;
	wire [16-1:0] node11365;
	wire [16-1:0] node11366;
	wire [16-1:0] node11367;
	wire [16-1:0] node11370;
	wire [16-1:0] node11373;
	wire [16-1:0] node11374;
	wire [16-1:0] node11377;
	wire [16-1:0] node11380;
	wire [16-1:0] node11381;
	wire [16-1:0] node11382;
	wire [16-1:0] node11385;
	wire [16-1:0] node11388;
	wire [16-1:0] node11389;
	wire [16-1:0] node11392;
	wire [16-1:0] node11395;
	wire [16-1:0] node11396;
	wire [16-1:0] node11397;
	wire [16-1:0] node11398;
	wire [16-1:0] node11401;
	wire [16-1:0] node11404;
	wire [16-1:0] node11405;
	wire [16-1:0] node11409;
	wire [16-1:0] node11410;
	wire [16-1:0] node11411;
	wire [16-1:0] node11414;
	wire [16-1:0] node11417;
	wire [16-1:0] node11418;
	wire [16-1:0] node11421;
	wire [16-1:0] node11424;
	wire [16-1:0] node11425;
	wire [16-1:0] node11426;
	wire [16-1:0] node11427;
	wire [16-1:0] node11428;
	wire [16-1:0] node11429;
	wire [16-1:0] node11430;
	wire [16-1:0] node11434;
	wire [16-1:0] node11435;
	wire [16-1:0] node11438;
	wire [16-1:0] node11441;
	wire [16-1:0] node11442;
	wire [16-1:0] node11443;
	wire [16-1:0] node11446;
	wire [16-1:0] node11449;
	wire [16-1:0] node11450;
	wire [16-1:0] node11453;
	wire [16-1:0] node11456;
	wire [16-1:0] node11457;
	wire [16-1:0] node11458;
	wire [16-1:0] node11459;
	wire [16-1:0] node11462;
	wire [16-1:0] node11465;
	wire [16-1:0] node11466;
	wire [16-1:0] node11469;
	wire [16-1:0] node11472;
	wire [16-1:0] node11473;
	wire [16-1:0] node11476;
	wire [16-1:0] node11477;
	wire [16-1:0] node11481;
	wire [16-1:0] node11482;
	wire [16-1:0] node11483;
	wire [16-1:0] node11484;
	wire [16-1:0] node11485;
	wire [16-1:0] node11488;
	wire [16-1:0] node11491;
	wire [16-1:0] node11492;
	wire [16-1:0] node11495;
	wire [16-1:0] node11498;
	wire [16-1:0] node11499;
	wire [16-1:0] node11500;
	wire [16-1:0] node11503;
	wire [16-1:0] node11506;
	wire [16-1:0] node11507;
	wire [16-1:0] node11510;
	wire [16-1:0] node11513;
	wire [16-1:0] node11514;
	wire [16-1:0] node11515;
	wire [16-1:0] node11516;
	wire [16-1:0] node11519;
	wire [16-1:0] node11522;
	wire [16-1:0] node11524;
	wire [16-1:0] node11527;
	wire [16-1:0] node11528;
	wire [16-1:0] node11529;
	wire [16-1:0] node11532;
	wire [16-1:0] node11535;
	wire [16-1:0] node11536;
	wire [16-1:0] node11539;
	wire [16-1:0] node11542;
	wire [16-1:0] node11543;
	wire [16-1:0] node11544;
	wire [16-1:0] node11545;
	wire [16-1:0] node11546;
	wire [16-1:0] node11547;
	wire [16-1:0] node11550;
	wire [16-1:0] node11553;
	wire [16-1:0] node11554;
	wire [16-1:0] node11557;
	wire [16-1:0] node11560;
	wire [16-1:0] node11561;
	wire [16-1:0] node11562;
	wire [16-1:0] node11565;
	wire [16-1:0] node11568;
	wire [16-1:0] node11569;
	wire [16-1:0] node11572;
	wire [16-1:0] node11575;
	wire [16-1:0] node11576;
	wire [16-1:0] node11577;
	wire [16-1:0] node11578;
	wire [16-1:0] node11582;
	wire [16-1:0] node11583;
	wire [16-1:0] node11587;
	wire [16-1:0] node11588;
	wire [16-1:0] node11589;
	wire [16-1:0] node11592;
	wire [16-1:0] node11595;
	wire [16-1:0] node11596;
	wire [16-1:0] node11599;
	wire [16-1:0] node11602;
	wire [16-1:0] node11603;
	wire [16-1:0] node11604;
	wire [16-1:0] node11605;
	wire [16-1:0] node11606;
	wire [16-1:0] node11609;
	wire [16-1:0] node11612;
	wire [16-1:0] node11613;
	wire [16-1:0] node11616;
	wire [16-1:0] node11619;
	wire [16-1:0] node11620;
	wire [16-1:0] node11621;
	wire [16-1:0] node11624;
	wire [16-1:0] node11627;
	wire [16-1:0] node11628;
	wire [16-1:0] node11631;
	wire [16-1:0] node11634;
	wire [16-1:0] node11635;
	wire [16-1:0] node11636;
	wire [16-1:0] node11637;
	wire [16-1:0] node11640;
	wire [16-1:0] node11643;
	wire [16-1:0] node11644;
	wire [16-1:0] node11647;
	wire [16-1:0] node11650;
	wire [16-1:0] node11651;
	wire [16-1:0] node11652;
	wire [16-1:0] node11655;
	wire [16-1:0] node11658;
	wire [16-1:0] node11659;
	wire [16-1:0] node11662;
	wire [16-1:0] node11665;
	wire [16-1:0] node11666;
	wire [16-1:0] node11667;
	wire [16-1:0] node11668;
	wire [16-1:0] node11669;
	wire [16-1:0] node11670;
	wire [16-1:0] node11671;
	wire [16-1:0] node11672;
	wire [16-1:0] node11673;
	wire [16-1:0] node11674;
	wire [16-1:0] node11675;
	wire [16-1:0] node11679;
	wire [16-1:0] node11680;
	wire [16-1:0] node11683;
	wire [16-1:0] node11686;
	wire [16-1:0] node11687;
	wire [16-1:0] node11688;
	wire [16-1:0] node11691;
	wire [16-1:0] node11694;
	wire [16-1:0] node11695;
	wire [16-1:0] node11698;
	wire [16-1:0] node11701;
	wire [16-1:0] node11702;
	wire [16-1:0] node11703;
	wire [16-1:0] node11704;
	wire [16-1:0] node11707;
	wire [16-1:0] node11710;
	wire [16-1:0] node11711;
	wire [16-1:0] node11714;
	wire [16-1:0] node11717;
	wire [16-1:0] node11718;
	wire [16-1:0] node11719;
	wire [16-1:0] node11722;
	wire [16-1:0] node11725;
	wire [16-1:0] node11726;
	wire [16-1:0] node11729;
	wire [16-1:0] node11732;
	wire [16-1:0] node11733;
	wire [16-1:0] node11734;
	wire [16-1:0] node11735;
	wire [16-1:0] node11736;
	wire [16-1:0] node11739;
	wire [16-1:0] node11742;
	wire [16-1:0] node11743;
	wire [16-1:0] node11746;
	wire [16-1:0] node11749;
	wire [16-1:0] node11750;
	wire [16-1:0] node11752;
	wire [16-1:0] node11755;
	wire [16-1:0] node11756;
	wire [16-1:0] node11759;
	wire [16-1:0] node11762;
	wire [16-1:0] node11763;
	wire [16-1:0] node11764;
	wire [16-1:0] node11765;
	wire [16-1:0] node11768;
	wire [16-1:0] node11771;
	wire [16-1:0] node11772;
	wire [16-1:0] node11775;
	wire [16-1:0] node11778;
	wire [16-1:0] node11779;
	wire [16-1:0] node11780;
	wire [16-1:0] node11783;
	wire [16-1:0] node11786;
	wire [16-1:0] node11787;
	wire [16-1:0] node11790;
	wire [16-1:0] node11793;
	wire [16-1:0] node11794;
	wire [16-1:0] node11795;
	wire [16-1:0] node11796;
	wire [16-1:0] node11797;
	wire [16-1:0] node11798;
	wire [16-1:0] node11801;
	wire [16-1:0] node11804;
	wire [16-1:0] node11805;
	wire [16-1:0] node11808;
	wire [16-1:0] node11811;
	wire [16-1:0] node11812;
	wire [16-1:0] node11813;
	wire [16-1:0] node11816;
	wire [16-1:0] node11819;
	wire [16-1:0] node11820;
	wire [16-1:0] node11823;
	wire [16-1:0] node11826;
	wire [16-1:0] node11827;
	wire [16-1:0] node11828;
	wire [16-1:0] node11829;
	wire [16-1:0] node11832;
	wire [16-1:0] node11835;
	wire [16-1:0] node11836;
	wire [16-1:0] node11839;
	wire [16-1:0] node11842;
	wire [16-1:0] node11843;
	wire [16-1:0] node11844;
	wire [16-1:0] node11847;
	wire [16-1:0] node11850;
	wire [16-1:0] node11851;
	wire [16-1:0] node11854;
	wire [16-1:0] node11857;
	wire [16-1:0] node11858;
	wire [16-1:0] node11859;
	wire [16-1:0] node11860;
	wire [16-1:0] node11861;
	wire [16-1:0] node11864;
	wire [16-1:0] node11867;
	wire [16-1:0] node11868;
	wire [16-1:0] node11871;
	wire [16-1:0] node11874;
	wire [16-1:0] node11875;
	wire [16-1:0] node11876;
	wire [16-1:0] node11880;
	wire [16-1:0] node11881;
	wire [16-1:0] node11884;
	wire [16-1:0] node11887;
	wire [16-1:0] node11888;
	wire [16-1:0] node11889;
	wire [16-1:0] node11890;
	wire [16-1:0] node11893;
	wire [16-1:0] node11896;
	wire [16-1:0] node11897;
	wire [16-1:0] node11900;
	wire [16-1:0] node11903;
	wire [16-1:0] node11904;
	wire [16-1:0] node11905;
	wire [16-1:0] node11908;
	wire [16-1:0] node11911;
	wire [16-1:0] node11912;
	wire [16-1:0] node11915;
	wire [16-1:0] node11918;
	wire [16-1:0] node11919;
	wire [16-1:0] node11920;
	wire [16-1:0] node11921;
	wire [16-1:0] node11922;
	wire [16-1:0] node11923;
	wire [16-1:0] node11924;
	wire [16-1:0] node11927;
	wire [16-1:0] node11930;
	wire [16-1:0] node11931;
	wire [16-1:0] node11935;
	wire [16-1:0] node11936;
	wire [16-1:0] node11938;
	wire [16-1:0] node11941;
	wire [16-1:0] node11942;
	wire [16-1:0] node11945;
	wire [16-1:0] node11948;
	wire [16-1:0] node11949;
	wire [16-1:0] node11950;
	wire [16-1:0] node11951;
	wire [16-1:0] node11954;
	wire [16-1:0] node11957;
	wire [16-1:0] node11958;
	wire [16-1:0] node11961;
	wire [16-1:0] node11964;
	wire [16-1:0] node11965;
	wire [16-1:0] node11966;
	wire [16-1:0] node11969;
	wire [16-1:0] node11972;
	wire [16-1:0] node11973;
	wire [16-1:0] node11976;
	wire [16-1:0] node11979;
	wire [16-1:0] node11980;
	wire [16-1:0] node11981;
	wire [16-1:0] node11982;
	wire [16-1:0] node11983;
	wire [16-1:0] node11986;
	wire [16-1:0] node11989;
	wire [16-1:0] node11990;
	wire [16-1:0] node11993;
	wire [16-1:0] node11996;
	wire [16-1:0] node11997;
	wire [16-1:0] node11998;
	wire [16-1:0] node12001;
	wire [16-1:0] node12004;
	wire [16-1:0] node12005;
	wire [16-1:0] node12008;
	wire [16-1:0] node12011;
	wire [16-1:0] node12012;
	wire [16-1:0] node12013;
	wire [16-1:0] node12014;
	wire [16-1:0] node12017;
	wire [16-1:0] node12020;
	wire [16-1:0] node12021;
	wire [16-1:0] node12024;
	wire [16-1:0] node12027;
	wire [16-1:0] node12028;
	wire [16-1:0] node12030;
	wire [16-1:0] node12033;
	wire [16-1:0] node12035;
	wire [16-1:0] node12038;
	wire [16-1:0] node12039;
	wire [16-1:0] node12040;
	wire [16-1:0] node12041;
	wire [16-1:0] node12042;
	wire [16-1:0] node12043;
	wire [16-1:0] node12046;
	wire [16-1:0] node12049;
	wire [16-1:0] node12052;
	wire [16-1:0] node12053;
	wire [16-1:0] node12054;
	wire [16-1:0] node12057;
	wire [16-1:0] node12060;
	wire [16-1:0] node12061;
	wire [16-1:0] node12064;
	wire [16-1:0] node12067;
	wire [16-1:0] node12068;
	wire [16-1:0] node12069;
	wire [16-1:0] node12070;
	wire [16-1:0] node12073;
	wire [16-1:0] node12076;
	wire [16-1:0] node12077;
	wire [16-1:0] node12080;
	wire [16-1:0] node12083;
	wire [16-1:0] node12084;
	wire [16-1:0] node12085;
	wire [16-1:0] node12088;
	wire [16-1:0] node12091;
	wire [16-1:0] node12092;
	wire [16-1:0] node12095;
	wire [16-1:0] node12098;
	wire [16-1:0] node12099;
	wire [16-1:0] node12100;
	wire [16-1:0] node12101;
	wire [16-1:0] node12103;
	wire [16-1:0] node12106;
	wire [16-1:0] node12107;
	wire [16-1:0] node12110;
	wire [16-1:0] node12113;
	wire [16-1:0] node12114;
	wire [16-1:0] node12115;
	wire [16-1:0] node12118;
	wire [16-1:0] node12121;
	wire [16-1:0] node12123;
	wire [16-1:0] node12126;
	wire [16-1:0] node12127;
	wire [16-1:0] node12128;
	wire [16-1:0] node12129;
	wire [16-1:0] node12132;
	wire [16-1:0] node12135;
	wire [16-1:0] node12136;
	wire [16-1:0] node12139;
	wire [16-1:0] node12142;
	wire [16-1:0] node12143;
	wire [16-1:0] node12144;
	wire [16-1:0] node12147;
	wire [16-1:0] node12150;
	wire [16-1:0] node12151;
	wire [16-1:0] node12154;
	wire [16-1:0] node12157;
	wire [16-1:0] node12158;
	wire [16-1:0] node12159;
	wire [16-1:0] node12160;
	wire [16-1:0] node12161;
	wire [16-1:0] node12162;
	wire [16-1:0] node12163;
	wire [16-1:0] node12164;
	wire [16-1:0] node12167;
	wire [16-1:0] node12170;
	wire [16-1:0] node12171;
	wire [16-1:0] node12174;
	wire [16-1:0] node12177;
	wire [16-1:0] node12178;
	wire [16-1:0] node12179;
	wire [16-1:0] node12182;
	wire [16-1:0] node12185;
	wire [16-1:0] node12186;
	wire [16-1:0] node12189;
	wire [16-1:0] node12192;
	wire [16-1:0] node12193;
	wire [16-1:0] node12194;
	wire [16-1:0] node12195;
	wire [16-1:0] node12198;
	wire [16-1:0] node12201;
	wire [16-1:0] node12202;
	wire [16-1:0] node12206;
	wire [16-1:0] node12207;
	wire [16-1:0] node12208;
	wire [16-1:0] node12212;
	wire [16-1:0] node12213;
	wire [16-1:0] node12216;
	wire [16-1:0] node12219;
	wire [16-1:0] node12220;
	wire [16-1:0] node12221;
	wire [16-1:0] node12222;
	wire [16-1:0] node12224;
	wire [16-1:0] node12227;
	wire [16-1:0] node12228;
	wire [16-1:0] node12231;
	wire [16-1:0] node12234;
	wire [16-1:0] node12235;
	wire [16-1:0] node12236;
	wire [16-1:0] node12239;
	wire [16-1:0] node12242;
	wire [16-1:0] node12243;
	wire [16-1:0] node12246;
	wire [16-1:0] node12249;
	wire [16-1:0] node12250;
	wire [16-1:0] node12251;
	wire [16-1:0] node12252;
	wire [16-1:0] node12255;
	wire [16-1:0] node12258;
	wire [16-1:0] node12259;
	wire [16-1:0] node12263;
	wire [16-1:0] node12264;
	wire [16-1:0] node12265;
	wire [16-1:0] node12268;
	wire [16-1:0] node12271;
	wire [16-1:0] node12272;
	wire [16-1:0] node12275;
	wire [16-1:0] node12278;
	wire [16-1:0] node12279;
	wire [16-1:0] node12280;
	wire [16-1:0] node12281;
	wire [16-1:0] node12282;
	wire [16-1:0] node12283;
	wire [16-1:0] node12286;
	wire [16-1:0] node12290;
	wire [16-1:0] node12291;
	wire [16-1:0] node12292;
	wire [16-1:0] node12295;
	wire [16-1:0] node12298;
	wire [16-1:0] node12299;
	wire [16-1:0] node12302;
	wire [16-1:0] node12305;
	wire [16-1:0] node12306;
	wire [16-1:0] node12307;
	wire [16-1:0] node12308;
	wire [16-1:0] node12311;
	wire [16-1:0] node12314;
	wire [16-1:0] node12315;
	wire [16-1:0] node12318;
	wire [16-1:0] node12321;
	wire [16-1:0] node12322;
	wire [16-1:0] node12323;
	wire [16-1:0] node12326;
	wire [16-1:0] node12329;
	wire [16-1:0] node12331;
	wire [16-1:0] node12334;
	wire [16-1:0] node12335;
	wire [16-1:0] node12336;
	wire [16-1:0] node12337;
	wire [16-1:0] node12338;
	wire [16-1:0] node12341;
	wire [16-1:0] node12344;
	wire [16-1:0] node12345;
	wire [16-1:0] node12348;
	wire [16-1:0] node12351;
	wire [16-1:0] node12352;
	wire [16-1:0] node12353;
	wire [16-1:0] node12356;
	wire [16-1:0] node12359;
	wire [16-1:0] node12360;
	wire [16-1:0] node12363;
	wire [16-1:0] node12366;
	wire [16-1:0] node12367;
	wire [16-1:0] node12368;
	wire [16-1:0] node12369;
	wire [16-1:0] node12372;
	wire [16-1:0] node12375;
	wire [16-1:0] node12377;
	wire [16-1:0] node12380;
	wire [16-1:0] node12381;
	wire [16-1:0] node12382;
	wire [16-1:0] node12385;
	wire [16-1:0] node12388;
	wire [16-1:0] node12390;
	wire [16-1:0] node12393;
	wire [16-1:0] node12394;
	wire [16-1:0] node12395;
	wire [16-1:0] node12396;
	wire [16-1:0] node12397;
	wire [16-1:0] node12398;
	wire [16-1:0] node12400;
	wire [16-1:0] node12403;
	wire [16-1:0] node12404;
	wire [16-1:0] node12407;
	wire [16-1:0] node12410;
	wire [16-1:0] node12411;
	wire [16-1:0] node12412;
	wire [16-1:0] node12415;
	wire [16-1:0] node12418;
	wire [16-1:0] node12419;
	wire [16-1:0] node12422;
	wire [16-1:0] node12425;
	wire [16-1:0] node12426;
	wire [16-1:0] node12427;
	wire [16-1:0] node12428;
	wire [16-1:0] node12431;
	wire [16-1:0] node12434;
	wire [16-1:0] node12435;
	wire [16-1:0] node12439;
	wire [16-1:0] node12440;
	wire [16-1:0] node12442;
	wire [16-1:0] node12445;
	wire [16-1:0] node12446;
	wire [16-1:0] node12450;
	wire [16-1:0] node12451;
	wire [16-1:0] node12452;
	wire [16-1:0] node12453;
	wire [16-1:0] node12454;
	wire [16-1:0] node12458;
	wire [16-1:0] node12459;
	wire [16-1:0] node12462;
	wire [16-1:0] node12465;
	wire [16-1:0] node12466;
	wire [16-1:0] node12467;
	wire [16-1:0] node12470;
	wire [16-1:0] node12473;
	wire [16-1:0] node12474;
	wire [16-1:0] node12477;
	wire [16-1:0] node12480;
	wire [16-1:0] node12481;
	wire [16-1:0] node12482;
	wire [16-1:0] node12483;
	wire [16-1:0] node12486;
	wire [16-1:0] node12489;
	wire [16-1:0] node12490;
	wire [16-1:0] node12493;
	wire [16-1:0] node12496;
	wire [16-1:0] node12497;
	wire [16-1:0] node12499;
	wire [16-1:0] node12502;
	wire [16-1:0] node12503;
	wire [16-1:0] node12506;
	wire [16-1:0] node12509;
	wire [16-1:0] node12510;
	wire [16-1:0] node12511;
	wire [16-1:0] node12512;
	wire [16-1:0] node12513;
	wire [16-1:0] node12514;
	wire [16-1:0] node12517;
	wire [16-1:0] node12520;
	wire [16-1:0] node12521;
	wire [16-1:0] node12524;
	wire [16-1:0] node12527;
	wire [16-1:0] node12528;
	wire [16-1:0] node12529;
	wire [16-1:0] node12532;
	wire [16-1:0] node12535;
	wire [16-1:0] node12536;
	wire [16-1:0] node12539;
	wire [16-1:0] node12542;
	wire [16-1:0] node12543;
	wire [16-1:0] node12544;
	wire [16-1:0] node12546;
	wire [16-1:0] node12549;
	wire [16-1:0] node12550;
	wire [16-1:0] node12553;
	wire [16-1:0] node12556;
	wire [16-1:0] node12557;
	wire [16-1:0] node12558;
	wire [16-1:0] node12561;
	wire [16-1:0] node12564;
	wire [16-1:0] node12565;
	wire [16-1:0] node12568;
	wire [16-1:0] node12571;
	wire [16-1:0] node12572;
	wire [16-1:0] node12573;
	wire [16-1:0] node12574;
	wire [16-1:0] node12575;
	wire [16-1:0] node12578;
	wire [16-1:0] node12581;
	wire [16-1:0] node12582;
	wire [16-1:0] node12585;
	wire [16-1:0] node12588;
	wire [16-1:0] node12589;
	wire [16-1:0] node12590;
	wire [16-1:0] node12593;
	wire [16-1:0] node12596;
	wire [16-1:0] node12597;
	wire [16-1:0] node12600;
	wire [16-1:0] node12603;
	wire [16-1:0] node12604;
	wire [16-1:0] node12605;
	wire [16-1:0] node12606;
	wire [16-1:0] node12610;
	wire [16-1:0] node12611;
	wire [16-1:0] node12614;
	wire [16-1:0] node12617;
	wire [16-1:0] node12618;
	wire [16-1:0] node12619;
	wire [16-1:0] node12623;
	wire [16-1:0] node12624;
	wire [16-1:0] node12627;
	wire [16-1:0] node12630;
	wire [16-1:0] node12631;
	wire [16-1:0] node12632;
	wire [16-1:0] node12633;
	wire [16-1:0] node12634;
	wire [16-1:0] node12635;
	wire [16-1:0] node12636;
	wire [16-1:0] node12637;
	wire [16-1:0] node12638;
	wire [16-1:0] node12641;
	wire [16-1:0] node12644;
	wire [16-1:0] node12645;
	wire [16-1:0] node12648;
	wire [16-1:0] node12651;
	wire [16-1:0] node12652;
	wire [16-1:0] node12653;
	wire [16-1:0] node12656;
	wire [16-1:0] node12659;
	wire [16-1:0] node12660;
	wire [16-1:0] node12663;
	wire [16-1:0] node12666;
	wire [16-1:0] node12667;
	wire [16-1:0] node12668;
	wire [16-1:0] node12669;
	wire [16-1:0] node12672;
	wire [16-1:0] node12675;
	wire [16-1:0] node12676;
	wire [16-1:0] node12679;
	wire [16-1:0] node12682;
	wire [16-1:0] node12683;
	wire [16-1:0] node12684;
	wire [16-1:0] node12687;
	wire [16-1:0] node12690;
	wire [16-1:0] node12691;
	wire [16-1:0] node12694;
	wire [16-1:0] node12697;
	wire [16-1:0] node12698;
	wire [16-1:0] node12699;
	wire [16-1:0] node12700;
	wire [16-1:0] node12701;
	wire [16-1:0] node12704;
	wire [16-1:0] node12707;
	wire [16-1:0] node12708;
	wire [16-1:0] node12712;
	wire [16-1:0] node12713;
	wire [16-1:0] node12714;
	wire [16-1:0] node12717;
	wire [16-1:0] node12720;
	wire [16-1:0] node12721;
	wire [16-1:0] node12724;
	wire [16-1:0] node12727;
	wire [16-1:0] node12728;
	wire [16-1:0] node12729;
	wire [16-1:0] node12730;
	wire [16-1:0] node12733;
	wire [16-1:0] node12736;
	wire [16-1:0] node12737;
	wire [16-1:0] node12740;
	wire [16-1:0] node12743;
	wire [16-1:0] node12744;
	wire [16-1:0] node12746;
	wire [16-1:0] node12749;
	wire [16-1:0] node12750;
	wire [16-1:0] node12753;
	wire [16-1:0] node12756;
	wire [16-1:0] node12757;
	wire [16-1:0] node12758;
	wire [16-1:0] node12759;
	wire [16-1:0] node12760;
	wire [16-1:0] node12761;
	wire [16-1:0] node12764;
	wire [16-1:0] node12767;
	wire [16-1:0] node12768;
	wire [16-1:0] node12771;
	wire [16-1:0] node12774;
	wire [16-1:0] node12775;
	wire [16-1:0] node12776;
	wire [16-1:0] node12779;
	wire [16-1:0] node12782;
	wire [16-1:0] node12783;
	wire [16-1:0] node12786;
	wire [16-1:0] node12789;
	wire [16-1:0] node12790;
	wire [16-1:0] node12791;
	wire [16-1:0] node12792;
	wire [16-1:0] node12795;
	wire [16-1:0] node12798;
	wire [16-1:0] node12799;
	wire [16-1:0] node12802;
	wire [16-1:0] node12805;
	wire [16-1:0] node12806;
	wire [16-1:0] node12807;
	wire [16-1:0] node12810;
	wire [16-1:0] node12813;
	wire [16-1:0] node12814;
	wire [16-1:0] node12817;
	wire [16-1:0] node12820;
	wire [16-1:0] node12821;
	wire [16-1:0] node12822;
	wire [16-1:0] node12823;
	wire [16-1:0] node12824;
	wire [16-1:0] node12827;
	wire [16-1:0] node12830;
	wire [16-1:0] node12831;
	wire [16-1:0] node12834;
	wire [16-1:0] node12837;
	wire [16-1:0] node12838;
	wire [16-1:0] node12839;
	wire [16-1:0] node12842;
	wire [16-1:0] node12845;
	wire [16-1:0] node12846;
	wire [16-1:0] node12849;
	wire [16-1:0] node12852;
	wire [16-1:0] node12853;
	wire [16-1:0] node12854;
	wire [16-1:0] node12855;
	wire [16-1:0] node12858;
	wire [16-1:0] node12861;
	wire [16-1:0] node12862;
	wire [16-1:0] node12865;
	wire [16-1:0] node12868;
	wire [16-1:0] node12869;
	wire [16-1:0] node12870;
	wire [16-1:0] node12873;
	wire [16-1:0] node12876;
	wire [16-1:0] node12877;
	wire [16-1:0] node12880;
	wire [16-1:0] node12883;
	wire [16-1:0] node12884;
	wire [16-1:0] node12885;
	wire [16-1:0] node12886;
	wire [16-1:0] node12887;
	wire [16-1:0] node12888;
	wire [16-1:0] node12889;
	wire [16-1:0] node12892;
	wire [16-1:0] node12895;
	wire [16-1:0] node12896;
	wire [16-1:0] node12899;
	wire [16-1:0] node12902;
	wire [16-1:0] node12903;
	wire [16-1:0] node12904;
	wire [16-1:0] node12907;
	wire [16-1:0] node12910;
	wire [16-1:0] node12911;
	wire [16-1:0] node12914;
	wire [16-1:0] node12917;
	wire [16-1:0] node12918;
	wire [16-1:0] node12919;
	wire [16-1:0] node12920;
	wire [16-1:0] node12923;
	wire [16-1:0] node12926;
	wire [16-1:0] node12927;
	wire [16-1:0] node12930;
	wire [16-1:0] node12933;
	wire [16-1:0] node12934;
	wire [16-1:0] node12935;
	wire [16-1:0] node12939;
	wire [16-1:0] node12940;
	wire [16-1:0] node12943;
	wire [16-1:0] node12946;
	wire [16-1:0] node12947;
	wire [16-1:0] node12948;
	wire [16-1:0] node12949;
	wire [16-1:0] node12950;
	wire [16-1:0] node12953;
	wire [16-1:0] node12956;
	wire [16-1:0] node12957;
	wire [16-1:0] node12960;
	wire [16-1:0] node12963;
	wire [16-1:0] node12964;
	wire [16-1:0] node12965;
	wire [16-1:0] node12968;
	wire [16-1:0] node12971;
	wire [16-1:0] node12972;
	wire [16-1:0] node12975;
	wire [16-1:0] node12978;
	wire [16-1:0] node12979;
	wire [16-1:0] node12980;
	wire [16-1:0] node12981;
	wire [16-1:0] node12984;
	wire [16-1:0] node12987;
	wire [16-1:0] node12988;
	wire [16-1:0] node12991;
	wire [16-1:0] node12994;
	wire [16-1:0] node12995;
	wire [16-1:0] node12996;
	wire [16-1:0] node12999;
	wire [16-1:0] node13002;
	wire [16-1:0] node13003;
	wire [16-1:0] node13006;
	wire [16-1:0] node13009;
	wire [16-1:0] node13010;
	wire [16-1:0] node13011;
	wire [16-1:0] node13012;
	wire [16-1:0] node13013;
	wire [16-1:0] node13014;
	wire [16-1:0] node13017;
	wire [16-1:0] node13020;
	wire [16-1:0] node13021;
	wire [16-1:0] node13024;
	wire [16-1:0] node13027;
	wire [16-1:0] node13028;
	wire [16-1:0] node13029;
	wire [16-1:0] node13032;
	wire [16-1:0] node13035;
	wire [16-1:0] node13036;
	wire [16-1:0] node13039;
	wire [16-1:0] node13042;
	wire [16-1:0] node13043;
	wire [16-1:0] node13044;
	wire [16-1:0] node13045;
	wire [16-1:0] node13048;
	wire [16-1:0] node13051;
	wire [16-1:0] node13052;
	wire [16-1:0] node13055;
	wire [16-1:0] node13058;
	wire [16-1:0] node13059;
	wire [16-1:0] node13060;
	wire [16-1:0] node13063;
	wire [16-1:0] node13066;
	wire [16-1:0] node13067;
	wire [16-1:0] node13070;
	wire [16-1:0] node13073;
	wire [16-1:0] node13074;
	wire [16-1:0] node13075;
	wire [16-1:0] node13076;
	wire [16-1:0] node13077;
	wire [16-1:0] node13081;
	wire [16-1:0] node13082;
	wire [16-1:0] node13085;
	wire [16-1:0] node13088;
	wire [16-1:0] node13089;
	wire [16-1:0] node13091;
	wire [16-1:0] node13094;
	wire [16-1:0] node13095;
	wire [16-1:0] node13098;
	wire [16-1:0] node13101;
	wire [16-1:0] node13102;
	wire [16-1:0] node13103;
	wire [16-1:0] node13104;
	wire [16-1:0] node13107;
	wire [16-1:0] node13110;
	wire [16-1:0] node13111;
	wire [16-1:0] node13114;
	wire [16-1:0] node13117;
	wire [16-1:0] node13118;
	wire [16-1:0] node13119;
	wire [16-1:0] node13122;
	wire [16-1:0] node13125;
	wire [16-1:0] node13126;
	wire [16-1:0] node13129;
	wire [16-1:0] node13132;
	wire [16-1:0] node13133;
	wire [16-1:0] node13134;
	wire [16-1:0] node13135;
	wire [16-1:0] node13136;
	wire [16-1:0] node13137;
	wire [16-1:0] node13138;
	wire [16-1:0] node13139;
	wire [16-1:0] node13142;
	wire [16-1:0] node13145;
	wire [16-1:0] node13146;
	wire [16-1:0] node13150;
	wire [16-1:0] node13151;
	wire [16-1:0] node13152;
	wire [16-1:0] node13155;
	wire [16-1:0] node13158;
	wire [16-1:0] node13159;
	wire [16-1:0] node13162;
	wire [16-1:0] node13165;
	wire [16-1:0] node13166;
	wire [16-1:0] node13167;
	wire [16-1:0] node13168;
	wire [16-1:0] node13171;
	wire [16-1:0] node13174;
	wire [16-1:0] node13175;
	wire [16-1:0] node13178;
	wire [16-1:0] node13181;
	wire [16-1:0] node13182;
	wire [16-1:0] node13183;
	wire [16-1:0] node13187;
	wire [16-1:0] node13188;
	wire [16-1:0] node13191;
	wire [16-1:0] node13194;
	wire [16-1:0] node13195;
	wire [16-1:0] node13196;
	wire [16-1:0] node13197;
	wire [16-1:0] node13198;
	wire [16-1:0] node13201;
	wire [16-1:0] node13204;
	wire [16-1:0] node13205;
	wire [16-1:0] node13208;
	wire [16-1:0] node13211;
	wire [16-1:0] node13212;
	wire [16-1:0] node13213;
	wire [16-1:0] node13216;
	wire [16-1:0] node13219;
	wire [16-1:0] node13221;
	wire [16-1:0] node13224;
	wire [16-1:0] node13225;
	wire [16-1:0] node13226;
	wire [16-1:0] node13228;
	wire [16-1:0] node13231;
	wire [16-1:0] node13232;
	wire [16-1:0] node13235;
	wire [16-1:0] node13238;
	wire [16-1:0] node13239;
	wire [16-1:0] node13240;
	wire [16-1:0] node13243;
	wire [16-1:0] node13246;
	wire [16-1:0] node13247;
	wire [16-1:0] node13250;
	wire [16-1:0] node13253;
	wire [16-1:0] node13254;
	wire [16-1:0] node13255;
	wire [16-1:0] node13256;
	wire [16-1:0] node13257;
	wire [16-1:0] node13259;
	wire [16-1:0] node13262;
	wire [16-1:0] node13264;
	wire [16-1:0] node13267;
	wire [16-1:0] node13268;
	wire [16-1:0] node13269;
	wire [16-1:0] node13272;
	wire [16-1:0] node13275;
	wire [16-1:0] node13276;
	wire [16-1:0] node13279;
	wire [16-1:0] node13282;
	wire [16-1:0] node13283;
	wire [16-1:0] node13284;
	wire [16-1:0] node13285;
	wire [16-1:0] node13288;
	wire [16-1:0] node13291;
	wire [16-1:0] node13292;
	wire [16-1:0] node13295;
	wire [16-1:0] node13298;
	wire [16-1:0] node13299;
	wire [16-1:0] node13300;
	wire [16-1:0] node13303;
	wire [16-1:0] node13306;
	wire [16-1:0] node13307;
	wire [16-1:0] node13310;
	wire [16-1:0] node13313;
	wire [16-1:0] node13314;
	wire [16-1:0] node13315;
	wire [16-1:0] node13316;
	wire [16-1:0] node13317;
	wire [16-1:0] node13320;
	wire [16-1:0] node13323;
	wire [16-1:0] node13324;
	wire [16-1:0] node13328;
	wire [16-1:0] node13329;
	wire [16-1:0] node13330;
	wire [16-1:0] node13333;
	wire [16-1:0] node13336;
	wire [16-1:0] node13337;
	wire [16-1:0] node13340;
	wire [16-1:0] node13343;
	wire [16-1:0] node13344;
	wire [16-1:0] node13345;
	wire [16-1:0] node13346;
	wire [16-1:0] node13349;
	wire [16-1:0] node13352;
	wire [16-1:0] node13353;
	wire [16-1:0] node13356;
	wire [16-1:0] node13359;
	wire [16-1:0] node13360;
	wire [16-1:0] node13361;
	wire [16-1:0] node13364;
	wire [16-1:0] node13367;
	wire [16-1:0] node13368;
	wire [16-1:0] node13371;
	wire [16-1:0] node13374;
	wire [16-1:0] node13375;
	wire [16-1:0] node13376;
	wire [16-1:0] node13377;
	wire [16-1:0] node13378;
	wire [16-1:0] node13379;
	wire [16-1:0] node13381;
	wire [16-1:0] node13384;
	wire [16-1:0] node13385;
	wire [16-1:0] node13388;
	wire [16-1:0] node13391;
	wire [16-1:0] node13393;
	wire [16-1:0] node13394;
	wire [16-1:0] node13397;
	wire [16-1:0] node13400;
	wire [16-1:0] node13401;
	wire [16-1:0] node13402;
	wire [16-1:0] node13403;
	wire [16-1:0] node13406;
	wire [16-1:0] node13409;
	wire [16-1:0] node13410;
	wire [16-1:0] node13413;
	wire [16-1:0] node13416;
	wire [16-1:0] node13417;
	wire [16-1:0] node13418;
	wire [16-1:0] node13421;
	wire [16-1:0] node13424;
	wire [16-1:0] node13425;
	wire [16-1:0] node13428;
	wire [16-1:0] node13431;
	wire [16-1:0] node13432;
	wire [16-1:0] node13433;
	wire [16-1:0] node13434;
	wire [16-1:0] node13436;
	wire [16-1:0] node13439;
	wire [16-1:0] node13440;
	wire [16-1:0] node13444;
	wire [16-1:0] node13445;
	wire [16-1:0] node13446;
	wire [16-1:0] node13450;
	wire [16-1:0] node13451;
	wire [16-1:0] node13454;
	wire [16-1:0] node13457;
	wire [16-1:0] node13458;
	wire [16-1:0] node13459;
	wire [16-1:0] node13461;
	wire [16-1:0] node13465;
	wire [16-1:0] node13466;
	wire [16-1:0] node13467;
	wire [16-1:0] node13470;
	wire [16-1:0] node13473;
	wire [16-1:0] node13474;
	wire [16-1:0] node13478;
	wire [16-1:0] node13479;
	wire [16-1:0] node13480;
	wire [16-1:0] node13481;
	wire [16-1:0] node13482;
	wire [16-1:0] node13483;
	wire [16-1:0] node13486;
	wire [16-1:0] node13489;
	wire [16-1:0] node13490;
	wire [16-1:0] node13494;
	wire [16-1:0] node13495;
	wire [16-1:0] node13496;
	wire [16-1:0] node13499;
	wire [16-1:0] node13502;
	wire [16-1:0] node13503;
	wire [16-1:0] node13506;
	wire [16-1:0] node13509;
	wire [16-1:0] node13510;
	wire [16-1:0] node13511;
	wire [16-1:0] node13512;
	wire [16-1:0] node13515;
	wire [16-1:0] node13518;
	wire [16-1:0] node13520;
	wire [16-1:0] node13523;
	wire [16-1:0] node13524;
	wire [16-1:0] node13527;
	wire [16-1:0] node13529;
	wire [16-1:0] node13532;
	wire [16-1:0] node13533;
	wire [16-1:0] node13534;
	wire [16-1:0] node13535;
	wire [16-1:0] node13536;
	wire [16-1:0] node13539;
	wire [16-1:0] node13542;
	wire [16-1:0] node13543;
	wire [16-1:0] node13546;
	wire [16-1:0] node13549;
	wire [16-1:0] node13550;
	wire [16-1:0] node13551;
	wire [16-1:0] node13554;
	wire [16-1:0] node13557;
	wire [16-1:0] node13558;
	wire [16-1:0] node13561;
	wire [16-1:0] node13564;
	wire [16-1:0] node13565;
	wire [16-1:0] node13566;
	wire [16-1:0] node13567;
	wire [16-1:0] node13570;
	wire [16-1:0] node13573;
	wire [16-1:0] node13574;
	wire [16-1:0] node13577;
	wire [16-1:0] node13580;
	wire [16-1:0] node13581;
	wire [16-1:0] node13582;
	wire [16-1:0] node13585;
	wire [16-1:0] node13588;
	wire [16-1:0] node13589;
	wire [16-1:0] node13592;
	wire [16-1:0] node13595;
	wire [16-1:0] node13596;
	wire [16-1:0] node13597;
	wire [16-1:0] node13598;
	wire [16-1:0] node13599;
	wire [16-1:0] node13600;
	wire [16-1:0] node13601;
	wire [16-1:0] node13602;
	wire [16-1:0] node13603;
	wire [16-1:0] node13604;
	wire [16-1:0] node13607;
	wire [16-1:0] node13610;
	wire [16-1:0] node13611;
	wire [16-1:0] node13615;
	wire [16-1:0] node13616;
	wire [16-1:0] node13617;
	wire [16-1:0] node13620;
	wire [16-1:0] node13623;
	wire [16-1:0] node13624;
	wire [16-1:0] node13627;
	wire [16-1:0] node13630;
	wire [16-1:0] node13631;
	wire [16-1:0] node13632;
	wire [16-1:0] node13633;
	wire [16-1:0] node13636;
	wire [16-1:0] node13639;
	wire [16-1:0] node13640;
	wire [16-1:0] node13643;
	wire [16-1:0] node13646;
	wire [16-1:0] node13647;
	wire [16-1:0] node13648;
	wire [16-1:0] node13652;
	wire [16-1:0] node13653;
	wire [16-1:0] node13656;
	wire [16-1:0] node13659;
	wire [16-1:0] node13660;
	wire [16-1:0] node13661;
	wire [16-1:0] node13662;
	wire [16-1:0] node13663;
	wire [16-1:0] node13666;
	wire [16-1:0] node13669;
	wire [16-1:0] node13670;
	wire [16-1:0] node13673;
	wire [16-1:0] node13676;
	wire [16-1:0] node13677;
	wire [16-1:0] node13678;
	wire [16-1:0] node13681;
	wire [16-1:0] node13684;
	wire [16-1:0] node13685;
	wire [16-1:0] node13688;
	wire [16-1:0] node13691;
	wire [16-1:0] node13692;
	wire [16-1:0] node13693;
	wire [16-1:0] node13694;
	wire [16-1:0] node13697;
	wire [16-1:0] node13700;
	wire [16-1:0] node13702;
	wire [16-1:0] node13705;
	wire [16-1:0] node13706;
	wire [16-1:0] node13707;
	wire [16-1:0] node13710;
	wire [16-1:0] node13713;
	wire [16-1:0] node13714;
	wire [16-1:0] node13717;
	wire [16-1:0] node13720;
	wire [16-1:0] node13721;
	wire [16-1:0] node13722;
	wire [16-1:0] node13723;
	wire [16-1:0] node13724;
	wire [16-1:0] node13725;
	wire [16-1:0] node13728;
	wire [16-1:0] node13731;
	wire [16-1:0] node13732;
	wire [16-1:0] node13735;
	wire [16-1:0] node13738;
	wire [16-1:0] node13739;
	wire [16-1:0] node13740;
	wire [16-1:0] node13743;
	wire [16-1:0] node13746;
	wire [16-1:0] node13747;
	wire [16-1:0] node13750;
	wire [16-1:0] node13753;
	wire [16-1:0] node13754;
	wire [16-1:0] node13755;
	wire [16-1:0] node13756;
	wire [16-1:0] node13759;
	wire [16-1:0] node13762;
	wire [16-1:0] node13763;
	wire [16-1:0] node13766;
	wire [16-1:0] node13769;
	wire [16-1:0] node13770;
	wire [16-1:0] node13771;
	wire [16-1:0] node13774;
	wire [16-1:0] node13777;
	wire [16-1:0] node13778;
	wire [16-1:0] node13781;
	wire [16-1:0] node13784;
	wire [16-1:0] node13785;
	wire [16-1:0] node13786;
	wire [16-1:0] node13787;
	wire [16-1:0] node13788;
	wire [16-1:0] node13791;
	wire [16-1:0] node13794;
	wire [16-1:0] node13795;
	wire [16-1:0] node13798;
	wire [16-1:0] node13801;
	wire [16-1:0] node13802;
	wire [16-1:0] node13803;
	wire [16-1:0] node13806;
	wire [16-1:0] node13809;
	wire [16-1:0] node13810;
	wire [16-1:0] node13813;
	wire [16-1:0] node13816;
	wire [16-1:0] node13817;
	wire [16-1:0] node13818;
	wire [16-1:0] node13820;
	wire [16-1:0] node13823;
	wire [16-1:0] node13824;
	wire [16-1:0] node13827;
	wire [16-1:0] node13830;
	wire [16-1:0] node13831;
	wire [16-1:0] node13832;
	wire [16-1:0] node13835;
	wire [16-1:0] node13838;
	wire [16-1:0] node13839;
	wire [16-1:0] node13842;
	wire [16-1:0] node13845;
	wire [16-1:0] node13846;
	wire [16-1:0] node13847;
	wire [16-1:0] node13848;
	wire [16-1:0] node13849;
	wire [16-1:0] node13850;
	wire [16-1:0] node13851;
	wire [16-1:0] node13855;
	wire [16-1:0] node13856;
	wire [16-1:0] node13859;
	wire [16-1:0] node13862;
	wire [16-1:0] node13863;
	wire [16-1:0] node13864;
	wire [16-1:0] node13867;
	wire [16-1:0] node13870;
	wire [16-1:0] node13871;
	wire [16-1:0] node13875;
	wire [16-1:0] node13876;
	wire [16-1:0] node13877;
	wire [16-1:0] node13878;
	wire [16-1:0] node13881;
	wire [16-1:0] node13884;
	wire [16-1:0] node13885;
	wire [16-1:0] node13889;
	wire [16-1:0] node13890;
	wire [16-1:0] node13891;
	wire [16-1:0] node13894;
	wire [16-1:0] node13897;
	wire [16-1:0] node13899;
	wire [16-1:0] node13902;
	wire [16-1:0] node13903;
	wire [16-1:0] node13904;
	wire [16-1:0] node13905;
	wire [16-1:0] node13906;
	wire [16-1:0] node13909;
	wire [16-1:0] node13912;
	wire [16-1:0] node13913;
	wire [16-1:0] node13916;
	wire [16-1:0] node13919;
	wire [16-1:0] node13920;
	wire [16-1:0] node13921;
	wire [16-1:0] node13924;
	wire [16-1:0] node13927;
	wire [16-1:0] node13928;
	wire [16-1:0] node13931;
	wire [16-1:0] node13934;
	wire [16-1:0] node13935;
	wire [16-1:0] node13936;
	wire [16-1:0] node13937;
	wire [16-1:0] node13940;
	wire [16-1:0] node13943;
	wire [16-1:0] node13944;
	wire [16-1:0] node13947;
	wire [16-1:0] node13950;
	wire [16-1:0] node13951;
	wire [16-1:0] node13952;
	wire [16-1:0] node13955;
	wire [16-1:0] node13958;
	wire [16-1:0] node13959;
	wire [16-1:0] node13962;
	wire [16-1:0] node13965;
	wire [16-1:0] node13966;
	wire [16-1:0] node13967;
	wire [16-1:0] node13968;
	wire [16-1:0] node13969;
	wire [16-1:0] node13970;
	wire [16-1:0] node13973;
	wire [16-1:0] node13976;
	wire [16-1:0] node13977;
	wire [16-1:0] node13980;
	wire [16-1:0] node13983;
	wire [16-1:0] node13984;
	wire [16-1:0] node13985;
	wire [16-1:0] node13988;
	wire [16-1:0] node13991;
	wire [16-1:0] node13992;
	wire [16-1:0] node13996;
	wire [16-1:0] node13997;
	wire [16-1:0] node13998;
	wire [16-1:0] node13999;
	wire [16-1:0] node14002;
	wire [16-1:0] node14005;
	wire [16-1:0] node14006;
	wire [16-1:0] node14009;
	wire [16-1:0] node14012;
	wire [16-1:0] node14013;
	wire [16-1:0] node14016;
	wire [16-1:0] node14017;
	wire [16-1:0] node14020;
	wire [16-1:0] node14023;
	wire [16-1:0] node14024;
	wire [16-1:0] node14025;
	wire [16-1:0] node14026;
	wire [16-1:0] node14027;
	wire [16-1:0] node14030;
	wire [16-1:0] node14033;
	wire [16-1:0] node14034;
	wire [16-1:0] node14037;
	wire [16-1:0] node14040;
	wire [16-1:0] node14041;
	wire [16-1:0] node14042;
	wire [16-1:0] node14045;
	wire [16-1:0] node14048;
	wire [16-1:0] node14049;
	wire [16-1:0] node14052;
	wire [16-1:0] node14055;
	wire [16-1:0] node14056;
	wire [16-1:0] node14057;
	wire [16-1:0] node14058;
	wire [16-1:0] node14061;
	wire [16-1:0] node14064;
	wire [16-1:0] node14066;
	wire [16-1:0] node14069;
	wire [16-1:0] node14070;
	wire [16-1:0] node14071;
	wire [16-1:0] node14074;
	wire [16-1:0] node14077;
	wire [16-1:0] node14078;
	wire [16-1:0] node14081;
	wire [16-1:0] node14084;
	wire [16-1:0] node14085;
	wire [16-1:0] node14086;
	wire [16-1:0] node14087;
	wire [16-1:0] node14088;
	wire [16-1:0] node14089;
	wire [16-1:0] node14090;
	wire [16-1:0] node14091;
	wire [16-1:0] node14094;
	wire [16-1:0] node14097;
	wire [16-1:0] node14098;
	wire [16-1:0] node14102;
	wire [16-1:0] node14103;
	wire [16-1:0] node14104;
	wire [16-1:0] node14107;
	wire [16-1:0] node14110;
	wire [16-1:0] node14111;
	wire [16-1:0] node14115;
	wire [16-1:0] node14116;
	wire [16-1:0] node14117;
	wire [16-1:0] node14118;
	wire [16-1:0] node14121;
	wire [16-1:0] node14124;
	wire [16-1:0] node14125;
	wire [16-1:0] node14128;
	wire [16-1:0] node14131;
	wire [16-1:0] node14132;
	wire [16-1:0] node14133;
	wire [16-1:0] node14136;
	wire [16-1:0] node14139;
	wire [16-1:0] node14140;
	wire [16-1:0] node14143;
	wire [16-1:0] node14146;
	wire [16-1:0] node14147;
	wire [16-1:0] node14148;
	wire [16-1:0] node14149;
	wire [16-1:0] node14150;
	wire [16-1:0] node14153;
	wire [16-1:0] node14156;
	wire [16-1:0] node14157;
	wire [16-1:0] node14160;
	wire [16-1:0] node14163;
	wire [16-1:0] node14164;
	wire [16-1:0] node14165;
	wire [16-1:0] node14168;
	wire [16-1:0] node14171;
	wire [16-1:0] node14172;
	wire [16-1:0] node14176;
	wire [16-1:0] node14177;
	wire [16-1:0] node14178;
	wire [16-1:0] node14179;
	wire [16-1:0] node14182;
	wire [16-1:0] node14185;
	wire [16-1:0] node14186;
	wire [16-1:0] node14189;
	wire [16-1:0] node14192;
	wire [16-1:0] node14193;
	wire [16-1:0] node14194;
	wire [16-1:0] node14197;
	wire [16-1:0] node14200;
	wire [16-1:0] node14201;
	wire [16-1:0] node14204;
	wire [16-1:0] node14207;
	wire [16-1:0] node14208;
	wire [16-1:0] node14209;
	wire [16-1:0] node14210;
	wire [16-1:0] node14211;
	wire [16-1:0] node14212;
	wire [16-1:0] node14215;
	wire [16-1:0] node14218;
	wire [16-1:0] node14219;
	wire [16-1:0] node14222;
	wire [16-1:0] node14225;
	wire [16-1:0] node14226;
	wire [16-1:0] node14227;
	wire [16-1:0] node14230;
	wire [16-1:0] node14233;
	wire [16-1:0] node14234;
	wire [16-1:0] node14237;
	wire [16-1:0] node14240;
	wire [16-1:0] node14241;
	wire [16-1:0] node14242;
	wire [16-1:0] node14243;
	wire [16-1:0] node14246;
	wire [16-1:0] node14249;
	wire [16-1:0] node14250;
	wire [16-1:0] node14253;
	wire [16-1:0] node14256;
	wire [16-1:0] node14257;
	wire [16-1:0] node14258;
	wire [16-1:0] node14261;
	wire [16-1:0] node14264;
	wire [16-1:0] node14265;
	wire [16-1:0] node14268;
	wire [16-1:0] node14271;
	wire [16-1:0] node14272;
	wire [16-1:0] node14273;
	wire [16-1:0] node14274;
	wire [16-1:0] node14275;
	wire [16-1:0] node14278;
	wire [16-1:0] node14281;
	wire [16-1:0] node14282;
	wire [16-1:0] node14285;
	wire [16-1:0] node14288;
	wire [16-1:0] node14289;
	wire [16-1:0] node14290;
	wire [16-1:0] node14293;
	wire [16-1:0] node14296;
	wire [16-1:0] node14298;
	wire [16-1:0] node14301;
	wire [16-1:0] node14302;
	wire [16-1:0] node14303;
	wire [16-1:0] node14305;
	wire [16-1:0] node14308;
	wire [16-1:0] node14309;
	wire [16-1:0] node14312;
	wire [16-1:0] node14315;
	wire [16-1:0] node14316;
	wire [16-1:0] node14317;
	wire [16-1:0] node14320;
	wire [16-1:0] node14323;
	wire [16-1:0] node14324;
	wire [16-1:0] node14327;
	wire [16-1:0] node14330;
	wire [16-1:0] node14331;
	wire [16-1:0] node14332;
	wire [16-1:0] node14333;
	wire [16-1:0] node14334;
	wire [16-1:0] node14335;
	wire [16-1:0] node14336;
	wire [16-1:0] node14339;
	wire [16-1:0] node14342;
	wire [16-1:0] node14343;
	wire [16-1:0] node14346;
	wire [16-1:0] node14349;
	wire [16-1:0] node14350;
	wire [16-1:0] node14351;
	wire [16-1:0] node14354;
	wire [16-1:0] node14357;
	wire [16-1:0] node14358;
	wire [16-1:0] node14361;
	wire [16-1:0] node14364;
	wire [16-1:0] node14365;
	wire [16-1:0] node14366;
	wire [16-1:0] node14367;
	wire [16-1:0] node14370;
	wire [16-1:0] node14373;
	wire [16-1:0] node14374;
	wire [16-1:0] node14377;
	wire [16-1:0] node14380;
	wire [16-1:0] node14381;
	wire [16-1:0] node14383;
	wire [16-1:0] node14386;
	wire [16-1:0] node14387;
	wire [16-1:0] node14390;
	wire [16-1:0] node14393;
	wire [16-1:0] node14394;
	wire [16-1:0] node14395;
	wire [16-1:0] node14396;
	wire [16-1:0] node14397;
	wire [16-1:0] node14400;
	wire [16-1:0] node14403;
	wire [16-1:0] node14404;
	wire [16-1:0] node14407;
	wire [16-1:0] node14410;
	wire [16-1:0] node14411;
	wire [16-1:0] node14412;
	wire [16-1:0] node14415;
	wire [16-1:0] node14418;
	wire [16-1:0] node14419;
	wire [16-1:0] node14422;
	wire [16-1:0] node14425;
	wire [16-1:0] node14426;
	wire [16-1:0] node14427;
	wire [16-1:0] node14428;
	wire [16-1:0] node14431;
	wire [16-1:0] node14434;
	wire [16-1:0] node14435;
	wire [16-1:0] node14438;
	wire [16-1:0] node14441;
	wire [16-1:0] node14442;
	wire [16-1:0] node14444;
	wire [16-1:0] node14447;
	wire [16-1:0] node14448;
	wire [16-1:0] node14451;
	wire [16-1:0] node14454;
	wire [16-1:0] node14455;
	wire [16-1:0] node14456;
	wire [16-1:0] node14457;
	wire [16-1:0] node14458;
	wire [16-1:0] node14459;
	wire [16-1:0] node14462;
	wire [16-1:0] node14465;
	wire [16-1:0] node14466;
	wire [16-1:0] node14470;
	wire [16-1:0] node14471;
	wire [16-1:0] node14473;
	wire [16-1:0] node14476;
	wire [16-1:0] node14477;
	wire [16-1:0] node14480;
	wire [16-1:0] node14483;
	wire [16-1:0] node14484;
	wire [16-1:0] node14485;
	wire [16-1:0] node14486;
	wire [16-1:0] node14489;
	wire [16-1:0] node14492;
	wire [16-1:0] node14493;
	wire [16-1:0] node14496;
	wire [16-1:0] node14499;
	wire [16-1:0] node14500;
	wire [16-1:0] node14501;
	wire [16-1:0] node14504;
	wire [16-1:0] node14507;
	wire [16-1:0] node14508;
	wire [16-1:0] node14511;
	wire [16-1:0] node14514;
	wire [16-1:0] node14515;
	wire [16-1:0] node14516;
	wire [16-1:0] node14517;
	wire [16-1:0] node14518;
	wire [16-1:0] node14521;
	wire [16-1:0] node14524;
	wire [16-1:0] node14525;
	wire [16-1:0] node14528;
	wire [16-1:0] node14531;
	wire [16-1:0] node14532;
	wire [16-1:0] node14533;
	wire [16-1:0] node14536;
	wire [16-1:0] node14539;
	wire [16-1:0] node14540;
	wire [16-1:0] node14543;
	wire [16-1:0] node14546;
	wire [16-1:0] node14547;
	wire [16-1:0] node14548;
	wire [16-1:0] node14549;
	wire [16-1:0] node14553;
	wire [16-1:0] node14554;
	wire [16-1:0] node14557;
	wire [16-1:0] node14560;
	wire [16-1:0] node14561;
	wire [16-1:0] node14562;
	wire [16-1:0] node14565;
	wire [16-1:0] node14568;
	wire [16-1:0] node14569;
	wire [16-1:0] node14572;
	wire [16-1:0] node14575;
	wire [16-1:0] node14576;
	wire [16-1:0] node14577;
	wire [16-1:0] node14578;
	wire [16-1:0] node14579;
	wire [16-1:0] node14580;
	wire [16-1:0] node14581;
	wire [16-1:0] node14582;
	wire [16-1:0] node14583;
	wire [16-1:0] node14587;
	wire [16-1:0] node14588;
	wire [16-1:0] node14591;
	wire [16-1:0] node14594;
	wire [16-1:0] node14595;
	wire [16-1:0] node14596;
	wire [16-1:0] node14599;
	wire [16-1:0] node14602;
	wire [16-1:0] node14603;
	wire [16-1:0] node14606;
	wire [16-1:0] node14609;
	wire [16-1:0] node14610;
	wire [16-1:0] node14611;
	wire [16-1:0] node14612;
	wire [16-1:0] node14615;
	wire [16-1:0] node14618;
	wire [16-1:0] node14619;
	wire [16-1:0] node14622;
	wire [16-1:0] node14625;
	wire [16-1:0] node14626;
	wire [16-1:0] node14627;
	wire [16-1:0] node14630;
	wire [16-1:0] node14633;
	wire [16-1:0] node14635;
	wire [16-1:0] node14638;
	wire [16-1:0] node14639;
	wire [16-1:0] node14640;
	wire [16-1:0] node14641;
	wire [16-1:0] node14642;
	wire [16-1:0] node14645;
	wire [16-1:0] node14648;
	wire [16-1:0] node14649;
	wire [16-1:0] node14652;
	wire [16-1:0] node14655;
	wire [16-1:0] node14656;
	wire [16-1:0] node14657;
	wire [16-1:0] node14661;
	wire [16-1:0] node14662;
	wire [16-1:0] node14665;
	wire [16-1:0] node14668;
	wire [16-1:0] node14669;
	wire [16-1:0] node14670;
	wire [16-1:0] node14671;
	wire [16-1:0] node14674;
	wire [16-1:0] node14677;
	wire [16-1:0] node14678;
	wire [16-1:0] node14681;
	wire [16-1:0] node14684;
	wire [16-1:0] node14685;
	wire [16-1:0] node14686;
	wire [16-1:0] node14689;
	wire [16-1:0] node14692;
	wire [16-1:0] node14693;
	wire [16-1:0] node14696;
	wire [16-1:0] node14699;
	wire [16-1:0] node14700;
	wire [16-1:0] node14701;
	wire [16-1:0] node14702;
	wire [16-1:0] node14703;
	wire [16-1:0] node14704;
	wire [16-1:0] node14707;
	wire [16-1:0] node14710;
	wire [16-1:0] node14711;
	wire [16-1:0] node14714;
	wire [16-1:0] node14717;
	wire [16-1:0] node14718;
	wire [16-1:0] node14719;
	wire [16-1:0] node14722;
	wire [16-1:0] node14725;
	wire [16-1:0] node14726;
	wire [16-1:0] node14729;
	wire [16-1:0] node14732;
	wire [16-1:0] node14733;
	wire [16-1:0] node14734;
	wire [16-1:0] node14735;
	wire [16-1:0] node14738;
	wire [16-1:0] node14741;
	wire [16-1:0] node14742;
	wire [16-1:0] node14745;
	wire [16-1:0] node14748;
	wire [16-1:0] node14749;
	wire [16-1:0] node14751;
	wire [16-1:0] node14754;
	wire [16-1:0] node14755;
	wire [16-1:0] node14758;
	wire [16-1:0] node14761;
	wire [16-1:0] node14762;
	wire [16-1:0] node14763;
	wire [16-1:0] node14764;
	wire [16-1:0] node14765;
	wire [16-1:0] node14768;
	wire [16-1:0] node14771;
	wire [16-1:0] node14772;
	wire [16-1:0] node14775;
	wire [16-1:0] node14778;
	wire [16-1:0] node14779;
	wire [16-1:0] node14780;
	wire [16-1:0] node14783;
	wire [16-1:0] node14786;
	wire [16-1:0] node14787;
	wire [16-1:0] node14790;
	wire [16-1:0] node14793;
	wire [16-1:0] node14794;
	wire [16-1:0] node14795;
	wire [16-1:0] node14796;
	wire [16-1:0] node14799;
	wire [16-1:0] node14802;
	wire [16-1:0] node14803;
	wire [16-1:0] node14806;
	wire [16-1:0] node14809;
	wire [16-1:0] node14810;
	wire [16-1:0] node14811;
	wire [16-1:0] node14814;
	wire [16-1:0] node14817;
	wire [16-1:0] node14818;
	wire [16-1:0] node14821;
	wire [16-1:0] node14824;
	wire [16-1:0] node14825;
	wire [16-1:0] node14826;
	wire [16-1:0] node14827;
	wire [16-1:0] node14828;
	wire [16-1:0] node14829;
	wire [16-1:0] node14830;
	wire [16-1:0] node14833;
	wire [16-1:0] node14836;
	wire [16-1:0] node14837;
	wire [16-1:0] node14841;
	wire [16-1:0] node14842;
	wire [16-1:0] node14843;
	wire [16-1:0] node14846;
	wire [16-1:0] node14849;
	wire [16-1:0] node14850;
	wire [16-1:0] node14853;
	wire [16-1:0] node14856;
	wire [16-1:0] node14857;
	wire [16-1:0] node14858;
	wire [16-1:0] node14859;
	wire [16-1:0] node14862;
	wire [16-1:0] node14865;
	wire [16-1:0] node14866;
	wire [16-1:0] node14869;
	wire [16-1:0] node14872;
	wire [16-1:0] node14873;
	wire [16-1:0] node14874;
	wire [16-1:0] node14877;
	wire [16-1:0] node14880;
	wire [16-1:0] node14882;
	wire [16-1:0] node14885;
	wire [16-1:0] node14886;
	wire [16-1:0] node14887;
	wire [16-1:0] node14888;
	wire [16-1:0] node14889;
	wire [16-1:0] node14892;
	wire [16-1:0] node14895;
	wire [16-1:0] node14896;
	wire [16-1:0] node14899;
	wire [16-1:0] node14902;
	wire [16-1:0] node14903;
	wire [16-1:0] node14904;
	wire [16-1:0] node14907;
	wire [16-1:0] node14910;
	wire [16-1:0] node14911;
	wire [16-1:0] node14914;
	wire [16-1:0] node14917;
	wire [16-1:0] node14918;
	wire [16-1:0] node14919;
	wire [16-1:0] node14921;
	wire [16-1:0] node14924;
	wire [16-1:0] node14925;
	wire [16-1:0] node14928;
	wire [16-1:0] node14931;
	wire [16-1:0] node14932;
	wire [16-1:0] node14933;
	wire [16-1:0] node14936;
	wire [16-1:0] node14939;
	wire [16-1:0] node14940;
	wire [16-1:0] node14943;
	wire [16-1:0] node14946;
	wire [16-1:0] node14947;
	wire [16-1:0] node14948;
	wire [16-1:0] node14949;
	wire [16-1:0] node14950;
	wire [16-1:0] node14951;
	wire [16-1:0] node14954;
	wire [16-1:0] node14957;
	wire [16-1:0] node14958;
	wire [16-1:0] node14961;
	wire [16-1:0] node14964;
	wire [16-1:0] node14965;
	wire [16-1:0] node14966;
	wire [16-1:0] node14969;
	wire [16-1:0] node14972;
	wire [16-1:0] node14973;
	wire [16-1:0] node14977;
	wire [16-1:0] node14978;
	wire [16-1:0] node14979;
	wire [16-1:0] node14980;
	wire [16-1:0] node14983;
	wire [16-1:0] node14986;
	wire [16-1:0] node14987;
	wire [16-1:0] node14990;
	wire [16-1:0] node14993;
	wire [16-1:0] node14994;
	wire [16-1:0] node14995;
	wire [16-1:0] node14998;
	wire [16-1:0] node15001;
	wire [16-1:0] node15002;
	wire [16-1:0] node15005;
	wire [16-1:0] node15008;
	wire [16-1:0] node15009;
	wire [16-1:0] node15010;
	wire [16-1:0] node15011;
	wire [16-1:0] node15012;
	wire [16-1:0] node15015;
	wire [16-1:0] node15018;
	wire [16-1:0] node15019;
	wire [16-1:0] node15022;
	wire [16-1:0] node15025;
	wire [16-1:0] node15026;
	wire [16-1:0] node15027;
	wire [16-1:0] node15030;
	wire [16-1:0] node15033;
	wire [16-1:0] node15034;
	wire [16-1:0] node15037;
	wire [16-1:0] node15040;
	wire [16-1:0] node15041;
	wire [16-1:0] node15042;
	wire [16-1:0] node15043;
	wire [16-1:0] node15046;
	wire [16-1:0] node15049;
	wire [16-1:0] node15050;
	wire [16-1:0] node15053;
	wire [16-1:0] node15056;
	wire [16-1:0] node15057;
	wire [16-1:0] node15059;
	wire [16-1:0] node15062;
	wire [16-1:0] node15063;
	wire [16-1:0] node15066;
	wire [16-1:0] node15069;
	wire [16-1:0] node15070;
	wire [16-1:0] node15071;
	wire [16-1:0] node15072;
	wire [16-1:0] node15073;
	wire [16-1:0] node15074;
	wire [16-1:0] node15075;
	wire [16-1:0] node15076;
	wire [16-1:0] node15079;
	wire [16-1:0] node15082;
	wire [16-1:0] node15083;
	wire [16-1:0] node15086;
	wire [16-1:0] node15089;
	wire [16-1:0] node15090;
	wire [16-1:0] node15091;
	wire [16-1:0] node15094;
	wire [16-1:0] node15097;
	wire [16-1:0] node15098;
	wire [16-1:0] node15101;
	wire [16-1:0] node15104;
	wire [16-1:0] node15105;
	wire [16-1:0] node15106;
	wire [16-1:0] node15108;
	wire [16-1:0] node15111;
	wire [16-1:0] node15112;
	wire [16-1:0] node15115;
	wire [16-1:0] node15118;
	wire [16-1:0] node15119;
	wire [16-1:0] node15120;
	wire [16-1:0] node15123;
	wire [16-1:0] node15126;
	wire [16-1:0] node15127;
	wire [16-1:0] node15130;
	wire [16-1:0] node15133;
	wire [16-1:0] node15134;
	wire [16-1:0] node15135;
	wire [16-1:0] node15136;
	wire [16-1:0] node15137;
	wire [16-1:0] node15140;
	wire [16-1:0] node15143;
	wire [16-1:0] node15144;
	wire [16-1:0] node15147;
	wire [16-1:0] node15150;
	wire [16-1:0] node15151;
	wire [16-1:0] node15153;
	wire [16-1:0] node15156;
	wire [16-1:0] node15157;
	wire [16-1:0] node15160;
	wire [16-1:0] node15163;
	wire [16-1:0] node15164;
	wire [16-1:0] node15165;
	wire [16-1:0] node15166;
	wire [16-1:0] node15169;
	wire [16-1:0] node15172;
	wire [16-1:0] node15173;
	wire [16-1:0] node15176;
	wire [16-1:0] node15179;
	wire [16-1:0] node15180;
	wire [16-1:0] node15181;
	wire [16-1:0] node15184;
	wire [16-1:0] node15187;
	wire [16-1:0] node15189;
	wire [16-1:0] node15192;
	wire [16-1:0] node15193;
	wire [16-1:0] node15194;
	wire [16-1:0] node15195;
	wire [16-1:0] node15196;
	wire [16-1:0] node15198;
	wire [16-1:0] node15201;
	wire [16-1:0] node15202;
	wire [16-1:0] node15205;
	wire [16-1:0] node15208;
	wire [16-1:0] node15209;
	wire [16-1:0] node15210;
	wire [16-1:0] node15213;
	wire [16-1:0] node15216;
	wire [16-1:0] node15217;
	wire [16-1:0] node15220;
	wire [16-1:0] node15223;
	wire [16-1:0] node15224;
	wire [16-1:0] node15225;
	wire [16-1:0] node15226;
	wire [16-1:0] node15229;
	wire [16-1:0] node15232;
	wire [16-1:0] node15233;
	wire [16-1:0] node15236;
	wire [16-1:0] node15239;
	wire [16-1:0] node15240;
	wire [16-1:0] node15241;
	wire [16-1:0] node15244;
	wire [16-1:0] node15247;
	wire [16-1:0] node15248;
	wire [16-1:0] node15251;
	wire [16-1:0] node15254;
	wire [16-1:0] node15255;
	wire [16-1:0] node15256;
	wire [16-1:0] node15257;
	wire [16-1:0] node15259;
	wire [16-1:0] node15262;
	wire [16-1:0] node15263;
	wire [16-1:0] node15266;
	wire [16-1:0] node15269;
	wire [16-1:0] node15270;
	wire [16-1:0] node15271;
	wire [16-1:0] node15274;
	wire [16-1:0] node15277;
	wire [16-1:0] node15278;
	wire [16-1:0] node15281;
	wire [16-1:0] node15284;
	wire [16-1:0] node15285;
	wire [16-1:0] node15286;
	wire [16-1:0] node15287;
	wire [16-1:0] node15290;
	wire [16-1:0] node15293;
	wire [16-1:0] node15294;
	wire [16-1:0] node15297;
	wire [16-1:0] node15300;
	wire [16-1:0] node15301;
	wire [16-1:0] node15303;
	wire [16-1:0] node15306;
	wire [16-1:0] node15307;
	wire [16-1:0] node15310;
	wire [16-1:0] node15313;
	wire [16-1:0] node15314;
	wire [16-1:0] node15315;
	wire [16-1:0] node15316;
	wire [16-1:0] node15317;
	wire [16-1:0] node15318;
	wire [16-1:0] node15319;
	wire [16-1:0] node15322;
	wire [16-1:0] node15325;
	wire [16-1:0] node15326;
	wire [16-1:0] node15329;
	wire [16-1:0] node15332;
	wire [16-1:0] node15333;
	wire [16-1:0] node15334;
	wire [16-1:0] node15337;
	wire [16-1:0] node15340;
	wire [16-1:0] node15341;
	wire [16-1:0] node15344;
	wire [16-1:0] node15347;
	wire [16-1:0] node15348;
	wire [16-1:0] node15349;
	wire [16-1:0] node15350;
	wire [16-1:0] node15353;
	wire [16-1:0] node15356;
	wire [16-1:0] node15357;
	wire [16-1:0] node15360;
	wire [16-1:0] node15363;
	wire [16-1:0] node15364;
	wire [16-1:0] node15365;
	wire [16-1:0] node15368;
	wire [16-1:0] node15371;
	wire [16-1:0] node15372;
	wire [16-1:0] node15375;
	wire [16-1:0] node15378;
	wire [16-1:0] node15379;
	wire [16-1:0] node15380;
	wire [16-1:0] node15381;
	wire [16-1:0] node15382;
	wire [16-1:0] node15385;
	wire [16-1:0] node15388;
	wire [16-1:0] node15389;
	wire [16-1:0] node15392;
	wire [16-1:0] node15395;
	wire [16-1:0] node15396;
	wire [16-1:0] node15398;
	wire [16-1:0] node15401;
	wire [16-1:0] node15402;
	wire [16-1:0] node15405;
	wire [16-1:0] node15408;
	wire [16-1:0] node15409;
	wire [16-1:0] node15410;
	wire [16-1:0] node15411;
	wire [16-1:0] node15414;
	wire [16-1:0] node15417;
	wire [16-1:0] node15418;
	wire [16-1:0] node15421;
	wire [16-1:0] node15424;
	wire [16-1:0] node15425;
	wire [16-1:0] node15426;
	wire [16-1:0] node15429;
	wire [16-1:0] node15432;
	wire [16-1:0] node15433;
	wire [16-1:0] node15436;
	wire [16-1:0] node15439;
	wire [16-1:0] node15440;
	wire [16-1:0] node15441;
	wire [16-1:0] node15442;
	wire [16-1:0] node15443;
	wire [16-1:0] node15444;
	wire [16-1:0] node15447;
	wire [16-1:0] node15450;
	wire [16-1:0] node15451;
	wire [16-1:0] node15454;
	wire [16-1:0] node15457;
	wire [16-1:0] node15458;
	wire [16-1:0] node15459;
	wire [16-1:0] node15462;
	wire [16-1:0] node15465;
	wire [16-1:0] node15466;
	wire [16-1:0] node15469;
	wire [16-1:0] node15472;
	wire [16-1:0] node15473;
	wire [16-1:0] node15474;
	wire [16-1:0] node15475;
	wire [16-1:0] node15478;
	wire [16-1:0] node15481;
	wire [16-1:0] node15482;
	wire [16-1:0] node15485;
	wire [16-1:0] node15488;
	wire [16-1:0] node15489;
	wire [16-1:0] node15490;
	wire [16-1:0] node15493;
	wire [16-1:0] node15496;
	wire [16-1:0] node15497;
	wire [16-1:0] node15500;
	wire [16-1:0] node15503;
	wire [16-1:0] node15504;
	wire [16-1:0] node15505;
	wire [16-1:0] node15506;
	wire [16-1:0] node15508;
	wire [16-1:0] node15511;
	wire [16-1:0] node15512;
	wire [16-1:0] node15515;
	wire [16-1:0] node15518;
	wire [16-1:0] node15519;
	wire [16-1:0] node15520;
	wire [16-1:0] node15523;
	wire [16-1:0] node15526;
	wire [16-1:0] node15528;
	wire [16-1:0] node15531;
	wire [16-1:0] node15532;
	wire [16-1:0] node15533;
	wire [16-1:0] node15535;
	wire [16-1:0] node15538;
	wire [16-1:0] node15539;
	wire [16-1:0] node15542;
	wire [16-1:0] node15545;
	wire [16-1:0] node15546;
	wire [16-1:0] node15547;
	wire [16-1:0] node15550;
	wire [16-1:0] node15553;
	wire [16-1:0] node15555;
	wire [16-1:0] node15558;
	wire [16-1:0] node15559;
	wire [16-1:0] node15560;
	wire [16-1:0] node15561;
	wire [16-1:0] node15562;
	wire [16-1:0] node15563;
	wire [16-1:0] node15564;
	wire [16-1:0] node15565;
	wire [16-1:0] node15566;
	wire [16-1:0] node15567;
	wire [16-1:0] node15568;
	wire [16-1:0] node15569;
	wire [16-1:0] node15570;
	wire [16-1:0] node15573;
	wire [16-1:0] node15576;
	wire [16-1:0] node15577;
	wire [16-1:0] node15580;
	wire [16-1:0] node15583;
	wire [16-1:0] node15584;
	wire [16-1:0] node15585;
	wire [16-1:0] node15588;
	wire [16-1:0] node15591;
	wire [16-1:0] node15592;
	wire [16-1:0] node15596;
	wire [16-1:0] node15597;
	wire [16-1:0] node15598;
	wire [16-1:0] node15599;
	wire [16-1:0] node15603;
	wire [16-1:0] node15604;
	wire [16-1:0] node15607;
	wire [16-1:0] node15610;
	wire [16-1:0] node15611;
	wire [16-1:0] node15612;
	wire [16-1:0] node15615;
	wire [16-1:0] node15618;
	wire [16-1:0] node15619;
	wire [16-1:0] node15623;
	wire [16-1:0] node15624;
	wire [16-1:0] node15625;
	wire [16-1:0] node15626;
	wire [16-1:0] node15627;
	wire [16-1:0] node15631;
	wire [16-1:0] node15632;
	wire [16-1:0] node15635;
	wire [16-1:0] node15638;
	wire [16-1:0] node15639;
	wire [16-1:0] node15640;
	wire [16-1:0] node15643;
	wire [16-1:0] node15646;
	wire [16-1:0] node15647;
	wire [16-1:0] node15650;
	wire [16-1:0] node15653;
	wire [16-1:0] node15654;
	wire [16-1:0] node15655;
	wire [16-1:0] node15657;
	wire [16-1:0] node15660;
	wire [16-1:0] node15661;
	wire [16-1:0] node15664;
	wire [16-1:0] node15667;
	wire [16-1:0] node15668;
	wire [16-1:0] node15669;
	wire [16-1:0] node15672;
	wire [16-1:0] node15675;
	wire [16-1:0] node15676;
	wire [16-1:0] node15679;
	wire [16-1:0] node15682;
	wire [16-1:0] node15683;
	wire [16-1:0] node15684;
	wire [16-1:0] node15685;
	wire [16-1:0] node15686;
	wire [16-1:0] node15687;
	wire [16-1:0] node15690;
	wire [16-1:0] node15693;
	wire [16-1:0] node15694;
	wire [16-1:0] node15697;
	wire [16-1:0] node15700;
	wire [16-1:0] node15701;
	wire [16-1:0] node15702;
	wire [16-1:0] node15705;
	wire [16-1:0] node15708;
	wire [16-1:0] node15709;
	wire [16-1:0] node15712;
	wire [16-1:0] node15715;
	wire [16-1:0] node15716;
	wire [16-1:0] node15717;
	wire [16-1:0] node15718;
	wire [16-1:0] node15722;
	wire [16-1:0] node15723;
	wire [16-1:0] node15726;
	wire [16-1:0] node15729;
	wire [16-1:0] node15730;
	wire [16-1:0] node15732;
	wire [16-1:0] node15735;
	wire [16-1:0] node15736;
	wire [16-1:0] node15739;
	wire [16-1:0] node15742;
	wire [16-1:0] node15743;
	wire [16-1:0] node15744;
	wire [16-1:0] node15745;
	wire [16-1:0] node15746;
	wire [16-1:0] node15749;
	wire [16-1:0] node15752;
	wire [16-1:0] node15753;
	wire [16-1:0] node15756;
	wire [16-1:0] node15759;
	wire [16-1:0] node15760;
	wire [16-1:0] node15761;
	wire [16-1:0] node15764;
	wire [16-1:0] node15767;
	wire [16-1:0] node15768;
	wire [16-1:0] node15771;
	wire [16-1:0] node15774;
	wire [16-1:0] node15775;
	wire [16-1:0] node15776;
	wire [16-1:0] node15777;
	wire [16-1:0] node15780;
	wire [16-1:0] node15783;
	wire [16-1:0] node15784;
	wire [16-1:0] node15787;
	wire [16-1:0] node15790;
	wire [16-1:0] node15791;
	wire [16-1:0] node15792;
	wire [16-1:0] node15795;
	wire [16-1:0] node15798;
	wire [16-1:0] node15800;
	wire [16-1:0] node15803;
	wire [16-1:0] node15804;
	wire [16-1:0] node15805;
	wire [16-1:0] node15806;
	wire [16-1:0] node15807;
	wire [16-1:0] node15808;
	wire [16-1:0] node15810;
	wire [16-1:0] node15813;
	wire [16-1:0] node15814;
	wire [16-1:0] node15817;
	wire [16-1:0] node15820;
	wire [16-1:0] node15821;
	wire [16-1:0] node15822;
	wire [16-1:0] node15825;
	wire [16-1:0] node15828;
	wire [16-1:0] node15829;
	wire [16-1:0] node15832;
	wire [16-1:0] node15835;
	wire [16-1:0] node15836;
	wire [16-1:0] node15837;
	wire [16-1:0] node15838;
	wire [16-1:0] node15841;
	wire [16-1:0] node15844;
	wire [16-1:0] node15845;
	wire [16-1:0] node15848;
	wire [16-1:0] node15851;
	wire [16-1:0] node15852;
	wire [16-1:0] node15853;
	wire [16-1:0] node15856;
	wire [16-1:0] node15859;
	wire [16-1:0] node15860;
	wire [16-1:0] node15864;
	wire [16-1:0] node15865;
	wire [16-1:0] node15866;
	wire [16-1:0] node15867;
	wire [16-1:0] node15868;
	wire [16-1:0] node15871;
	wire [16-1:0] node15874;
	wire [16-1:0] node15875;
	wire [16-1:0] node15878;
	wire [16-1:0] node15881;
	wire [16-1:0] node15882;
	wire [16-1:0] node15883;
	wire [16-1:0] node15886;
	wire [16-1:0] node15889;
	wire [16-1:0] node15890;
	wire [16-1:0] node15893;
	wire [16-1:0] node15896;
	wire [16-1:0] node15897;
	wire [16-1:0] node15898;
	wire [16-1:0] node15899;
	wire [16-1:0] node15902;
	wire [16-1:0] node15905;
	wire [16-1:0] node15906;
	wire [16-1:0] node15909;
	wire [16-1:0] node15912;
	wire [16-1:0] node15913;
	wire [16-1:0] node15914;
	wire [16-1:0] node15917;
	wire [16-1:0] node15920;
	wire [16-1:0] node15921;
	wire [16-1:0] node15924;
	wire [16-1:0] node15927;
	wire [16-1:0] node15928;
	wire [16-1:0] node15929;
	wire [16-1:0] node15930;
	wire [16-1:0] node15931;
	wire [16-1:0] node15932;
	wire [16-1:0] node15935;
	wire [16-1:0] node15938;
	wire [16-1:0] node15939;
	wire [16-1:0] node15942;
	wire [16-1:0] node15945;
	wire [16-1:0] node15946;
	wire [16-1:0] node15947;
	wire [16-1:0] node15950;
	wire [16-1:0] node15953;
	wire [16-1:0] node15954;
	wire [16-1:0] node15957;
	wire [16-1:0] node15960;
	wire [16-1:0] node15961;
	wire [16-1:0] node15962;
	wire [16-1:0] node15963;
	wire [16-1:0] node15966;
	wire [16-1:0] node15969;
	wire [16-1:0] node15970;
	wire [16-1:0] node15973;
	wire [16-1:0] node15976;
	wire [16-1:0] node15977;
	wire [16-1:0] node15978;
	wire [16-1:0] node15981;
	wire [16-1:0] node15984;
	wire [16-1:0] node15985;
	wire [16-1:0] node15988;
	wire [16-1:0] node15991;
	wire [16-1:0] node15992;
	wire [16-1:0] node15993;
	wire [16-1:0] node15994;
	wire [16-1:0] node15995;
	wire [16-1:0] node15998;
	wire [16-1:0] node16001;
	wire [16-1:0] node16003;
	wire [16-1:0] node16006;
	wire [16-1:0] node16007;
	wire [16-1:0] node16008;
	wire [16-1:0] node16011;
	wire [16-1:0] node16014;
	wire [16-1:0] node16015;
	wire [16-1:0] node16019;
	wire [16-1:0] node16020;
	wire [16-1:0] node16021;
	wire [16-1:0] node16022;
	wire [16-1:0] node16025;
	wire [16-1:0] node16028;
	wire [16-1:0] node16029;
	wire [16-1:0] node16032;
	wire [16-1:0] node16035;
	wire [16-1:0] node16036;
	wire [16-1:0] node16037;
	wire [16-1:0] node16040;
	wire [16-1:0] node16043;
	wire [16-1:0] node16044;
	wire [16-1:0] node16047;
	wire [16-1:0] node16050;
	wire [16-1:0] node16051;
	wire [16-1:0] node16052;
	wire [16-1:0] node16053;
	wire [16-1:0] node16054;
	wire [16-1:0] node16055;
	wire [16-1:0] node16056;
	wire [16-1:0] node16057;
	wire [16-1:0] node16060;
	wire [16-1:0] node16063;
	wire [16-1:0] node16064;
	wire [16-1:0] node16067;
	wire [16-1:0] node16070;
	wire [16-1:0] node16071;
	wire [16-1:0] node16072;
	wire [16-1:0] node16075;
	wire [16-1:0] node16078;
	wire [16-1:0] node16079;
	wire [16-1:0] node16083;
	wire [16-1:0] node16084;
	wire [16-1:0] node16085;
	wire [16-1:0] node16086;
	wire [16-1:0] node16089;
	wire [16-1:0] node16092;
	wire [16-1:0] node16093;
	wire [16-1:0] node16096;
	wire [16-1:0] node16099;
	wire [16-1:0] node16100;
	wire [16-1:0] node16101;
	wire [16-1:0] node16104;
	wire [16-1:0] node16107;
	wire [16-1:0] node16108;
	wire [16-1:0] node16111;
	wire [16-1:0] node16114;
	wire [16-1:0] node16115;
	wire [16-1:0] node16116;
	wire [16-1:0] node16117;
	wire [16-1:0] node16118;
	wire [16-1:0] node16121;
	wire [16-1:0] node16124;
	wire [16-1:0] node16125;
	wire [16-1:0] node16128;
	wire [16-1:0] node16131;
	wire [16-1:0] node16132;
	wire [16-1:0] node16133;
	wire [16-1:0] node16136;
	wire [16-1:0] node16139;
	wire [16-1:0] node16140;
	wire [16-1:0] node16143;
	wire [16-1:0] node16146;
	wire [16-1:0] node16147;
	wire [16-1:0] node16148;
	wire [16-1:0] node16149;
	wire [16-1:0] node16152;
	wire [16-1:0] node16155;
	wire [16-1:0] node16156;
	wire [16-1:0] node16159;
	wire [16-1:0] node16162;
	wire [16-1:0] node16163;
	wire [16-1:0] node16165;
	wire [16-1:0] node16168;
	wire [16-1:0] node16169;
	wire [16-1:0] node16172;
	wire [16-1:0] node16175;
	wire [16-1:0] node16176;
	wire [16-1:0] node16177;
	wire [16-1:0] node16178;
	wire [16-1:0] node16179;
	wire [16-1:0] node16180;
	wire [16-1:0] node16183;
	wire [16-1:0] node16186;
	wire [16-1:0] node16187;
	wire [16-1:0] node16190;
	wire [16-1:0] node16193;
	wire [16-1:0] node16194;
	wire [16-1:0] node16195;
	wire [16-1:0] node16198;
	wire [16-1:0] node16201;
	wire [16-1:0] node16202;
	wire [16-1:0] node16206;
	wire [16-1:0] node16207;
	wire [16-1:0] node16208;
	wire [16-1:0] node16209;
	wire [16-1:0] node16212;
	wire [16-1:0] node16215;
	wire [16-1:0] node16216;
	wire [16-1:0] node16219;
	wire [16-1:0] node16222;
	wire [16-1:0] node16223;
	wire [16-1:0] node16224;
	wire [16-1:0] node16228;
	wire [16-1:0] node16229;
	wire [16-1:0] node16232;
	wire [16-1:0] node16235;
	wire [16-1:0] node16236;
	wire [16-1:0] node16237;
	wire [16-1:0] node16238;
	wire [16-1:0] node16239;
	wire [16-1:0] node16242;
	wire [16-1:0] node16245;
	wire [16-1:0] node16246;
	wire [16-1:0] node16249;
	wire [16-1:0] node16252;
	wire [16-1:0] node16253;
	wire [16-1:0] node16254;
	wire [16-1:0] node16257;
	wire [16-1:0] node16260;
	wire [16-1:0] node16261;
	wire [16-1:0] node16264;
	wire [16-1:0] node16267;
	wire [16-1:0] node16268;
	wire [16-1:0] node16269;
	wire [16-1:0] node16270;
	wire [16-1:0] node16273;
	wire [16-1:0] node16276;
	wire [16-1:0] node16277;
	wire [16-1:0] node16281;
	wire [16-1:0] node16282;
	wire [16-1:0] node16284;
	wire [16-1:0] node16287;
	wire [16-1:0] node16288;
	wire [16-1:0] node16291;
	wire [16-1:0] node16294;
	wire [16-1:0] node16295;
	wire [16-1:0] node16296;
	wire [16-1:0] node16297;
	wire [16-1:0] node16298;
	wire [16-1:0] node16299;
	wire [16-1:0] node16300;
	wire [16-1:0] node16303;
	wire [16-1:0] node16306;
	wire [16-1:0] node16307;
	wire [16-1:0] node16311;
	wire [16-1:0] node16312;
	wire [16-1:0] node16313;
	wire [16-1:0] node16316;
	wire [16-1:0] node16319;
	wire [16-1:0] node16320;
	wire [16-1:0] node16323;
	wire [16-1:0] node16326;
	wire [16-1:0] node16327;
	wire [16-1:0] node16328;
	wire [16-1:0] node16329;
	wire [16-1:0] node16332;
	wire [16-1:0] node16335;
	wire [16-1:0] node16336;
	wire [16-1:0] node16340;
	wire [16-1:0] node16341;
	wire [16-1:0] node16342;
	wire [16-1:0] node16345;
	wire [16-1:0] node16348;
	wire [16-1:0] node16349;
	wire [16-1:0] node16352;
	wire [16-1:0] node16355;
	wire [16-1:0] node16356;
	wire [16-1:0] node16357;
	wire [16-1:0] node16358;
	wire [16-1:0] node16359;
	wire [16-1:0] node16362;
	wire [16-1:0] node16365;
	wire [16-1:0] node16366;
	wire [16-1:0] node16370;
	wire [16-1:0] node16371;
	wire [16-1:0] node16372;
	wire [16-1:0] node16375;
	wire [16-1:0] node16378;
	wire [16-1:0] node16379;
	wire [16-1:0] node16382;
	wire [16-1:0] node16385;
	wire [16-1:0] node16386;
	wire [16-1:0] node16387;
	wire [16-1:0] node16388;
	wire [16-1:0] node16391;
	wire [16-1:0] node16394;
	wire [16-1:0] node16395;
	wire [16-1:0] node16398;
	wire [16-1:0] node16401;
	wire [16-1:0] node16402;
	wire [16-1:0] node16403;
	wire [16-1:0] node16406;
	wire [16-1:0] node16409;
	wire [16-1:0] node16410;
	wire [16-1:0] node16413;
	wire [16-1:0] node16416;
	wire [16-1:0] node16417;
	wire [16-1:0] node16418;
	wire [16-1:0] node16419;
	wire [16-1:0] node16420;
	wire [16-1:0] node16421;
	wire [16-1:0] node16424;
	wire [16-1:0] node16427;
	wire [16-1:0] node16428;
	wire [16-1:0] node16431;
	wire [16-1:0] node16434;
	wire [16-1:0] node16435;
	wire [16-1:0] node16436;
	wire [16-1:0] node16439;
	wire [16-1:0] node16442;
	wire [16-1:0] node16443;
	wire [16-1:0] node16447;
	wire [16-1:0] node16448;
	wire [16-1:0] node16449;
	wire [16-1:0] node16450;
	wire [16-1:0] node16453;
	wire [16-1:0] node16456;
	wire [16-1:0] node16457;
	wire [16-1:0] node16460;
	wire [16-1:0] node16463;
	wire [16-1:0] node16464;
	wire [16-1:0] node16465;
	wire [16-1:0] node16468;
	wire [16-1:0] node16471;
	wire [16-1:0] node16472;
	wire [16-1:0] node16475;
	wire [16-1:0] node16478;
	wire [16-1:0] node16479;
	wire [16-1:0] node16480;
	wire [16-1:0] node16481;
	wire [16-1:0] node16482;
	wire [16-1:0] node16486;
	wire [16-1:0] node16487;
	wire [16-1:0] node16491;
	wire [16-1:0] node16492;
	wire [16-1:0] node16493;
	wire [16-1:0] node16496;
	wire [16-1:0] node16499;
	wire [16-1:0] node16500;
	wire [16-1:0] node16503;
	wire [16-1:0] node16506;
	wire [16-1:0] node16507;
	wire [16-1:0] node16508;
	wire [16-1:0] node16509;
	wire [16-1:0] node16512;
	wire [16-1:0] node16515;
	wire [16-1:0] node16516;
	wire [16-1:0] node16519;
	wire [16-1:0] node16522;
	wire [16-1:0] node16523;
	wire [16-1:0] node16524;
	wire [16-1:0] node16527;
	wire [16-1:0] node16530;
	wire [16-1:0] node16531;
	wire [16-1:0] node16534;
	wire [16-1:0] node16537;
	wire [16-1:0] node16538;
	wire [16-1:0] node16539;
	wire [16-1:0] node16540;
	wire [16-1:0] node16541;
	wire [16-1:0] node16542;
	wire [16-1:0] node16543;
	wire [16-1:0] node16544;
	wire [16-1:0] node16545;
	wire [16-1:0] node16548;
	wire [16-1:0] node16551;
	wire [16-1:0] node16552;
	wire [16-1:0] node16555;
	wire [16-1:0] node16558;
	wire [16-1:0] node16559;
	wire [16-1:0] node16560;
	wire [16-1:0] node16564;
	wire [16-1:0] node16565;
	wire [16-1:0] node16568;
	wire [16-1:0] node16571;
	wire [16-1:0] node16572;
	wire [16-1:0] node16573;
	wire [16-1:0] node16574;
	wire [16-1:0] node16577;
	wire [16-1:0] node16580;
	wire [16-1:0] node16581;
	wire [16-1:0] node16584;
	wire [16-1:0] node16587;
	wire [16-1:0] node16588;
	wire [16-1:0] node16589;
	wire [16-1:0] node16592;
	wire [16-1:0] node16595;
	wire [16-1:0] node16597;
	wire [16-1:0] node16600;
	wire [16-1:0] node16601;
	wire [16-1:0] node16602;
	wire [16-1:0] node16603;
	wire [16-1:0] node16604;
	wire [16-1:0] node16607;
	wire [16-1:0] node16610;
	wire [16-1:0] node16611;
	wire [16-1:0] node16614;
	wire [16-1:0] node16617;
	wire [16-1:0] node16618;
	wire [16-1:0] node16619;
	wire [16-1:0] node16622;
	wire [16-1:0] node16625;
	wire [16-1:0] node16626;
	wire [16-1:0] node16629;
	wire [16-1:0] node16632;
	wire [16-1:0] node16633;
	wire [16-1:0] node16634;
	wire [16-1:0] node16635;
	wire [16-1:0] node16638;
	wire [16-1:0] node16641;
	wire [16-1:0] node16642;
	wire [16-1:0] node16645;
	wire [16-1:0] node16648;
	wire [16-1:0] node16649;
	wire [16-1:0] node16650;
	wire [16-1:0] node16653;
	wire [16-1:0] node16656;
	wire [16-1:0] node16657;
	wire [16-1:0] node16661;
	wire [16-1:0] node16662;
	wire [16-1:0] node16663;
	wire [16-1:0] node16664;
	wire [16-1:0] node16665;
	wire [16-1:0] node16666;
	wire [16-1:0] node16670;
	wire [16-1:0] node16671;
	wire [16-1:0] node16674;
	wire [16-1:0] node16677;
	wire [16-1:0] node16678;
	wire [16-1:0] node16679;
	wire [16-1:0] node16682;
	wire [16-1:0] node16685;
	wire [16-1:0] node16686;
	wire [16-1:0] node16689;
	wire [16-1:0] node16692;
	wire [16-1:0] node16693;
	wire [16-1:0] node16694;
	wire [16-1:0] node16695;
	wire [16-1:0] node16698;
	wire [16-1:0] node16701;
	wire [16-1:0] node16702;
	wire [16-1:0] node16705;
	wire [16-1:0] node16708;
	wire [16-1:0] node16709;
	wire [16-1:0] node16710;
	wire [16-1:0] node16713;
	wire [16-1:0] node16716;
	wire [16-1:0] node16718;
	wire [16-1:0] node16721;
	wire [16-1:0] node16722;
	wire [16-1:0] node16723;
	wire [16-1:0] node16724;
	wire [16-1:0] node16725;
	wire [16-1:0] node16728;
	wire [16-1:0] node16731;
	wire [16-1:0] node16732;
	wire [16-1:0] node16735;
	wire [16-1:0] node16738;
	wire [16-1:0] node16739;
	wire [16-1:0] node16741;
	wire [16-1:0] node16744;
	wire [16-1:0] node16745;
	wire [16-1:0] node16748;
	wire [16-1:0] node16751;
	wire [16-1:0] node16752;
	wire [16-1:0] node16753;
	wire [16-1:0] node16754;
	wire [16-1:0] node16758;
	wire [16-1:0] node16759;
	wire [16-1:0] node16762;
	wire [16-1:0] node16765;
	wire [16-1:0] node16766;
	wire [16-1:0] node16767;
	wire [16-1:0] node16770;
	wire [16-1:0] node16773;
	wire [16-1:0] node16774;
	wire [16-1:0] node16777;
	wire [16-1:0] node16780;
	wire [16-1:0] node16781;
	wire [16-1:0] node16782;
	wire [16-1:0] node16783;
	wire [16-1:0] node16784;
	wire [16-1:0] node16785;
	wire [16-1:0] node16786;
	wire [16-1:0] node16789;
	wire [16-1:0] node16792;
	wire [16-1:0] node16793;
	wire [16-1:0] node16796;
	wire [16-1:0] node16799;
	wire [16-1:0] node16800;
	wire [16-1:0] node16801;
	wire [16-1:0] node16804;
	wire [16-1:0] node16807;
	wire [16-1:0] node16808;
	wire [16-1:0] node16811;
	wire [16-1:0] node16814;
	wire [16-1:0] node16815;
	wire [16-1:0] node16816;
	wire [16-1:0] node16817;
	wire [16-1:0] node16820;
	wire [16-1:0] node16823;
	wire [16-1:0] node16824;
	wire [16-1:0] node16827;
	wire [16-1:0] node16830;
	wire [16-1:0] node16831;
	wire [16-1:0] node16832;
	wire [16-1:0] node16835;
	wire [16-1:0] node16838;
	wire [16-1:0] node16839;
	wire [16-1:0] node16842;
	wire [16-1:0] node16845;
	wire [16-1:0] node16846;
	wire [16-1:0] node16847;
	wire [16-1:0] node16848;
	wire [16-1:0] node16849;
	wire [16-1:0] node16852;
	wire [16-1:0] node16855;
	wire [16-1:0] node16856;
	wire [16-1:0] node16859;
	wire [16-1:0] node16862;
	wire [16-1:0] node16863;
	wire [16-1:0] node16864;
	wire [16-1:0] node16867;
	wire [16-1:0] node16870;
	wire [16-1:0] node16871;
	wire [16-1:0] node16874;
	wire [16-1:0] node16877;
	wire [16-1:0] node16878;
	wire [16-1:0] node16879;
	wire [16-1:0] node16880;
	wire [16-1:0] node16883;
	wire [16-1:0] node16886;
	wire [16-1:0] node16887;
	wire [16-1:0] node16891;
	wire [16-1:0] node16892;
	wire [16-1:0] node16893;
	wire [16-1:0] node16896;
	wire [16-1:0] node16899;
	wire [16-1:0] node16901;
	wire [16-1:0] node16904;
	wire [16-1:0] node16905;
	wire [16-1:0] node16906;
	wire [16-1:0] node16907;
	wire [16-1:0] node16908;
	wire [16-1:0] node16909;
	wire [16-1:0] node16912;
	wire [16-1:0] node16915;
	wire [16-1:0] node16916;
	wire [16-1:0] node16919;
	wire [16-1:0] node16922;
	wire [16-1:0] node16923;
	wire [16-1:0] node16924;
	wire [16-1:0] node16927;
	wire [16-1:0] node16930;
	wire [16-1:0] node16931;
	wire [16-1:0] node16935;
	wire [16-1:0] node16936;
	wire [16-1:0] node16937;
	wire [16-1:0] node16939;
	wire [16-1:0] node16942;
	wire [16-1:0] node16943;
	wire [16-1:0] node16946;
	wire [16-1:0] node16949;
	wire [16-1:0] node16950;
	wire [16-1:0] node16951;
	wire [16-1:0] node16954;
	wire [16-1:0] node16957;
	wire [16-1:0] node16958;
	wire [16-1:0] node16961;
	wire [16-1:0] node16964;
	wire [16-1:0] node16965;
	wire [16-1:0] node16966;
	wire [16-1:0] node16967;
	wire [16-1:0] node16968;
	wire [16-1:0] node16971;
	wire [16-1:0] node16974;
	wire [16-1:0] node16975;
	wire [16-1:0] node16978;
	wire [16-1:0] node16981;
	wire [16-1:0] node16982;
	wire [16-1:0] node16983;
	wire [16-1:0] node16986;
	wire [16-1:0] node16989;
	wire [16-1:0] node16990;
	wire [16-1:0] node16993;
	wire [16-1:0] node16996;
	wire [16-1:0] node16997;
	wire [16-1:0] node16998;
	wire [16-1:0] node16999;
	wire [16-1:0] node17002;
	wire [16-1:0] node17005;
	wire [16-1:0] node17006;
	wire [16-1:0] node17009;
	wire [16-1:0] node17012;
	wire [16-1:0] node17013;
	wire [16-1:0] node17014;
	wire [16-1:0] node17017;
	wire [16-1:0] node17020;
	wire [16-1:0] node17022;
	wire [16-1:0] node17025;
	wire [16-1:0] node17026;
	wire [16-1:0] node17027;
	wire [16-1:0] node17028;
	wire [16-1:0] node17029;
	wire [16-1:0] node17030;
	wire [16-1:0] node17031;
	wire [16-1:0] node17032;
	wire [16-1:0] node17035;
	wire [16-1:0] node17038;
	wire [16-1:0] node17039;
	wire [16-1:0] node17042;
	wire [16-1:0] node17045;
	wire [16-1:0] node17046;
	wire [16-1:0] node17047;
	wire [16-1:0] node17050;
	wire [16-1:0] node17053;
	wire [16-1:0] node17054;
	wire [16-1:0] node17057;
	wire [16-1:0] node17060;
	wire [16-1:0] node17061;
	wire [16-1:0] node17062;
	wire [16-1:0] node17063;
	wire [16-1:0] node17066;
	wire [16-1:0] node17069;
	wire [16-1:0] node17070;
	wire [16-1:0] node17073;
	wire [16-1:0] node17076;
	wire [16-1:0] node17077;
	wire [16-1:0] node17078;
	wire [16-1:0] node17081;
	wire [16-1:0] node17084;
	wire [16-1:0] node17085;
	wire [16-1:0] node17088;
	wire [16-1:0] node17091;
	wire [16-1:0] node17092;
	wire [16-1:0] node17093;
	wire [16-1:0] node17094;
	wire [16-1:0] node17095;
	wire [16-1:0] node17098;
	wire [16-1:0] node17101;
	wire [16-1:0] node17102;
	wire [16-1:0] node17105;
	wire [16-1:0] node17108;
	wire [16-1:0] node17109;
	wire [16-1:0] node17110;
	wire [16-1:0] node17113;
	wire [16-1:0] node17116;
	wire [16-1:0] node17117;
	wire [16-1:0] node17121;
	wire [16-1:0] node17122;
	wire [16-1:0] node17123;
	wire [16-1:0] node17124;
	wire [16-1:0] node17127;
	wire [16-1:0] node17130;
	wire [16-1:0] node17131;
	wire [16-1:0] node17134;
	wire [16-1:0] node17137;
	wire [16-1:0] node17138;
	wire [16-1:0] node17140;
	wire [16-1:0] node17143;
	wire [16-1:0] node17144;
	wire [16-1:0] node17148;
	wire [16-1:0] node17149;
	wire [16-1:0] node17150;
	wire [16-1:0] node17151;
	wire [16-1:0] node17152;
	wire [16-1:0] node17153;
	wire [16-1:0] node17156;
	wire [16-1:0] node17159;
	wire [16-1:0] node17160;
	wire [16-1:0] node17164;
	wire [16-1:0] node17165;
	wire [16-1:0] node17166;
	wire [16-1:0] node17170;
	wire [16-1:0] node17171;
	wire [16-1:0] node17174;
	wire [16-1:0] node17177;
	wire [16-1:0] node17178;
	wire [16-1:0] node17179;
	wire [16-1:0] node17180;
	wire [16-1:0] node17183;
	wire [16-1:0] node17186;
	wire [16-1:0] node17187;
	wire [16-1:0] node17190;
	wire [16-1:0] node17193;
	wire [16-1:0] node17194;
	wire [16-1:0] node17195;
	wire [16-1:0] node17198;
	wire [16-1:0] node17201;
	wire [16-1:0] node17202;
	wire [16-1:0] node17205;
	wire [16-1:0] node17208;
	wire [16-1:0] node17209;
	wire [16-1:0] node17210;
	wire [16-1:0] node17211;
	wire [16-1:0] node17212;
	wire [16-1:0] node17215;
	wire [16-1:0] node17218;
	wire [16-1:0] node17219;
	wire [16-1:0] node17222;
	wire [16-1:0] node17225;
	wire [16-1:0] node17226;
	wire [16-1:0] node17227;
	wire [16-1:0] node17230;
	wire [16-1:0] node17233;
	wire [16-1:0] node17234;
	wire [16-1:0] node17237;
	wire [16-1:0] node17240;
	wire [16-1:0] node17241;
	wire [16-1:0] node17242;
	wire [16-1:0] node17243;
	wire [16-1:0] node17246;
	wire [16-1:0] node17249;
	wire [16-1:0] node17250;
	wire [16-1:0] node17253;
	wire [16-1:0] node17256;
	wire [16-1:0] node17257;
	wire [16-1:0] node17258;
	wire [16-1:0] node17261;
	wire [16-1:0] node17264;
	wire [16-1:0] node17265;
	wire [16-1:0] node17268;
	wire [16-1:0] node17271;
	wire [16-1:0] node17272;
	wire [16-1:0] node17273;
	wire [16-1:0] node17274;
	wire [16-1:0] node17275;
	wire [16-1:0] node17276;
	wire [16-1:0] node17277;
	wire [16-1:0] node17280;
	wire [16-1:0] node17283;
	wire [16-1:0] node17286;
	wire [16-1:0] node17287;
	wire [16-1:0] node17288;
	wire [16-1:0] node17291;
	wire [16-1:0] node17294;
	wire [16-1:0] node17296;
	wire [16-1:0] node17299;
	wire [16-1:0] node17300;
	wire [16-1:0] node17301;
	wire [16-1:0] node17302;
	wire [16-1:0] node17305;
	wire [16-1:0] node17308;
	wire [16-1:0] node17309;
	wire [16-1:0] node17312;
	wire [16-1:0] node17315;
	wire [16-1:0] node17316;
	wire [16-1:0] node17317;
	wire [16-1:0] node17320;
	wire [16-1:0] node17323;
	wire [16-1:0] node17324;
	wire [16-1:0] node17327;
	wire [16-1:0] node17330;
	wire [16-1:0] node17331;
	wire [16-1:0] node17332;
	wire [16-1:0] node17333;
	wire [16-1:0] node17334;
	wire [16-1:0] node17337;
	wire [16-1:0] node17340;
	wire [16-1:0] node17341;
	wire [16-1:0] node17344;
	wire [16-1:0] node17347;
	wire [16-1:0] node17348;
	wire [16-1:0] node17349;
	wire [16-1:0] node17352;
	wire [16-1:0] node17355;
	wire [16-1:0] node17357;
	wire [16-1:0] node17360;
	wire [16-1:0] node17361;
	wire [16-1:0] node17362;
	wire [16-1:0] node17363;
	wire [16-1:0] node17366;
	wire [16-1:0] node17369;
	wire [16-1:0] node17370;
	wire [16-1:0] node17373;
	wire [16-1:0] node17376;
	wire [16-1:0] node17377;
	wire [16-1:0] node17378;
	wire [16-1:0] node17381;
	wire [16-1:0] node17384;
	wire [16-1:0] node17385;
	wire [16-1:0] node17388;
	wire [16-1:0] node17391;
	wire [16-1:0] node17392;
	wire [16-1:0] node17393;
	wire [16-1:0] node17394;
	wire [16-1:0] node17395;
	wire [16-1:0] node17397;
	wire [16-1:0] node17400;
	wire [16-1:0] node17401;
	wire [16-1:0] node17404;
	wire [16-1:0] node17407;
	wire [16-1:0] node17408;
	wire [16-1:0] node17409;
	wire [16-1:0] node17412;
	wire [16-1:0] node17415;
	wire [16-1:0] node17418;
	wire [16-1:0] node17419;
	wire [16-1:0] node17420;
	wire [16-1:0] node17421;
	wire [16-1:0] node17424;
	wire [16-1:0] node17427;
	wire [16-1:0] node17428;
	wire [16-1:0] node17431;
	wire [16-1:0] node17434;
	wire [16-1:0] node17435;
	wire [16-1:0] node17436;
	wire [16-1:0] node17439;
	wire [16-1:0] node17442;
	wire [16-1:0] node17443;
	wire [16-1:0] node17446;
	wire [16-1:0] node17449;
	wire [16-1:0] node17450;
	wire [16-1:0] node17451;
	wire [16-1:0] node17452;
	wire [16-1:0] node17453;
	wire [16-1:0] node17456;
	wire [16-1:0] node17459;
	wire [16-1:0] node17460;
	wire [16-1:0] node17463;
	wire [16-1:0] node17466;
	wire [16-1:0] node17467;
	wire [16-1:0] node17468;
	wire [16-1:0] node17471;
	wire [16-1:0] node17474;
	wire [16-1:0] node17475;
	wire [16-1:0] node17478;
	wire [16-1:0] node17481;
	wire [16-1:0] node17482;
	wire [16-1:0] node17483;
	wire [16-1:0] node17484;
	wire [16-1:0] node17487;
	wire [16-1:0] node17491;
	wire [16-1:0] node17492;
	wire [16-1:0] node17493;
	wire [16-1:0] node17496;
	wire [16-1:0] node17499;
	wire [16-1:0] node17500;
	wire [16-1:0] node17503;
	wire [16-1:0] node17506;
	wire [16-1:0] node17507;
	wire [16-1:0] node17508;
	wire [16-1:0] node17509;
	wire [16-1:0] node17510;
	wire [16-1:0] node17511;
	wire [16-1:0] node17512;
	wire [16-1:0] node17513;
	wire [16-1:0] node17514;
	wire [16-1:0] node17515;
	wire [16-1:0] node17518;
	wire [16-1:0] node17521;
	wire [16-1:0] node17522;
	wire [16-1:0] node17525;
	wire [16-1:0] node17528;
	wire [16-1:0] node17529;
	wire [16-1:0] node17530;
	wire [16-1:0] node17533;
	wire [16-1:0] node17536;
	wire [16-1:0] node17537;
	wire [16-1:0] node17540;
	wire [16-1:0] node17543;
	wire [16-1:0] node17544;
	wire [16-1:0] node17545;
	wire [16-1:0] node17546;
	wire [16-1:0] node17549;
	wire [16-1:0] node17552;
	wire [16-1:0] node17553;
	wire [16-1:0] node17556;
	wire [16-1:0] node17559;
	wire [16-1:0] node17560;
	wire [16-1:0] node17561;
	wire [16-1:0] node17564;
	wire [16-1:0] node17567;
	wire [16-1:0] node17568;
	wire [16-1:0] node17571;
	wire [16-1:0] node17574;
	wire [16-1:0] node17575;
	wire [16-1:0] node17576;
	wire [16-1:0] node17577;
	wire [16-1:0] node17578;
	wire [16-1:0] node17581;
	wire [16-1:0] node17584;
	wire [16-1:0] node17585;
	wire [16-1:0] node17588;
	wire [16-1:0] node17591;
	wire [16-1:0] node17592;
	wire [16-1:0] node17593;
	wire [16-1:0] node17596;
	wire [16-1:0] node17599;
	wire [16-1:0] node17600;
	wire [16-1:0] node17603;
	wire [16-1:0] node17606;
	wire [16-1:0] node17607;
	wire [16-1:0] node17608;
	wire [16-1:0] node17609;
	wire [16-1:0] node17612;
	wire [16-1:0] node17615;
	wire [16-1:0] node17616;
	wire [16-1:0] node17620;
	wire [16-1:0] node17621;
	wire [16-1:0] node17622;
	wire [16-1:0] node17625;
	wire [16-1:0] node17628;
	wire [16-1:0] node17629;
	wire [16-1:0] node17632;
	wire [16-1:0] node17635;
	wire [16-1:0] node17636;
	wire [16-1:0] node17637;
	wire [16-1:0] node17638;
	wire [16-1:0] node17639;
	wire [16-1:0] node17641;
	wire [16-1:0] node17644;
	wire [16-1:0] node17645;
	wire [16-1:0] node17648;
	wire [16-1:0] node17651;
	wire [16-1:0] node17652;
	wire [16-1:0] node17653;
	wire [16-1:0] node17656;
	wire [16-1:0] node17659;
	wire [16-1:0] node17660;
	wire [16-1:0] node17663;
	wire [16-1:0] node17666;
	wire [16-1:0] node17667;
	wire [16-1:0] node17668;
	wire [16-1:0] node17669;
	wire [16-1:0] node17672;
	wire [16-1:0] node17675;
	wire [16-1:0] node17676;
	wire [16-1:0] node17679;
	wire [16-1:0] node17682;
	wire [16-1:0] node17683;
	wire [16-1:0] node17684;
	wire [16-1:0] node17687;
	wire [16-1:0] node17690;
	wire [16-1:0] node17691;
	wire [16-1:0] node17694;
	wire [16-1:0] node17697;
	wire [16-1:0] node17698;
	wire [16-1:0] node17699;
	wire [16-1:0] node17700;
	wire [16-1:0] node17702;
	wire [16-1:0] node17705;
	wire [16-1:0] node17706;
	wire [16-1:0] node17709;
	wire [16-1:0] node17712;
	wire [16-1:0] node17713;
	wire [16-1:0] node17714;
	wire [16-1:0] node17717;
	wire [16-1:0] node17720;
	wire [16-1:0] node17722;
	wire [16-1:0] node17725;
	wire [16-1:0] node17726;
	wire [16-1:0] node17727;
	wire [16-1:0] node17728;
	wire [16-1:0] node17731;
	wire [16-1:0] node17734;
	wire [16-1:0] node17735;
	wire [16-1:0] node17739;
	wire [16-1:0] node17740;
	wire [16-1:0] node17741;
	wire [16-1:0] node17744;
	wire [16-1:0] node17747;
	wire [16-1:0] node17748;
	wire [16-1:0] node17752;
	wire [16-1:0] node17753;
	wire [16-1:0] node17754;
	wire [16-1:0] node17755;
	wire [16-1:0] node17756;
	wire [16-1:0] node17757;
	wire [16-1:0] node17758;
	wire [16-1:0] node17761;
	wire [16-1:0] node17764;
	wire [16-1:0] node17765;
	wire [16-1:0] node17768;
	wire [16-1:0] node17771;
	wire [16-1:0] node17772;
	wire [16-1:0] node17773;
	wire [16-1:0] node17776;
	wire [16-1:0] node17779;
	wire [16-1:0] node17780;
	wire [16-1:0] node17783;
	wire [16-1:0] node17786;
	wire [16-1:0] node17787;
	wire [16-1:0] node17788;
	wire [16-1:0] node17789;
	wire [16-1:0] node17792;
	wire [16-1:0] node17795;
	wire [16-1:0] node17796;
	wire [16-1:0] node17799;
	wire [16-1:0] node17802;
	wire [16-1:0] node17803;
	wire [16-1:0] node17804;
	wire [16-1:0] node17807;
	wire [16-1:0] node17810;
	wire [16-1:0] node17811;
	wire [16-1:0] node17814;
	wire [16-1:0] node17817;
	wire [16-1:0] node17818;
	wire [16-1:0] node17819;
	wire [16-1:0] node17820;
	wire [16-1:0] node17821;
	wire [16-1:0] node17824;
	wire [16-1:0] node17827;
	wire [16-1:0] node17828;
	wire [16-1:0] node17831;
	wire [16-1:0] node17834;
	wire [16-1:0] node17835;
	wire [16-1:0] node17836;
	wire [16-1:0] node17839;
	wire [16-1:0] node17842;
	wire [16-1:0] node17843;
	wire [16-1:0] node17846;
	wire [16-1:0] node17849;
	wire [16-1:0] node17850;
	wire [16-1:0] node17851;
	wire [16-1:0] node17852;
	wire [16-1:0] node17855;
	wire [16-1:0] node17858;
	wire [16-1:0] node17859;
	wire [16-1:0] node17862;
	wire [16-1:0] node17865;
	wire [16-1:0] node17866;
	wire [16-1:0] node17867;
	wire [16-1:0] node17870;
	wire [16-1:0] node17873;
	wire [16-1:0] node17874;
	wire [16-1:0] node17878;
	wire [16-1:0] node17879;
	wire [16-1:0] node17880;
	wire [16-1:0] node17881;
	wire [16-1:0] node17882;
	wire [16-1:0] node17883;
	wire [16-1:0] node17886;
	wire [16-1:0] node17889;
	wire [16-1:0] node17890;
	wire [16-1:0] node17893;
	wire [16-1:0] node17896;
	wire [16-1:0] node17897;
	wire [16-1:0] node17898;
	wire [16-1:0] node17901;
	wire [16-1:0] node17904;
	wire [16-1:0] node17905;
	wire [16-1:0] node17908;
	wire [16-1:0] node17911;
	wire [16-1:0] node17912;
	wire [16-1:0] node17913;
	wire [16-1:0] node17915;
	wire [16-1:0] node17918;
	wire [16-1:0] node17919;
	wire [16-1:0] node17922;
	wire [16-1:0] node17925;
	wire [16-1:0] node17926;
	wire [16-1:0] node17927;
	wire [16-1:0] node17930;
	wire [16-1:0] node17933;
	wire [16-1:0] node17935;
	wire [16-1:0] node17938;
	wire [16-1:0] node17939;
	wire [16-1:0] node17940;
	wire [16-1:0] node17941;
	wire [16-1:0] node17942;
	wire [16-1:0] node17945;
	wire [16-1:0] node17948;
	wire [16-1:0] node17949;
	wire [16-1:0] node17952;
	wire [16-1:0] node17955;
	wire [16-1:0] node17956;
	wire [16-1:0] node17957;
	wire [16-1:0] node17960;
	wire [16-1:0] node17963;
	wire [16-1:0] node17964;
	wire [16-1:0] node17967;
	wire [16-1:0] node17970;
	wire [16-1:0] node17971;
	wire [16-1:0] node17972;
	wire [16-1:0] node17973;
	wire [16-1:0] node17976;
	wire [16-1:0] node17979;
	wire [16-1:0] node17980;
	wire [16-1:0] node17983;
	wire [16-1:0] node17986;
	wire [16-1:0] node17987;
	wire [16-1:0] node17988;
	wire [16-1:0] node17991;
	wire [16-1:0] node17994;
	wire [16-1:0] node17995;
	wire [16-1:0] node17998;
	wire [16-1:0] node18001;
	wire [16-1:0] node18002;
	wire [16-1:0] node18003;
	wire [16-1:0] node18004;
	wire [16-1:0] node18005;
	wire [16-1:0] node18006;
	wire [16-1:0] node18007;
	wire [16-1:0] node18008;
	wire [16-1:0] node18011;
	wire [16-1:0] node18014;
	wire [16-1:0] node18015;
	wire [16-1:0] node18018;
	wire [16-1:0] node18021;
	wire [16-1:0] node18022;
	wire [16-1:0] node18023;
	wire [16-1:0] node18026;
	wire [16-1:0] node18029;
	wire [16-1:0] node18030;
	wire [16-1:0] node18033;
	wire [16-1:0] node18036;
	wire [16-1:0] node18037;
	wire [16-1:0] node18038;
	wire [16-1:0] node18039;
	wire [16-1:0] node18042;
	wire [16-1:0] node18045;
	wire [16-1:0] node18046;
	wire [16-1:0] node18049;
	wire [16-1:0] node18052;
	wire [16-1:0] node18053;
	wire [16-1:0] node18054;
	wire [16-1:0] node18057;
	wire [16-1:0] node18060;
	wire [16-1:0] node18061;
	wire [16-1:0] node18064;
	wire [16-1:0] node18067;
	wire [16-1:0] node18068;
	wire [16-1:0] node18069;
	wire [16-1:0] node18070;
	wire [16-1:0] node18071;
	wire [16-1:0] node18074;
	wire [16-1:0] node18077;
	wire [16-1:0] node18078;
	wire [16-1:0] node18081;
	wire [16-1:0] node18084;
	wire [16-1:0] node18085;
	wire [16-1:0] node18086;
	wire [16-1:0] node18089;
	wire [16-1:0] node18092;
	wire [16-1:0] node18094;
	wire [16-1:0] node18097;
	wire [16-1:0] node18098;
	wire [16-1:0] node18099;
	wire [16-1:0] node18100;
	wire [16-1:0] node18103;
	wire [16-1:0] node18106;
	wire [16-1:0] node18107;
	wire [16-1:0] node18110;
	wire [16-1:0] node18113;
	wire [16-1:0] node18114;
	wire [16-1:0] node18115;
	wire [16-1:0] node18119;
	wire [16-1:0] node18120;
	wire [16-1:0] node18123;
	wire [16-1:0] node18126;
	wire [16-1:0] node18127;
	wire [16-1:0] node18128;
	wire [16-1:0] node18129;
	wire [16-1:0] node18130;
	wire [16-1:0] node18131;
	wire [16-1:0] node18134;
	wire [16-1:0] node18137;
	wire [16-1:0] node18138;
	wire [16-1:0] node18141;
	wire [16-1:0] node18144;
	wire [16-1:0] node18145;
	wire [16-1:0] node18146;
	wire [16-1:0] node18149;
	wire [16-1:0] node18152;
	wire [16-1:0] node18153;
	wire [16-1:0] node18156;
	wire [16-1:0] node18159;
	wire [16-1:0] node18160;
	wire [16-1:0] node18161;
	wire [16-1:0] node18162;
	wire [16-1:0] node18165;
	wire [16-1:0] node18168;
	wire [16-1:0] node18169;
	wire [16-1:0] node18172;
	wire [16-1:0] node18175;
	wire [16-1:0] node18176;
	wire [16-1:0] node18178;
	wire [16-1:0] node18181;
	wire [16-1:0] node18183;
	wire [16-1:0] node18186;
	wire [16-1:0] node18187;
	wire [16-1:0] node18188;
	wire [16-1:0] node18189;
	wire [16-1:0] node18191;
	wire [16-1:0] node18194;
	wire [16-1:0] node18195;
	wire [16-1:0] node18199;
	wire [16-1:0] node18200;
	wire [16-1:0] node18201;
	wire [16-1:0] node18204;
	wire [16-1:0] node18207;
	wire [16-1:0] node18208;
	wire [16-1:0] node18211;
	wire [16-1:0] node18214;
	wire [16-1:0] node18215;
	wire [16-1:0] node18216;
	wire [16-1:0] node18217;
	wire [16-1:0] node18220;
	wire [16-1:0] node18223;
	wire [16-1:0] node18224;
	wire [16-1:0] node18227;
	wire [16-1:0] node18230;
	wire [16-1:0] node18231;
	wire [16-1:0] node18232;
	wire [16-1:0] node18235;
	wire [16-1:0] node18238;
	wire [16-1:0] node18239;
	wire [16-1:0] node18242;
	wire [16-1:0] node18245;
	wire [16-1:0] node18246;
	wire [16-1:0] node18247;
	wire [16-1:0] node18248;
	wire [16-1:0] node18249;
	wire [16-1:0] node18250;
	wire [16-1:0] node18251;
	wire [16-1:0] node18255;
	wire [16-1:0] node18256;
	wire [16-1:0] node18259;
	wire [16-1:0] node18262;
	wire [16-1:0] node18263;
	wire [16-1:0] node18264;
	wire [16-1:0] node18267;
	wire [16-1:0] node18270;
	wire [16-1:0] node18271;
	wire [16-1:0] node18274;
	wire [16-1:0] node18277;
	wire [16-1:0] node18278;
	wire [16-1:0] node18279;
	wire [16-1:0] node18280;
	wire [16-1:0] node18283;
	wire [16-1:0] node18286;
	wire [16-1:0] node18287;
	wire [16-1:0] node18290;
	wire [16-1:0] node18293;
	wire [16-1:0] node18294;
	wire [16-1:0] node18295;
	wire [16-1:0] node18298;
	wire [16-1:0] node18301;
	wire [16-1:0] node18302;
	wire [16-1:0] node18305;
	wire [16-1:0] node18308;
	wire [16-1:0] node18309;
	wire [16-1:0] node18310;
	wire [16-1:0] node18311;
	wire [16-1:0] node18312;
	wire [16-1:0] node18315;
	wire [16-1:0] node18318;
	wire [16-1:0] node18319;
	wire [16-1:0] node18322;
	wire [16-1:0] node18325;
	wire [16-1:0] node18326;
	wire [16-1:0] node18327;
	wire [16-1:0] node18330;
	wire [16-1:0] node18333;
	wire [16-1:0] node18334;
	wire [16-1:0] node18337;
	wire [16-1:0] node18340;
	wire [16-1:0] node18341;
	wire [16-1:0] node18342;
	wire [16-1:0] node18343;
	wire [16-1:0] node18347;
	wire [16-1:0] node18348;
	wire [16-1:0] node18351;
	wire [16-1:0] node18354;
	wire [16-1:0] node18355;
	wire [16-1:0] node18356;
	wire [16-1:0] node18359;
	wire [16-1:0] node18362;
	wire [16-1:0] node18363;
	wire [16-1:0] node18366;
	wire [16-1:0] node18369;
	wire [16-1:0] node18370;
	wire [16-1:0] node18371;
	wire [16-1:0] node18372;
	wire [16-1:0] node18373;
	wire [16-1:0] node18374;
	wire [16-1:0] node18377;
	wire [16-1:0] node18380;
	wire [16-1:0] node18381;
	wire [16-1:0] node18384;
	wire [16-1:0] node18387;
	wire [16-1:0] node18388;
	wire [16-1:0] node18389;
	wire [16-1:0] node18392;
	wire [16-1:0] node18395;
	wire [16-1:0] node18396;
	wire [16-1:0] node18399;
	wire [16-1:0] node18402;
	wire [16-1:0] node18403;
	wire [16-1:0] node18404;
	wire [16-1:0] node18405;
	wire [16-1:0] node18408;
	wire [16-1:0] node18411;
	wire [16-1:0] node18412;
	wire [16-1:0] node18415;
	wire [16-1:0] node18418;
	wire [16-1:0] node18419;
	wire [16-1:0] node18420;
	wire [16-1:0] node18423;
	wire [16-1:0] node18426;
	wire [16-1:0] node18427;
	wire [16-1:0] node18430;
	wire [16-1:0] node18433;
	wire [16-1:0] node18434;
	wire [16-1:0] node18435;
	wire [16-1:0] node18436;
	wire [16-1:0] node18437;
	wire [16-1:0] node18440;
	wire [16-1:0] node18443;
	wire [16-1:0] node18444;
	wire [16-1:0] node18447;
	wire [16-1:0] node18450;
	wire [16-1:0] node18451;
	wire [16-1:0] node18452;
	wire [16-1:0] node18455;
	wire [16-1:0] node18458;
	wire [16-1:0] node18459;
	wire [16-1:0] node18462;
	wire [16-1:0] node18465;
	wire [16-1:0] node18466;
	wire [16-1:0] node18467;
	wire [16-1:0] node18469;
	wire [16-1:0] node18472;
	wire [16-1:0] node18473;
	wire [16-1:0] node18476;
	wire [16-1:0] node18479;
	wire [16-1:0] node18480;
	wire [16-1:0] node18481;
	wire [16-1:0] node18484;
	wire [16-1:0] node18487;
	wire [16-1:0] node18488;
	wire [16-1:0] node18491;
	wire [16-1:0] node18494;
	wire [16-1:0] node18495;
	wire [16-1:0] node18496;
	wire [16-1:0] node18497;
	wire [16-1:0] node18498;
	wire [16-1:0] node18499;
	wire [16-1:0] node18500;
	wire [16-1:0] node18501;
	wire [16-1:0] node18502;
	wire [16-1:0] node18505;
	wire [16-1:0] node18508;
	wire [16-1:0] node18509;
	wire [16-1:0] node18512;
	wire [16-1:0] node18515;
	wire [16-1:0] node18516;
	wire [16-1:0] node18517;
	wire [16-1:0] node18520;
	wire [16-1:0] node18523;
	wire [16-1:0] node18524;
	wire [16-1:0] node18527;
	wire [16-1:0] node18530;
	wire [16-1:0] node18531;
	wire [16-1:0] node18532;
	wire [16-1:0] node18533;
	wire [16-1:0] node18536;
	wire [16-1:0] node18539;
	wire [16-1:0] node18540;
	wire [16-1:0] node18543;
	wire [16-1:0] node18546;
	wire [16-1:0] node18547;
	wire [16-1:0] node18548;
	wire [16-1:0] node18551;
	wire [16-1:0] node18554;
	wire [16-1:0] node18555;
	wire [16-1:0] node18559;
	wire [16-1:0] node18560;
	wire [16-1:0] node18561;
	wire [16-1:0] node18562;
	wire [16-1:0] node18563;
	wire [16-1:0] node18566;
	wire [16-1:0] node18569;
	wire [16-1:0] node18570;
	wire [16-1:0] node18573;
	wire [16-1:0] node18576;
	wire [16-1:0] node18577;
	wire [16-1:0] node18578;
	wire [16-1:0] node18581;
	wire [16-1:0] node18584;
	wire [16-1:0] node18585;
	wire [16-1:0] node18588;
	wire [16-1:0] node18591;
	wire [16-1:0] node18592;
	wire [16-1:0] node18593;
	wire [16-1:0] node18594;
	wire [16-1:0] node18597;
	wire [16-1:0] node18600;
	wire [16-1:0] node18601;
	wire [16-1:0] node18604;
	wire [16-1:0] node18607;
	wire [16-1:0] node18608;
	wire [16-1:0] node18609;
	wire [16-1:0] node18612;
	wire [16-1:0] node18615;
	wire [16-1:0] node18616;
	wire [16-1:0] node18619;
	wire [16-1:0] node18622;
	wire [16-1:0] node18623;
	wire [16-1:0] node18624;
	wire [16-1:0] node18625;
	wire [16-1:0] node18626;
	wire [16-1:0] node18628;
	wire [16-1:0] node18631;
	wire [16-1:0] node18632;
	wire [16-1:0] node18635;
	wire [16-1:0] node18638;
	wire [16-1:0] node18639;
	wire [16-1:0] node18640;
	wire [16-1:0] node18643;
	wire [16-1:0] node18646;
	wire [16-1:0] node18647;
	wire [16-1:0] node18650;
	wire [16-1:0] node18653;
	wire [16-1:0] node18654;
	wire [16-1:0] node18655;
	wire [16-1:0] node18656;
	wire [16-1:0] node18659;
	wire [16-1:0] node18662;
	wire [16-1:0] node18663;
	wire [16-1:0] node18666;
	wire [16-1:0] node18669;
	wire [16-1:0] node18670;
	wire [16-1:0] node18671;
	wire [16-1:0] node18674;
	wire [16-1:0] node18677;
	wire [16-1:0] node18678;
	wire [16-1:0] node18682;
	wire [16-1:0] node18683;
	wire [16-1:0] node18684;
	wire [16-1:0] node18685;
	wire [16-1:0] node18686;
	wire [16-1:0] node18689;
	wire [16-1:0] node18692;
	wire [16-1:0] node18693;
	wire [16-1:0] node18696;
	wire [16-1:0] node18699;
	wire [16-1:0] node18700;
	wire [16-1:0] node18702;
	wire [16-1:0] node18705;
	wire [16-1:0] node18707;
	wire [16-1:0] node18710;
	wire [16-1:0] node18711;
	wire [16-1:0] node18712;
	wire [16-1:0] node18713;
	wire [16-1:0] node18716;
	wire [16-1:0] node18719;
	wire [16-1:0] node18720;
	wire [16-1:0] node18723;
	wire [16-1:0] node18726;
	wire [16-1:0] node18727;
	wire [16-1:0] node18728;
	wire [16-1:0] node18731;
	wire [16-1:0] node18734;
	wire [16-1:0] node18735;
	wire [16-1:0] node18738;
	wire [16-1:0] node18741;
	wire [16-1:0] node18742;
	wire [16-1:0] node18743;
	wire [16-1:0] node18744;
	wire [16-1:0] node18745;
	wire [16-1:0] node18746;
	wire [16-1:0] node18747;
	wire [16-1:0] node18750;
	wire [16-1:0] node18753;
	wire [16-1:0] node18754;
	wire [16-1:0] node18757;
	wire [16-1:0] node18760;
	wire [16-1:0] node18761;
	wire [16-1:0] node18762;
	wire [16-1:0] node18765;
	wire [16-1:0] node18768;
	wire [16-1:0] node18769;
	wire [16-1:0] node18772;
	wire [16-1:0] node18775;
	wire [16-1:0] node18776;
	wire [16-1:0] node18777;
	wire [16-1:0] node18778;
	wire [16-1:0] node18781;
	wire [16-1:0] node18784;
	wire [16-1:0] node18785;
	wire [16-1:0] node18788;
	wire [16-1:0] node18791;
	wire [16-1:0] node18792;
	wire [16-1:0] node18793;
	wire [16-1:0] node18796;
	wire [16-1:0] node18799;
	wire [16-1:0] node18800;
	wire [16-1:0] node18803;
	wire [16-1:0] node18806;
	wire [16-1:0] node18807;
	wire [16-1:0] node18808;
	wire [16-1:0] node18809;
	wire [16-1:0] node18810;
	wire [16-1:0] node18813;
	wire [16-1:0] node18816;
	wire [16-1:0] node18817;
	wire [16-1:0] node18820;
	wire [16-1:0] node18823;
	wire [16-1:0] node18824;
	wire [16-1:0] node18826;
	wire [16-1:0] node18829;
	wire [16-1:0] node18830;
	wire [16-1:0] node18833;
	wire [16-1:0] node18836;
	wire [16-1:0] node18837;
	wire [16-1:0] node18838;
	wire [16-1:0] node18839;
	wire [16-1:0] node18842;
	wire [16-1:0] node18845;
	wire [16-1:0] node18846;
	wire [16-1:0] node18849;
	wire [16-1:0] node18852;
	wire [16-1:0] node18853;
	wire [16-1:0] node18854;
	wire [16-1:0] node18857;
	wire [16-1:0] node18860;
	wire [16-1:0] node18861;
	wire [16-1:0] node18864;
	wire [16-1:0] node18867;
	wire [16-1:0] node18868;
	wire [16-1:0] node18869;
	wire [16-1:0] node18870;
	wire [16-1:0] node18871;
	wire [16-1:0] node18872;
	wire [16-1:0] node18875;
	wire [16-1:0] node18878;
	wire [16-1:0] node18879;
	wire [16-1:0] node18882;
	wire [16-1:0] node18885;
	wire [16-1:0] node18886;
	wire [16-1:0] node18887;
	wire [16-1:0] node18890;
	wire [16-1:0] node18893;
	wire [16-1:0] node18894;
	wire [16-1:0] node18898;
	wire [16-1:0] node18899;
	wire [16-1:0] node18900;
	wire [16-1:0] node18901;
	wire [16-1:0] node18904;
	wire [16-1:0] node18907;
	wire [16-1:0] node18908;
	wire [16-1:0] node18911;
	wire [16-1:0] node18914;
	wire [16-1:0] node18915;
	wire [16-1:0] node18916;
	wire [16-1:0] node18919;
	wire [16-1:0] node18922;
	wire [16-1:0] node18924;
	wire [16-1:0] node18927;
	wire [16-1:0] node18928;
	wire [16-1:0] node18929;
	wire [16-1:0] node18930;
	wire [16-1:0] node18931;
	wire [16-1:0] node18934;
	wire [16-1:0] node18937;
	wire [16-1:0] node18938;
	wire [16-1:0] node18941;
	wire [16-1:0] node18944;
	wire [16-1:0] node18945;
	wire [16-1:0] node18946;
	wire [16-1:0] node18949;
	wire [16-1:0] node18952;
	wire [16-1:0] node18954;
	wire [16-1:0] node18957;
	wire [16-1:0] node18958;
	wire [16-1:0] node18959;
	wire [16-1:0] node18960;
	wire [16-1:0] node18963;
	wire [16-1:0] node18966;
	wire [16-1:0] node18967;
	wire [16-1:0] node18970;
	wire [16-1:0] node18973;
	wire [16-1:0] node18974;
	wire [16-1:0] node18975;
	wire [16-1:0] node18978;
	wire [16-1:0] node18981;
	wire [16-1:0] node18982;
	wire [16-1:0] node18985;
	wire [16-1:0] node18988;
	wire [16-1:0] node18989;
	wire [16-1:0] node18990;
	wire [16-1:0] node18991;
	wire [16-1:0] node18992;
	wire [16-1:0] node18993;
	wire [16-1:0] node18994;
	wire [16-1:0] node18995;
	wire [16-1:0] node18998;
	wire [16-1:0] node19001;
	wire [16-1:0] node19002;
	wire [16-1:0] node19005;
	wire [16-1:0] node19008;
	wire [16-1:0] node19009;
	wire [16-1:0] node19010;
	wire [16-1:0] node19013;
	wire [16-1:0] node19016;
	wire [16-1:0] node19017;
	wire [16-1:0] node19020;
	wire [16-1:0] node19023;
	wire [16-1:0] node19024;
	wire [16-1:0] node19025;
	wire [16-1:0] node19026;
	wire [16-1:0] node19029;
	wire [16-1:0] node19032;
	wire [16-1:0] node19033;
	wire [16-1:0] node19036;
	wire [16-1:0] node19039;
	wire [16-1:0] node19040;
	wire [16-1:0] node19041;
	wire [16-1:0] node19044;
	wire [16-1:0] node19047;
	wire [16-1:0] node19048;
	wire [16-1:0] node19051;
	wire [16-1:0] node19054;
	wire [16-1:0] node19055;
	wire [16-1:0] node19056;
	wire [16-1:0] node19057;
	wire [16-1:0] node19058;
	wire [16-1:0] node19061;
	wire [16-1:0] node19064;
	wire [16-1:0] node19065;
	wire [16-1:0] node19069;
	wire [16-1:0] node19070;
	wire [16-1:0] node19071;
	wire [16-1:0] node19074;
	wire [16-1:0] node19077;
	wire [16-1:0] node19078;
	wire [16-1:0] node19081;
	wire [16-1:0] node19084;
	wire [16-1:0] node19085;
	wire [16-1:0] node19086;
	wire [16-1:0] node19088;
	wire [16-1:0] node19091;
	wire [16-1:0] node19092;
	wire [16-1:0] node19095;
	wire [16-1:0] node19098;
	wire [16-1:0] node19099;
	wire [16-1:0] node19100;
	wire [16-1:0] node19103;
	wire [16-1:0] node19106;
	wire [16-1:0] node19107;
	wire [16-1:0] node19110;
	wire [16-1:0] node19113;
	wire [16-1:0] node19114;
	wire [16-1:0] node19115;
	wire [16-1:0] node19116;
	wire [16-1:0] node19117;
	wire [16-1:0] node19118;
	wire [16-1:0] node19121;
	wire [16-1:0] node19124;
	wire [16-1:0] node19125;
	wire [16-1:0] node19128;
	wire [16-1:0] node19131;
	wire [16-1:0] node19132;
	wire [16-1:0] node19133;
	wire [16-1:0] node19136;
	wire [16-1:0] node19139;
	wire [16-1:0] node19140;
	wire [16-1:0] node19143;
	wire [16-1:0] node19146;
	wire [16-1:0] node19147;
	wire [16-1:0] node19148;
	wire [16-1:0] node19149;
	wire [16-1:0] node19152;
	wire [16-1:0] node19155;
	wire [16-1:0] node19156;
	wire [16-1:0] node19159;
	wire [16-1:0] node19162;
	wire [16-1:0] node19163;
	wire [16-1:0] node19164;
	wire [16-1:0] node19167;
	wire [16-1:0] node19170;
	wire [16-1:0] node19171;
	wire [16-1:0] node19174;
	wire [16-1:0] node19177;
	wire [16-1:0] node19178;
	wire [16-1:0] node19179;
	wire [16-1:0] node19180;
	wire [16-1:0] node19181;
	wire [16-1:0] node19184;
	wire [16-1:0] node19187;
	wire [16-1:0] node19188;
	wire [16-1:0] node19191;
	wire [16-1:0] node19194;
	wire [16-1:0] node19195;
	wire [16-1:0] node19197;
	wire [16-1:0] node19200;
	wire [16-1:0] node19201;
	wire [16-1:0] node19204;
	wire [16-1:0] node19207;
	wire [16-1:0] node19208;
	wire [16-1:0] node19209;
	wire [16-1:0] node19210;
	wire [16-1:0] node19213;
	wire [16-1:0] node19216;
	wire [16-1:0] node19217;
	wire [16-1:0] node19220;
	wire [16-1:0] node19223;
	wire [16-1:0] node19224;
	wire [16-1:0] node19225;
	wire [16-1:0] node19228;
	wire [16-1:0] node19231;
	wire [16-1:0] node19233;
	wire [16-1:0] node19236;
	wire [16-1:0] node19237;
	wire [16-1:0] node19238;
	wire [16-1:0] node19239;
	wire [16-1:0] node19240;
	wire [16-1:0] node19241;
	wire [16-1:0] node19242;
	wire [16-1:0] node19245;
	wire [16-1:0] node19248;
	wire [16-1:0] node19249;
	wire [16-1:0] node19252;
	wire [16-1:0] node19255;
	wire [16-1:0] node19256;
	wire [16-1:0] node19257;
	wire [16-1:0] node19260;
	wire [16-1:0] node19263;
	wire [16-1:0] node19264;
	wire [16-1:0] node19267;
	wire [16-1:0] node19270;
	wire [16-1:0] node19271;
	wire [16-1:0] node19272;
	wire [16-1:0] node19273;
	wire [16-1:0] node19276;
	wire [16-1:0] node19279;
	wire [16-1:0] node19280;
	wire [16-1:0] node19283;
	wire [16-1:0] node19286;
	wire [16-1:0] node19287;
	wire [16-1:0] node19288;
	wire [16-1:0] node19292;
	wire [16-1:0] node19293;
	wire [16-1:0] node19296;
	wire [16-1:0] node19299;
	wire [16-1:0] node19300;
	wire [16-1:0] node19301;
	wire [16-1:0] node19302;
	wire [16-1:0] node19303;
	wire [16-1:0] node19306;
	wire [16-1:0] node19309;
	wire [16-1:0] node19310;
	wire [16-1:0] node19313;
	wire [16-1:0] node19316;
	wire [16-1:0] node19317;
	wire [16-1:0] node19318;
	wire [16-1:0] node19321;
	wire [16-1:0] node19324;
	wire [16-1:0] node19325;
	wire [16-1:0] node19328;
	wire [16-1:0] node19331;
	wire [16-1:0] node19332;
	wire [16-1:0] node19333;
	wire [16-1:0] node19334;
	wire [16-1:0] node19338;
	wire [16-1:0] node19339;
	wire [16-1:0] node19342;
	wire [16-1:0] node19345;
	wire [16-1:0] node19346;
	wire [16-1:0] node19348;
	wire [16-1:0] node19351;
	wire [16-1:0] node19352;
	wire [16-1:0] node19355;
	wire [16-1:0] node19358;
	wire [16-1:0] node19359;
	wire [16-1:0] node19360;
	wire [16-1:0] node19361;
	wire [16-1:0] node19362;
	wire [16-1:0] node19363;
	wire [16-1:0] node19367;
	wire [16-1:0] node19368;
	wire [16-1:0] node19371;
	wire [16-1:0] node19374;
	wire [16-1:0] node19375;
	wire [16-1:0] node19376;
	wire [16-1:0] node19379;
	wire [16-1:0] node19382;
	wire [16-1:0] node19383;
	wire [16-1:0] node19387;
	wire [16-1:0] node19388;
	wire [16-1:0] node19389;
	wire [16-1:0] node19390;
	wire [16-1:0] node19393;
	wire [16-1:0] node19396;
	wire [16-1:0] node19397;
	wire [16-1:0] node19400;
	wire [16-1:0] node19403;
	wire [16-1:0] node19404;
	wire [16-1:0] node19405;
	wire [16-1:0] node19408;
	wire [16-1:0] node19411;
	wire [16-1:0] node19412;
	wire [16-1:0] node19415;
	wire [16-1:0] node19418;
	wire [16-1:0] node19419;
	wire [16-1:0] node19420;
	wire [16-1:0] node19421;
	wire [16-1:0] node19422;
	wire [16-1:0] node19425;
	wire [16-1:0] node19428;
	wire [16-1:0] node19429;
	wire [16-1:0] node19432;
	wire [16-1:0] node19435;
	wire [16-1:0] node19436;
	wire [16-1:0] node19438;
	wire [16-1:0] node19441;
	wire [16-1:0] node19442;
	wire [16-1:0] node19445;
	wire [16-1:0] node19448;
	wire [16-1:0] node19449;
	wire [16-1:0] node19450;
	wire [16-1:0] node19451;
	wire [16-1:0] node19454;
	wire [16-1:0] node19457;
	wire [16-1:0] node19458;
	wire [16-1:0] node19461;
	wire [16-1:0] node19464;
	wire [16-1:0] node19465;
	wire [16-1:0] node19466;
	wire [16-1:0] node19469;
	wire [16-1:0] node19472;
	wire [16-1:0] node19473;
	wire [16-1:0] node19476;
	wire [16-1:0] node19479;
	wire [16-1:0] node19480;
	wire [16-1:0] node19481;
	wire [16-1:0] node19482;
	wire [16-1:0] node19483;
	wire [16-1:0] node19484;
	wire [16-1:0] node19485;
	wire [16-1:0] node19486;
	wire [16-1:0] node19487;
	wire [16-1:0] node19488;
	wire [16-1:0] node19489;
	wire [16-1:0] node19492;
	wire [16-1:0] node19495;
	wire [16-1:0] node19496;
	wire [16-1:0] node19499;
	wire [16-1:0] node19502;
	wire [16-1:0] node19503;
	wire [16-1:0] node19504;
	wire [16-1:0] node19507;
	wire [16-1:0] node19510;
	wire [16-1:0] node19511;
	wire [16-1:0] node19515;
	wire [16-1:0] node19516;
	wire [16-1:0] node19517;
	wire [16-1:0] node19518;
	wire [16-1:0] node19522;
	wire [16-1:0] node19523;
	wire [16-1:0] node19526;
	wire [16-1:0] node19529;
	wire [16-1:0] node19530;
	wire [16-1:0] node19531;
	wire [16-1:0] node19534;
	wire [16-1:0] node19537;
	wire [16-1:0] node19538;
	wire [16-1:0] node19541;
	wire [16-1:0] node19544;
	wire [16-1:0] node19545;
	wire [16-1:0] node19546;
	wire [16-1:0] node19547;
	wire [16-1:0] node19548;
	wire [16-1:0] node19551;
	wire [16-1:0] node19554;
	wire [16-1:0] node19556;
	wire [16-1:0] node19559;
	wire [16-1:0] node19560;
	wire [16-1:0] node19561;
	wire [16-1:0] node19564;
	wire [16-1:0] node19567;
	wire [16-1:0] node19568;
	wire [16-1:0] node19571;
	wire [16-1:0] node19574;
	wire [16-1:0] node19575;
	wire [16-1:0] node19576;
	wire [16-1:0] node19577;
	wire [16-1:0] node19580;
	wire [16-1:0] node19583;
	wire [16-1:0] node19584;
	wire [16-1:0] node19587;
	wire [16-1:0] node19590;
	wire [16-1:0] node19591;
	wire [16-1:0] node19592;
	wire [16-1:0] node19595;
	wire [16-1:0] node19598;
	wire [16-1:0] node19599;
	wire [16-1:0] node19602;
	wire [16-1:0] node19605;
	wire [16-1:0] node19606;
	wire [16-1:0] node19607;
	wire [16-1:0] node19608;
	wire [16-1:0] node19609;
	wire [16-1:0] node19610;
	wire [16-1:0] node19613;
	wire [16-1:0] node19616;
	wire [16-1:0] node19617;
	wire [16-1:0] node19620;
	wire [16-1:0] node19623;
	wire [16-1:0] node19624;
	wire [16-1:0] node19625;
	wire [16-1:0] node19628;
	wire [16-1:0] node19631;
	wire [16-1:0] node19632;
	wire [16-1:0] node19636;
	wire [16-1:0] node19637;
	wire [16-1:0] node19638;
	wire [16-1:0] node19639;
	wire [16-1:0] node19642;
	wire [16-1:0] node19645;
	wire [16-1:0] node19646;
	wire [16-1:0] node19649;
	wire [16-1:0] node19652;
	wire [16-1:0] node19653;
	wire [16-1:0] node19654;
	wire [16-1:0] node19657;
	wire [16-1:0] node19660;
	wire [16-1:0] node19661;
	wire [16-1:0] node19664;
	wire [16-1:0] node19667;
	wire [16-1:0] node19668;
	wire [16-1:0] node19669;
	wire [16-1:0] node19670;
	wire [16-1:0] node19671;
	wire [16-1:0] node19674;
	wire [16-1:0] node19677;
	wire [16-1:0] node19678;
	wire [16-1:0] node19681;
	wire [16-1:0] node19684;
	wire [16-1:0] node19685;
	wire [16-1:0] node19686;
	wire [16-1:0] node19689;
	wire [16-1:0] node19692;
	wire [16-1:0] node19693;
	wire [16-1:0] node19696;
	wire [16-1:0] node19699;
	wire [16-1:0] node19700;
	wire [16-1:0] node19701;
	wire [16-1:0] node19702;
	wire [16-1:0] node19705;
	wire [16-1:0] node19708;
	wire [16-1:0] node19709;
	wire [16-1:0] node19712;
	wire [16-1:0] node19715;
	wire [16-1:0] node19716;
	wire [16-1:0] node19717;
	wire [16-1:0] node19720;
	wire [16-1:0] node19723;
	wire [16-1:0] node19724;
	wire [16-1:0] node19727;
	wire [16-1:0] node19730;
	wire [16-1:0] node19731;
	wire [16-1:0] node19732;
	wire [16-1:0] node19733;
	wire [16-1:0] node19734;
	wire [16-1:0] node19735;
	wire [16-1:0] node19736;
	wire [16-1:0] node19739;
	wire [16-1:0] node19742;
	wire [16-1:0] node19743;
	wire [16-1:0] node19747;
	wire [16-1:0] node19748;
	wire [16-1:0] node19749;
	wire [16-1:0] node19752;
	wire [16-1:0] node19755;
	wire [16-1:0] node19756;
	wire [16-1:0] node19759;
	wire [16-1:0] node19762;
	wire [16-1:0] node19763;
	wire [16-1:0] node19764;
	wire [16-1:0] node19765;
	wire [16-1:0] node19768;
	wire [16-1:0] node19771;
	wire [16-1:0] node19772;
	wire [16-1:0] node19775;
	wire [16-1:0] node19778;
	wire [16-1:0] node19779;
	wire [16-1:0] node19780;
	wire [16-1:0] node19783;
	wire [16-1:0] node19786;
	wire [16-1:0] node19787;
	wire [16-1:0] node19790;
	wire [16-1:0] node19793;
	wire [16-1:0] node19794;
	wire [16-1:0] node19795;
	wire [16-1:0] node19796;
	wire [16-1:0] node19797;
	wire [16-1:0] node19800;
	wire [16-1:0] node19803;
	wire [16-1:0] node19804;
	wire [16-1:0] node19807;
	wire [16-1:0] node19810;
	wire [16-1:0] node19811;
	wire [16-1:0] node19812;
	wire [16-1:0] node19815;
	wire [16-1:0] node19818;
	wire [16-1:0] node19819;
	wire [16-1:0] node19823;
	wire [16-1:0] node19824;
	wire [16-1:0] node19825;
	wire [16-1:0] node19826;
	wire [16-1:0] node19829;
	wire [16-1:0] node19832;
	wire [16-1:0] node19833;
	wire [16-1:0] node19836;
	wire [16-1:0] node19839;
	wire [16-1:0] node19840;
	wire [16-1:0] node19841;
	wire [16-1:0] node19844;
	wire [16-1:0] node19847;
	wire [16-1:0] node19848;
	wire [16-1:0] node19851;
	wire [16-1:0] node19854;
	wire [16-1:0] node19855;
	wire [16-1:0] node19856;
	wire [16-1:0] node19857;
	wire [16-1:0] node19858;
	wire [16-1:0] node19859;
	wire [16-1:0] node19862;
	wire [16-1:0] node19865;
	wire [16-1:0] node19866;
	wire [16-1:0] node19869;
	wire [16-1:0] node19872;
	wire [16-1:0] node19873;
	wire [16-1:0] node19876;
	wire [16-1:0] node19877;
	wire [16-1:0] node19880;
	wire [16-1:0] node19883;
	wire [16-1:0] node19884;
	wire [16-1:0] node19885;
	wire [16-1:0] node19886;
	wire [16-1:0] node19889;
	wire [16-1:0] node19892;
	wire [16-1:0] node19893;
	wire [16-1:0] node19897;
	wire [16-1:0] node19898;
	wire [16-1:0] node19899;
	wire [16-1:0] node19903;
	wire [16-1:0] node19904;
	wire [16-1:0] node19907;
	wire [16-1:0] node19910;
	wire [16-1:0] node19911;
	wire [16-1:0] node19912;
	wire [16-1:0] node19913;
	wire [16-1:0] node19914;
	wire [16-1:0] node19917;
	wire [16-1:0] node19920;
	wire [16-1:0] node19921;
	wire [16-1:0] node19924;
	wire [16-1:0] node19927;
	wire [16-1:0] node19928;
	wire [16-1:0] node19929;
	wire [16-1:0] node19932;
	wire [16-1:0] node19935;
	wire [16-1:0] node19936;
	wire [16-1:0] node19939;
	wire [16-1:0] node19942;
	wire [16-1:0] node19943;
	wire [16-1:0] node19944;
	wire [16-1:0] node19945;
	wire [16-1:0] node19948;
	wire [16-1:0] node19951;
	wire [16-1:0] node19952;
	wire [16-1:0] node19955;
	wire [16-1:0] node19958;
	wire [16-1:0] node19959;
	wire [16-1:0] node19960;
	wire [16-1:0] node19963;
	wire [16-1:0] node19966;
	wire [16-1:0] node19967;
	wire [16-1:0] node19970;
	wire [16-1:0] node19973;
	wire [16-1:0] node19974;
	wire [16-1:0] node19975;
	wire [16-1:0] node19976;
	wire [16-1:0] node19977;
	wire [16-1:0] node19978;
	wire [16-1:0] node19979;
	wire [16-1:0] node19980;
	wire [16-1:0] node19983;
	wire [16-1:0] node19986;
	wire [16-1:0] node19987;
	wire [16-1:0] node19990;
	wire [16-1:0] node19993;
	wire [16-1:0] node19994;
	wire [16-1:0] node19995;
	wire [16-1:0] node19998;
	wire [16-1:0] node20001;
	wire [16-1:0] node20002;
	wire [16-1:0] node20005;
	wire [16-1:0] node20008;
	wire [16-1:0] node20009;
	wire [16-1:0] node20010;
	wire [16-1:0] node20011;
	wire [16-1:0] node20014;
	wire [16-1:0] node20017;
	wire [16-1:0] node20018;
	wire [16-1:0] node20021;
	wire [16-1:0] node20024;
	wire [16-1:0] node20025;
	wire [16-1:0] node20026;
	wire [16-1:0] node20030;
	wire [16-1:0] node20031;
	wire [16-1:0] node20034;
	wire [16-1:0] node20037;
	wire [16-1:0] node20038;
	wire [16-1:0] node20039;
	wire [16-1:0] node20040;
	wire [16-1:0] node20041;
	wire [16-1:0] node20044;
	wire [16-1:0] node20047;
	wire [16-1:0] node20048;
	wire [16-1:0] node20051;
	wire [16-1:0] node20054;
	wire [16-1:0] node20055;
	wire [16-1:0] node20056;
	wire [16-1:0] node20059;
	wire [16-1:0] node20062;
	wire [16-1:0] node20064;
	wire [16-1:0] node20067;
	wire [16-1:0] node20068;
	wire [16-1:0] node20069;
	wire [16-1:0] node20070;
	wire [16-1:0] node20073;
	wire [16-1:0] node20076;
	wire [16-1:0] node20077;
	wire [16-1:0] node20080;
	wire [16-1:0] node20083;
	wire [16-1:0] node20084;
	wire [16-1:0] node20085;
	wire [16-1:0] node20088;
	wire [16-1:0] node20091;
	wire [16-1:0] node20092;
	wire [16-1:0] node20095;
	wire [16-1:0] node20098;
	wire [16-1:0] node20099;
	wire [16-1:0] node20100;
	wire [16-1:0] node20101;
	wire [16-1:0] node20102;
	wire [16-1:0] node20103;
	wire [16-1:0] node20106;
	wire [16-1:0] node20109;
	wire [16-1:0] node20110;
	wire [16-1:0] node20113;
	wire [16-1:0] node20116;
	wire [16-1:0] node20117;
	wire [16-1:0] node20118;
	wire [16-1:0] node20121;
	wire [16-1:0] node20124;
	wire [16-1:0] node20125;
	wire [16-1:0] node20129;
	wire [16-1:0] node20130;
	wire [16-1:0] node20131;
	wire [16-1:0] node20132;
	wire [16-1:0] node20136;
	wire [16-1:0] node20137;
	wire [16-1:0] node20141;
	wire [16-1:0] node20142;
	wire [16-1:0] node20143;
	wire [16-1:0] node20146;
	wire [16-1:0] node20149;
	wire [16-1:0] node20150;
	wire [16-1:0] node20153;
	wire [16-1:0] node20156;
	wire [16-1:0] node20157;
	wire [16-1:0] node20158;
	wire [16-1:0] node20159;
	wire [16-1:0] node20160;
	wire [16-1:0] node20163;
	wire [16-1:0] node20166;
	wire [16-1:0] node20167;
	wire [16-1:0] node20170;
	wire [16-1:0] node20173;
	wire [16-1:0] node20174;
	wire [16-1:0] node20175;
	wire [16-1:0] node20178;
	wire [16-1:0] node20181;
	wire [16-1:0] node20183;
	wire [16-1:0] node20186;
	wire [16-1:0] node20187;
	wire [16-1:0] node20188;
	wire [16-1:0] node20189;
	wire [16-1:0] node20192;
	wire [16-1:0] node20195;
	wire [16-1:0] node20196;
	wire [16-1:0] node20199;
	wire [16-1:0] node20202;
	wire [16-1:0] node20203;
	wire [16-1:0] node20204;
	wire [16-1:0] node20207;
	wire [16-1:0] node20210;
	wire [16-1:0] node20211;
	wire [16-1:0] node20214;
	wire [16-1:0] node20217;
	wire [16-1:0] node20218;
	wire [16-1:0] node20219;
	wire [16-1:0] node20220;
	wire [16-1:0] node20221;
	wire [16-1:0] node20222;
	wire [16-1:0] node20223;
	wire [16-1:0] node20227;
	wire [16-1:0] node20228;
	wire [16-1:0] node20231;
	wire [16-1:0] node20234;
	wire [16-1:0] node20235;
	wire [16-1:0] node20236;
	wire [16-1:0] node20239;
	wire [16-1:0] node20242;
	wire [16-1:0] node20243;
	wire [16-1:0] node20246;
	wire [16-1:0] node20249;
	wire [16-1:0] node20250;
	wire [16-1:0] node20251;
	wire [16-1:0] node20252;
	wire [16-1:0] node20255;
	wire [16-1:0] node20258;
	wire [16-1:0] node20259;
	wire [16-1:0] node20262;
	wire [16-1:0] node20265;
	wire [16-1:0] node20266;
	wire [16-1:0] node20267;
	wire [16-1:0] node20270;
	wire [16-1:0] node20273;
	wire [16-1:0] node20274;
	wire [16-1:0] node20277;
	wire [16-1:0] node20280;
	wire [16-1:0] node20281;
	wire [16-1:0] node20282;
	wire [16-1:0] node20283;
	wire [16-1:0] node20284;
	wire [16-1:0] node20287;
	wire [16-1:0] node20290;
	wire [16-1:0] node20291;
	wire [16-1:0] node20294;
	wire [16-1:0] node20297;
	wire [16-1:0] node20298;
	wire [16-1:0] node20299;
	wire [16-1:0] node20302;
	wire [16-1:0] node20305;
	wire [16-1:0] node20306;
	wire [16-1:0] node20309;
	wire [16-1:0] node20312;
	wire [16-1:0] node20313;
	wire [16-1:0] node20314;
	wire [16-1:0] node20315;
	wire [16-1:0] node20318;
	wire [16-1:0] node20321;
	wire [16-1:0] node20322;
	wire [16-1:0] node20325;
	wire [16-1:0] node20328;
	wire [16-1:0] node20329;
	wire [16-1:0] node20330;
	wire [16-1:0] node20333;
	wire [16-1:0] node20336;
	wire [16-1:0] node20337;
	wire [16-1:0] node20340;
	wire [16-1:0] node20343;
	wire [16-1:0] node20344;
	wire [16-1:0] node20345;
	wire [16-1:0] node20346;
	wire [16-1:0] node20347;
	wire [16-1:0] node20348;
	wire [16-1:0] node20351;
	wire [16-1:0] node20354;
	wire [16-1:0] node20355;
	wire [16-1:0] node20358;
	wire [16-1:0] node20361;
	wire [16-1:0] node20362;
	wire [16-1:0] node20363;
	wire [16-1:0] node20366;
	wire [16-1:0] node20369;
	wire [16-1:0] node20370;
	wire [16-1:0] node20373;
	wire [16-1:0] node20376;
	wire [16-1:0] node20377;
	wire [16-1:0] node20378;
	wire [16-1:0] node20379;
	wire [16-1:0] node20382;
	wire [16-1:0] node20385;
	wire [16-1:0] node20386;
	wire [16-1:0] node20389;
	wire [16-1:0] node20392;
	wire [16-1:0] node20393;
	wire [16-1:0] node20394;
	wire [16-1:0] node20397;
	wire [16-1:0] node20400;
	wire [16-1:0] node20401;
	wire [16-1:0] node20404;
	wire [16-1:0] node20407;
	wire [16-1:0] node20408;
	wire [16-1:0] node20409;
	wire [16-1:0] node20410;
	wire [16-1:0] node20411;
	wire [16-1:0] node20414;
	wire [16-1:0] node20418;
	wire [16-1:0] node20419;
	wire [16-1:0] node20420;
	wire [16-1:0] node20423;
	wire [16-1:0] node20426;
	wire [16-1:0] node20427;
	wire [16-1:0] node20430;
	wire [16-1:0] node20433;
	wire [16-1:0] node20434;
	wire [16-1:0] node20435;
	wire [16-1:0] node20436;
	wire [16-1:0] node20439;
	wire [16-1:0] node20442;
	wire [16-1:0] node20443;
	wire [16-1:0] node20446;
	wire [16-1:0] node20449;
	wire [16-1:0] node20450;
	wire [16-1:0] node20451;
	wire [16-1:0] node20454;
	wire [16-1:0] node20457;
	wire [16-1:0] node20459;
	wire [16-1:0] node20462;
	wire [16-1:0] node20463;
	wire [16-1:0] node20464;
	wire [16-1:0] node20465;
	wire [16-1:0] node20466;
	wire [16-1:0] node20467;
	wire [16-1:0] node20468;
	wire [16-1:0] node20469;
	wire [16-1:0] node20470;
	wire [16-1:0] node20473;
	wire [16-1:0] node20476;
	wire [16-1:0] node20477;
	wire [16-1:0] node20480;
	wire [16-1:0] node20483;
	wire [16-1:0] node20484;
	wire [16-1:0] node20485;
	wire [16-1:0] node20488;
	wire [16-1:0] node20491;
	wire [16-1:0] node20492;
	wire [16-1:0] node20495;
	wire [16-1:0] node20498;
	wire [16-1:0] node20499;
	wire [16-1:0] node20500;
	wire [16-1:0] node20501;
	wire [16-1:0] node20504;
	wire [16-1:0] node20507;
	wire [16-1:0] node20508;
	wire [16-1:0] node20511;
	wire [16-1:0] node20514;
	wire [16-1:0] node20515;
	wire [16-1:0] node20516;
	wire [16-1:0] node20519;
	wire [16-1:0] node20522;
	wire [16-1:0] node20523;
	wire [16-1:0] node20527;
	wire [16-1:0] node20528;
	wire [16-1:0] node20529;
	wire [16-1:0] node20530;
	wire [16-1:0] node20531;
	wire [16-1:0] node20534;
	wire [16-1:0] node20537;
	wire [16-1:0] node20538;
	wire [16-1:0] node20541;
	wire [16-1:0] node20544;
	wire [16-1:0] node20545;
	wire [16-1:0] node20546;
	wire [16-1:0] node20549;
	wire [16-1:0] node20552;
	wire [16-1:0] node20553;
	wire [16-1:0] node20556;
	wire [16-1:0] node20559;
	wire [16-1:0] node20560;
	wire [16-1:0] node20561;
	wire [16-1:0] node20562;
	wire [16-1:0] node20566;
	wire [16-1:0] node20567;
	wire [16-1:0] node20570;
	wire [16-1:0] node20573;
	wire [16-1:0] node20574;
	wire [16-1:0] node20575;
	wire [16-1:0] node20578;
	wire [16-1:0] node20581;
	wire [16-1:0] node20582;
	wire [16-1:0] node20585;
	wire [16-1:0] node20588;
	wire [16-1:0] node20589;
	wire [16-1:0] node20590;
	wire [16-1:0] node20591;
	wire [16-1:0] node20592;
	wire [16-1:0] node20593;
	wire [16-1:0] node20596;
	wire [16-1:0] node20600;
	wire [16-1:0] node20601;
	wire [16-1:0] node20602;
	wire [16-1:0] node20605;
	wire [16-1:0] node20608;
	wire [16-1:0] node20609;
	wire [16-1:0] node20612;
	wire [16-1:0] node20615;
	wire [16-1:0] node20616;
	wire [16-1:0] node20617;
	wire [16-1:0] node20618;
	wire [16-1:0] node20621;
	wire [16-1:0] node20624;
	wire [16-1:0] node20625;
	wire [16-1:0] node20628;
	wire [16-1:0] node20631;
	wire [16-1:0] node20632;
	wire [16-1:0] node20633;
	wire [16-1:0] node20636;
	wire [16-1:0] node20639;
	wire [16-1:0] node20640;
	wire [16-1:0] node20643;
	wire [16-1:0] node20646;
	wire [16-1:0] node20647;
	wire [16-1:0] node20648;
	wire [16-1:0] node20649;
	wire [16-1:0] node20650;
	wire [16-1:0] node20654;
	wire [16-1:0] node20655;
	wire [16-1:0] node20659;
	wire [16-1:0] node20660;
	wire [16-1:0] node20661;
	wire [16-1:0] node20664;
	wire [16-1:0] node20667;
	wire [16-1:0] node20668;
	wire [16-1:0] node20671;
	wire [16-1:0] node20674;
	wire [16-1:0] node20675;
	wire [16-1:0] node20676;
	wire [16-1:0] node20677;
	wire [16-1:0] node20680;
	wire [16-1:0] node20683;
	wire [16-1:0] node20684;
	wire [16-1:0] node20687;
	wire [16-1:0] node20690;
	wire [16-1:0] node20691;
	wire [16-1:0] node20692;
	wire [16-1:0] node20695;
	wire [16-1:0] node20698;
	wire [16-1:0] node20699;
	wire [16-1:0] node20702;
	wire [16-1:0] node20705;
	wire [16-1:0] node20706;
	wire [16-1:0] node20707;
	wire [16-1:0] node20708;
	wire [16-1:0] node20709;
	wire [16-1:0] node20710;
	wire [16-1:0] node20712;
	wire [16-1:0] node20715;
	wire [16-1:0] node20716;
	wire [16-1:0] node20719;
	wire [16-1:0] node20722;
	wire [16-1:0] node20723;
	wire [16-1:0] node20724;
	wire [16-1:0] node20727;
	wire [16-1:0] node20730;
	wire [16-1:0] node20731;
	wire [16-1:0] node20734;
	wire [16-1:0] node20737;
	wire [16-1:0] node20738;
	wire [16-1:0] node20739;
	wire [16-1:0] node20741;
	wire [16-1:0] node20744;
	wire [16-1:0] node20745;
	wire [16-1:0] node20748;
	wire [16-1:0] node20751;
	wire [16-1:0] node20752;
	wire [16-1:0] node20753;
	wire [16-1:0] node20756;
	wire [16-1:0] node20759;
	wire [16-1:0] node20760;
	wire [16-1:0] node20763;
	wire [16-1:0] node20766;
	wire [16-1:0] node20767;
	wire [16-1:0] node20768;
	wire [16-1:0] node20769;
	wire [16-1:0] node20770;
	wire [16-1:0] node20773;
	wire [16-1:0] node20776;
	wire [16-1:0] node20777;
	wire [16-1:0] node20780;
	wire [16-1:0] node20783;
	wire [16-1:0] node20784;
	wire [16-1:0] node20785;
	wire [16-1:0] node20788;
	wire [16-1:0] node20791;
	wire [16-1:0] node20792;
	wire [16-1:0] node20795;
	wire [16-1:0] node20798;
	wire [16-1:0] node20799;
	wire [16-1:0] node20800;
	wire [16-1:0] node20801;
	wire [16-1:0] node20804;
	wire [16-1:0] node20807;
	wire [16-1:0] node20808;
	wire [16-1:0] node20811;
	wire [16-1:0] node20814;
	wire [16-1:0] node20815;
	wire [16-1:0] node20816;
	wire [16-1:0] node20819;
	wire [16-1:0] node20822;
	wire [16-1:0] node20824;
	wire [16-1:0] node20827;
	wire [16-1:0] node20828;
	wire [16-1:0] node20829;
	wire [16-1:0] node20830;
	wire [16-1:0] node20831;
	wire [16-1:0] node20832;
	wire [16-1:0] node20835;
	wire [16-1:0] node20838;
	wire [16-1:0] node20840;
	wire [16-1:0] node20843;
	wire [16-1:0] node20844;
	wire [16-1:0] node20845;
	wire [16-1:0] node20848;
	wire [16-1:0] node20851;
	wire [16-1:0] node20852;
	wire [16-1:0] node20855;
	wire [16-1:0] node20858;
	wire [16-1:0] node20859;
	wire [16-1:0] node20860;
	wire [16-1:0] node20861;
	wire [16-1:0] node20864;
	wire [16-1:0] node20867;
	wire [16-1:0] node20868;
	wire [16-1:0] node20871;
	wire [16-1:0] node20874;
	wire [16-1:0] node20875;
	wire [16-1:0] node20876;
	wire [16-1:0] node20879;
	wire [16-1:0] node20882;
	wire [16-1:0] node20884;
	wire [16-1:0] node20887;
	wire [16-1:0] node20888;
	wire [16-1:0] node20889;
	wire [16-1:0] node20890;
	wire [16-1:0] node20891;
	wire [16-1:0] node20895;
	wire [16-1:0] node20896;
	wire [16-1:0] node20900;
	wire [16-1:0] node20901;
	wire [16-1:0] node20903;
	wire [16-1:0] node20906;
	wire [16-1:0] node20907;
	wire [16-1:0] node20910;
	wire [16-1:0] node20913;
	wire [16-1:0] node20914;
	wire [16-1:0] node20915;
	wire [16-1:0] node20917;
	wire [16-1:0] node20920;
	wire [16-1:0] node20921;
	wire [16-1:0] node20924;
	wire [16-1:0] node20927;
	wire [16-1:0] node20928;
	wire [16-1:0] node20929;
	wire [16-1:0] node20932;
	wire [16-1:0] node20935;
	wire [16-1:0] node20936;
	wire [16-1:0] node20939;
	wire [16-1:0] node20942;
	wire [16-1:0] node20943;
	wire [16-1:0] node20944;
	wire [16-1:0] node20945;
	wire [16-1:0] node20946;
	wire [16-1:0] node20947;
	wire [16-1:0] node20948;
	wire [16-1:0] node20949;
	wire [16-1:0] node20952;
	wire [16-1:0] node20955;
	wire [16-1:0] node20956;
	wire [16-1:0] node20959;
	wire [16-1:0] node20962;
	wire [16-1:0] node20963;
	wire [16-1:0] node20964;
	wire [16-1:0] node20967;
	wire [16-1:0] node20970;
	wire [16-1:0] node20971;
	wire [16-1:0] node20974;
	wire [16-1:0] node20977;
	wire [16-1:0] node20978;
	wire [16-1:0] node20979;
	wire [16-1:0] node20980;
	wire [16-1:0] node20983;
	wire [16-1:0] node20986;
	wire [16-1:0] node20988;
	wire [16-1:0] node20991;
	wire [16-1:0] node20992;
	wire [16-1:0] node20994;
	wire [16-1:0] node20997;
	wire [16-1:0] node20998;
	wire [16-1:0] node21001;
	wire [16-1:0] node21004;
	wire [16-1:0] node21005;
	wire [16-1:0] node21006;
	wire [16-1:0] node21007;
	wire [16-1:0] node21008;
	wire [16-1:0] node21011;
	wire [16-1:0] node21014;
	wire [16-1:0] node21015;
	wire [16-1:0] node21018;
	wire [16-1:0] node21021;
	wire [16-1:0] node21022;
	wire [16-1:0] node21023;
	wire [16-1:0] node21027;
	wire [16-1:0] node21028;
	wire [16-1:0] node21031;
	wire [16-1:0] node21034;
	wire [16-1:0] node21035;
	wire [16-1:0] node21036;
	wire [16-1:0] node21037;
	wire [16-1:0] node21040;
	wire [16-1:0] node21043;
	wire [16-1:0] node21044;
	wire [16-1:0] node21047;
	wire [16-1:0] node21050;
	wire [16-1:0] node21051;
	wire [16-1:0] node21052;
	wire [16-1:0] node21055;
	wire [16-1:0] node21058;
	wire [16-1:0] node21059;
	wire [16-1:0] node21062;
	wire [16-1:0] node21065;
	wire [16-1:0] node21066;
	wire [16-1:0] node21067;
	wire [16-1:0] node21068;
	wire [16-1:0] node21069;
	wire [16-1:0] node21070;
	wire [16-1:0] node21073;
	wire [16-1:0] node21076;
	wire [16-1:0] node21077;
	wire [16-1:0] node21080;
	wire [16-1:0] node21083;
	wire [16-1:0] node21084;
	wire [16-1:0] node21085;
	wire [16-1:0] node21089;
	wire [16-1:0] node21090;
	wire [16-1:0] node21093;
	wire [16-1:0] node21096;
	wire [16-1:0] node21097;
	wire [16-1:0] node21098;
	wire [16-1:0] node21099;
	wire [16-1:0] node21102;
	wire [16-1:0] node21105;
	wire [16-1:0] node21106;
	wire [16-1:0] node21109;
	wire [16-1:0] node21112;
	wire [16-1:0] node21113;
	wire [16-1:0] node21114;
	wire [16-1:0] node21117;
	wire [16-1:0] node21120;
	wire [16-1:0] node21121;
	wire [16-1:0] node21124;
	wire [16-1:0] node21127;
	wire [16-1:0] node21128;
	wire [16-1:0] node21129;
	wire [16-1:0] node21130;
	wire [16-1:0] node21131;
	wire [16-1:0] node21134;
	wire [16-1:0] node21137;
	wire [16-1:0] node21139;
	wire [16-1:0] node21142;
	wire [16-1:0] node21143;
	wire [16-1:0] node21144;
	wire [16-1:0] node21147;
	wire [16-1:0] node21150;
	wire [16-1:0] node21151;
	wire [16-1:0] node21154;
	wire [16-1:0] node21157;
	wire [16-1:0] node21158;
	wire [16-1:0] node21159;
	wire [16-1:0] node21160;
	wire [16-1:0] node21163;
	wire [16-1:0] node21166;
	wire [16-1:0] node21168;
	wire [16-1:0] node21171;
	wire [16-1:0] node21172;
	wire [16-1:0] node21174;
	wire [16-1:0] node21177;
	wire [16-1:0] node21178;
	wire [16-1:0] node21182;
	wire [16-1:0] node21183;
	wire [16-1:0] node21184;
	wire [16-1:0] node21185;
	wire [16-1:0] node21186;
	wire [16-1:0] node21187;
	wire [16-1:0] node21188;
	wire [16-1:0] node21191;
	wire [16-1:0] node21194;
	wire [16-1:0] node21195;
	wire [16-1:0] node21199;
	wire [16-1:0] node21200;
	wire [16-1:0] node21202;
	wire [16-1:0] node21205;
	wire [16-1:0] node21206;
	wire [16-1:0] node21210;
	wire [16-1:0] node21211;
	wire [16-1:0] node21212;
	wire [16-1:0] node21213;
	wire [16-1:0] node21216;
	wire [16-1:0] node21219;
	wire [16-1:0] node21220;
	wire [16-1:0] node21224;
	wire [16-1:0] node21225;
	wire [16-1:0] node21226;
	wire [16-1:0] node21229;
	wire [16-1:0] node21232;
	wire [16-1:0] node21233;
	wire [16-1:0] node21237;
	wire [16-1:0] node21238;
	wire [16-1:0] node21239;
	wire [16-1:0] node21240;
	wire [16-1:0] node21241;
	wire [16-1:0] node21244;
	wire [16-1:0] node21247;
	wire [16-1:0] node21248;
	wire [16-1:0] node21251;
	wire [16-1:0] node21254;
	wire [16-1:0] node21255;
	wire [16-1:0] node21256;
	wire [16-1:0] node21259;
	wire [16-1:0] node21262;
	wire [16-1:0] node21263;
	wire [16-1:0] node21266;
	wire [16-1:0] node21269;
	wire [16-1:0] node21270;
	wire [16-1:0] node21271;
	wire [16-1:0] node21272;
	wire [16-1:0] node21275;
	wire [16-1:0] node21278;
	wire [16-1:0] node21279;
	wire [16-1:0] node21282;
	wire [16-1:0] node21285;
	wire [16-1:0] node21286;
	wire [16-1:0] node21287;
	wire [16-1:0] node21290;
	wire [16-1:0] node21293;
	wire [16-1:0] node21294;
	wire [16-1:0] node21297;
	wire [16-1:0] node21300;
	wire [16-1:0] node21301;
	wire [16-1:0] node21302;
	wire [16-1:0] node21303;
	wire [16-1:0] node21304;
	wire [16-1:0] node21305;
	wire [16-1:0] node21308;
	wire [16-1:0] node21311;
	wire [16-1:0] node21312;
	wire [16-1:0] node21315;
	wire [16-1:0] node21318;
	wire [16-1:0] node21319;
	wire [16-1:0] node21320;
	wire [16-1:0] node21323;
	wire [16-1:0] node21326;
	wire [16-1:0] node21327;
	wire [16-1:0] node21330;
	wire [16-1:0] node21333;
	wire [16-1:0] node21334;
	wire [16-1:0] node21335;
	wire [16-1:0] node21336;
	wire [16-1:0] node21339;
	wire [16-1:0] node21342;
	wire [16-1:0] node21343;
	wire [16-1:0] node21346;
	wire [16-1:0] node21349;
	wire [16-1:0] node21350;
	wire [16-1:0] node21352;
	wire [16-1:0] node21355;
	wire [16-1:0] node21357;
	wire [16-1:0] node21360;
	wire [16-1:0] node21361;
	wire [16-1:0] node21362;
	wire [16-1:0] node21363;
	wire [16-1:0] node21364;
	wire [16-1:0] node21367;
	wire [16-1:0] node21370;
	wire [16-1:0] node21372;
	wire [16-1:0] node21375;
	wire [16-1:0] node21376;
	wire [16-1:0] node21377;
	wire [16-1:0] node21380;
	wire [16-1:0] node21383;
	wire [16-1:0] node21384;
	wire [16-1:0] node21387;
	wire [16-1:0] node21390;
	wire [16-1:0] node21391;
	wire [16-1:0] node21392;
	wire [16-1:0] node21394;
	wire [16-1:0] node21397;
	wire [16-1:0] node21398;
	wire [16-1:0] node21401;
	wire [16-1:0] node21404;
	wire [16-1:0] node21405;
	wire [16-1:0] node21406;
	wire [16-1:0] node21409;
	wire [16-1:0] node21412;
	wire [16-1:0] node21413;
	wire [16-1:0] node21416;
	wire [16-1:0] node21419;
	wire [16-1:0] node21420;
	wire [16-1:0] node21421;
	wire [16-1:0] node21422;
	wire [16-1:0] node21423;
	wire [16-1:0] node21424;
	wire [16-1:0] node21425;
	wire [16-1:0] node21426;
	wire [16-1:0] node21427;
	wire [16-1:0] node21428;
	wire [16-1:0] node21431;
	wire [16-1:0] node21434;
	wire [16-1:0] node21435;
	wire [16-1:0] node21439;
	wire [16-1:0] node21440;
	wire [16-1:0] node21441;
	wire [16-1:0] node21444;
	wire [16-1:0] node21447;
	wire [16-1:0] node21449;
	wire [16-1:0] node21452;
	wire [16-1:0] node21453;
	wire [16-1:0] node21454;
	wire [16-1:0] node21455;
	wire [16-1:0] node21458;
	wire [16-1:0] node21461;
	wire [16-1:0] node21462;
	wire [16-1:0] node21465;
	wire [16-1:0] node21468;
	wire [16-1:0] node21469;
	wire [16-1:0] node21470;
	wire [16-1:0] node21473;
	wire [16-1:0] node21476;
	wire [16-1:0] node21478;
	wire [16-1:0] node21481;
	wire [16-1:0] node21482;
	wire [16-1:0] node21483;
	wire [16-1:0] node21484;
	wire [16-1:0] node21485;
	wire [16-1:0] node21488;
	wire [16-1:0] node21491;
	wire [16-1:0] node21492;
	wire [16-1:0] node21495;
	wire [16-1:0] node21498;
	wire [16-1:0] node21499;
	wire [16-1:0] node21500;
	wire [16-1:0] node21503;
	wire [16-1:0] node21506;
	wire [16-1:0] node21507;
	wire [16-1:0] node21510;
	wire [16-1:0] node21513;
	wire [16-1:0] node21514;
	wire [16-1:0] node21515;
	wire [16-1:0] node21516;
	wire [16-1:0] node21519;
	wire [16-1:0] node21522;
	wire [16-1:0] node21523;
	wire [16-1:0] node21526;
	wire [16-1:0] node21529;
	wire [16-1:0] node21530;
	wire [16-1:0] node21531;
	wire [16-1:0] node21534;
	wire [16-1:0] node21537;
	wire [16-1:0] node21538;
	wire [16-1:0] node21541;
	wire [16-1:0] node21544;
	wire [16-1:0] node21545;
	wire [16-1:0] node21546;
	wire [16-1:0] node21547;
	wire [16-1:0] node21548;
	wire [16-1:0] node21549;
	wire [16-1:0] node21552;
	wire [16-1:0] node21555;
	wire [16-1:0] node21556;
	wire [16-1:0] node21559;
	wire [16-1:0] node21562;
	wire [16-1:0] node21563;
	wire [16-1:0] node21564;
	wire [16-1:0] node21567;
	wire [16-1:0] node21570;
	wire [16-1:0] node21571;
	wire [16-1:0] node21574;
	wire [16-1:0] node21577;
	wire [16-1:0] node21578;
	wire [16-1:0] node21579;
	wire [16-1:0] node21581;
	wire [16-1:0] node21584;
	wire [16-1:0] node21585;
	wire [16-1:0] node21588;
	wire [16-1:0] node21591;
	wire [16-1:0] node21592;
	wire [16-1:0] node21593;
	wire [16-1:0] node21596;
	wire [16-1:0] node21599;
	wire [16-1:0] node21600;
	wire [16-1:0] node21603;
	wire [16-1:0] node21606;
	wire [16-1:0] node21607;
	wire [16-1:0] node21608;
	wire [16-1:0] node21609;
	wire [16-1:0] node21610;
	wire [16-1:0] node21614;
	wire [16-1:0] node21615;
	wire [16-1:0] node21618;
	wire [16-1:0] node21621;
	wire [16-1:0] node21622;
	wire [16-1:0] node21623;
	wire [16-1:0] node21626;
	wire [16-1:0] node21629;
	wire [16-1:0] node21630;
	wire [16-1:0] node21633;
	wire [16-1:0] node21636;
	wire [16-1:0] node21637;
	wire [16-1:0] node21638;
	wire [16-1:0] node21639;
	wire [16-1:0] node21642;
	wire [16-1:0] node21645;
	wire [16-1:0] node21646;
	wire [16-1:0] node21649;
	wire [16-1:0] node21652;
	wire [16-1:0] node21653;
	wire [16-1:0] node21654;
	wire [16-1:0] node21657;
	wire [16-1:0] node21660;
	wire [16-1:0] node21663;
	wire [16-1:0] node21664;
	wire [16-1:0] node21665;
	wire [16-1:0] node21666;
	wire [16-1:0] node21667;
	wire [16-1:0] node21668;
	wire [16-1:0] node21669;
	wire [16-1:0] node21672;
	wire [16-1:0] node21675;
	wire [16-1:0] node21676;
	wire [16-1:0] node21679;
	wire [16-1:0] node21682;
	wire [16-1:0] node21683;
	wire [16-1:0] node21684;
	wire [16-1:0] node21687;
	wire [16-1:0] node21690;
	wire [16-1:0] node21691;
	wire [16-1:0] node21694;
	wire [16-1:0] node21697;
	wire [16-1:0] node21698;
	wire [16-1:0] node21699;
	wire [16-1:0] node21700;
	wire [16-1:0] node21703;
	wire [16-1:0] node21706;
	wire [16-1:0] node21707;
	wire [16-1:0] node21710;
	wire [16-1:0] node21713;
	wire [16-1:0] node21714;
	wire [16-1:0] node21715;
	wire [16-1:0] node21718;
	wire [16-1:0] node21721;
	wire [16-1:0] node21722;
	wire [16-1:0] node21726;
	wire [16-1:0] node21727;
	wire [16-1:0] node21728;
	wire [16-1:0] node21729;
	wire [16-1:0] node21730;
	wire [16-1:0] node21733;
	wire [16-1:0] node21736;
	wire [16-1:0] node21737;
	wire [16-1:0] node21741;
	wire [16-1:0] node21742;
	wire [16-1:0] node21743;
	wire [16-1:0] node21746;
	wire [16-1:0] node21749;
	wire [16-1:0] node21750;
	wire [16-1:0] node21753;
	wire [16-1:0] node21756;
	wire [16-1:0] node21757;
	wire [16-1:0] node21758;
	wire [16-1:0] node21759;
	wire [16-1:0] node21762;
	wire [16-1:0] node21765;
	wire [16-1:0] node21766;
	wire [16-1:0] node21769;
	wire [16-1:0] node21772;
	wire [16-1:0] node21773;
	wire [16-1:0] node21774;
	wire [16-1:0] node21777;
	wire [16-1:0] node21780;
	wire [16-1:0] node21781;
	wire [16-1:0] node21784;
	wire [16-1:0] node21787;
	wire [16-1:0] node21788;
	wire [16-1:0] node21789;
	wire [16-1:0] node21790;
	wire [16-1:0] node21791;
	wire [16-1:0] node21792;
	wire [16-1:0] node21796;
	wire [16-1:0] node21797;
	wire [16-1:0] node21800;
	wire [16-1:0] node21803;
	wire [16-1:0] node21804;
	wire [16-1:0] node21806;
	wire [16-1:0] node21809;
	wire [16-1:0] node21810;
	wire [16-1:0] node21813;
	wire [16-1:0] node21816;
	wire [16-1:0] node21817;
	wire [16-1:0] node21818;
	wire [16-1:0] node21819;
	wire [16-1:0] node21822;
	wire [16-1:0] node21825;
	wire [16-1:0] node21826;
	wire [16-1:0] node21829;
	wire [16-1:0] node21832;
	wire [16-1:0] node21833;
	wire [16-1:0] node21834;
	wire [16-1:0] node21837;
	wire [16-1:0] node21840;
	wire [16-1:0] node21842;
	wire [16-1:0] node21845;
	wire [16-1:0] node21846;
	wire [16-1:0] node21847;
	wire [16-1:0] node21848;
	wire [16-1:0] node21849;
	wire [16-1:0] node21852;
	wire [16-1:0] node21855;
	wire [16-1:0] node21856;
	wire [16-1:0] node21859;
	wire [16-1:0] node21862;
	wire [16-1:0] node21863;
	wire [16-1:0] node21864;
	wire [16-1:0] node21867;
	wire [16-1:0] node21870;
	wire [16-1:0] node21871;
	wire [16-1:0] node21874;
	wire [16-1:0] node21877;
	wire [16-1:0] node21878;
	wire [16-1:0] node21879;
	wire [16-1:0] node21880;
	wire [16-1:0] node21883;
	wire [16-1:0] node21886;
	wire [16-1:0] node21887;
	wire [16-1:0] node21890;
	wire [16-1:0] node21893;
	wire [16-1:0] node21894;
	wire [16-1:0] node21896;
	wire [16-1:0] node21899;
	wire [16-1:0] node21900;
	wire [16-1:0] node21903;
	wire [16-1:0] node21906;
	wire [16-1:0] node21907;
	wire [16-1:0] node21908;
	wire [16-1:0] node21909;
	wire [16-1:0] node21910;
	wire [16-1:0] node21911;
	wire [16-1:0] node21912;
	wire [16-1:0] node21913;
	wire [16-1:0] node21916;
	wire [16-1:0] node21919;
	wire [16-1:0] node21920;
	wire [16-1:0] node21924;
	wire [16-1:0] node21925;
	wire [16-1:0] node21926;
	wire [16-1:0] node21929;
	wire [16-1:0] node21932;
	wire [16-1:0] node21933;
	wire [16-1:0] node21936;
	wire [16-1:0] node21939;
	wire [16-1:0] node21940;
	wire [16-1:0] node21941;
	wire [16-1:0] node21942;
	wire [16-1:0] node21945;
	wire [16-1:0] node21948;
	wire [16-1:0] node21949;
	wire [16-1:0] node21952;
	wire [16-1:0] node21955;
	wire [16-1:0] node21956;
	wire [16-1:0] node21957;
	wire [16-1:0] node21960;
	wire [16-1:0] node21963;
	wire [16-1:0] node21964;
	wire [16-1:0] node21968;
	wire [16-1:0] node21969;
	wire [16-1:0] node21970;
	wire [16-1:0] node21971;
	wire [16-1:0] node21972;
	wire [16-1:0] node21975;
	wire [16-1:0] node21978;
	wire [16-1:0] node21979;
	wire [16-1:0] node21982;
	wire [16-1:0] node21985;
	wire [16-1:0] node21986;
	wire [16-1:0] node21987;
	wire [16-1:0] node21990;
	wire [16-1:0] node21993;
	wire [16-1:0] node21994;
	wire [16-1:0] node21997;
	wire [16-1:0] node22000;
	wire [16-1:0] node22001;
	wire [16-1:0] node22002;
	wire [16-1:0] node22003;
	wire [16-1:0] node22006;
	wire [16-1:0] node22009;
	wire [16-1:0] node22010;
	wire [16-1:0] node22013;
	wire [16-1:0] node22016;
	wire [16-1:0] node22017;
	wire [16-1:0] node22018;
	wire [16-1:0] node22021;
	wire [16-1:0] node22024;
	wire [16-1:0] node22025;
	wire [16-1:0] node22028;
	wire [16-1:0] node22031;
	wire [16-1:0] node22032;
	wire [16-1:0] node22033;
	wire [16-1:0] node22034;
	wire [16-1:0] node22035;
	wire [16-1:0] node22036;
	wire [16-1:0] node22039;
	wire [16-1:0] node22042;
	wire [16-1:0] node22043;
	wire [16-1:0] node22046;
	wire [16-1:0] node22049;
	wire [16-1:0] node22050;
	wire [16-1:0] node22051;
	wire [16-1:0] node22054;
	wire [16-1:0] node22057;
	wire [16-1:0] node22058;
	wire [16-1:0] node22061;
	wire [16-1:0] node22064;
	wire [16-1:0] node22065;
	wire [16-1:0] node22066;
	wire [16-1:0] node22067;
	wire [16-1:0] node22070;
	wire [16-1:0] node22073;
	wire [16-1:0] node22074;
	wire [16-1:0] node22077;
	wire [16-1:0] node22080;
	wire [16-1:0] node22081;
	wire [16-1:0] node22082;
	wire [16-1:0] node22085;
	wire [16-1:0] node22088;
	wire [16-1:0] node22089;
	wire [16-1:0] node22092;
	wire [16-1:0] node22095;
	wire [16-1:0] node22096;
	wire [16-1:0] node22097;
	wire [16-1:0] node22098;
	wire [16-1:0] node22099;
	wire [16-1:0] node22102;
	wire [16-1:0] node22105;
	wire [16-1:0] node22106;
	wire [16-1:0] node22110;
	wire [16-1:0] node22111;
	wire [16-1:0] node22112;
	wire [16-1:0] node22115;
	wire [16-1:0] node22118;
	wire [16-1:0] node22119;
	wire [16-1:0] node22122;
	wire [16-1:0] node22125;
	wire [16-1:0] node22126;
	wire [16-1:0] node22127;
	wire [16-1:0] node22128;
	wire [16-1:0] node22131;
	wire [16-1:0] node22134;
	wire [16-1:0] node22135;
	wire [16-1:0] node22138;
	wire [16-1:0] node22141;
	wire [16-1:0] node22142;
	wire [16-1:0] node22143;
	wire [16-1:0] node22146;
	wire [16-1:0] node22149;
	wire [16-1:0] node22150;
	wire [16-1:0] node22153;
	wire [16-1:0] node22156;
	wire [16-1:0] node22157;
	wire [16-1:0] node22158;
	wire [16-1:0] node22159;
	wire [16-1:0] node22160;
	wire [16-1:0] node22161;
	wire [16-1:0] node22162;
	wire [16-1:0] node22165;
	wire [16-1:0] node22168;
	wire [16-1:0] node22170;
	wire [16-1:0] node22173;
	wire [16-1:0] node22174;
	wire [16-1:0] node22175;
	wire [16-1:0] node22178;
	wire [16-1:0] node22181;
	wire [16-1:0] node22183;
	wire [16-1:0] node22186;
	wire [16-1:0] node22187;
	wire [16-1:0] node22188;
	wire [16-1:0] node22189;
	wire [16-1:0] node22192;
	wire [16-1:0] node22195;
	wire [16-1:0] node22196;
	wire [16-1:0] node22199;
	wire [16-1:0] node22202;
	wire [16-1:0] node22203;
	wire [16-1:0] node22204;
	wire [16-1:0] node22207;
	wire [16-1:0] node22210;
	wire [16-1:0] node22211;
	wire [16-1:0] node22214;
	wire [16-1:0] node22217;
	wire [16-1:0] node22218;
	wire [16-1:0] node22219;
	wire [16-1:0] node22220;
	wire [16-1:0] node22221;
	wire [16-1:0] node22224;
	wire [16-1:0] node22227;
	wire [16-1:0] node22228;
	wire [16-1:0] node22231;
	wire [16-1:0] node22234;
	wire [16-1:0] node22235;
	wire [16-1:0] node22236;
	wire [16-1:0] node22239;
	wire [16-1:0] node22242;
	wire [16-1:0] node22243;
	wire [16-1:0] node22247;
	wire [16-1:0] node22248;
	wire [16-1:0] node22249;
	wire [16-1:0] node22250;
	wire [16-1:0] node22253;
	wire [16-1:0] node22256;
	wire [16-1:0] node22257;
	wire [16-1:0] node22260;
	wire [16-1:0] node22263;
	wire [16-1:0] node22264;
	wire [16-1:0] node22265;
	wire [16-1:0] node22268;
	wire [16-1:0] node22271;
	wire [16-1:0] node22272;
	wire [16-1:0] node22275;
	wire [16-1:0] node22278;
	wire [16-1:0] node22279;
	wire [16-1:0] node22280;
	wire [16-1:0] node22281;
	wire [16-1:0] node22282;
	wire [16-1:0] node22283;
	wire [16-1:0] node22286;
	wire [16-1:0] node22289;
	wire [16-1:0] node22290;
	wire [16-1:0] node22293;
	wire [16-1:0] node22296;
	wire [16-1:0] node22297;
	wire [16-1:0] node22298;
	wire [16-1:0] node22301;
	wire [16-1:0] node22304;
	wire [16-1:0] node22305;
	wire [16-1:0] node22308;
	wire [16-1:0] node22311;
	wire [16-1:0] node22312;
	wire [16-1:0] node22313;
	wire [16-1:0] node22314;
	wire [16-1:0] node22317;
	wire [16-1:0] node22320;
	wire [16-1:0] node22321;
	wire [16-1:0] node22324;
	wire [16-1:0] node22327;
	wire [16-1:0] node22328;
	wire [16-1:0] node22329;
	wire [16-1:0] node22332;
	wire [16-1:0] node22335;
	wire [16-1:0] node22336;
	wire [16-1:0] node22339;
	wire [16-1:0] node22342;
	wire [16-1:0] node22343;
	wire [16-1:0] node22344;
	wire [16-1:0] node22345;
	wire [16-1:0] node22347;
	wire [16-1:0] node22350;
	wire [16-1:0] node22351;
	wire [16-1:0] node22354;
	wire [16-1:0] node22357;
	wire [16-1:0] node22358;
	wire [16-1:0] node22359;
	wire [16-1:0] node22362;
	wire [16-1:0] node22365;
	wire [16-1:0] node22366;
	wire [16-1:0] node22369;
	wire [16-1:0] node22372;
	wire [16-1:0] node22373;
	wire [16-1:0] node22374;
	wire [16-1:0] node22375;
	wire [16-1:0] node22378;
	wire [16-1:0] node22381;
	wire [16-1:0] node22382;
	wire [16-1:0] node22385;
	wire [16-1:0] node22388;
	wire [16-1:0] node22389;
	wire [16-1:0] node22390;
	wire [16-1:0] node22393;
	wire [16-1:0] node22396;
	wire [16-1:0] node22397;
	wire [16-1:0] node22400;
	wire [16-1:0] node22403;
	wire [16-1:0] node22404;
	wire [16-1:0] node22405;
	wire [16-1:0] node22406;
	wire [16-1:0] node22407;
	wire [16-1:0] node22408;
	wire [16-1:0] node22409;
	wire [16-1:0] node22410;
	wire [16-1:0] node22411;
	wire [16-1:0] node22414;
	wire [16-1:0] node22417;
	wire [16-1:0] node22418;
	wire [16-1:0] node22421;
	wire [16-1:0] node22424;
	wire [16-1:0] node22425;
	wire [16-1:0] node22426;
	wire [16-1:0] node22429;
	wire [16-1:0] node22432;
	wire [16-1:0] node22433;
	wire [16-1:0] node22437;
	wire [16-1:0] node22438;
	wire [16-1:0] node22439;
	wire [16-1:0] node22440;
	wire [16-1:0] node22443;
	wire [16-1:0] node22446;
	wire [16-1:0] node22447;
	wire [16-1:0] node22450;
	wire [16-1:0] node22453;
	wire [16-1:0] node22454;
	wire [16-1:0] node22455;
	wire [16-1:0] node22458;
	wire [16-1:0] node22461;
	wire [16-1:0] node22462;
	wire [16-1:0] node22465;
	wire [16-1:0] node22468;
	wire [16-1:0] node22469;
	wire [16-1:0] node22470;
	wire [16-1:0] node22471;
	wire [16-1:0] node22472;
	wire [16-1:0] node22475;
	wire [16-1:0] node22478;
	wire [16-1:0] node22479;
	wire [16-1:0] node22482;
	wire [16-1:0] node22485;
	wire [16-1:0] node22486;
	wire [16-1:0] node22487;
	wire [16-1:0] node22490;
	wire [16-1:0] node22493;
	wire [16-1:0] node22494;
	wire [16-1:0] node22497;
	wire [16-1:0] node22500;
	wire [16-1:0] node22501;
	wire [16-1:0] node22502;
	wire [16-1:0] node22503;
	wire [16-1:0] node22506;
	wire [16-1:0] node22509;
	wire [16-1:0] node22510;
	wire [16-1:0] node22513;
	wire [16-1:0] node22516;
	wire [16-1:0] node22517;
	wire [16-1:0] node22518;
	wire [16-1:0] node22521;
	wire [16-1:0] node22524;
	wire [16-1:0] node22525;
	wire [16-1:0] node22528;
	wire [16-1:0] node22531;
	wire [16-1:0] node22532;
	wire [16-1:0] node22533;
	wire [16-1:0] node22534;
	wire [16-1:0] node22535;
	wire [16-1:0] node22536;
	wire [16-1:0] node22540;
	wire [16-1:0] node22541;
	wire [16-1:0] node22544;
	wire [16-1:0] node22547;
	wire [16-1:0] node22548;
	wire [16-1:0] node22549;
	wire [16-1:0] node22552;
	wire [16-1:0] node22555;
	wire [16-1:0] node22556;
	wire [16-1:0] node22559;
	wire [16-1:0] node22562;
	wire [16-1:0] node22563;
	wire [16-1:0] node22564;
	wire [16-1:0] node22565;
	wire [16-1:0] node22569;
	wire [16-1:0] node22570;
	wire [16-1:0] node22573;
	wire [16-1:0] node22576;
	wire [16-1:0] node22577;
	wire [16-1:0] node22578;
	wire [16-1:0] node22581;
	wire [16-1:0] node22584;
	wire [16-1:0] node22585;
	wire [16-1:0] node22588;
	wire [16-1:0] node22591;
	wire [16-1:0] node22592;
	wire [16-1:0] node22593;
	wire [16-1:0] node22594;
	wire [16-1:0] node22595;
	wire [16-1:0] node22598;
	wire [16-1:0] node22601;
	wire [16-1:0] node22602;
	wire [16-1:0] node22605;
	wire [16-1:0] node22608;
	wire [16-1:0] node22609;
	wire [16-1:0] node22611;
	wire [16-1:0] node22614;
	wire [16-1:0] node22615;
	wire [16-1:0] node22618;
	wire [16-1:0] node22621;
	wire [16-1:0] node22622;
	wire [16-1:0] node22623;
	wire [16-1:0] node22624;
	wire [16-1:0] node22627;
	wire [16-1:0] node22630;
	wire [16-1:0] node22631;
	wire [16-1:0] node22634;
	wire [16-1:0] node22637;
	wire [16-1:0] node22638;
	wire [16-1:0] node22640;
	wire [16-1:0] node22643;
	wire [16-1:0] node22644;
	wire [16-1:0] node22647;
	wire [16-1:0] node22650;
	wire [16-1:0] node22651;
	wire [16-1:0] node22652;
	wire [16-1:0] node22653;
	wire [16-1:0] node22654;
	wire [16-1:0] node22655;
	wire [16-1:0] node22657;
	wire [16-1:0] node22660;
	wire [16-1:0] node22661;
	wire [16-1:0] node22664;
	wire [16-1:0] node22667;
	wire [16-1:0] node22668;
	wire [16-1:0] node22669;
	wire [16-1:0] node22672;
	wire [16-1:0] node22675;
	wire [16-1:0] node22676;
	wire [16-1:0] node22679;
	wire [16-1:0] node22682;
	wire [16-1:0] node22683;
	wire [16-1:0] node22684;
	wire [16-1:0] node22685;
	wire [16-1:0] node22688;
	wire [16-1:0] node22691;
	wire [16-1:0] node22692;
	wire [16-1:0] node22695;
	wire [16-1:0] node22698;
	wire [16-1:0] node22699;
	wire [16-1:0] node22701;
	wire [16-1:0] node22704;
	wire [16-1:0] node22705;
	wire [16-1:0] node22709;
	wire [16-1:0] node22710;
	wire [16-1:0] node22711;
	wire [16-1:0] node22712;
	wire [16-1:0] node22713;
	wire [16-1:0] node22716;
	wire [16-1:0] node22719;
	wire [16-1:0] node22720;
	wire [16-1:0] node22723;
	wire [16-1:0] node22726;
	wire [16-1:0] node22727;
	wire [16-1:0] node22728;
	wire [16-1:0] node22731;
	wire [16-1:0] node22734;
	wire [16-1:0] node22735;
	wire [16-1:0] node22738;
	wire [16-1:0] node22741;
	wire [16-1:0] node22742;
	wire [16-1:0] node22743;
	wire [16-1:0] node22744;
	wire [16-1:0] node22747;
	wire [16-1:0] node22750;
	wire [16-1:0] node22751;
	wire [16-1:0] node22754;
	wire [16-1:0] node22757;
	wire [16-1:0] node22758;
	wire [16-1:0] node22759;
	wire [16-1:0] node22762;
	wire [16-1:0] node22765;
	wire [16-1:0] node22766;
	wire [16-1:0] node22769;
	wire [16-1:0] node22772;
	wire [16-1:0] node22773;
	wire [16-1:0] node22774;
	wire [16-1:0] node22775;
	wire [16-1:0] node22776;
	wire [16-1:0] node22777;
	wire [16-1:0] node22780;
	wire [16-1:0] node22783;
	wire [16-1:0] node22784;
	wire [16-1:0] node22787;
	wire [16-1:0] node22790;
	wire [16-1:0] node22791;
	wire [16-1:0] node22792;
	wire [16-1:0] node22795;
	wire [16-1:0] node22798;
	wire [16-1:0] node22799;
	wire [16-1:0] node22802;
	wire [16-1:0] node22805;
	wire [16-1:0] node22806;
	wire [16-1:0] node22807;
	wire [16-1:0] node22808;
	wire [16-1:0] node22811;
	wire [16-1:0] node22814;
	wire [16-1:0] node22815;
	wire [16-1:0] node22818;
	wire [16-1:0] node22821;
	wire [16-1:0] node22822;
	wire [16-1:0] node22823;
	wire [16-1:0] node22826;
	wire [16-1:0] node22829;
	wire [16-1:0] node22830;
	wire [16-1:0] node22833;
	wire [16-1:0] node22836;
	wire [16-1:0] node22837;
	wire [16-1:0] node22838;
	wire [16-1:0] node22839;
	wire [16-1:0] node22840;
	wire [16-1:0] node22843;
	wire [16-1:0] node22846;
	wire [16-1:0] node22847;
	wire [16-1:0] node22850;
	wire [16-1:0] node22853;
	wire [16-1:0] node22854;
	wire [16-1:0] node22855;
	wire [16-1:0] node22858;
	wire [16-1:0] node22861;
	wire [16-1:0] node22862;
	wire [16-1:0] node22865;
	wire [16-1:0] node22868;
	wire [16-1:0] node22869;
	wire [16-1:0] node22870;
	wire [16-1:0] node22872;
	wire [16-1:0] node22875;
	wire [16-1:0] node22876;
	wire [16-1:0] node22879;
	wire [16-1:0] node22882;
	wire [16-1:0] node22883;
	wire [16-1:0] node22884;
	wire [16-1:0] node22887;
	wire [16-1:0] node22890;
	wire [16-1:0] node22891;
	wire [16-1:0] node22894;
	wire [16-1:0] node22897;
	wire [16-1:0] node22898;
	wire [16-1:0] node22899;
	wire [16-1:0] node22900;
	wire [16-1:0] node22901;
	wire [16-1:0] node22902;
	wire [16-1:0] node22903;
	wire [16-1:0] node22904;
	wire [16-1:0] node22907;
	wire [16-1:0] node22910;
	wire [16-1:0] node22911;
	wire [16-1:0] node22914;
	wire [16-1:0] node22917;
	wire [16-1:0] node22918;
	wire [16-1:0] node22919;
	wire [16-1:0] node22923;
	wire [16-1:0] node22924;
	wire [16-1:0] node22927;
	wire [16-1:0] node22930;
	wire [16-1:0] node22931;
	wire [16-1:0] node22932;
	wire [16-1:0] node22933;
	wire [16-1:0] node22936;
	wire [16-1:0] node22939;
	wire [16-1:0] node22940;
	wire [16-1:0] node22943;
	wire [16-1:0] node22946;
	wire [16-1:0] node22947;
	wire [16-1:0] node22948;
	wire [16-1:0] node22952;
	wire [16-1:0] node22954;
	wire [16-1:0] node22957;
	wire [16-1:0] node22958;
	wire [16-1:0] node22959;
	wire [16-1:0] node22960;
	wire [16-1:0] node22961;
	wire [16-1:0] node22964;
	wire [16-1:0] node22967;
	wire [16-1:0] node22968;
	wire [16-1:0] node22971;
	wire [16-1:0] node22974;
	wire [16-1:0] node22975;
	wire [16-1:0] node22976;
	wire [16-1:0] node22979;
	wire [16-1:0] node22982;
	wire [16-1:0] node22983;
	wire [16-1:0] node22986;
	wire [16-1:0] node22989;
	wire [16-1:0] node22990;
	wire [16-1:0] node22991;
	wire [16-1:0] node22992;
	wire [16-1:0] node22995;
	wire [16-1:0] node22998;
	wire [16-1:0] node22999;
	wire [16-1:0] node23002;
	wire [16-1:0] node23005;
	wire [16-1:0] node23006;
	wire [16-1:0] node23007;
	wire [16-1:0] node23011;
	wire [16-1:0] node23012;
	wire [16-1:0] node23015;
	wire [16-1:0] node23018;
	wire [16-1:0] node23019;
	wire [16-1:0] node23020;
	wire [16-1:0] node23021;
	wire [16-1:0] node23022;
	wire [16-1:0] node23023;
	wire [16-1:0] node23026;
	wire [16-1:0] node23029;
	wire [16-1:0] node23030;
	wire [16-1:0] node23033;
	wire [16-1:0] node23036;
	wire [16-1:0] node23037;
	wire [16-1:0] node23038;
	wire [16-1:0] node23041;
	wire [16-1:0] node23044;
	wire [16-1:0] node23045;
	wire [16-1:0] node23048;
	wire [16-1:0] node23051;
	wire [16-1:0] node23052;
	wire [16-1:0] node23053;
	wire [16-1:0] node23054;
	wire [16-1:0] node23057;
	wire [16-1:0] node23060;
	wire [16-1:0] node23061;
	wire [16-1:0] node23064;
	wire [16-1:0] node23067;
	wire [16-1:0] node23068;
	wire [16-1:0] node23069;
	wire [16-1:0] node23072;
	wire [16-1:0] node23075;
	wire [16-1:0] node23076;
	wire [16-1:0] node23079;
	wire [16-1:0] node23082;
	wire [16-1:0] node23083;
	wire [16-1:0] node23084;
	wire [16-1:0] node23085;
	wire [16-1:0] node23087;
	wire [16-1:0] node23090;
	wire [16-1:0] node23091;
	wire [16-1:0] node23094;
	wire [16-1:0] node23097;
	wire [16-1:0] node23098;
	wire [16-1:0] node23099;
	wire [16-1:0] node23102;
	wire [16-1:0] node23105;
	wire [16-1:0] node23106;
	wire [16-1:0] node23109;
	wire [16-1:0] node23112;
	wire [16-1:0] node23113;
	wire [16-1:0] node23114;
	wire [16-1:0] node23115;
	wire [16-1:0] node23118;
	wire [16-1:0] node23121;
	wire [16-1:0] node23122;
	wire [16-1:0] node23125;
	wire [16-1:0] node23128;
	wire [16-1:0] node23129;
	wire [16-1:0] node23130;
	wire [16-1:0] node23133;
	wire [16-1:0] node23136;
	wire [16-1:0] node23137;
	wire [16-1:0] node23140;
	wire [16-1:0] node23143;
	wire [16-1:0] node23144;
	wire [16-1:0] node23145;
	wire [16-1:0] node23146;
	wire [16-1:0] node23147;
	wire [16-1:0] node23148;
	wire [16-1:0] node23149;
	wire [16-1:0] node23152;
	wire [16-1:0] node23155;
	wire [16-1:0] node23156;
	wire [16-1:0] node23159;
	wire [16-1:0] node23162;
	wire [16-1:0] node23163;
	wire [16-1:0] node23164;
	wire [16-1:0] node23167;
	wire [16-1:0] node23170;
	wire [16-1:0] node23171;
	wire [16-1:0] node23174;
	wire [16-1:0] node23177;
	wire [16-1:0] node23178;
	wire [16-1:0] node23179;
	wire [16-1:0] node23180;
	wire [16-1:0] node23183;
	wire [16-1:0] node23186;
	wire [16-1:0] node23187;
	wire [16-1:0] node23190;
	wire [16-1:0] node23193;
	wire [16-1:0] node23194;
	wire [16-1:0] node23195;
	wire [16-1:0] node23198;
	wire [16-1:0] node23201;
	wire [16-1:0] node23202;
	wire [16-1:0] node23205;
	wire [16-1:0] node23208;
	wire [16-1:0] node23209;
	wire [16-1:0] node23210;
	wire [16-1:0] node23211;
	wire [16-1:0] node23213;
	wire [16-1:0] node23216;
	wire [16-1:0] node23217;
	wire [16-1:0] node23220;
	wire [16-1:0] node23223;
	wire [16-1:0] node23224;
	wire [16-1:0] node23225;
	wire [16-1:0] node23228;
	wire [16-1:0] node23231;
	wire [16-1:0] node23232;
	wire [16-1:0] node23235;
	wire [16-1:0] node23238;
	wire [16-1:0] node23239;
	wire [16-1:0] node23240;
	wire [16-1:0] node23242;
	wire [16-1:0] node23245;
	wire [16-1:0] node23247;
	wire [16-1:0] node23250;
	wire [16-1:0] node23251;
	wire [16-1:0] node23252;
	wire [16-1:0] node23255;
	wire [16-1:0] node23258;
	wire [16-1:0] node23259;
	wire [16-1:0] node23262;
	wire [16-1:0] node23265;
	wire [16-1:0] node23266;
	wire [16-1:0] node23267;
	wire [16-1:0] node23268;
	wire [16-1:0] node23269;
	wire [16-1:0] node23271;
	wire [16-1:0] node23274;
	wire [16-1:0] node23275;
	wire [16-1:0] node23278;
	wire [16-1:0] node23281;
	wire [16-1:0] node23282;
	wire [16-1:0] node23283;
	wire [16-1:0] node23286;
	wire [16-1:0] node23289;
	wire [16-1:0] node23290;
	wire [16-1:0] node23293;
	wire [16-1:0] node23296;
	wire [16-1:0] node23297;
	wire [16-1:0] node23298;
	wire [16-1:0] node23299;
	wire [16-1:0] node23302;
	wire [16-1:0] node23305;
	wire [16-1:0] node23306;
	wire [16-1:0] node23309;
	wire [16-1:0] node23312;
	wire [16-1:0] node23313;
	wire [16-1:0] node23315;
	wire [16-1:0] node23318;
	wire [16-1:0] node23319;
	wire [16-1:0] node23322;
	wire [16-1:0] node23325;
	wire [16-1:0] node23326;
	wire [16-1:0] node23327;
	wire [16-1:0] node23328;
	wire [16-1:0] node23329;
	wire [16-1:0] node23332;
	wire [16-1:0] node23335;
	wire [16-1:0] node23336;
	wire [16-1:0] node23339;
	wire [16-1:0] node23342;
	wire [16-1:0] node23343;
	wire [16-1:0] node23344;
	wire [16-1:0] node23347;
	wire [16-1:0] node23350;
	wire [16-1:0] node23351;
	wire [16-1:0] node23354;
	wire [16-1:0] node23357;
	wire [16-1:0] node23358;
	wire [16-1:0] node23359;
	wire [16-1:0] node23360;
	wire [16-1:0] node23363;
	wire [16-1:0] node23366;
	wire [16-1:0] node23367;
	wire [16-1:0] node23370;
	wire [16-1:0] node23373;
	wire [16-1:0] node23374;
	wire [16-1:0] node23375;
	wire [16-1:0] node23378;
	wire [16-1:0] node23381;
	wire [16-1:0] node23382;
	wire [16-1:0] node23385;
	wire [16-1:0] node23388;
	wire [16-1:0] node23389;
	wire [16-1:0] node23390;
	wire [16-1:0] node23391;
	wire [16-1:0] node23392;
	wire [16-1:0] node23393;
	wire [16-1:0] node23394;
	wire [16-1:0] node23395;
	wire [16-1:0] node23396;
	wire [16-1:0] node23397;
	wire [16-1:0] node23398;
	wire [16-1:0] node23399;
	wire [16-1:0] node23402;
	wire [16-1:0] node23405;
	wire [16-1:0] node23406;
	wire [16-1:0] node23409;
	wire [16-1:0] node23412;
	wire [16-1:0] node23413;
	wire [16-1:0] node23414;
	wire [16-1:0] node23417;
	wire [16-1:0] node23420;
	wire [16-1:0] node23421;
	wire [16-1:0] node23424;
	wire [16-1:0] node23427;
	wire [16-1:0] node23428;
	wire [16-1:0] node23429;
	wire [16-1:0] node23430;
	wire [16-1:0] node23433;
	wire [16-1:0] node23436;
	wire [16-1:0] node23437;
	wire [16-1:0] node23440;
	wire [16-1:0] node23443;
	wire [16-1:0] node23444;
	wire [16-1:0] node23445;
	wire [16-1:0] node23448;
	wire [16-1:0] node23451;
	wire [16-1:0] node23453;
	wire [16-1:0] node23456;
	wire [16-1:0] node23457;
	wire [16-1:0] node23458;
	wire [16-1:0] node23459;
	wire [16-1:0] node23462;
	wire [16-1:0] node23463;
	wire [16-1:0] node23466;
	wire [16-1:0] node23469;
	wire [16-1:0] node23470;
	wire [16-1:0] node23471;
	wire [16-1:0] node23474;
	wire [16-1:0] node23477;
	wire [16-1:0] node23478;
	wire [16-1:0] node23481;
	wire [16-1:0] node23484;
	wire [16-1:0] node23485;
	wire [16-1:0] node23486;
	wire [16-1:0] node23487;
	wire [16-1:0] node23490;
	wire [16-1:0] node23493;
	wire [16-1:0] node23494;
	wire [16-1:0] node23497;
	wire [16-1:0] node23500;
	wire [16-1:0] node23501;
	wire [16-1:0] node23502;
	wire [16-1:0] node23505;
	wire [16-1:0] node23508;
	wire [16-1:0] node23510;
	wire [16-1:0] node23513;
	wire [16-1:0] node23514;
	wire [16-1:0] node23515;
	wire [16-1:0] node23516;
	wire [16-1:0] node23517;
	wire [16-1:0] node23518;
	wire [16-1:0] node23521;
	wire [16-1:0] node23524;
	wire [16-1:0] node23525;
	wire [16-1:0] node23528;
	wire [16-1:0] node23531;
	wire [16-1:0] node23532;
	wire [16-1:0] node23533;
	wire [16-1:0] node23537;
	wire [16-1:0] node23538;
	wire [16-1:0] node23541;
	wire [16-1:0] node23544;
	wire [16-1:0] node23545;
	wire [16-1:0] node23546;
	wire [16-1:0] node23547;
	wire [16-1:0] node23550;
	wire [16-1:0] node23553;
	wire [16-1:0] node23554;
	wire [16-1:0] node23557;
	wire [16-1:0] node23560;
	wire [16-1:0] node23561;
	wire [16-1:0] node23562;
	wire [16-1:0] node23565;
	wire [16-1:0] node23568;
	wire [16-1:0] node23569;
	wire [16-1:0] node23572;
	wire [16-1:0] node23575;
	wire [16-1:0] node23576;
	wire [16-1:0] node23577;
	wire [16-1:0] node23578;
	wire [16-1:0] node23579;
	wire [16-1:0] node23582;
	wire [16-1:0] node23585;
	wire [16-1:0] node23586;
	wire [16-1:0] node23589;
	wire [16-1:0] node23592;
	wire [16-1:0] node23593;
	wire [16-1:0] node23594;
	wire [16-1:0] node23597;
	wire [16-1:0] node23600;
	wire [16-1:0] node23601;
	wire [16-1:0] node23604;
	wire [16-1:0] node23607;
	wire [16-1:0] node23608;
	wire [16-1:0] node23609;
	wire [16-1:0] node23610;
	wire [16-1:0] node23613;
	wire [16-1:0] node23616;
	wire [16-1:0] node23617;
	wire [16-1:0] node23620;
	wire [16-1:0] node23623;
	wire [16-1:0] node23624;
	wire [16-1:0] node23625;
	wire [16-1:0] node23629;
	wire [16-1:0] node23630;
	wire [16-1:0] node23634;
	wire [16-1:0] node23635;
	wire [16-1:0] node23636;
	wire [16-1:0] node23637;
	wire [16-1:0] node23638;
	wire [16-1:0] node23639;
	wire [16-1:0] node23640;
	wire [16-1:0] node23643;
	wire [16-1:0] node23647;
	wire [16-1:0] node23648;
	wire [16-1:0] node23649;
	wire [16-1:0] node23652;
	wire [16-1:0] node23655;
	wire [16-1:0] node23656;
	wire [16-1:0] node23659;
	wire [16-1:0] node23662;
	wire [16-1:0] node23663;
	wire [16-1:0] node23664;
	wire [16-1:0] node23665;
	wire [16-1:0] node23668;
	wire [16-1:0] node23671;
	wire [16-1:0] node23672;
	wire [16-1:0] node23675;
	wire [16-1:0] node23678;
	wire [16-1:0] node23680;
	wire [16-1:0] node23681;
	wire [16-1:0] node23684;
	wire [16-1:0] node23687;
	wire [16-1:0] node23688;
	wire [16-1:0] node23689;
	wire [16-1:0] node23690;
	wire [16-1:0] node23691;
	wire [16-1:0] node23694;
	wire [16-1:0] node23697;
	wire [16-1:0] node23698;
	wire [16-1:0] node23701;
	wire [16-1:0] node23704;
	wire [16-1:0] node23705;
	wire [16-1:0] node23706;
	wire [16-1:0] node23709;
	wire [16-1:0] node23712;
	wire [16-1:0] node23713;
	wire [16-1:0] node23716;
	wire [16-1:0] node23719;
	wire [16-1:0] node23720;
	wire [16-1:0] node23721;
	wire [16-1:0] node23722;
	wire [16-1:0] node23725;
	wire [16-1:0] node23728;
	wire [16-1:0] node23729;
	wire [16-1:0] node23732;
	wire [16-1:0] node23735;
	wire [16-1:0] node23736;
	wire [16-1:0] node23737;
	wire [16-1:0] node23740;
	wire [16-1:0] node23743;
	wire [16-1:0] node23745;
	wire [16-1:0] node23748;
	wire [16-1:0] node23749;
	wire [16-1:0] node23750;
	wire [16-1:0] node23751;
	wire [16-1:0] node23752;
	wire [16-1:0] node23753;
	wire [16-1:0] node23756;
	wire [16-1:0] node23759;
	wire [16-1:0] node23760;
	wire [16-1:0] node23763;
	wire [16-1:0] node23766;
	wire [16-1:0] node23767;
	wire [16-1:0] node23768;
	wire [16-1:0] node23771;
	wire [16-1:0] node23774;
	wire [16-1:0] node23775;
	wire [16-1:0] node23778;
	wire [16-1:0] node23781;
	wire [16-1:0] node23782;
	wire [16-1:0] node23783;
	wire [16-1:0] node23784;
	wire [16-1:0] node23787;
	wire [16-1:0] node23790;
	wire [16-1:0] node23791;
	wire [16-1:0] node23795;
	wire [16-1:0] node23796;
	wire [16-1:0] node23797;
	wire [16-1:0] node23800;
	wire [16-1:0] node23803;
	wire [16-1:0] node23804;
	wire [16-1:0] node23807;
	wire [16-1:0] node23810;
	wire [16-1:0] node23811;
	wire [16-1:0] node23812;
	wire [16-1:0] node23813;
	wire [16-1:0] node23814;
	wire [16-1:0] node23817;
	wire [16-1:0] node23820;
	wire [16-1:0] node23821;
	wire [16-1:0] node23824;
	wire [16-1:0] node23827;
	wire [16-1:0] node23828;
	wire [16-1:0] node23829;
	wire [16-1:0] node23832;
	wire [16-1:0] node23835;
	wire [16-1:0] node23836;
	wire [16-1:0] node23839;
	wire [16-1:0] node23842;
	wire [16-1:0] node23843;
	wire [16-1:0] node23844;
	wire [16-1:0] node23845;
	wire [16-1:0] node23848;
	wire [16-1:0] node23851;
	wire [16-1:0] node23852;
	wire [16-1:0] node23855;
	wire [16-1:0] node23858;
	wire [16-1:0] node23859;
	wire [16-1:0] node23860;
	wire [16-1:0] node23863;
	wire [16-1:0] node23866;
	wire [16-1:0] node23867;
	wire [16-1:0] node23870;
	wire [16-1:0] node23873;
	wire [16-1:0] node23874;
	wire [16-1:0] node23875;
	wire [16-1:0] node23876;
	wire [16-1:0] node23877;
	wire [16-1:0] node23878;
	wire [16-1:0] node23879;
	wire [16-1:0] node23880;
	wire [16-1:0] node23883;
	wire [16-1:0] node23886;
	wire [16-1:0] node23887;
	wire [16-1:0] node23890;
	wire [16-1:0] node23893;
	wire [16-1:0] node23894;
	wire [16-1:0] node23895;
	wire [16-1:0] node23898;
	wire [16-1:0] node23901;
	wire [16-1:0] node23902;
	wire [16-1:0] node23906;
	wire [16-1:0] node23907;
	wire [16-1:0] node23908;
	wire [16-1:0] node23909;
	wire [16-1:0] node23912;
	wire [16-1:0] node23915;
	wire [16-1:0] node23916;
	wire [16-1:0] node23919;
	wire [16-1:0] node23922;
	wire [16-1:0] node23923;
	wire [16-1:0] node23924;
	wire [16-1:0] node23927;
	wire [16-1:0] node23930;
	wire [16-1:0] node23931;
	wire [16-1:0] node23934;
	wire [16-1:0] node23937;
	wire [16-1:0] node23938;
	wire [16-1:0] node23939;
	wire [16-1:0] node23940;
	wire [16-1:0] node23941;
	wire [16-1:0] node23944;
	wire [16-1:0] node23947;
	wire [16-1:0] node23948;
	wire [16-1:0] node23951;
	wire [16-1:0] node23954;
	wire [16-1:0] node23955;
	wire [16-1:0] node23956;
	wire [16-1:0] node23959;
	wire [16-1:0] node23962;
	wire [16-1:0] node23964;
	wire [16-1:0] node23967;
	wire [16-1:0] node23968;
	wire [16-1:0] node23970;
	wire [16-1:0] node23971;
	wire [16-1:0] node23974;
	wire [16-1:0] node23977;
	wire [16-1:0] node23978;
	wire [16-1:0] node23979;
	wire [16-1:0] node23982;
	wire [16-1:0] node23985;
	wire [16-1:0] node23986;
	wire [16-1:0] node23989;
	wire [16-1:0] node23992;
	wire [16-1:0] node23993;
	wire [16-1:0] node23994;
	wire [16-1:0] node23995;
	wire [16-1:0] node23996;
	wire [16-1:0] node23997;
	wire [16-1:0] node24000;
	wire [16-1:0] node24003;
	wire [16-1:0] node24004;
	wire [16-1:0] node24008;
	wire [16-1:0] node24009;
	wire [16-1:0] node24010;
	wire [16-1:0] node24013;
	wire [16-1:0] node24016;
	wire [16-1:0] node24017;
	wire [16-1:0] node24021;
	wire [16-1:0] node24022;
	wire [16-1:0] node24023;
	wire [16-1:0] node24024;
	wire [16-1:0] node24027;
	wire [16-1:0] node24030;
	wire [16-1:0] node24031;
	wire [16-1:0] node24034;
	wire [16-1:0] node24037;
	wire [16-1:0] node24038;
	wire [16-1:0] node24039;
	wire [16-1:0] node24042;
	wire [16-1:0] node24045;
	wire [16-1:0] node24046;
	wire [16-1:0] node24050;
	wire [16-1:0] node24051;
	wire [16-1:0] node24052;
	wire [16-1:0] node24053;
	wire [16-1:0] node24054;
	wire [16-1:0] node24057;
	wire [16-1:0] node24060;
	wire [16-1:0] node24062;
	wire [16-1:0] node24065;
	wire [16-1:0] node24066;
	wire [16-1:0] node24067;
	wire [16-1:0] node24070;
	wire [16-1:0] node24073;
	wire [16-1:0] node24075;
	wire [16-1:0] node24078;
	wire [16-1:0] node24079;
	wire [16-1:0] node24080;
	wire [16-1:0] node24081;
	wire [16-1:0] node24084;
	wire [16-1:0] node24087;
	wire [16-1:0] node24088;
	wire [16-1:0] node24091;
	wire [16-1:0] node24094;
	wire [16-1:0] node24095;
	wire [16-1:0] node24096;
	wire [16-1:0] node24100;
	wire [16-1:0] node24101;
	wire [16-1:0] node24104;
	wire [16-1:0] node24107;
	wire [16-1:0] node24108;
	wire [16-1:0] node24109;
	wire [16-1:0] node24110;
	wire [16-1:0] node24111;
	wire [16-1:0] node24112;
	wire [16-1:0] node24113;
	wire [16-1:0] node24116;
	wire [16-1:0] node24119;
	wire [16-1:0] node24120;
	wire [16-1:0] node24123;
	wire [16-1:0] node24126;
	wire [16-1:0] node24127;
	wire [16-1:0] node24128;
	wire [16-1:0] node24131;
	wire [16-1:0] node24134;
	wire [16-1:0] node24135;
	wire [16-1:0] node24138;
	wire [16-1:0] node24141;
	wire [16-1:0] node24142;
	wire [16-1:0] node24143;
	wire [16-1:0] node24144;
	wire [16-1:0] node24148;
	wire [16-1:0] node24149;
	wire [16-1:0] node24152;
	wire [16-1:0] node24155;
	wire [16-1:0] node24156;
	wire [16-1:0] node24157;
	wire [16-1:0] node24161;
	wire [16-1:0] node24162;
	wire [16-1:0] node24165;
	wire [16-1:0] node24168;
	wire [16-1:0] node24169;
	wire [16-1:0] node24170;
	wire [16-1:0] node24171;
	wire [16-1:0] node24172;
	wire [16-1:0] node24175;
	wire [16-1:0] node24178;
	wire [16-1:0] node24179;
	wire [16-1:0] node24182;
	wire [16-1:0] node24185;
	wire [16-1:0] node24186;
	wire [16-1:0] node24187;
	wire [16-1:0] node24190;
	wire [16-1:0] node24193;
	wire [16-1:0] node24195;
	wire [16-1:0] node24198;
	wire [16-1:0] node24199;
	wire [16-1:0] node24200;
	wire [16-1:0] node24202;
	wire [16-1:0] node24205;
	wire [16-1:0] node24206;
	wire [16-1:0] node24209;
	wire [16-1:0] node24212;
	wire [16-1:0] node24213;
	wire [16-1:0] node24215;
	wire [16-1:0] node24218;
	wire [16-1:0] node24219;
	wire [16-1:0] node24223;
	wire [16-1:0] node24224;
	wire [16-1:0] node24225;
	wire [16-1:0] node24226;
	wire [16-1:0] node24227;
	wire [16-1:0] node24229;
	wire [16-1:0] node24232;
	wire [16-1:0] node24233;
	wire [16-1:0] node24237;
	wire [16-1:0] node24238;
	wire [16-1:0] node24239;
	wire [16-1:0] node24242;
	wire [16-1:0] node24245;
	wire [16-1:0] node24246;
	wire [16-1:0] node24250;
	wire [16-1:0] node24251;
	wire [16-1:0] node24252;
	wire [16-1:0] node24253;
	wire [16-1:0] node24256;
	wire [16-1:0] node24259;
	wire [16-1:0] node24260;
	wire [16-1:0] node24263;
	wire [16-1:0] node24266;
	wire [16-1:0] node24267;
	wire [16-1:0] node24268;
	wire [16-1:0] node24271;
	wire [16-1:0] node24274;
	wire [16-1:0] node24276;
	wire [16-1:0] node24279;
	wire [16-1:0] node24280;
	wire [16-1:0] node24281;
	wire [16-1:0] node24282;
	wire [16-1:0] node24283;
	wire [16-1:0] node24287;
	wire [16-1:0] node24288;
	wire [16-1:0] node24291;
	wire [16-1:0] node24294;
	wire [16-1:0] node24295;
	wire [16-1:0] node24296;
	wire [16-1:0] node24299;
	wire [16-1:0] node24302;
	wire [16-1:0] node24303;
	wire [16-1:0] node24306;
	wire [16-1:0] node24309;
	wire [16-1:0] node24310;
	wire [16-1:0] node24311;
	wire [16-1:0] node24313;
	wire [16-1:0] node24316;
	wire [16-1:0] node24317;
	wire [16-1:0] node24320;
	wire [16-1:0] node24323;
	wire [16-1:0] node24324;
	wire [16-1:0] node24325;
	wire [16-1:0] node24329;
	wire [16-1:0] node24330;
	wire [16-1:0] node24333;
	wire [16-1:0] node24336;
	wire [16-1:0] node24337;
	wire [16-1:0] node24338;
	wire [16-1:0] node24339;
	wire [16-1:0] node24340;
	wire [16-1:0] node24341;
	wire [16-1:0] node24342;
	wire [16-1:0] node24343;
	wire [16-1:0] node24344;
	wire [16-1:0] node24347;
	wire [16-1:0] node24350;
	wire [16-1:0] node24351;
	wire [16-1:0] node24354;
	wire [16-1:0] node24357;
	wire [16-1:0] node24358;
	wire [16-1:0] node24359;
	wire [16-1:0] node24362;
	wire [16-1:0] node24365;
	wire [16-1:0] node24366;
	wire [16-1:0] node24370;
	wire [16-1:0] node24371;
	wire [16-1:0] node24372;
	wire [16-1:0] node24373;
	wire [16-1:0] node24376;
	wire [16-1:0] node24379;
	wire [16-1:0] node24380;
	wire [16-1:0] node24383;
	wire [16-1:0] node24386;
	wire [16-1:0] node24387;
	wire [16-1:0] node24388;
	wire [16-1:0] node24391;
	wire [16-1:0] node24394;
	wire [16-1:0] node24395;
	wire [16-1:0] node24398;
	wire [16-1:0] node24401;
	wire [16-1:0] node24402;
	wire [16-1:0] node24403;
	wire [16-1:0] node24404;
	wire [16-1:0] node24405;
	wire [16-1:0] node24408;
	wire [16-1:0] node24411;
	wire [16-1:0] node24412;
	wire [16-1:0] node24416;
	wire [16-1:0] node24417;
	wire [16-1:0] node24418;
	wire [16-1:0] node24421;
	wire [16-1:0] node24424;
	wire [16-1:0] node24425;
	wire [16-1:0] node24428;
	wire [16-1:0] node24431;
	wire [16-1:0] node24432;
	wire [16-1:0] node24433;
	wire [16-1:0] node24434;
	wire [16-1:0] node24437;
	wire [16-1:0] node24440;
	wire [16-1:0] node24441;
	wire [16-1:0] node24444;
	wire [16-1:0] node24447;
	wire [16-1:0] node24448;
	wire [16-1:0] node24449;
	wire [16-1:0] node24452;
	wire [16-1:0] node24455;
	wire [16-1:0] node24457;
	wire [16-1:0] node24460;
	wire [16-1:0] node24461;
	wire [16-1:0] node24462;
	wire [16-1:0] node24463;
	wire [16-1:0] node24464;
	wire [16-1:0] node24465;
	wire [16-1:0] node24468;
	wire [16-1:0] node24471;
	wire [16-1:0] node24472;
	wire [16-1:0] node24475;
	wire [16-1:0] node24478;
	wire [16-1:0] node24479;
	wire [16-1:0] node24481;
	wire [16-1:0] node24484;
	wire [16-1:0] node24485;
	wire [16-1:0] node24488;
	wire [16-1:0] node24491;
	wire [16-1:0] node24492;
	wire [16-1:0] node24494;
	wire [16-1:0] node24495;
	wire [16-1:0] node24498;
	wire [16-1:0] node24501;
	wire [16-1:0] node24502;
	wire [16-1:0] node24503;
	wire [16-1:0] node24506;
	wire [16-1:0] node24509;
	wire [16-1:0] node24510;
	wire [16-1:0] node24513;
	wire [16-1:0] node24516;
	wire [16-1:0] node24517;
	wire [16-1:0] node24518;
	wire [16-1:0] node24519;
	wire [16-1:0] node24520;
	wire [16-1:0] node24523;
	wire [16-1:0] node24526;
	wire [16-1:0] node24527;
	wire [16-1:0] node24530;
	wire [16-1:0] node24533;
	wire [16-1:0] node24534;
	wire [16-1:0] node24535;
	wire [16-1:0] node24538;
	wire [16-1:0] node24541;
	wire [16-1:0] node24542;
	wire [16-1:0] node24545;
	wire [16-1:0] node24548;
	wire [16-1:0] node24549;
	wire [16-1:0] node24550;
	wire [16-1:0] node24551;
	wire [16-1:0] node24554;
	wire [16-1:0] node24557;
	wire [16-1:0] node24558;
	wire [16-1:0] node24561;
	wire [16-1:0] node24564;
	wire [16-1:0] node24565;
	wire [16-1:0] node24566;
	wire [16-1:0] node24569;
	wire [16-1:0] node24572;
	wire [16-1:0] node24573;
	wire [16-1:0] node24576;
	wire [16-1:0] node24579;
	wire [16-1:0] node24580;
	wire [16-1:0] node24581;
	wire [16-1:0] node24582;
	wire [16-1:0] node24583;
	wire [16-1:0] node24584;
	wire [16-1:0] node24585;
	wire [16-1:0] node24588;
	wire [16-1:0] node24591;
	wire [16-1:0] node24592;
	wire [16-1:0] node24595;
	wire [16-1:0] node24598;
	wire [16-1:0] node24599;
	wire [16-1:0] node24600;
	wire [16-1:0] node24603;
	wire [16-1:0] node24606;
	wire [16-1:0] node24607;
	wire [16-1:0] node24610;
	wire [16-1:0] node24613;
	wire [16-1:0] node24614;
	wire [16-1:0] node24615;
	wire [16-1:0] node24616;
	wire [16-1:0] node24619;
	wire [16-1:0] node24622;
	wire [16-1:0] node24623;
	wire [16-1:0] node24626;
	wire [16-1:0] node24629;
	wire [16-1:0] node24630;
	wire [16-1:0] node24631;
	wire [16-1:0] node24634;
	wire [16-1:0] node24637;
	wire [16-1:0] node24639;
	wire [16-1:0] node24642;
	wire [16-1:0] node24643;
	wire [16-1:0] node24644;
	wire [16-1:0] node24645;
	wire [16-1:0] node24646;
	wire [16-1:0] node24649;
	wire [16-1:0] node24652;
	wire [16-1:0] node24653;
	wire [16-1:0] node24656;
	wire [16-1:0] node24659;
	wire [16-1:0] node24660;
	wire [16-1:0] node24661;
	wire [16-1:0] node24664;
	wire [16-1:0] node24667;
	wire [16-1:0] node24668;
	wire [16-1:0] node24671;
	wire [16-1:0] node24674;
	wire [16-1:0] node24675;
	wire [16-1:0] node24676;
	wire [16-1:0] node24677;
	wire [16-1:0] node24680;
	wire [16-1:0] node24683;
	wire [16-1:0] node24684;
	wire [16-1:0] node24687;
	wire [16-1:0] node24690;
	wire [16-1:0] node24691;
	wire [16-1:0] node24692;
	wire [16-1:0] node24695;
	wire [16-1:0] node24698;
	wire [16-1:0] node24699;
	wire [16-1:0] node24702;
	wire [16-1:0] node24705;
	wire [16-1:0] node24706;
	wire [16-1:0] node24707;
	wire [16-1:0] node24708;
	wire [16-1:0] node24709;
	wire [16-1:0] node24710;
	wire [16-1:0] node24713;
	wire [16-1:0] node24716;
	wire [16-1:0] node24717;
	wire [16-1:0] node24720;
	wire [16-1:0] node24723;
	wire [16-1:0] node24724;
	wire [16-1:0] node24726;
	wire [16-1:0] node24729;
	wire [16-1:0] node24730;
	wire [16-1:0] node24733;
	wire [16-1:0] node24736;
	wire [16-1:0] node24737;
	wire [16-1:0] node24738;
	wire [16-1:0] node24739;
	wire [16-1:0] node24742;
	wire [16-1:0] node24745;
	wire [16-1:0] node24746;
	wire [16-1:0] node24749;
	wire [16-1:0] node24752;
	wire [16-1:0] node24753;
	wire [16-1:0] node24754;
	wire [16-1:0] node24757;
	wire [16-1:0] node24760;
	wire [16-1:0] node24761;
	wire [16-1:0] node24764;
	wire [16-1:0] node24767;
	wire [16-1:0] node24768;
	wire [16-1:0] node24769;
	wire [16-1:0] node24770;
	wire [16-1:0] node24771;
	wire [16-1:0] node24774;
	wire [16-1:0] node24777;
	wire [16-1:0] node24778;
	wire [16-1:0] node24782;
	wire [16-1:0] node24783;
	wire [16-1:0] node24784;
	wire [16-1:0] node24787;
	wire [16-1:0] node24790;
	wire [16-1:0] node24791;
	wire [16-1:0] node24794;
	wire [16-1:0] node24797;
	wire [16-1:0] node24798;
	wire [16-1:0] node24799;
	wire [16-1:0] node24800;
	wire [16-1:0] node24803;
	wire [16-1:0] node24806;
	wire [16-1:0] node24807;
	wire [16-1:0] node24810;
	wire [16-1:0] node24813;
	wire [16-1:0] node24814;
	wire [16-1:0] node24816;
	wire [16-1:0] node24819;
	wire [16-1:0] node24821;
	wire [16-1:0] node24824;
	wire [16-1:0] node24825;
	wire [16-1:0] node24826;
	wire [16-1:0] node24827;
	wire [16-1:0] node24828;
	wire [16-1:0] node24829;
	wire [16-1:0] node24830;
	wire [16-1:0] node24831;
	wire [16-1:0] node24835;
	wire [16-1:0] node24836;
	wire [16-1:0] node24840;
	wire [16-1:0] node24841;
	wire [16-1:0] node24842;
	wire [16-1:0] node24845;
	wire [16-1:0] node24848;
	wire [16-1:0] node24849;
	wire [16-1:0] node24853;
	wire [16-1:0] node24854;
	wire [16-1:0] node24855;
	wire [16-1:0] node24856;
	wire [16-1:0] node24859;
	wire [16-1:0] node24862;
	wire [16-1:0] node24863;
	wire [16-1:0] node24866;
	wire [16-1:0] node24869;
	wire [16-1:0] node24870;
	wire [16-1:0] node24871;
	wire [16-1:0] node24874;
	wire [16-1:0] node24877;
	wire [16-1:0] node24878;
	wire [16-1:0] node24882;
	wire [16-1:0] node24883;
	wire [16-1:0] node24884;
	wire [16-1:0] node24885;
	wire [16-1:0] node24887;
	wire [16-1:0] node24890;
	wire [16-1:0] node24891;
	wire [16-1:0] node24894;
	wire [16-1:0] node24897;
	wire [16-1:0] node24898;
	wire [16-1:0] node24899;
	wire [16-1:0] node24902;
	wire [16-1:0] node24905;
	wire [16-1:0] node24907;
	wire [16-1:0] node24910;
	wire [16-1:0] node24911;
	wire [16-1:0] node24912;
	wire [16-1:0] node24913;
	wire [16-1:0] node24916;
	wire [16-1:0] node24919;
	wire [16-1:0] node24920;
	wire [16-1:0] node24923;
	wire [16-1:0] node24926;
	wire [16-1:0] node24927;
	wire [16-1:0] node24928;
	wire [16-1:0] node24932;
	wire [16-1:0] node24933;
	wire [16-1:0] node24937;
	wire [16-1:0] node24938;
	wire [16-1:0] node24939;
	wire [16-1:0] node24940;
	wire [16-1:0] node24941;
	wire [16-1:0] node24942;
	wire [16-1:0] node24945;
	wire [16-1:0] node24948;
	wire [16-1:0] node24949;
	wire [16-1:0] node24952;
	wire [16-1:0] node24955;
	wire [16-1:0] node24956;
	wire [16-1:0] node24957;
	wire [16-1:0] node24960;
	wire [16-1:0] node24963;
	wire [16-1:0] node24964;
	wire [16-1:0] node24967;
	wire [16-1:0] node24970;
	wire [16-1:0] node24971;
	wire [16-1:0] node24972;
	wire [16-1:0] node24973;
	wire [16-1:0] node24976;
	wire [16-1:0] node24979;
	wire [16-1:0] node24980;
	wire [16-1:0] node24983;
	wire [16-1:0] node24986;
	wire [16-1:0] node24987;
	wire [16-1:0] node24988;
	wire [16-1:0] node24991;
	wire [16-1:0] node24994;
	wire [16-1:0] node24995;
	wire [16-1:0] node24998;
	wire [16-1:0] node25001;
	wire [16-1:0] node25002;
	wire [16-1:0] node25003;
	wire [16-1:0] node25004;
	wire [16-1:0] node25007;
	wire [16-1:0] node25008;
	wire [16-1:0] node25011;
	wire [16-1:0] node25014;
	wire [16-1:0] node25015;
	wire [16-1:0] node25017;
	wire [16-1:0] node25020;
	wire [16-1:0] node25021;
	wire [16-1:0] node25024;
	wire [16-1:0] node25027;
	wire [16-1:0] node25028;
	wire [16-1:0] node25029;
	wire [16-1:0] node25031;
	wire [16-1:0] node25034;
	wire [16-1:0] node25035;
	wire [16-1:0] node25038;
	wire [16-1:0] node25041;
	wire [16-1:0] node25042;
	wire [16-1:0] node25043;
	wire [16-1:0] node25046;
	wire [16-1:0] node25049;
	wire [16-1:0] node25050;
	wire [16-1:0] node25054;
	wire [16-1:0] node25055;
	wire [16-1:0] node25056;
	wire [16-1:0] node25057;
	wire [16-1:0] node25058;
	wire [16-1:0] node25059;
	wire [16-1:0] node25060;
	wire [16-1:0] node25064;
	wire [16-1:0] node25065;
	wire [16-1:0] node25068;
	wire [16-1:0] node25071;
	wire [16-1:0] node25072;
	wire [16-1:0] node25073;
	wire [16-1:0] node25076;
	wire [16-1:0] node25079;
	wire [16-1:0] node25080;
	wire [16-1:0] node25084;
	wire [16-1:0] node25085;
	wire [16-1:0] node25086;
	wire [16-1:0] node25087;
	wire [16-1:0] node25090;
	wire [16-1:0] node25093;
	wire [16-1:0] node25094;
	wire [16-1:0] node25097;
	wire [16-1:0] node25100;
	wire [16-1:0] node25101;
	wire [16-1:0] node25102;
	wire [16-1:0] node25105;
	wire [16-1:0] node25108;
	wire [16-1:0] node25109;
	wire [16-1:0] node25112;
	wire [16-1:0] node25115;
	wire [16-1:0] node25116;
	wire [16-1:0] node25117;
	wire [16-1:0] node25118;
	wire [16-1:0] node25119;
	wire [16-1:0] node25122;
	wire [16-1:0] node25125;
	wire [16-1:0] node25126;
	wire [16-1:0] node25129;
	wire [16-1:0] node25132;
	wire [16-1:0] node25133;
	wire [16-1:0] node25134;
	wire [16-1:0] node25138;
	wire [16-1:0] node25139;
	wire [16-1:0] node25142;
	wire [16-1:0] node25145;
	wire [16-1:0] node25146;
	wire [16-1:0] node25147;
	wire [16-1:0] node25148;
	wire [16-1:0] node25151;
	wire [16-1:0] node25154;
	wire [16-1:0] node25155;
	wire [16-1:0] node25158;
	wire [16-1:0] node25161;
	wire [16-1:0] node25162;
	wire [16-1:0] node25163;
	wire [16-1:0] node25166;
	wire [16-1:0] node25169;
	wire [16-1:0] node25171;
	wire [16-1:0] node25174;
	wire [16-1:0] node25175;
	wire [16-1:0] node25176;
	wire [16-1:0] node25177;
	wire [16-1:0] node25178;
	wire [16-1:0] node25179;
	wire [16-1:0] node25182;
	wire [16-1:0] node25185;
	wire [16-1:0] node25186;
	wire [16-1:0] node25189;
	wire [16-1:0] node25192;
	wire [16-1:0] node25193;
	wire [16-1:0] node25194;
	wire [16-1:0] node25197;
	wire [16-1:0] node25200;
	wire [16-1:0] node25201;
	wire [16-1:0] node25204;
	wire [16-1:0] node25207;
	wire [16-1:0] node25208;
	wire [16-1:0] node25209;
	wire [16-1:0] node25211;
	wire [16-1:0] node25214;
	wire [16-1:0] node25215;
	wire [16-1:0] node25218;
	wire [16-1:0] node25221;
	wire [16-1:0] node25222;
	wire [16-1:0] node25223;
	wire [16-1:0] node25226;
	wire [16-1:0] node25229;
	wire [16-1:0] node25230;
	wire [16-1:0] node25233;
	wire [16-1:0] node25236;
	wire [16-1:0] node25237;
	wire [16-1:0] node25238;
	wire [16-1:0] node25239;
	wire [16-1:0] node25240;
	wire [16-1:0] node25243;
	wire [16-1:0] node25246;
	wire [16-1:0] node25247;
	wire [16-1:0] node25251;
	wire [16-1:0] node25252;
	wire [16-1:0] node25254;
	wire [16-1:0] node25257;
	wire [16-1:0] node25258;
	wire [16-1:0] node25262;
	wire [16-1:0] node25263;
	wire [16-1:0] node25264;
	wire [16-1:0] node25265;
	wire [16-1:0] node25268;
	wire [16-1:0] node25271;
	wire [16-1:0] node25272;
	wire [16-1:0] node25275;
	wire [16-1:0] node25278;
	wire [16-1:0] node25279;
	wire [16-1:0] node25280;
	wire [16-1:0] node25283;
	wire [16-1:0] node25286;
	wire [16-1:0] node25287;
	wire [16-1:0] node25290;
	wire [16-1:0] node25293;
	wire [16-1:0] node25294;
	wire [16-1:0] node25295;
	wire [16-1:0] node25296;
	wire [16-1:0] node25297;
	wire [16-1:0] node25298;
	wire [16-1:0] node25299;
	wire [16-1:0] node25300;
	wire [16-1:0] node25301;
	wire [16-1:0] node25302;
	wire [16-1:0] node25305;
	wire [16-1:0] node25308;
	wire [16-1:0] node25309;
	wire [16-1:0] node25312;
	wire [16-1:0] node25315;
	wire [16-1:0] node25316;
	wire [16-1:0] node25317;
	wire [16-1:0] node25321;
	wire [16-1:0] node25322;
	wire [16-1:0] node25326;
	wire [16-1:0] node25327;
	wire [16-1:0] node25328;
	wire [16-1:0] node25330;
	wire [16-1:0] node25333;
	wire [16-1:0] node25334;
	wire [16-1:0] node25337;
	wire [16-1:0] node25340;
	wire [16-1:0] node25341;
	wire [16-1:0] node25342;
	wire [16-1:0] node25345;
	wire [16-1:0] node25348;
	wire [16-1:0] node25349;
	wire [16-1:0] node25352;
	wire [16-1:0] node25355;
	wire [16-1:0] node25356;
	wire [16-1:0] node25357;
	wire [16-1:0] node25358;
	wire [16-1:0] node25359;
	wire [16-1:0] node25362;
	wire [16-1:0] node25365;
	wire [16-1:0] node25366;
	wire [16-1:0] node25369;
	wire [16-1:0] node25372;
	wire [16-1:0] node25373;
	wire [16-1:0] node25374;
	wire [16-1:0] node25377;
	wire [16-1:0] node25380;
	wire [16-1:0] node25382;
	wire [16-1:0] node25385;
	wire [16-1:0] node25386;
	wire [16-1:0] node25387;
	wire [16-1:0] node25388;
	wire [16-1:0] node25391;
	wire [16-1:0] node25394;
	wire [16-1:0] node25395;
	wire [16-1:0] node25398;
	wire [16-1:0] node25401;
	wire [16-1:0] node25402;
	wire [16-1:0] node25403;
	wire [16-1:0] node25406;
	wire [16-1:0] node25409;
	wire [16-1:0] node25410;
	wire [16-1:0] node25414;
	wire [16-1:0] node25415;
	wire [16-1:0] node25416;
	wire [16-1:0] node25417;
	wire [16-1:0] node25418;
	wire [16-1:0] node25419;
	wire [16-1:0] node25422;
	wire [16-1:0] node25425;
	wire [16-1:0] node25426;
	wire [16-1:0] node25430;
	wire [16-1:0] node25431;
	wire [16-1:0] node25432;
	wire [16-1:0] node25435;
	wire [16-1:0] node25438;
	wire [16-1:0] node25439;
	wire [16-1:0] node25442;
	wire [16-1:0] node25445;
	wire [16-1:0] node25446;
	wire [16-1:0] node25447;
	wire [16-1:0] node25448;
	wire [16-1:0] node25451;
	wire [16-1:0] node25454;
	wire [16-1:0] node25455;
	wire [16-1:0] node25458;
	wire [16-1:0] node25461;
	wire [16-1:0] node25462;
	wire [16-1:0] node25463;
	wire [16-1:0] node25466;
	wire [16-1:0] node25469;
	wire [16-1:0] node25470;
	wire [16-1:0] node25473;
	wire [16-1:0] node25476;
	wire [16-1:0] node25477;
	wire [16-1:0] node25478;
	wire [16-1:0] node25479;
	wire [16-1:0] node25480;
	wire [16-1:0] node25483;
	wire [16-1:0] node25486;
	wire [16-1:0] node25487;
	wire [16-1:0] node25490;
	wire [16-1:0] node25493;
	wire [16-1:0] node25494;
	wire [16-1:0] node25495;
	wire [16-1:0] node25498;
	wire [16-1:0] node25501;
	wire [16-1:0] node25502;
	wire [16-1:0] node25505;
	wire [16-1:0] node25508;
	wire [16-1:0] node25509;
	wire [16-1:0] node25510;
	wire [16-1:0] node25512;
	wire [16-1:0] node25515;
	wire [16-1:0] node25516;
	wire [16-1:0] node25520;
	wire [16-1:0] node25521;
	wire [16-1:0] node25522;
	wire [16-1:0] node25525;
	wire [16-1:0] node25528;
	wire [16-1:0] node25529;
	wire [16-1:0] node25532;
	wire [16-1:0] node25535;
	wire [16-1:0] node25536;
	wire [16-1:0] node25537;
	wire [16-1:0] node25538;
	wire [16-1:0] node25539;
	wire [16-1:0] node25540;
	wire [16-1:0] node25541;
	wire [16-1:0] node25544;
	wire [16-1:0] node25547;
	wire [16-1:0] node25548;
	wire [16-1:0] node25552;
	wire [16-1:0] node25553;
	wire [16-1:0] node25554;
	wire [16-1:0] node25558;
	wire [16-1:0] node25559;
	wire [16-1:0] node25562;
	wire [16-1:0] node25565;
	wire [16-1:0] node25566;
	wire [16-1:0] node25567;
	wire [16-1:0] node25568;
	wire [16-1:0] node25571;
	wire [16-1:0] node25574;
	wire [16-1:0] node25575;
	wire [16-1:0] node25578;
	wire [16-1:0] node25581;
	wire [16-1:0] node25582;
	wire [16-1:0] node25583;
	wire [16-1:0] node25586;
	wire [16-1:0] node25589;
	wire [16-1:0] node25590;
	wire [16-1:0] node25593;
	wire [16-1:0] node25596;
	wire [16-1:0] node25597;
	wire [16-1:0] node25598;
	wire [16-1:0] node25599;
	wire [16-1:0] node25600;
	wire [16-1:0] node25603;
	wire [16-1:0] node25606;
	wire [16-1:0] node25607;
	wire [16-1:0] node25610;
	wire [16-1:0] node25613;
	wire [16-1:0] node25614;
	wire [16-1:0] node25615;
	wire [16-1:0] node25619;
	wire [16-1:0] node25620;
	wire [16-1:0] node25623;
	wire [16-1:0] node25626;
	wire [16-1:0] node25627;
	wire [16-1:0] node25629;
	wire [16-1:0] node25630;
	wire [16-1:0] node25633;
	wire [16-1:0] node25636;
	wire [16-1:0] node25637;
	wire [16-1:0] node25638;
	wire [16-1:0] node25641;
	wire [16-1:0] node25644;
	wire [16-1:0] node25645;
	wire [16-1:0] node25648;
	wire [16-1:0] node25651;
	wire [16-1:0] node25652;
	wire [16-1:0] node25653;
	wire [16-1:0] node25654;
	wire [16-1:0] node25655;
	wire [16-1:0] node25656;
	wire [16-1:0] node25659;
	wire [16-1:0] node25662;
	wire [16-1:0] node25664;
	wire [16-1:0] node25667;
	wire [16-1:0] node25668;
	wire [16-1:0] node25669;
	wire [16-1:0] node25672;
	wire [16-1:0] node25675;
	wire [16-1:0] node25676;
	wire [16-1:0] node25679;
	wire [16-1:0] node25682;
	wire [16-1:0] node25683;
	wire [16-1:0] node25684;
	wire [16-1:0] node25685;
	wire [16-1:0] node25688;
	wire [16-1:0] node25691;
	wire [16-1:0] node25692;
	wire [16-1:0] node25695;
	wire [16-1:0] node25698;
	wire [16-1:0] node25699;
	wire [16-1:0] node25700;
	wire [16-1:0] node25703;
	wire [16-1:0] node25706;
	wire [16-1:0] node25707;
	wire [16-1:0] node25710;
	wire [16-1:0] node25713;
	wire [16-1:0] node25714;
	wire [16-1:0] node25715;
	wire [16-1:0] node25716;
	wire [16-1:0] node25717;
	wire [16-1:0] node25720;
	wire [16-1:0] node25723;
	wire [16-1:0] node25724;
	wire [16-1:0] node25727;
	wire [16-1:0] node25730;
	wire [16-1:0] node25731;
	wire [16-1:0] node25732;
	wire [16-1:0] node25735;
	wire [16-1:0] node25738;
	wire [16-1:0] node25739;
	wire [16-1:0] node25742;
	wire [16-1:0] node25745;
	wire [16-1:0] node25746;
	wire [16-1:0] node25747;
	wire [16-1:0] node25748;
	wire [16-1:0] node25751;
	wire [16-1:0] node25754;
	wire [16-1:0] node25755;
	wire [16-1:0] node25758;
	wire [16-1:0] node25761;
	wire [16-1:0] node25762;
	wire [16-1:0] node25763;
	wire [16-1:0] node25766;
	wire [16-1:0] node25769;
	wire [16-1:0] node25770;
	wire [16-1:0] node25773;
	wire [16-1:0] node25776;
	wire [16-1:0] node25777;
	wire [16-1:0] node25778;
	wire [16-1:0] node25779;
	wire [16-1:0] node25780;
	wire [16-1:0] node25781;
	wire [16-1:0] node25782;
	wire [16-1:0] node25783;
	wire [16-1:0] node25786;
	wire [16-1:0] node25789;
	wire [16-1:0] node25790;
	wire [16-1:0] node25793;
	wire [16-1:0] node25796;
	wire [16-1:0] node25797;
	wire [16-1:0] node25798;
	wire [16-1:0] node25801;
	wire [16-1:0] node25804;
	wire [16-1:0] node25806;
	wire [16-1:0] node25809;
	wire [16-1:0] node25810;
	wire [16-1:0] node25811;
	wire [16-1:0] node25812;
	wire [16-1:0] node25815;
	wire [16-1:0] node25818;
	wire [16-1:0] node25819;
	wire [16-1:0] node25822;
	wire [16-1:0] node25825;
	wire [16-1:0] node25827;
	wire [16-1:0] node25828;
	wire [16-1:0] node25832;
	wire [16-1:0] node25833;
	wire [16-1:0] node25834;
	wire [16-1:0] node25835;
	wire [16-1:0] node25836;
	wire [16-1:0] node25839;
	wire [16-1:0] node25842;
	wire [16-1:0] node25843;
	wire [16-1:0] node25846;
	wire [16-1:0] node25849;
	wire [16-1:0] node25850;
	wire [16-1:0] node25851;
	wire [16-1:0] node25854;
	wire [16-1:0] node25857;
	wire [16-1:0] node25858;
	wire [16-1:0] node25861;
	wire [16-1:0] node25864;
	wire [16-1:0] node25865;
	wire [16-1:0] node25866;
	wire [16-1:0] node25867;
	wire [16-1:0] node25870;
	wire [16-1:0] node25873;
	wire [16-1:0] node25874;
	wire [16-1:0] node25877;
	wire [16-1:0] node25880;
	wire [16-1:0] node25881;
	wire [16-1:0] node25882;
	wire [16-1:0] node25885;
	wire [16-1:0] node25888;
	wire [16-1:0] node25890;
	wire [16-1:0] node25893;
	wire [16-1:0] node25894;
	wire [16-1:0] node25895;
	wire [16-1:0] node25896;
	wire [16-1:0] node25897;
	wire [16-1:0] node25899;
	wire [16-1:0] node25902;
	wire [16-1:0] node25903;
	wire [16-1:0] node25906;
	wire [16-1:0] node25909;
	wire [16-1:0] node25910;
	wire [16-1:0] node25912;
	wire [16-1:0] node25915;
	wire [16-1:0] node25916;
	wire [16-1:0] node25919;
	wire [16-1:0] node25922;
	wire [16-1:0] node25923;
	wire [16-1:0] node25924;
	wire [16-1:0] node25925;
	wire [16-1:0] node25928;
	wire [16-1:0] node25931;
	wire [16-1:0] node25932;
	wire [16-1:0] node25935;
	wire [16-1:0] node25938;
	wire [16-1:0] node25939;
	wire [16-1:0] node25940;
	wire [16-1:0] node25943;
	wire [16-1:0] node25946;
	wire [16-1:0] node25947;
	wire [16-1:0] node25950;
	wire [16-1:0] node25953;
	wire [16-1:0] node25954;
	wire [16-1:0] node25955;
	wire [16-1:0] node25956;
	wire [16-1:0] node25957;
	wire [16-1:0] node25960;
	wire [16-1:0] node25963;
	wire [16-1:0] node25964;
	wire [16-1:0] node25967;
	wire [16-1:0] node25970;
	wire [16-1:0] node25971;
	wire [16-1:0] node25972;
	wire [16-1:0] node25975;
	wire [16-1:0] node25978;
	wire [16-1:0] node25979;
	wire [16-1:0] node25982;
	wire [16-1:0] node25985;
	wire [16-1:0] node25986;
	wire [16-1:0] node25987;
	wire [16-1:0] node25988;
	wire [16-1:0] node25991;
	wire [16-1:0] node25994;
	wire [16-1:0] node25995;
	wire [16-1:0] node25998;
	wire [16-1:0] node26001;
	wire [16-1:0] node26002;
	wire [16-1:0] node26003;
	wire [16-1:0] node26006;
	wire [16-1:0] node26009;
	wire [16-1:0] node26011;
	wire [16-1:0] node26014;
	wire [16-1:0] node26015;
	wire [16-1:0] node26016;
	wire [16-1:0] node26017;
	wire [16-1:0] node26018;
	wire [16-1:0] node26019;
	wire [16-1:0] node26020;
	wire [16-1:0] node26023;
	wire [16-1:0] node26026;
	wire [16-1:0] node26027;
	wire [16-1:0] node26031;
	wire [16-1:0] node26032;
	wire [16-1:0] node26033;
	wire [16-1:0] node26036;
	wire [16-1:0] node26039;
	wire [16-1:0] node26041;
	wire [16-1:0] node26044;
	wire [16-1:0] node26045;
	wire [16-1:0] node26046;
	wire [16-1:0] node26047;
	wire [16-1:0] node26050;
	wire [16-1:0] node26053;
	wire [16-1:0] node26054;
	wire [16-1:0] node26057;
	wire [16-1:0] node26060;
	wire [16-1:0] node26061;
	wire [16-1:0] node26062;
	wire [16-1:0] node26065;
	wire [16-1:0] node26068;
	wire [16-1:0] node26069;
	wire [16-1:0] node26072;
	wire [16-1:0] node26075;
	wire [16-1:0] node26076;
	wire [16-1:0] node26077;
	wire [16-1:0] node26078;
	wire [16-1:0] node26079;
	wire [16-1:0] node26082;
	wire [16-1:0] node26085;
	wire [16-1:0] node26086;
	wire [16-1:0] node26089;
	wire [16-1:0] node26092;
	wire [16-1:0] node26093;
	wire [16-1:0] node26094;
	wire [16-1:0] node26097;
	wire [16-1:0] node26100;
	wire [16-1:0] node26101;
	wire [16-1:0] node26104;
	wire [16-1:0] node26107;
	wire [16-1:0] node26108;
	wire [16-1:0] node26109;
	wire [16-1:0] node26110;
	wire [16-1:0] node26113;
	wire [16-1:0] node26116;
	wire [16-1:0] node26117;
	wire [16-1:0] node26120;
	wire [16-1:0] node26123;
	wire [16-1:0] node26124;
	wire [16-1:0] node26126;
	wire [16-1:0] node26129;
	wire [16-1:0] node26130;
	wire [16-1:0] node26134;
	wire [16-1:0] node26135;
	wire [16-1:0] node26136;
	wire [16-1:0] node26137;
	wire [16-1:0] node26138;
	wire [16-1:0] node26139;
	wire [16-1:0] node26142;
	wire [16-1:0] node26145;
	wire [16-1:0] node26147;
	wire [16-1:0] node26150;
	wire [16-1:0] node26151;
	wire [16-1:0] node26152;
	wire [16-1:0] node26155;
	wire [16-1:0] node26158;
	wire [16-1:0] node26159;
	wire [16-1:0] node26162;
	wire [16-1:0] node26165;
	wire [16-1:0] node26166;
	wire [16-1:0] node26167;
	wire [16-1:0] node26168;
	wire [16-1:0] node26172;
	wire [16-1:0] node26173;
	wire [16-1:0] node26176;
	wire [16-1:0] node26179;
	wire [16-1:0] node26180;
	wire [16-1:0] node26181;
	wire [16-1:0] node26184;
	wire [16-1:0] node26187;
	wire [16-1:0] node26188;
	wire [16-1:0] node26191;
	wire [16-1:0] node26194;
	wire [16-1:0] node26195;
	wire [16-1:0] node26196;
	wire [16-1:0] node26197;
	wire [16-1:0] node26198;
	wire [16-1:0] node26201;
	wire [16-1:0] node26204;
	wire [16-1:0] node26205;
	wire [16-1:0] node26208;
	wire [16-1:0] node26211;
	wire [16-1:0] node26212;
	wire [16-1:0] node26213;
	wire [16-1:0] node26216;
	wire [16-1:0] node26219;
	wire [16-1:0] node26220;
	wire [16-1:0] node26223;
	wire [16-1:0] node26226;
	wire [16-1:0] node26227;
	wire [16-1:0] node26228;
	wire [16-1:0] node26229;
	wire [16-1:0] node26232;
	wire [16-1:0] node26235;
	wire [16-1:0] node26237;
	wire [16-1:0] node26240;
	wire [16-1:0] node26241;
	wire [16-1:0] node26243;
	wire [16-1:0] node26246;
	wire [16-1:0] node26247;
	wire [16-1:0] node26250;
	wire [16-1:0] node26253;
	wire [16-1:0] node26254;
	wire [16-1:0] node26255;
	wire [16-1:0] node26256;
	wire [16-1:0] node26257;
	wire [16-1:0] node26258;
	wire [16-1:0] node26259;
	wire [16-1:0] node26260;
	wire [16-1:0] node26261;
	wire [16-1:0] node26264;
	wire [16-1:0] node26267;
	wire [16-1:0] node26268;
	wire [16-1:0] node26272;
	wire [16-1:0] node26273;
	wire [16-1:0] node26274;
	wire [16-1:0] node26277;
	wire [16-1:0] node26280;
	wire [16-1:0] node26281;
	wire [16-1:0] node26284;
	wire [16-1:0] node26287;
	wire [16-1:0] node26288;
	wire [16-1:0] node26289;
	wire [16-1:0] node26290;
	wire [16-1:0] node26293;
	wire [16-1:0] node26296;
	wire [16-1:0] node26297;
	wire [16-1:0] node26301;
	wire [16-1:0] node26302;
	wire [16-1:0] node26303;
	wire [16-1:0] node26306;
	wire [16-1:0] node26309;
	wire [16-1:0] node26310;
	wire [16-1:0] node26313;
	wire [16-1:0] node26316;
	wire [16-1:0] node26317;
	wire [16-1:0] node26318;
	wire [16-1:0] node26319;
	wire [16-1:0] node26320;
	wire [16-1:0] node26323;
	wire [16-1:0] node26326;
	wire [16-1:0] node26327;
	wire [16-1:0] node26330;
	wire [16-1:0] node26333;
	wire [16-1:0] node26334;
	wire [16-1:0] node26335;
	wire [16-1:0] node26338;
	wire [16-1:0] node26342;
	wire [16-1:0] node26343;
	wire [16-1:0] node26344;
	wire [16-1:0] node26346;
	wire [16-1:0] node26349;
	wire [16-1:0] node26350;
	wire [16-1:0] node26353;
	wire [16-1:0] node26356;
	wire [16-1:0] node26357;
	wire [16-1:0] node26358;
	wire [16-1:0] node26362;
	wire [16-1:0] node26363;
	wire [16-1:0] node26366;
	wire [16-1:0] node26369;
	wire [16-1:0] node26370;
	wire [16-1:0] node26371;
	wire [16-1:0] node26372;
	wire [16-1:0] node26373;
	wire [16-1:0] node26374;
	wire [16-1:0] node26377;
	wire [16-1:0] node26380;
	wire [16-1:0] node26381;
	wire [16-1:0] node26384;
	wire [16-1:0] node26387;
	wire [16-1:0] node26388;
	wire [16-1:0] node26389;
	wire [16-1:0] node26392;
	wire [16-1:0] node26395;
	wire [16-1:0] node26396;
	wire [16-1:0] node26400;
	wire [16-1:0] node26401;
	wire [16-1:0] node26402;
	wire [16-1:0] node26403;
	wire [16-1:0] node26406;
	wire [16-1:0] node26409;
	wire [16-1:0] node26410;
	wire [16-1:0] node26413;
	wire [16-1:0] node26416;
	wire [16-1:0] node26417;
	wire [16-1:0] node26418;
	wire [16-1:0] node26421;
	wire [16-1:0] node26424;
	wire [16-1:0] node26425;
	wire [16-1:0] node26428;
	wire [16-1:0] node26431;
	wire [16-1:0] node26432;
	wire [16-1:0] node26433;
	wire [16-1:0] node26434;
	wire [16-1:0] node26435;
	wire [16-1:0] node26438;
	wire [16-1:0] node26441;
	wire [16-1:0] node26442;
	wire [16-1:0] node26446;
	wire [16-1:0] node26447;
	wire [16-1:0] node26449;
	wire [16-1:0] node26452;
	wire [16-1:0] node26453;
	wire [16-1:0] node26457;
	wire [16-1:0] node26458;
	wire [16-1:0] node26459;
	wire [16-1:0] node26460;
	wire [16-1:0] node26464;
	wire [16-1:0] node26465;
	wire [16-1:0] node26468;
	wire [16-1:0] node26471;
	wire [16-1:0] node26472;
	wire [16-1:0] node26473;
	wire [16-1:0] node26476;
	wire [16-1:0] node26479;
	wire [16-1:0] node26480;
	wire [16-1:0] node26483;
	wire [16-1:0] node26486;
	wire [16-1:0] node26487;
	wire [16-1:0] node26488;
	wire [16-1:0] node26489;
	wire [16-1:0] node26490;
	wire [16-1:0] node26491;
	wire [16-1:0] node26492;
	wire [16-1:0] node26495;
	wire [16-1:0] node26498;
	wire [16-1:0] node26499;
	wire [16-1:0] node26502;
	wire [16-1:0] node26505;
	wire [16-1:0] node26506;
	wire [16-1:0] node26507;
	wire [16-1:0] node26510;
	wire [16-1:0] node26513;
	wire [16-1:0] node26514;
	wire [16-1:0] node26517;
	wire [16-1:0] node26520;
	wire [16-1:0] node26521;
	wire [16-1:0] node26522;
	wire [16-1:0] node26523;
	wire [16-1:0] node26526;
	wire [16-1:0] node26529;
	wire [16-1:0] node26530;
	wire [16-1:0] node26534;
	wire [16-1:0] node26535;
	wire [16-1:0] node26536;
	wire [16-1:0] node26539;
	wire [16-1:0] node26542;
	wire [16-1:0] node26543;
	wire [16-1:0] node26546;
	wire [16-1:0] node26549;
	wire [16-1:0] node26550;
	wire [16-1:0] node26551;
	wire [16-1:0] node26552;
	wire [16-1:0] node26553;
	wire [16-1:0] node26557;
	wire [16-1:0] node26558;
	wire [16-1:0] node26561;
	wire [16-1:0] node26564;
	wire [16-1:0] node26565;
	wire [16-1:0] node26566;
	wire [16-1:0] node26569;
	wire [16-1:0] node26572;
	wire [16-1:0] node26573;
	wire [16-1:0] node26576;
	wire [16-1:0] node26579;
	wire [16-1:0] node26580;
	wire [16-1:0] node26581;
	wire [16-1:0] node26582;
	wire [16-1:0] node26585;
	wire [16-1:0] node26588;
	wire [16-1:0] node26589;
	wire [16-1:0] node26593;
	wire [16-1:0] node26594;
	wire [16-1:0] node26595;
	wire [16-1:0] node26598;
	wire [16-1:0] node26601;
	wire [16-1:0] node26603;
	wire [16-1:0] node26606;
	wire [16-1:0] node26607;
	wire [16-1:0] node26608;
	wire [16-1:0] node26609;
	wire [16-1:0] node26610;
	wire [16-1:0] node26611;
	wire [16-1:0] node26614;
	wire [16-1:0] node26617;
	wire [16-1:0] node26618;
	wire [16-1:0] node26621;
	wire [16-1:0] node26624;
	wire [16-1:0] node26625;
	wire [16-1:0] node26626;
	wire [16-1:0] node26629;
	wire [16-1:0] node26632;
	wire [16-1:0] node26633;
	wire [16-1:0] node26637;
	wire [16-1:0] node26638;
	wire [16-1:0] node26639;
	wire [16-1:0] node26640;
	wire [16-1:0] node26644;
	wire [16-1:0] node26645;
	wire [16-1:0] node26648;
	wire [16-1:0] node26651;
	wire [16-1:0] node26652;
	wire [16-1:0] node26653;
	wire [16-1:0] node26656;
	wire [16-1:0] node26659;
	wire [16-1:0] node26660;
	wire [16-1:0] node26663;
	wire [16-1:0] node26666;
	wire [16-1:0] node26667;
	wire [16-1:0] node26668;
	wire [16-1:0] node26669;
	wire [16-1:0] node26670;
	wire [16-1:0] node26674;
	wire [16-1:0] node26675;
	wire [16-1:0] node26678;
	wire [16-1:0] node26681;
	wire [16-1:0] node26682;
	wire [16-1:0] node26683;
	wire [16-1:0] node26686;
	wire [16-1:0] node26689;
	wire [16-1:0] node26690;
	wire [16-1:0] node26693;
	wire [16-1:0] node26696;
	wire [16-1:0] node26697;
	wire [16-1:0] node26698;
	wire [16-1:0] node26699;
	wire [16-1:0] node26702;
	wire [16-1:0] node26705;
	wire [16-1:0] node26706;
	wire [16-1:0] node26709;
	wire [16-1:0] node26712;
	wire [16-1:0] node26713;
	wire [16-1:0] node26714;
	wire [16-1:0] node26717;
	wire [16-1:0] node26720;
	wire [16-1:0] node26721;
	wire [16-1:0] node26724;
	wire [16-1:0] node26727;
	wire [16-1:0] node26728;
	wire [16-1:0] node26729;
	wire [16-1:0] node26730;
	wire [16-1:0] node26731;
	wire [16-1:0] node26732;
	wire [16-1:0] node26733;
	wire [16-1:0] node26734;
	wire [16-1:0] node26737;
	wire [16-1:0] node26740;
	wire [16-1:0] node26741;
	wire [16-1:0] node26744;
	wire [16-1:0] node26747;
	wire [16-1:0] node26748;
	wire [16-1:0] node26749;
	wire [16-1:0] node26752;
	wire [16-1:0] node26755;
	wire [16-1:0] node26756;
	wire [16-1:0] node26759;
	wire [16-1:0] node26762;
	wire [16-1:0] node26763;
	wire [16-1:0] node26764;
	wire [16-1:0] node26765;
	wire [16-1:0] node26768;
	wire [16-1:0] node26771;
	wire [16-1:0] node26772;
	wire [16-1:0] node26776;
	wire [16-1:0] node26777;
	wire [16-1:0] node26778;
	wire [16-1:0] node26781;
	wire [16-1:0] node26784;
	wire [16-1:0] node26785;
	wire [16-1:0] node26788;
	wire [16-1:0] node26791;
	wire [16-1:0] node26792;
	wire [16-1:0] node26793;
	wire [16-1:0] node26794;
	wire [16-1:0] node26795;
	wire [16-1:0] node26798;
	wire [16-1:0] node26801;
	wire [16-1:0] node26802;
	wire [16-1:0] node26805;
	wire [16-1:0] node26808;
	wire [16-1:0] node26809;
	wire [16-1:0] node26811;
	wire [16-1:0] node26814;
	wire [16-1:0] node26815;
	wire [16-1:0] node26818;
	wire [16-1:0] node26821;
	wire [16-1:0] node26822;
	wire [16-1:0] node26823;
	wire [16-1:0] node26824;
	wire [16-1:0] node26827;
	wire [16-1:0] node26830;
	wire [16-1:0] node26831;
	wire [16-1:0] node26834;
	wire [16-1:0] node26837;
	wire [16-1:0] node26838;
	wire [16-1:0] node26839;
	wire [16-1:0] node26842;
	wire [16-1:0] node26845;
	wire [16-1:0] node26846;
	wire [16-1:0] node26849;
	wire [16-1:0] node26852;
	wire [16-1:0] node26853;
	wire [16-1:0] node26854;
	wire [16-1:0] node26855;
	wire [16-1:0] node26856;
	wire [16-1:0] node26857;
	wire [16-1:0] node26860;
	wire [16-1:0] node26863;
	wire [16-1:0] node26864;
	wire [16-1:0] node26867;
	wire [16-1:0] node26870;
	wire [16-1:0] node26871;
	wire [16-1:0] node26872;
	wire [16-1:0] node26875;
	wire [16-1:0] node26878;
	wire [16-1:0] node26879;
	wire [16-1:0] node26882;
	wire [16-1:0] node26885;
	wire [16-1:0] node26886;
	wire [16-1:0] node26887;
	wire [16-1:0] node26888;
	wire [16-1:0] node26891;
	wire [16-1:0] node26894;
	wire [16-1:0] node26895;
	wire [16-1:0] node26898;
	wire [16-1:0] node26901;
	wire [16-1:0] node26902;
	wire [16-1:0] node26903;
	wire [16-1:0] node26906;
	wire [16-1:0] node26909;
	wire [16-1:0] node26910;
	wire [16-1:0] node26913;
	wire [16-1:0] node26916;
	wire [16-1:0] node26917;
	wire [16-1:0] node26918;
	wire [16-1:0] node26919;
	wire [16-1:0] node26920;
	wire [16-1:0] node26923;
	wire [16-1:0] node26926;
	wire [16-1:0] node26928;
	wire [16-1:0] node26931;
	wire [16-1:0] node26932;
	wire [16-1:0] node26934;
	wire [16-1:0] node26937;
	wire [16-1:0] node26938;
	wire [16-1:0] node26941;
	wire [16-1:0] node26944;
	wire [16-1:0] node26945;
	wire [16-1:0] node26946;
	wire [16-1:0] node26947;
	wire [16-1:0] node26950;
	wire [16-1:0] node26953;
	wire [16-1:0] node26954;
	wire [16-1:0] node26957;
	wire [16-1:0] node26960;
	wire [16-1:0] node26961;
	wire [16-1:0] node26963;
	wire [16-1:0] node26966;
	wire [16-1:0] node26967;
	wire [16-1:0] node26970;
	wire [16-1:0] node26973;
	wire [16-1:0] node26974;
	wire [16-1:0] node26975;
	wire [16-1:0] node26976;
	wire [16-1:0] node26977;
	wire [16-1:0] node26978;
	wire [16-1:0] node26979;
	wire [16-1:0] node26982;
	wire [16-1:0] node26985;
	wire [16-1:0] node26986;
	wire [16-1:0] node26989;
	wire [16-1:0] node26992;
	wire [16-1:0] node26993;
	wire [16-1:0] node26994;
	wire [16-1:0] node26997;
	wire [16-1:0] node27000;
	wire [16-1:0] node27001;
	wire [16-1:0] node27005;
	wire [16-1:0] node27006;
	wire [16-1:0] node27007;
	wire [16-1:0] node27008;
	wire [16-1:0] node27011;
	wire [16-1:0] node27014;
	wire [16-1:0] node27015;
	wire [16-1:0] node27019;
	wire [16-1:0] node27020;
	wire [16-1:0] node27021;
	wire [16-1:0] node27024;
	wire [16-1:0] node27027;
	wire [16-1:0] node27028;
	wire [16-1:0] node27031;
	wire [16-1:0] node27034;
	wire [16-1:0] node27035;
	wire [16-1:0] node27036;
	wire [16-1:0] node27037;
	wire [16-1:0] node27038;
	wire [16-1:0] node27042;
	wire [16-1:0] node27043;
	wire [16-1:0] node27047;
	wire [16-1:0] node27048;
	wire [16-1:0] node27050;
	wire [16-1:0] node27053;
	wire [16-1:0] node27054;
	wire [16-1:0] node27058;
	wire [16-1:0] node27059;
	wire [16-1:0] node27060;
	wire [16-1:0] node27061;
	wire [16-1:0] node27064;
	wire [16-1:0] node27067;
	wire [16-1:0] node27068;
	wire [16-1:0] node27071;
	wire [16-1:0] node27074;
	wire [16-1:0] node27075;
	wire [16-1:0] node27076;
	wire [16-1:0] node27080;
	wire [16-1:0] node27081;
	wire [16-1:0] node27084;
	wire [16-1:0] node27087;
	wire [16-1:0] node27088;
	wire [16-1:0] node27089;
	wire [16-1:0] node27090;
	wire [16-1:0] node27091;
	wire [16-1:0] node27092;
	wire [16-1:0] node27096;
	wire [16-1:0] node27097;
	wire [16-1:0] node27100;
	wire [16-1:0] node27103;
	wire [16-1:0] node27104;
	wire [16-1:0] node27105;
	wire [16-1:0] node27108;
	wire [16-1:0] node27111;
	wire [16-1:0] node27112;
	wire [16-1:0] node27115;
	wire [16-1:0] node27118;
	wire [16-1:0] node27119;
	wire [16-1:0] node27120;
	wire [16-1:0] node27121;
	wire [16-1:0] node27124;
	wire [16-1:0] node27127;
	wire [16-1:0] node27128;
	wire [16-1:0] node27131;
	wire [16-1:0] node27134;
	wire [16-1:0] node27135;
	wire [16-1:0] node27136;
	wire [16-1:0] node27139;
	wire [16-1:0] node27142;
	wire [16-1:0] node27143;
	wire [16-1:0] node27146;
	wire [16-1:0] node27149;
	wire [16-1:0] node27150;
	wire [16-1:0] node27151;
	wire [16-1:0] node27152;
	wire [16-1:0] node27153;
	wire [16-1:0] node27156;
	wire [16-1:0] node27159;
	wire [16-1:0] node27160;
	wire [16-1:0] node27163;
	wire [16-1:0] node27166;
	wire [16-1:0] node27167;
	wire [16-1:0] node27168;
	wire [16-1:0] node27171;
	wire [16-1:0] node27174;
	wire [16-1:0] node27175;
	wire [16-1:0] node27178;
	wire [16-1:0] node27181;
	wire [16-1:0] node27182;
	wire [16-1:0] node27183;
	wire [16-1:0] node27185;
	wire [16-1:0] node27188;
	wire [16-1:0] node27189;
	wire [16-1:0] node27192;
	wire [16-1:0] node27195;
	wire [16-1:0] node27196;
	wire [16-1:0] node27197;
	wire [16-1:0] node27200;
	wire [16-1:0] node27203;
	wire [16-1:0] node27205;
	wire [16-1:0] node27208;
	wire [16-1:0] node27209;
	wire [16-1:0] node27210;
	wire [16-1:0] node27211;
	wire [16-1:0] node27212;
	wire [16-1:0] node27213;
	wire [16-1:0] node27214;
	wire [16-1:0] node27215;
	wire [16-1:0] node27216;
	wire [16-1:0] node27217;
	wire [16-1:0] node27218;
	wire [16-1:0] node27221;
	wire [16-1:0] node27224;
	wire [16-1:0] node27225;
	wire [16-1:0] node27228;
	wire [16-1:0] node27231;
	wire [16-1:0] node27232;
	wire [16-1:0] node27233;
	wire [16-1:0] node27236;
	wire [16-1:0] node27239;
	wire [16-1:0] node27240;
	wire [16-1:0] node27243;
	wire [16-1:0] node27246;
	wire [16-1:0] node27247;
	wire [16-1:0] node27248;
	wire [16-1:0] node27249;
	wire [16-1:0] node27252;
	wire [16-1:0] node27255;
	wire [16-1:0] node27257;
	wire [16-1:0] node27260;
	wire [16-1:0] node27261;
	wire [16-1:0] node27262;
	wire [16-1:0] node27265;
	wire [16-1:0] node27268;
	wire [16-1:0] node27269;
	wire [16-1:0] node27272;
	wire [16-1:0] node27275;
	wire [16-1:0] node27276;
	wire [16-1:0] node27277;
	wire [16-1:0] node27278;
	wire [16-1:0] node27279;
	wire [16-1:0] node27282;
	wire [16-1:0] node27285;
	wire [16-1:0] node27286;
	wire [16-1:0] node27290;
	wire [16-1:0] node27291;
	wire [16-1:0] node27293;
	wire [16-1:0] node27296;
	wire [16-1:0] node27297;
	wire [16-1:0] node27301;
	wire [16-1:0] node27302;
	wire [16-1:0] node27303;
	wire [16-1:0] node27304;
	wire [16-1:0] node27307;
	wire [16-1:0] node27310;
	wire [16-1:0] node27311;
	wire [16-1:0] node27314;
	wire [16-1:0] node27317;
	wire [16-1:0] node27318;
	wire [16-1:0] node27319;
	wire [16-1:0] node27322;
	wire [16-1:0] node27325;
	wire [16-1:0] node27326;
	wire [16-1:0] node27330;
	wire [16-1:0] node27331;
	wire [16-1:0] node27332;
	wire [16-1:0] node27333;
	wire [16-1:0] node27334;
	wire [16-1:0] node27335;
	wire [16-1:0] node27338;
	wire [16-1:0] node27341;
	wire [16-1:0] node27342;
	wire [16-1:0] node27345;
	wire [16-1:0] node27348;
	wire [16-1:0] node27349;
	wire [16-1:0] node27350;
	wire [16-1:0] node27354;
	wire [16-1:0] node27355;
	wire [16-1:0] node27358;
	wire [16-1:0] node27361;
	wire [16-1:0] node27362;
	wire [16-1:0] node27363;
	wire [16-1:0] node27365;
	wire [16-1:0] node27368;
	wire [16-1:0] node27369;
	wire [16-1:0] node27372;
	wire [16-1:0] node27375;
	wire [16-1:0] node27376;
	wire [16-1:0] node27377;
	wire [16-1:0] node27380;
	wire [16-1:0] node27383;
	wire [16-1:0] node27384;
	wire [16-1:0] node27387;
	wire [16-1:0] node27390;
	wire [16-1:0] node27391;
	wire [16-1:0] node27392;
	wire [16-1:0] node27393;
	wire [16-1:0] node27394;
	wire [16-1:0] node27397;
	wire [16-1:0] node27400;
	wire [16-1:0] node27402;
	wire [16-1:0] node27405;
	wire [16-1:0] node27406;
	wire [16-1:0] node27407;
	wire [16-1:0] node27410;
	wire [16-1:0] node27413;
	wire [16-1:0] node27414;
	wire [16-1:0] node27417;
	wire [16-1:0] node27420;
	wire [16-1:0] node27421;
	wire [16-1:0] node27422;
	wire [16-1:0] node27423;
	wire [16-1:0] node27426;
	wire [16-1:0] node27429;
	wire [16-1:0] node27430;
	wire [16-1:0] node27433;
	wire [16-1:0] node27436;
	wire [16-1:0] node27437;
	wire [16-1:0] node27438;
	wire [16-1:0] node27441;
	wire [16-1:0] node27444;
	wire [16-1:0] node27445;
	wire [16-1:0] node27448;
	wire [16-1:0] node27451;
	wire [16-1:0] node27452;
	wire [16-1:0] node27453;
	wire [16-1:0] node27454;
	wire [16-1:0] node27455;
	wire [16-1:0] node27456;
	wire [16-1:0] node27457;
	wire [16-1:0] node27460;
	wire [16-1:0] node27463;
	wire [16-1:0] node27464;
	wire [16-1:0] node27468;
	wire [16-1:0] node27469;
	wire [16-1:0] node27470;
	wire [16-1:0] node27473;
	wire [16-1:0] node27476;
	wire [16-1:0] node27477;
	wire [16-1:0] node27480;
	wire [16-1:0] node27483;
	wire [16-1:0] node27484;
	wire [16-1:0] node27485;
	wire [16-1:0] node27486;
	wire [16-1:0] node27489;
	wire [16-1:0] node27492;
	wire [16-1:0] node27493;
	wire [16-1:0] node27496;
	wire [16-1:0] node27499;
	wire [16-1:0] node27500;
	wire [16-1:0] node27501;
	wire [16-1:0] node27504;
	wire [16-1:0] node27507;
	wire [16-1:0] node27508;
	wire [16-1:0] node27511;
	wire [16-1:0] node27514;
	wire [16-1:0] node27515;
	wire [16-1:0] node27516;
	wire [16-1:0] node27517;
	wire [16-1:0] node27518;
	wire [16-1:0] node27521;
	wire [16-1:0] node27524;
	wire [16-1:0] node27525;
	wire [16-1:0] node27528;
	wire [16-1:0] node27531;
	wire [16-1:0] node27532;
	wire [16-1:0] node27533;
	wire [16-1:0] node27536;
	wire [16-1:0] node27539;
	wire [16-1:0] node27540;
	wire [16-1:0] node27543;
	wire [16-1:0] node27546;
	wire [16-1:0] node27547;
	wire [16-1:0] node27548;
	wire [16-1:0] node27549;
	wire [16-1:0] node27552;
	wire [16-1:0] node27555;
	wire [16-1:0] node27556;
	wire [16-1:0] node27559;
	wire [16-1:0] node27562;
	wire [16-1:0] node27563;
	wire [16-1:0] node27565;
	wire [16-1:0] node27568;
	wire [16-1:0] node27569;
	wire [16-1:0] node27573;
	wire [16-1:0] node27574;
	wire [16-1:0] node27575;
	wire [16-1:0] node27576;
	wire [16-1:0] node27577;
	wire [16-1:0] node27578;
	wire [16-1:0] node27581;
	wire [16-1:0] node27584;
	wire [16-1:0] node27585;
	wire [16-1:0] node27588;
	wire [16-1:0] node27591;
	wire [16-1:0] node27592;
	wire [16-1:0] node27593;
	wire [16-1:0] node27596;
	wire [16-1:0] node27599;
	wire [16-1:0] node27600;
	wire [16-1:0] node27603;
	wire [16-1:0] node27606;
	wire [16-1:0] node27607;
	wire [16-1:0] node27608;
	wire [16-1:0] node27609;
	wire [16-1:0] node27612;
	wire [16-1:0] node27615;
	wire [16-1:0] node27616;
	wire [16-1:0] node27619;
	wire [16-1:0] node27622;
	wire [16-1:0] node27623;
	wire [16-1:0] node27624;
	wire [16-1:0] node27627;
	wire [16-1:0] node27630;
	wire [16-1:0] node27631;
	wire [16-1:0] node27634;
	wire [16-1:0] node27637;
	wire [16-1:0] node27638;
	wire [16-1:0] node27639;
	wire [16-1:0] node27640;
	wire [16-1:0] node27641;
	wire [16-1:0] node27644;
	wire [16-1:0] node27647;
	wire [16-1:0] node27649;
	wire [16-1:0] node27652;
	wire [16-1:0] node27653;
	wire [16-1:0] node27654;
	wire [16-1:0] node27657;
	wire [16-1:0] node27660;
	wire [16-1:0] node27661;
	wire [16-1:0] node27665;
	wire [16-1:0] node27666;
	wire [16-1:0] node27667;
	wire [16-1:0] node27669;
	wire [16-1:0] node27672;
	wire [16-1:0] node27674;
	wire [16-1:0] node27677;
	wire [16-1:0] node27678;
	wire [16-1:0] node27679;
	wire [16-1:0] node27682;
	wire [16-1:0] node27686;
	wire [16-1:0] node27687;
	wire [16-1:0] node27688;
	wire [16-1:0] node27689;
	wire [16-1:0] node27690;
	wire [16-1:0] node27691;
	wire [16-1:0] node27692;
	wire [16-1:0] node27693;
	wire [16-1:0] node27696;
	wire [16-1:0] node27699;
	wire [16-1:0] node27701;
	wire [16-1:0] node27704;
	wire [16-1:0] node27705;
	wire [16-1:0] node27707;
	wire [16-1:0] node27710;
	wire [16-1:0] node27711;
	wire [16-1:0] node27714;
	wire [16-1:0] node27717;
	wire [16-1:0] node27718;
	wire [16-1:0] node27719;
	wire [16-1:0] node27720;
	wire [16-1:0] node27724;
	wire [16-1:0] node27725;
	wire [16-1:0] node27728;
	wire [16-1:0] node27731;
	wire [16-1:0] node27732;
	wire [16-1:0] node27733;
	wire [16-1:0] node27736;
	wire [16-1:0] node27739;
	wire [16-1:0] node27741;
	wire [16-1:0] node27744;
	wire [16-1:0] node27745;
	wire [16-1:0] node27746;
	wire [16-1:0] node27747;
	wire [16-1:0] node27748;
	wire [16-1:0] node27751;
	wire [16-1:0] node27754;
	wire [16-1:0] node27755;
	wire [16-1:0] node27758;
	wire [16-1:0] node27761;
	wire [16-1:0] node27762;
	wire [16-1:0] node27763;
	wire [16-1:0] node27766;
	wire [16-1:0] node27769;
	wire [16-1:0] node27770;
	wire [16-1:0] node27773;
	wire [16-1:0] node27776;
	wire [16-1:0] node27777;
	wire [16-1:0] node27778;
	wire [16-1:0] node27779;
	wire [16-1:0] node27782;
	wire [16-1:0] node27785;
	wire [16-1:0] node27786;
	wire [16-1:0] node27790;
	wire [16-1:0] node27791;
	wire [16-1:0] node27792;
	wire [16-1:0] node27795;
	wire [16-1:0] node27798;
	wire [16-1:0] node27799;
	wire [16-1:0] node27803;
	wire [16-1:0] node27804;
	wire [16-1:0] node27805;
	wire [16-1:0] node27806;
	wire [16-1:0] node27807;
	wire [16-1:0] node27808;
	wire [16-1:0] node27811;
	wire [16-1:0] node27814;
	wire [16-1:0] node27815;
	wire [16-1:0] node27818;
	wire [16-1:0] node27821;
	wire [16-1:0] node27822;
	wire [16-1:0] node27823;
	wire [16-1:0] node27826;
	wire [16-1:0] node27829;
	wire [16-1:0] node27830;
	wire [16-1:0] node27833;
	wire [16-1:0] node27836;
	wire [16-1:0] node27837;
	wire [16-1:0] node27838;
	wire [16-1:0] node27839;
	wire [16-1:0] node27842;
	wire [16-1:0] node27845;
	wire [16-1:0] node27846;
	wire [16-1:0] node27849;
	wire [16-1:0] node27852;
	wire [16-1:0] node27853;
	wire [16-1:0] node27854;
	wire [16-1:0] node27857;
	wire [16-1:0] node27860;
	wire [16-1:0] node27861;
	wire [16-1:0] node27864;
	wire [16-1:0] node27867;
	wire [16-1:0] node27868;
	wire [16-1:0] node27869;
	wire [16-1:0] node27870;
	wire [16-1:0] node27871;
	wire [16-1:0] node27875;
	wire [16-1:0] node27876;
	wire [16-1:0] node27879;
	wire [16-1:0] node27882;
	wire [16-1:0] node27883;
	wire [16-1:0] node27884;
	wire [16-1:0] node27887;
	wire [16-1:0] node27890;
	wire [16-1:0] node27891;
	wire [16-1:0] node27895;
	wire [16-1:0] node27896;
	wire [16-1:0] node27897;
	wire [16-1:0] node27898;
	wire [16-1:0] node27901;
	wire [16-1:0] node27904;
	wire [16-1:0] node27905;
	wire [16-1:0] node27908;
	wire [16-1:0] node27911;
	wire [16-1:0] node27912;
	wire [16-1:0] node27913;
	wire [16-1:0] node27916;
	wire [16-1:0] node27919;
	wire [16-1:0] node27920;
	wire [16-1:0] node27923;
	wire [16-1:0] node27926;
	wire [16-1:0] node27927;
	wire [16-1:0] node27928;
	wire [16-1:0] node27929;
	wire [16-1:0] node27930;
	wire [16-1:0] node27931;
	wire [16-1:0] node27932;
	wire [16-1:0] node27935;
	wire [16-1:0] node27938;
	wire [16-1:0] node27939;
	wire [16-1:0] node27942;
	wire [16-1:0] node27945;
	wire [16-1:0] node27946;
	wire [16-1:0] node27948;
	wire [16-1:0] node27951;
	wire [16-1:0] node27952;
	wire [16-1:0] node27955;
	wire [16-1:0] node27958;
	wire [16-1:0] node27959;
	wire [16-1:0] node27960;
	wire [16-1:0] node27961;
	wire [16-1:0] node27964;
	wire [16-1:0] node27967;
	wire [16-1:0] node27968;
	wire [16-1:0] node27971;
	wire [16-1:0] node27974;
	wire [16-1:0] node27975;
	wire [16-1:0] node27976;
	wire [16-1:0] node27979;
	wire [16-1:0] node27982;
	wire [16-1:0] node27983;
	wire [16-1:0] node27986;
	wire [16-1:0] node27989;
	wire [16-1:0] node27990;
	wire [16-1:0] node27991;
	wire [16-1:0] node27992;
	wire [16-1:0] node27994;
	wire [16-1:0] node27997;
	wire [16-1:0] node27998;
	wire [16-1:0] node28001;
	wire [16-1:0] node28004;
	wire [16-1:0] node28005;
	wire [16-1:0] node28006;
	wire [16-1:0] node28009;
	wire [16-1:0] node28012;
	wire [16-1:0] node28013;
	wire [16-1:0] node28016;
	wire [16-1:0] node28019;
	wire [16-1:0] node28020;
	wire [16-1:0] node28021;
	wire [16-1:0] node28022;
	wire [16-1:0] node28025;
	wire [16-1:0] node28028;
	wire [16-1:0] node28029;
	wire [16-1:0] node28032;
	wire [16-1:0] node28035;
	wire [16-1:0] node28036;
	wire [16-1:0] node28037;
	wire [16-1:0] node28040;
	wire [16-1:0] node28043;
	wire [16-1:0] node28045;
	wire [16-1:0] node28048;
	wire [16-1:0] node28049;
	wire [16-1:0] node28050;
	wire [16-1:0] node28051;
	wire [16-1:0] node28052;
	wire [16-1:0] node28053;
	wire [16-1:0] node28056;
	wire [16-1:0] node28059;
	wire [16-1:0] node28060;
	wire [16-1:0] node28063;
	wire [16-1:0] node28066;
	wire [16-1:0] node28067;
	wire [16-1:0] node28068;
	wire [16-1:0] node28071;
	wire [16-1:0] node28074;
	wire [16-1:0] node28075;
	wire [16-1:0] node28078;
	wire [16-1:0] node28081;
	wire [16-1:0] node28082;
	wire [16-1:0] node28083;
	wire [16-1:0] node28084;
	wire [16-1:0] node28087;
	wire [16-1:0] node28090;
	wire [16-1:0] node28091;
	wire [16-1:0] node28094;
	wire [16-1:0] node28097;
	wire [16-1:0] node28098;
	wire [16-1:0] node28099;
	wire [16-1:0] node28102;
	wire [16-1:0] node28105;
	wire [16-1:0] node28106;
	wire [16-1:0] node28109;
	wire [16-1:0] node28112;
	wire [16-1:0] node28113;
	wire [16-1:0] node28114;
	wire [16-1:0] node28115;
	wire [16-1:0] node28116;
	wire [16-1:0] node28119;
	wire [16-1:0] node28122;
	wire [16-1:0] node28123;
	wire [16-1:0] node28126;
	wire [16-1:0] node28129;
	wire [16-1:0] node28130;
	wire [16-1:0] node28131;
	wire [16-1:0] node28135;
	wire [16-1:0] node28137;
	wire [16-1:0] node28140;
	wire [16-1:0] node28141;
	wire [16-1:0] node28142;
	wire [16-1:0] node28143;
	wire [16-1:0] node28146;
	wire [16-1:0] node28149;
	wire [16-1:0] node28150;
	wire [16-1:0] node28153;
	wire [16-1:0] node28156;
	wire [16-1:0] node28157;
	wire [16-1:0] node28158;
	wire [16-1:0] node28161;
	wire [16-1:0] node28164;
	wire [16-1:0] node28165;
	wire [16-1:0] node28168;
	wire [16-1:0] node28171;
	wire [16-1:0] node28172;
	wire [16-1:0] node28173;
	wire [16-1:0] node28174;
	wire [16-1:0] node28175;
	wire [16-1:0] node28176;
	wire [16-1:0] node28177;
	wire [16-1:0] node28178;
	wire [16-1:0] node28179;
	wire [16-1:0] node28183;
	wire [16-1:0] node28184;
	wire [16-1:0] node28187;
	wire [16-1:0] node28190;
	wire [16-1:0] node28191;
	wire [16-1:0] node28192;
	wire [16-1:0] node28195;
	wire [16-1:0] node28198;
	wire [16-1:0] node28200;
	wire [16-1:0] node28203;
	wire [16-1:0] node28204;
	wire [16-1:0] node28205;
	wire [16-1:0] node28206;
	wire [16-1:0] node28209;
	wire [16-1:0] node28212;
	wire [16-1:0] node28213;
	wire [16-1:0] node28216;
	wire [16-1:0] node28219;
	wire [16-1:0] node28220;
	wire [16-1:0] node28221;
	wire [16-1:0] node28224;
	wire [16-1:0] node28227;
	wire [16-1:0] node28228;
	wire [16-1:0] node28231;
	wire [16-1:0] node28234;
	wire [16-1:0] node28235;
	wire [16-1:0] node28236;
	wire [16-1:0] node28237;
	wire [16-1:0] node28238;
	wire [16-1:0] node28242;
	wire [16-1:0] node28243;
	wire [16-1:0] node28246;
	wire [16-1:0] node28249;
	wire [16-1:0] node28250;
	wire [16-1:0] node28251;
	wire [16-1:0] node28254;
	wire [16-1:0] node28257;
	wire [16-1:0] node28258;
	wire [16-1:0] node28262;
	wire [16-1:0] node28263;
	wire [16-1:0] node28264;
	wire [16-1:0] node28265;
	wire [16-1:0] node28268;
	wire [16-1:0] node28271;
	wire [16-1:0] node28272;
	wire [16-1:0] node28276;
	wire [16-1:0] node28277;
	wire [16-1:0] node28278;
	wire [16-1:0] node28281;
	wire [16-1:0] node28284;
	wire [16-1:0] node28285;
	wire [16-1:0] node28289;
	wire [16-1:0] node28290;
	wire [16-1:0] node28291;
	wire [16-1:0] node28292;
	wire [16-1:0] node28293;
	wire [16-1:0] node28294;
	wire [16-1:0] node28297;
	wire [16-1:0] node28300;
	wire [16-1:0] node28302;
	wire [16-1:0] node28305;
	wire [16-1:0] node28306;
	wire [16-1:0] node28307;
	wire [16-1:0] node28310;
	wire [16-1:0] node28313;
	wire [16-1:0] node28314;
	wire [16-1:0] node28317;
	wire [16-1:0] node28320;
	wire [16-1:0] node28321;
	wire [16-1:0] node28322;
	wire [16-1:0] node28323;
	wire [16-1:0] node28326;
	wire [16-1:0] node28329;
	wire [16-1:0] node28331;
	wire [16-1:0] node28334;
	wire [16-1:0] node28335;
	wire [16-1:0] node28336;
	wire [16-1:0] node28339;
	wire [16-1:0] node28342;
	wire [16-1:0] node28343;
	wire [16-1:0] node28346;
	wire [16-1:0] node28349;
	wire [16-1:0] node28350;
	wire [16-1:0] node28351;
	wire [16-1:0] node28352;
	wire [16-1:0] node28353;
	wire [16-1:0] node28356;
	wire [16-1:0] node28359;
	wire [16-1:0] node28360;
	wire [16-1:0] node28364;
	wire [16-1:0] node28365;
	wire [16-1:0] node28366;
	wire [16-1:0] node28370;
	wire [16-1:0] node28371;
	wire [16-1:0] node28374;
	wire [16-1:0] node28377;
	wire [16-1:0] node28378;
	wire [16-1:0] node28379;
	wire [16-1:0] node28380;
	wire [16-1:0] node28383;
	wire [16-1:0] node28386;
	wire [16-1:0] node28388;
	wire [16-1:0] node28391;
	wire [16-1:0] node28392;
	wire [16-1:0] node28393;
	wire [16-1:0] node28396;
	wire [16-1:0] node28399;
	wire [16-1:0] node28400;
	wire [16-1:0] node28403;
	wire [16-1:0] node28406;
	wire [16-1:0] node28407;
	wire [16-1:0] node28408;
	wire [16-1:0] node28409;
	wire [16-1:0] node28410;
	wire [16-1:0] node28411;
	wire [16-1:0] node28412;
	wire [16-1:0] node28415;
	wire [16-1:0] node28418;
	wire [16-1:0] node28419;
	wire [16-1:0] node28422;
	wire [16-1:0] node28425;
	wire [16-1:0] node28426;
	wire [16-1:0] node28427;
	wire [16-1:0] node28430;
	wire [16-1:0] node28433;
	wire [16-1:0] node28434;
	wire [16-1:0] node28437;
	wire [16-1:0] node28440;
	wire [16-1:0] node28441;
	wire [16-1:0] node28442;
	wire [16-1:0] node28443;
	wire [16-1:0] node28446;
	wire [16-1:0] node28449;
	wire [16-1:0] node28450;
	wire [16-1:0] node28453;
	wire [16-1:0] node28456;
	wire [16-1:0] node28457;
	wire [16-1:0] node28458;
	wire [16-1:0] node28461;
	wire [16-1:0] node28464;
	wire [16-1:0] node28465;
	wire [16-1:0] node28468;
	wire [16-1:0] node28471;
	wire [16-1:0] node28472;
	wire [16-1:0] node28473;
	wire [16-1:0] node28474;
	wire [16-1:0] node28475;
	wire [16-1:0] node28478;
	wire [16-1:0] node28481;
	wire [16-1:0] node28482;
	wire [16-1:0] node28485;
	wire [16-1:0] node28488;
	wire [16-1:0] node28489;
	wire [16-1:0] node28490;
	wire [16-1:0] node28493;
	wire [16-1:0] node28496;
	wire [16-1:0] node28497;
	wire [16-1:0] node28500;
	wire [16-1:0] node28503;
	wire [16-1:0] node28504;
	wire [16-1:0] node28505;
	wire [16-1:0] node28506;
	wire [16-1:0] node28510;
	wire [16-1:0] node28511;
	wire [16-1:0] node28515;
	wire [16-1:0] node28516;
	wire [16-1:0] node28517;
	wire [16-1:0] node28521;
	wire [16-1:0] node28522;
	wire [16-1:0] node28525;
	wire [16-1:0] node28528;
	wire [16-1:0] node28529;
	wire [16-1:0] node28530;
	wire [16-1:0] node28531;
	wire [16-1:0] node28532;
	wire [16-1:0] node28533;
	wire [16-1:0] node28536;
	wire [16-1:0] node28539;
	wire [16-1:0] node28541;
	wire [16-1:0] node28544;
	wire [16-1:0] node28545;
	wire [16-1:0] node28546;
	wire [16-1:0] node28550;
	wire [16-1:0] node28551;
	wire [16-1:0] node28554;
	wire [16-1:0] node28557;
	wire [16-1:0] node28558;
	wire [16-1:0] node28559;
	wire [16-1:0] node28560;
	wire [16-1:0] node28563;
	wire [16-1:0] node28566;
	wire [16-1:0] node28567;
	wire [16-1:0] node28570;
	wire [16-1:0] node28573;
	wire [16-1:0] node28574;
	wire [16-1:0] node28575;
	wire [16-1:0] node28578;
	wire [16-1:0] node28581;
	wire [16-1:0] node28582;
	wire [16-1:0] node28585;
	wire [16-1:0] node28588;
	wire [16-1:0] node28589;
	wire [16-1:0] node28590;
	wire [16-1:0] node28591;
	wire [16-1:0] node28592;
	wire [16-1:0] node28595;
	wire [16-1:0] node28598;
	wire [16-1:0] node28599;
	wire [16-1:0] node28602;
	wire [16-1:0] node28605;
	wire [16-1:0] node28606;
	wire [16-1:0] node28607;
	wire [16-1:0] node28610;
	wire [16-1:0] node28613;
	wire [16-1:0] node28614;
	wire [16-1:0] node28617;
	wire [16-1:0] node28620;
	wire [16-1:0] node28621;
	wire [16-1:0] node28622;
	wire [16-1:0] node28623;
	wire [16-1:0] node28626;
	wire [16-1:0] node28629;
	wire [16-1:0] node28630;
	wire [16-1:0] node28633;
	wire [16-1:0] node28636;
	wire [16-1:0] node28637;
	wire [16-1:0] node28638;
	wire [16-1:0] node28641;
	wire [16-1:0] node28644;
	wire [16-1:0] node28645;
	wire [16-1:0] node28648;
	wire [16-1:0] node28651;
	wire [16-1:0] node28652;
	wire [16-1:0] node28653;
	wire [16-1:0] node28654;
	wire [16-1:0] node28655;
	wire [16-1:0] node28656;
	wire [16-1:0] node28657;
	wire [16-1:0] node28659;
	wire [16-1:0] node28662;
	wire [16-1:0] node28663;
	wire [16-1:0] node28666;
	wire [16-1:0] node28669;
	wire [16-1:0] node28670;
	wire [16-1:0] node28672;
	wire [16-1:0] node28675;
	wire [16-1:0] node28676;
	wire [16-1:0] node28679;
	wire [16-1:0] node28682;
	wire [16-1:0] node28683;
	wire [16-1:0] node28684;
	wire [16-1:0] node28685;
	wire [16-1:0] node28688;
	wire [16-1:0] node28691;
	wire [16-1:0] node28692;
	wire [16-1:0] node28696;
	wire [16-1:0] node28697;
	wire [16-1:0] node28698;
	wire [16-1:0] node28701;
	wire [16-1:0] node28704;
	wire [16-1:0] node28705;
	wire [16-1:0] node28708;
	wire [16-1:0] node28711;
	wire [16-1:0] node28712;
	wire [16-1:0] node28713;
	wire [16-1:0] node28714;
	wire [16-1:0] node28715;
	wire [16-1:0] node28718;
	wire [16-1:0] node28721;
	wire [16-1:0] node28722;
	wire [16-1:0] node28726;
	wire [16-1:0] node28727;
	wire [16-1:0] node28728;
	wire [16-1:0] node28731;
	wire [16-1:0] node28734;
	wire [16-1:0] node28735;
	wire [16-1:0] node28738;
	wire [16-1:0] node28741;
	wire [16-1:0] node28742;
	wire [16-1:0] node28743;
	wire [16-1:0] node28744;
	wire [16-1:0] node28747;
	wire [16-1:0] node28750;
	wire [16-1:0] node28751;
	wire [16-1:0] node28754;
	wire [16-1:0] node28757;
	wire [16-1:0] node28758;
	wire [16-1:0] node28760;
	wire [16-1:0] node28763;
	wire [16-1:0] node28764;
	wire [16-1:0] node28767;
	wire [16-1:0] node28770;
	wire [16-1:0] node28771;
	wire [16-1:0] node28772;
	wire [16-1:0] node28773;
	wire [16-1:0] node28774;
	wire [16-1:0] node28776;
	wire [16-1:0] node28779;
	wire [16-1:0] node28780;
	wire [16-1:0] node28783;
	wire [16-1:0] node28786;
	wire [16-1:0] node28787;
	wire [16-1:0] node28788;
	wire [16-1:0] node28791;
	wire [16-1:0] node28794;
	wire [16-1:0] node28795;
	wire [16-1:0] node28798;
	wire [16-1:0] node28801;
	wire [16-1:0] node28802;
	wire [16-1:0] node28803;
	wire [16-1:0] node28805;
	wire [16-1:0] node28808;
	wire [16-1:0] node28809;
	wire [16-1:0] node28812;
	wire [16-1:0] node28815;
	wire [16-1:0] node28816;
	wire [16-1:0] node28817;
	wire [16-1:0] node28820;
	wire [16-1:0] node28823;
	wire [16-1:0] node28824;
	wire [16-1:0] node28827;
	wire [16-1:0] node28830;
	wire [16-1:0] node28831;
	wire [16-1:0] node28832;
	wire [16-1:0] node28833;
	wire [16-1:0] node28835;
	wire [16-1:0] node28838;
	wire [16-1:0] node28839;
	wire [16-1:0] node28842;
	wire [16-1:0] node28845;
	wire [16-1:0] node28846;
	wire [16-1:0] node28847;
	wire [16-1:0] node28850;
	wire [16-1:0] node28853;
	wire [16-1:0] node28854;
	wire [16-1:0] node28857;
	wire [16-1:0] node28860;
	wire [16-1:0] node28861;
	wire [16-1:0] node28862;
	wire [16-1:0] node28863;
	wire [16-1:0] node28866;
	wire [16-1:0] node28869;
	wire [16-1:0] node28870;
	wire [16-1:0] node28873;
	wire [16-1:0] node28876;
	wire [16-1:0] node28877;
	wire [16-1:0] node28878;
	wire [16-1:0] node28881;
	wire [16-1:0] node28884;
	wire [16-1:0] node28885;
	wire [16-1:0] node28888;
	wire [16-1:0] node28891;
	wire [16-1:0] node28892;
	wire [16-1:0] node28893;
	wire [16-1:0] node28894;
	wire [16-1:0] node28895;
	wire [16-1:0] node28896;
	wire [16-1:0] node28897;
	wire [16-1:0] node28900;
	wire [16-1:0] node28903;
	wire [16-1:0] node28904;
	wire [16-1:0] node28907;
	wire [16-1:0] node28910;
	wire [16-1:0] node28911;
	wire [16-1:0] node28912;
	wire [16-1:0] node28915;
	wire [16-1:0] node28918;
	wire [16-1:0] node28919;
	wire [16-1:0] node28923;
	wire [16-1:0] node28924;
	wire [16-1:0] node28925;
	wire [16-1:0] node28926;
	wire [16-1:0] node28929;
	wire [16-1:0] node28932;
	wire [16-1:0] node28933;
	wire [16-1:0] node28937;
	wire [16-1:0] node28938;
	wire [16-1:0] node28939;
	wire [16-1:0] node28942;
	wire [16-1:0] node28945;
	wire [16-1:0] node28946;
	wire [16-1:0] node28949;
	wire [16-1:0] node28952;
	wire [16-1:0] node28953;
	wire [16-1:0] node28954;
	wire [16-1:0] node28955;
	wire [16-1:0] node28956;
	wire [16-1:0] node28959;
	wire [16-1:0] node28962;
	wire [16-1:0] node28963;
	wire [16-1:0] node28966;
	wire [16-1:0] node28969;
	wire [16-1:0] node28970;
	wire [16-1:0] node28971;
	wire [16-1:0] node28974;
	wire [16-1:0] node28977;
	wire [16-1:0] node28978;
	wire [16-1:0] node28981;
	wire [16-1:0] node28984;
	wire [16-1:0] node28985;
	wire [16-1:0] node28986;
	wire [16-1:0] node28987;
	wire [16-1:0] node28990;
	wire [16-1:0] node28993;
	wire [16-1:0] node28994;
	wire [16-1:0] node28998;
	wire [16-1:0] node28999;
	wire [16-1:0] node29000;
	wire [16-1:0] node29003;
	wire [16-1:0] node29006;
	wire [16-1:0] node29007;
	wire [16-1:0] node29010;
	wire [16-1:0] node29013;
	wire [16-1:0] node29014;
	wire [16-1:0] node29015;
	wire [16-1:0] node29016;
	wire [16-1:0] node29017;
	wire [16-1:0] node29018;
	wire [16-1:0] node29021;
	wire [16-1:0] node29024;
	wire [16-1:0] node29025;
	wire [16-1:0] node29028;
	wire [16-1:0] node29031;
	wire [16-1:0] node29032;
	wire [16-1:0] node29033;
	wire [16-1:0] node29036;
	wire [16-1:0] node29039;
	wire [16-1:0] node29041;
	wire [16-1:0] node29044;
	wire [16-1:0] node29045;
	wire [16-1:0] node29046;
	wire [16-1:0] node29047;
	wire [16-1:0] node29050;
	wire [16-1:0] node29053;
	wire [16-1:0] node29054;
	wire [16-1:0] node29057;
	wire [16-1:0] node29060;
	wire [16-1:0] node29061;
	wire [16-1:0] node29062;
	wire [16-1:0] node29065;
	wire [16-1:0] node29068;
	wire [16-1:0] node29069;
	wire [16-1:0] node29072;
	wire [16-1:0] node29075;
	wire [16-1:0] node29076;
	wire [16-1:0] node29077;
	wire [16-1:0] node29078;
	wire [16-1:0] node29079;
	wire [16-1:0] node29082;
	wire [16-1:0] node29085;
	wire [16-1:0] node29086;
	wire [16-1:0] node29090;
	wire [16-1:0] node29091;
	wire [16-1:0] node29092;
	wire [16-1:0] node29095;
	wire [16-1:0] node29098;
	wire [16-1:0] node29099;
	wire [16-1:0] node29102;
	wire [16-1:0] node29105;
	wire [16-1:0] node29106;
	wire [16-1:0] node29107;
	wire [16-1:0] node29108;
	wire [16-1:0] node29111;
	wire [16-1:0] node29114;
	wire [16-1:0] node29115;
	wire [16-1:0] node29118;
	wire [16-1:0] node29121;
	wire [16-1:0] node29122;
	wire [16-1:0] node29123;
	wire [16-1:0] node29126;
	wire [16-1:0] node29129;
	wire [16-1:0] node29130;
	wire [16-1:0] node29133;
	wire [16-1:0] node29136;
	wire [16-1:0] node29137;
	wire [16-1:0] node29138;
	wire [16-1:0] node29139;
	wire [16-1:0] node29140;
	wire [16-1:0] node29141;
	wire [16-1:0] node29142;
	wire [16-1:0] node29143;
	wire [16-1:0] node29144;
	wire [16-1:0] node29145;
	wire [16-1:0] node29148;
	wire [16-1:0] node29151;
	wire [16-1:0] node29152;
	wire [16-1:0] node29155;
	wire [16-1:0] node29158;
	wire [16-1:0] node29159;
	wire [16-1:0] node29160;
	wire [16-1:0] node29163;
	wire [16-1:0] node29166;
	wire [16-1:0] node29167;
	wire [16-1:0] node29170;
	wire [16-1:0] node29173;
	wire [16-1:0] node29174;
	wire [16-1:0] node29175;
	wire [16-1:0] node29176;
	wire [16-1:0] node29179;
	wire [16-1:0] node29182;
	wire [16-1:0] node29183;
	wire [16-1:0] node29186;
	wire [16-1:0] node29189;
	wire [16-1:0] node29190;
	wire [16-1:0] node29192;
	wire [16-1:0] node29195;
	wire [16-1:0] node29196;
	wire [16-1:0] node29200;
	wire [16-1:0] node29201;
	wire [16-1:0] node29202;
	wire [16-1:0] node29203;
	wire [16-1:0] node29204;
	wire [16-1:0] node29208;
	wire [16-1:0] node29209;
	wire [16-1:0] node29212;
	wire [16-1:0] node29215;
	wire [16-1:0] node29216;
	wire [16-1:0] node29218;
	wire [16-1:0] node29221;
	wire [16-1:0] node29222;
	wire [16-1:0] node29225;
	wire [16-1:0] node29228;
	wire [16-1:0] node29229;
	wire [16-1:0] node29230;
	wire [16-1:0] node29232;
	wire [16-1:0] node29235;
	wire [16-1:0] node29236;
	wire [16-1:0] node29239;
	wire [16-1:0] node29242;
	wire [16-1:0] node29243;
	wire [16-1:0] node29244;
	wire [16-1:0] node29247;
	wire [16-1:0] node29250;
	wire [16-1:0] node29251;
	wire [16-1:0] node29254;
	wire [16-1:0] node29257;
	wire [16-1:0] node29258;
	wire [16-1:0] node29259;
	wire [16-1:0] node29260;
	wire [16-1:0] node29261;
	wire [16-1:0] node29262;
	wire [16-1:0] node29265;
	wire [16-1:0] node29268;
	wire [16-1:0] node29269;
	wire [16-1:0] node29272;
	wire [16-1:0] node29275;
	wire [16-1:0] node29276;
	wire [16-1:0] node29277;
	wire [16-1:0] node29280;
	wire [16-1:0] node29283;
	wire [16-1:0] node29284;
	wire [16-1:0] node29287;
	wire [16-1:0] node29290;
	wire [16-1:0] node29291;
	wire [16-1:0] node29292;
	wire [16-1:0] node29294;
	wire [16-1:0] node29297;
	wire [16-1:0] node29298;
	wire [16-1:0] node29301;
	wire [16-1:0] node29304;
	wire [16-1:0] node29305;
	wire [16-1:0] node29306;
	wire [16-1:0] node29309;
	wire [16-1:0] node29312;
	wire [16-1:0] node29313;
	wire [16-1:0] node29316;
	wire [16-1:0] node29319;
	wire [16-1:0] node29320;
	wire [16-1:0] node29321;
	wire [16-1:0] node29322;
	wire [16-1:0] node29323;
	wire [16-1:0] node29326;
	wire [16-1:0] node29329;
	wire [16-1:0] node29330;
	wire [16-1:0] node29333;
	wire [16-1:0] node29336;
	wire [16-1:0] node29337;
	wire [16-1:0] node29338;
	wire [16-1:0] node29341;
	wire [16-1:0] node29344;
	wire [16-1:0] node29345;
	wire [16-1:0] node29348;
	wire [16-1:0] node29351;
	wire [16-1:0] node29352;
	wire [16-1:0] node29353;
	wire [16-1:0] node29354;
	wire [16-1:0] node29357;
	wire [16-1:0] node29360;
	wire [16-1:0] node29361;
	wire [16-1:0] node29364;
	wire [16-1:0] node29367;
	wire [16-1:0] node29368;
	wire [16-1:0] node29369;
	wire [16-1:0] node29372;
	wire [16-1:0] node29375;
	wire [16-1:0] node29376;
	wire [16-1:0] node29379;
	wire [16-1:0] node29382;
	wire [16-1:0] node29383;
	wire [16-1:0] node29384;
	wire [16-1:0] node29385;
	wire [16-1:0] node29386;
	wire [16-1:0] node29387;
	wire [16-1:0] node29388;
	wire [16-1:0] node29391;
	wire [16-1:0] node29394;
	wire [16-1:0] node29395;
	wire [16-1:0] node29399;
	wire [16-1:0] node29400;
	wire [16-1:0] node29401;
	wire [16-1:0] node29404;
	wire [16-1:0] node29407;
	wire [16-1:0] node29408;
	wire [16-1:0] node29411;
	wire [16-1:0] node29414;
	wire [16-1:0] node29415;
	wire [16-1:0] node29416;
	wire [16-1:0] node29417;
	wire [16-1:0] node29420;
	wire [16-1:0] node29423;
	wire [16-1:0] node29424;
	wire [16-1:0] node29427;
	wire [16-1:0] node29430;
	wire [16-1:0] node29431;
	wire [16-1:0] node29433;
	wire [16-1:0] node29436;
	wire [16-1:0] node29437;
	wire [16-1:0] node29441;
	wire [16-1:0] node29442;
	wire [16-1:0] node29443;
	wire [16-1:0] node29444;
	wire [16-1:0] node29446;
	wire [16-1:0] node29449;
	wire [16-1:0] node29450;
	wire [16-1:0] node29453;
	wire [16-1:0] node29456;
	wire [16-1:0] node29457;
	wire [16-1:0] node29458;
	wire [16-1:0] node29461;
	wire [16-1:0] node29464;
	wire [16-1:0] node29465;
	wire [16-1:0] node29468;
	wire [16-1:0] node29471;
	wire [16-1:0] node29472;
	wire [16-1:0] node29473;
	wire [16-1:0] node29474;
	wire [16-1:0] node29477;
	wire [16-1:0] node29480;
	wire [16-1:0] node29481;
	wire [16-1:0] node29484;
	wire [16-1:0] node29487;
	wire [16-1:0] node29488;
	wire [16-1:0] node29489;
	wire [16-1:0] node29492;
	wire [16-1:0] node29495;
	wire [16-1:0] node29496;
	wire [16-1:0] node29499;
	wire [16-1:0] node29502;
	wire [16-1:0] node29503;
	wire [16-1:0] node29504;
	wire [16-1:0] node29505;
	wire [16-1:0] node29506;
	wire [16-1:0] node29507;
	wire [16-1:0] node29510;
	wire [16-1:0] node29513;
	wire [16-1:0] node29514;
	wire [16-1:0] node29517;
	wire [16-1:0] node29520;
	wire [16-1:0] node29521;
	wire [16-1:0] node29522;
	wire [16-1:0] node29525;
	wire [16-1:0] node29528;
	wire [16-1:0] node29529;
	wire [16-1:0] node29532;
	wire [16-1:0] node29535;
	wire [16-1:0] node29536;
	wire [16-1:0] node29537;
	wire [16-1:0] node29538;
	wire [16-1:0] node29541;
	wire [16-1:0] node29544;
	wire [16-1:0] node29545;
	wire [16-1:0] node29548;
	wire [16-1:0] node29551;
	wire [16-1:0] node29552;
	wire [16-1:0] node29553;
	wire [16-1:0] node29556;
	wire [16-1:0] node29559;
	wire [16-1:0] node29560;
	wire [16-1:0] node29564;
	wire [16-1:0] node29565;
	wire [16-1:0] node29566;
	wire [16-1:0] node29567;
	wire [16-1:0] node29568;
	wire [16-1:0] node29571;
	wire [16-1:0] node29574;
	wire [16-1:0] node29575;
	wire [16-1:0] node29578;
	wire [16-1:0] node29581;
	wire [16-1:0] node29582;
	wire [16-1:0] node29583;
	wire [16-1:0] node29586;
	wire [16-1:0] node29589;
	wire [16-1:0] node29590;
	wire [16-1:0] node29593;
	wire [16-1:0] node29596;
	wire [16-1:0] node29597;
	wire [16-1:0] node29598;
	wire [16-1:0] node29599;
	wire [16-1:0] node29602;
	wire [16-1:0] node29605;
	wire [16-1:0] node29606;
	wire [16-1:0] node29609;
	wire [16-1:0] node29612;
	wire [16-1:0] node29613;
	wire [16-1:0] node29614;
	wire [16-1:0] node29618;
	wire [16-1:0] node29619;
	wire [16-1:0] node29622;
	wire [16-1:0] node29625;
	wire [16-1:0] node29626;
	wire [16-1:0] node29627;
	wire [16-1:0] node29628;
	wire [16-1:0] node29629;
	wire [16-1:0] node29630;
	wire [16-1:0] node29631;
	wire [16-1:0] node29632;
	wire [16-1:0] node29635;
	wire [16-1:0] node29638;
	wire [16-1:0] node29639;
	wire [16-1:0] node29642;
	wire [16-1:0] node29645;
	wire [16-1:0] node29646;
	wire [16-1:0] node29647;
	wire [16-1:0] node29650;
	wire [16-1:0] node29653;
	wire [16-1:0] node29656;
	wire [16-1:0] node29657;
	wire [16-1:0] node29658;
	wire [16-1:0] node29659;
	wire [16-1:0] node29662;
	wire [16-1:0] node29665;
	wire [16-1:0] node29666;
	wire [16-1:0] node29669;
	wire [16-1:0] node29672;
	wire [16-1:0] node29673;
	wire [16-1:0] node29674;
	wire [16-1:0] node29677;
	wire [16-1:0] node29680;
	wire [16-1:0] node29681;
	wire [16-1:0] node29684;
	wire [16-1:0] node29687;
	wire [16-1:0] node29688;
	wire [16-1:0] node29689;
	wire [16-1:0] node29690;
	wire [16-1:0] node29691;
	wire [16-1:0] node29694;
	wire [16-1:0] node29697;
	wire [16-1:0] node29699;
	wire [16-1:0] node29702;
	wire [16-1:0] node29703;
	wire [16-1:0] node29704;
	wire [16-1:0] node29707;
	wire [16-1:0] node29710;
	wire [16-1:0] node29711;
	wire [16-1:0] node29714;
	wire [16-1:0] node29717;
	wire [16-1:0] node29718;
	wire [16-1:0] node29719;
	wire [16-1:0] node29720;
	wire [16-1:0] node29723;
	wire [16-1:0] node29726;
	wire [16-1:0] node29727;
	wire [16-1:0] node29730;
	wire [16-1:0] node29733;
	wire [16-1:0] node29734;
	wire [16-1:0] node29735;
	wire [16-1:0] node29738;
	wire [16-1:0] node29741;
	wire [16-1:0] node29742;
	wire [16-1:0] node29745;
	wire [16-1:0] node29748;
	wire [16-1:0] node29749;
	wire [16-1:0] node29750;
	wire [16-1:0] node29751;
	wire [16-1:0] node29752;
	wire [16-1:0] node29753;
	wire [16-1:0] node29756;
	wire [16-1:0] node29759;
	wire [16-1:0] node29760;
	wire [16-1:0] node29763;
	wire [16-1:0] node29766;
	wire [16-1:0] node29767;
	wire [16-1:0] node29768;
	wire [16-1:0] node29771;
	wire [16-1:0] node29774;
	wire [16-1:0] node29775;
	wire [16-1:0] node29778;
	wire [16-1:0] node29781;
	wire [16-1:0] node29782;
	wire [16-1:0] node29783;
	wire [16-1:0] node29784;
	wire [16-1:0] node29787;
	wire [16-1:0] node29790;
	wire [16-1:0] node29791;
	wire [16-1:0] node29794;
	wire [16-1:0] node29797;
	wire [16-1:0] node29798;
	wire [16-1:0] node29799;
	wire [16-1:0] node29802;
	wire [16-1:0] node29805;
	wire [16-1:0] node29806;
	wire [16-1:0] node29809;
	wire [16-1:0] node29812;
	wire [16-1:0] node29813;
	wire [16-1:0] node29814;
	wire [16-1:0] node29815;
	wire [16-1:0] node29816;
	wire [16-1:0] node29819;
	wire [16-1:0] node29822;
	wire [16-1:0] node29823;
	wire [16-1:0] node29826;
	wire [16-1:0] node29829;
	wire [16-1:0] node29830;
	wire [16-1:0] node29831;
	wire [16-1:0] node29834;
	wire [16-1:0] node29837;
	wire [16-1:0] node29838;
	wire [16-1:0] node29841;
	wire [16-1:0] node29844;
	wire [16-1:0] node29845;
	wire [16-1:0] node29846;
	wire [16-1:0] node29849;
	wire [16-1:0] node29850;
	wire [16-1:0] node29853;
	wire [16-1:0] node29856;
	wire [16-1:0] node29857;
	wire [16-1:0] node29858;
	wire [16-1:0] node29862;
	wire [16-1:0] node29864;
	wire [16-1:0] node29867;
	wire [16-1:0] node29868;
	wire [16-1:0] node29869;
	wire [16-1:0] node29870;
	wire [16-1:0] node29871;
	wire [16-1:0] node29872;
	wire [16-1:0] node29873;
	wire [16-1:0] node29876;
	wire [16-1:0] node29879;
	wire [16-1:0] node29880;
	wire [16-1:0] node29883;
	wire [16-1:0] node29886;
	wire [16-1:0] node29887;
	wire [16-1:0] node29888;
	wire [16-1:0] node29891;
	wire [16-1:0] node29894;
	wire [16-1:0] node29895;
	wire [16-1:0] node29898;
	wire [16-1:0] node29901;
	wire [16-1:0] node29902;
	wire [16-1:0] node29903;
	wire [16-1:0] node29905;
	wire [16-1:0] node29908;
	wire [16-1:0] node29909;
	wire [16-1:0] node29912;
	wire [16-1:0] node29915;
	wire [16-1:0] node29916;
	wire [16-1:0] node29917;
	wire [16-1:0] node29920;
	wire [16-1:0] node29923;
	wire [16-1:0] node29924;
	wire [16-1:0] node29927;
	wire [16-1:0] node29930;
	wire [16-1:0] node29931;
	wire [16-1:0] node29932;
	wire [16-1:0] node29933;
	wire [16-1:0] node29934;
	wire [16-1:0] node29937;
	wire [16-1:0] node29940;
	wire [16-1:0] node29941;
	wire [16-1:0] node29944;
	wire [16-1:0] node29947;
	wire [16-1:0] node29948;
	wire [16-1:0] node29949;
	wire [16-1:0] node29952;
	wire [16-1:0] node29955;
	wire [16-1:0] node29957;
	wire [16-1:0] node29960;
	wire [16-1:0] node29961;
	wire [16-1:0] node29962;
	wire [16-1:0] node29963;
	wire [16-1:0] node29966;
	wire [16-1:0] node29969;
	wire [16-1:0] node29970;
	wire [16-1:0] node29973;
	wire [16-1:0] node29976;
	wire [16-1:0] node29977;
	wire [16-1:0] node29979;
	wire [16-1:0] node29982;
	wire [16-1:0] node29983;
	wire [16-1:0] node29986;
	wire [16-1:0] node29989;
	wire [16-1:0] node29990;
	wire [16-1:0] node29991;
	wire [16-1:0] node29992;
	wire [16-1:0] node29993;
	wire [16-1:0] node29994;
	wire [16-1:0] node29997;
	wire [16-1:0] node30000;
	wire [16-1:0] node30001;
	wire [16-1:0] node30004;
	wire [16-1:0] node30007;
	wire [16-1:0] node30008;
	wire [16-1:0] node30009;
	wire [16-1:0] node30012;
	wire [16-1:0] node30015;
	wire [16-1:0] node30016;
	wire [16-1:0] node30019;
	wire [16-1:0] node30022;
	wire [16-1:0] node30023;
	wire [16-1:0] node30024;
	wire [16-1:0] node30025;
	wire [16-1:0] node30028;
	wire [16-1:0] node30031;
	wire [16-1:0] node30032;
	wire [16-1:0] node30035;
	wire [16-1:0] node30038;
	wire [16-1:0] node30039;
	wire [16-1:0] node30040;
	wire [16-1:0] node30043;
	wire [16-1:0] node30046;
	wire [16-1:0] node30047;
	wire [16-1:0] node30050;
	wire [16-1:0] node30053;
	wire [16-1:0] node30054;
	wire [16-1:0] node30055;
	wire [16-1:0] node30056;
	wire [16-1:0] node30059;
	wire [16-1:0] node30060;
	wire [16-1:0] node30064;
	wire [16-1:0] node30065;
	wire [16-1:0] node30066;
	wire [16-1:0] node30069;
	wire [16-1:0] node30072;
	wire [16-1:0] node30073;
	wire [16-1:0] node30076;
	wire [16-1:0] node30079;
	wire [16-1:0] node30080;
	wire [16-1:0] node30081;
	wire [16-1:0] node30082;
	wire [16-1:0] node30085;
	wire [16-1:0] node30088;
	wire [16-1:0] node30089;
	wire [16-1:0] node30092;
	wire [16-1:0] node30095;
	wire [16-1:0] node30096;
	wire [16-1:0] node30097;
	wire [16-1:0] node30100;
	wire [16-1:0] node30103;
	wire [16-1:0] node30104;
	wire [16-1:0] node30107;
	wire [16-1:0] node30110;
	wire [16-1:0] node30111;
	wire [16-1:0] node30112;
	wire [16-1:0] node30113;
	wire [16-1:0] node30114;
	wire [16-1:0] node30115;
	wire [16-1:0] node30116;
	wire [16-1:0] node30117;
	wire [16-1:0] node30119;
	wire [16-1:0] node30122;
	wire [16-1:0] node30123;
	wire [16-1:0] node30127;
	wire [16-1:0] node30128;
	wire [16-1:0] node30129;
	wire [16-1:0] node30132;
	wire [16-1:0] node30135;
	wire [16-1:0] node30136;
	wire [16-1:0] node30139;
	wire [16-1:0] node30142;
	wire [16-1:0] node30143;
	wire [16-1:0] node30144;
	wire [16-1:0] node30145;
	wire [16-1:0] node30148;
	wire [16-1:0] node30151;
	wire [16-1:0] node30152;
	wire [16-1:0] node30155;
	wire [16-1:0] node30158;
	wire [16-1:0] node30159;
	wire [16-1:0] node30160;
	wire [16-1:0] node30163;
	wire [16-1:0] node30166;
	wire [16-1:0] node30167;
	wire [16-1:0] node30170;
	wire [16-1:0] node30173;
	wire [16-1:0] node30174;
	wire [16-1:0] node30175;
	wire [16-1:0] node30176;
	wire [16-1:0] node30177;
	wire [16-1:0] node30180;
	wire [16-1:0] node30183;
	wire [16-1:0] node30184;
	wire [16-1:0] node30187;
	wire [16-1:0] node30190;
	wire [16-1:0] node30191;
	wire [16-1:0] node30192;
	wire [16-1:0] node30195;
	wire [16-1:0] node30198;
	wire [16-1:0] node30200;
	wire [16-1:0] node30203;
	wire [16-1:0] node30204;
	wire [16-1:0] node30205;
	wire [16-1:0] node30207;
	wire [16-1:0] node30210;
	wire [16-1:0] node30211;
	wire [16-1:0] node30214;
	wire [16-1:0] node30217;
	wire [16-1:0] node30218;
	wire [16-1:0] node30220;
	wire [16-1:0] node30223;
	wire [16-1:0] node30225;
	wire [16-1:0] node30228;
	wire [16-1:0] node30229;
	wire [16-1:0] node30230;
	wire [16-1:0] node30231;
	wire [16-1:0] node30232;
	wire [16-1:0] node30233;
	wire [16-1:0] node30236;
	wire [16-1:0] node30239;
	wire [16-1:0] node30240;
	wire [16-1:0] node30243;
	wire [16-1:0] node30246;
	wire [16-1:0] node30247;
	wire [16-1:0] node30248;
	wire [16-1:0] node30251;
	wire [16-1:0] node30254;
	wire [16-1:0] node30255;
	wire [16-1:0] node30258;
	wire [16-1:0] node30261;
	wire [16-1:0] node30262;
	wire [16-1:0] node30263;
	wire [16-1:0] node30265;
	wire [16-1:0] node30268;
	wire [16-1:0] node30269;
	wire [16-1:0] node30272;
	wire [16-1:0] node30275;
	wire [16-1:0] node30276;
	wire [16-1:0] node30277;
	wire [16-1:0] node30280;
	wire [16-1:0] node30283;
	wire [16-1:0] node30284;
	wire [16-1:0] node30287;
	wire [16-1:0] node30290;
	wire [16-1:0] node30291;
	wire [16-1:0] node30292;
	wire [16-1:0] node30293;
	wire [16-1:0] node30294;
	wire [16-1:0] node30297;
	wire [16-1:0] node30300;
	wire [16-1:0] node30302;
	wire [16-1:0] node30305;
	wire [16-1:0] node30306;
	wire [16-1:0] node30307;
	wire [16-1:0] node30310;
	wire [16-1:0] node30313;
	wire [16-1:0] node30314;
	wire [16-1:0] node30317;
	wire [16-1:0] node30320;
	wire [16-1:0] node30321;
	wire [16-1:0] node30322;
	wire [16-1:0] node30323;
	wire [16-1:0] node30326;
	wire [16-1:0] node30329;
	wire [16-1:0] node30330;
	wire [16-1:0] node30333;
	wire [16-1:0] node30336;
	wire [16-1:0] node30337;
	wire [16-1:0] node30338;
	wire [16-1:0] node30341;
	wire [16-1:0] node30344;
	wire [16-1:0] node30345;
	wire [16-1:0] node30348;
	wire [16-1:0] node30351;
	wire [16-1:0] node30352;
	wire [16-1:0] node30353;
	wire [16-1:0] node30354;
	wire [16-1:0] node30355;
	wire [16-1:0] node30356;
	wire [16-1:0] node30357;
	wire [16-1:0] node30361;
	wire [16-1:0] node30363;
	wire [16-1:0] node30366;
	wire [16-1:0] node30367;
	wire [16-1:0] node30368;
	wire [16-1:0] node30371;
	wire [16-1:0] node30374;
	wire [16-1:0] node30375;
	wire [16-1:0] node30378;
	wire [16-1:0] node30381;
	wire [16-1:0] node30382;
	wire [16-1:0] node30383;
	wire [16-1:0] node30384;
	wire [16-1:0] node30387;
	wire [16-1:0] node30390;
	wire [16-1:0] node30391;
	wire [16-1:0] node30394;
	wire [16-1:0] node30397;
	wire [16-1:0] node30398;
	wire [16-1:0] node30399;
	wire [16-1:0] node30402;
	wire [16-1:0] node30405;
	wire [16-1:0] node30407;
	wire [16-1:0] node30410;
	wire [16-1:0] node30411;
	wire [16-1:0] node30412;
	wire [16-1:0] node30413;
	wire [16-1:0] node30414;
	wire [16-1:0] node30417;
	wire [16-1:0] node30420;
	wire [16-1:0] node30421;
	wire [16-1:0] node30424;
	wire [16-1:0] node30427;
	wire [16-1:0] node30428;
	wire [16-1:0] node30429;
	wire [16-1:0] node30432;
	wire [16-1:0] node30435;
	wire [16-1:0] node30436;
	wire [16-1:0] node30439;
	wire [16-1:0] node30442;
	wire [16-1:0] node30443;
	wire [16-1:0] node30444;
	wire [16-1:0] node30445;
	wire [16-1:0] node30448;
	wire [16-1:0] node30451;
	wire [16-1:0] node30452;
	wire [16-1:0] node30455;
	wire [16-1:0] node30458;
	wire [16-1:0] node30459;
	wire [16-1:0] node30461;
	wire [16-1:0] node30464;
	wire [16-1:0] node30465;
	wire [16-1:0] node30468;
	wire [16-1:0] node30471;
	wire [16-1:0] node30472;
	wire [16-1:0] node30473;
	wire [16-1:0] node30474;
	wire [16-1:0] node30476;
	wire [16-1:0] node30477;
	wire [16-1:0] node30480;
	wire [16-1:0] node30483;
	wire [16-1:0] node30484;
	wire [16-1:0] node30486;
	wire [16-1:0] node30489;
	wire [16-1:0] node30490;
	wire [16-1:0] node30493;
	wire [16-1:0] node30496;
	wire [16-1:0] node30497;
	wire [16-1:0] node30498;
	wire [16-1:0] node30499;
	wire [16-1:0] node30502;
	wire [16-1:0] node30505;
	wire [16-1:0] node30506;
	wire [16-1:0] node30509;
	wire [16-1:0] node30512;
	wire [16-1:0] node30513;
	wire [16-1:0] node30514;
	wire [16-1:0] node30517;
	wire [16-1:0] node30520;
	wire [16-1:0] node30521;
	wire [16-1:0] node30524;
	wire [16-1:0] node30527;
	wire [16-1:0] node30528;
	wire [16-1:0] node30529;
	wire [16-1:0] node30530;
	wire [16-1:0] node30532;
	wire [16-1:0] node30535;
	wire [16-1:0] node30536;
	wire [16-1:0] node30539;
	wire [16-1:0] node30542;
	wire [16-1:0] node30543;
	wire [16-1:0] node30544;
	wire [16-1:0] node30547;
	wire [16-1:0] node30550;
	wire [16-1:0] node30551;
	wire [16-1:0] node30554;
	wire [16-1:0] node30557;
	wire [16-1:0] node30558;
	wire [16-1:0] node30559;
	wire [16-1:0] node30560;
	wire [16-1:0] node30563;
	wire [16-1:0] node30566;
	wire [16-1:0] node30567;
	wire [16-1:0] node30570;
	wire [16-1:0] node30573;
	wire [16-1:0] node30574;
	wire [16-1:0] node30576;
	wire [16-1:0] node30579;
	wire [16-1:0] node30580;
	wire [16-1:0] node30583;
	wire [16-1:0] node30586;
	wire [16-1:0] node30587;
	wire [16-1:0] node30588;
	wire [16-1:0] node30589;
	wire [16-1:0] node30590;
	wire [16-1:0] node30591;
	wire [16-1:0] node30593;
	wire [16-1:0] node30594;
	wire [16-1:0] node30597;
	wire [16-1:0] node30600;
	wire [16-1:0] node30601;
	wire [16-1:0] node30602;
	wire [16-1:0] node30605;
	wire [16-1:0] node30608;
	wire [16-1:0] node30609;
	wire [16-1:0] node30612;
	wire [16-1:0] node30615;
	wire [16-1:0] node30616;
	wire [16-1:0] node30617;
	wire [16-1:0] node30618;
	wire [16-1:0] node30621;
	wire [16-1:0] node30624;
	wire [16-1:0] node30625;
	wire [16-1:0] node30628;
	wire [16-1:0] node30631;
	wire [16-1:0] node30632;
	wire [16-1:0] node30633;
	wire [16-1:0] node30636;
	wire [16-1:0] node30639;
	wire [16-1:0] node30640;
	wire [16-1:0] node30643;
	wire [16-1:0] node30646;
	wire [16-1:0] node30647;
	wire [16-1:0] node30648;
	wire [16-1:0] node30649;
	wire [16-1:0] node30650;
	wire [16-1:0] node30653;
	wire [16-1:0] node30656;
	wire [16-1:0] node30657;
	wire [16-1:0] node30660;
	wire [16-1:0] node30663;
	wire [16-1:0] node30664;
	wire [16-1:0] node30665;
	wire [16-1:0] node30668;
	wire [16-1:0] node30671;
	wire [16-1:0] node30672;
	wire [16-1:0] node30675;
	wire [16-1:0] node30678;
	wire [16-1:0] node30679;
	wire [16-1:0] node30680;
	wire [16-1:0] node30681;
	wire [16-1:0] node30684;
	wire [16-1:0] node30687;
	wire [16-1:0] node30688;
	wire [16-1:0] node30691;
	wire [16-1:0] node30694;
	wire [16-1:0] node30695;
	wire [16-1:0] node30696;
	wire [16-1:0] node30699;
	wire [16-1:0] node30702;
	wire [16-1:0] node30703;
	wire [16-1:0] node30706;
	wire [16-1:0] node30709;
	wire [16-1:0] node30710;
	wire [16-1:0] node30711;
	wire [16-1:0] node30712;
	wire [16-1:0] node30713;
	wire [16-1:0] node30714;
	wire [16-1:0] node30717;
	wire [16-1:0] node30720;
	wire [16-1:0] node30721;
	wire [16-1:0] node30724;
	wire [16-1:0] node30727;
	wire [16-1:0] node30728;
	wire [16-1:0] node30729;
	wire [16-1:0] node30732;
	wire [16-1:0] node30735;
	wire [16-1:0] node30736;
	wire [16-1:0] node30739;
	wire [16-1:0] node30742;
	wire [16-1:0] node30743;
	wire [16-1:0] node30744;
	wire [16-1:0] node30745;
	wire [16-1:0] node30748;
	wire [16-1:0] node30751;
	wire [16-1:0] node30753;
	wire [16-1:0] node30756;
	wire [16-1:0] node30758;
	wire [16-1:0] node30759;
	wire [16-1:0] node30762;
	wire [16-1:0] node30765;
	wire [16-1:0] node30766;
	wire [16-1:0] node30767;
	wire [16-1:0] node30768;
	wire [16-1:0] node30770;
	wire [16-1:0] node30773;
	wire [16-1:0] node30774;
	wire [16-1:0] node30778;
	wire [16-1:0] node30779;
	wire [16-1:0] node30780;
	wire [16-1:0] node30783;
	wire [16-1:0] node30786;
	wire [16-1:0] node30787;
	wire [16-1:0] node30790;
	wire [16-1:0] node30793;
	wire [16-1:0] node30794;
	wire [16-1:0] node30795;
	wire [16-1:0] node30796;
	wire [16-1:0] node30799;
	wire [16-1:0] node30802;
	wire [16-1:0] node30803;
	wire [16-1:0] node30806;
	wire [16-1:0] node30809;
	wire [16-1:0] node30810;
	wire [16-1:0] node30812;
	wire [16-1:0] node30815;
	wire [16-1:0] node30817;
	wire [16-1:0] node30820;
	wire [16-1:0] node30821;
	wire [16-1:0] node30822;
	wire [16-1:0] node30823;
	wire [16-1:0] node30824;
	wire [16-1:0] node30825;
	wire [16-1:0] node30828;
	wire [16-1:0] node30829;
	wire [16-1:0] node30832;
	wire [16-1:0] node30835;
	wire [16-1:0] node30836;
	wire [16-1:0] node30837;
	wire [16-1:0] node30840;
	wire [16-1:0] node30843;
	wire [16-1:0] node30844;
	wire [16-1:0] node30848;
	wire [16-1:0] node30849;
	wire [16-1:0] node30850;
	wire [16-1:0] node30851;
	wire [16-1:0] node30854;
	wire [16-1:0] node30857;
	wire [16-1:0] node30858;
	wire [16-1:0] node30861;
	wire [16-1:0] node30864;
	wire [16-1:0] node30865;
	wire [16-1:0] node30866;
	wire [16-1:0] node30869;
	wire [16-1:0] node30872;
	wire [16-1:0] node30873;
	wire [16-1:0] node30877;
	wire [16-1:0] node30878;
	wire [16-1:0] node30879;
	wire [16-1:0] node30880;
	wire [16-1:0] node30881;
	wire [16-1:0] node30884;
	wire [16-1:0] node30887;
	wire [16-1:0] node30888;
	wire [16-1:0] node30891;
	wire [16-1:0] node30894;
	wire [16-1:0] node30895;
	wire [16-1:0] node30896;
	wire [16-1:0] node30900;
	wire [16-1:0] node30901;
	wire [16-1:0] node30904;
	wire [16-1:0] node30907;
	wire [16-1:0] node30908;
	wire [16-1:0] node30909;
	wire [16-1:0] node30910;
	wire [16-1:0] node30913;
	wire [16-1:0] node30916;
	wire [16-1:0] node30917;
	wire [16-1:0] node30920;
	wire [16-1:0] node30923;
	wire [16-1:0] node30924;
	wire [16-1:0] node30925;
	wire [16-1:0] node30928;
	wire [16-1:0] node30931;
	wire [16-1:0] node30932;
	wire [16-1:0] node30935;
	wire [16-1:0] node30938;
	wire [16-1:0] node30939;
	wire [16-1:0] node30940;
	wire [16-1:0] node30941;
	wire [16-1:0] node30942;
	wire [16-1:0] node30943;
	wire [16-1:0] node30946;
	wire [16-1:0] node30949;
	wire [16-1:0] node30951;
	wire [16-1:0] node30954;
	wire [16-1:0] node30955;
	wire [16-1:0] node30956;
	wire [16-1:0] node30959;
	wire [16-1:0] node30962;
	wire [16-1:0] node30963;
	wire [16-1:0] node30966;
	wire [16-1:0] node30969;
	wire [16-1:0] node30970;
	wire [16-1:0] node30971;
	wire [16-1:0] node30972;
	wire [16-1:0] node30975;
	wire [16-1:0] node30978;
	wire [16-1:0] node30980;
	wire [16-1:0] node30983;
	wire [16-1:0] node30984;
	wire [16-1:0] node30985;
	wire [16-1:0] node30988;
	wire [16-1:0] node30991;
	wire [16-1:0] node30992;
	wire [16-1:0] node30995;
	wire [16-1:0] node30998;
	wire [16-1:0] node30999;
	wire [16-1:0] node31000;
	wire [16-1:0] node31001;
	wire [16-1:0] node31002;
	wire [16-1:0] node31005;
	wire [16-1:0] node31008;
	wire [16-1:0] node31009;
	wire [16-1:0] node31012;
	wire [16-1:0] node31015;
	wire [16-1:0] node31016;
	wire [16-1:0] node31017;
	wire [16-1:0] node31020;
	wire [16-1:0] node31023;
	wire [16-1:0] node31024;
	wire [16-1:0] node31027;
	wire [16-1:0] node31030;
	wire [16-1:0] node31031;
	wire [16-1:0] node31032;
	wire [16-1:0] node31034;
	wire [16-1:0] node31037;
	wire [16-1:0] node31038;
	wire [16-1:0] node31041;
	wire [16-1:0] node31044;
	wire [16-1:0] node31045;
	wire [16-1:0] node31046;
	wire [16-1:0] node31049;
	wire [16-1:0] node31052;
	wire [16-1:0] node31053;
	wire [16-1:0] node31056;

	assign outp = (inp[6]) ? node15558 : node1;
		assign node1 = (inp[1]) ? node7785 : node2;
			assign node2 = (inp[9]) ? node3888 : node3;
				assign node3 = (inp[13]) ? node1945 : node4;
					assign node4 = (inp[4]) ? node972 : node5;
						assign node5 = (inp[15]) ? node481 : node6;
							assign node6 = (inp[8]) ? node256 : node7;
								assign node7 = (inp[14]) ? node133 : node8;
									assign node8 = (inp[7]) ? node72 : node9;
										assign node9 = (inp[0]) ? node41 : node10;
											assign node10 = (inp[3]) ? node26 : node11;
												assign node11 = (inp[11]) ? node19 : node12;
													assign node12 = (inp[12]) ? node16 : node13;
														assign node13 = (inp[5]) ? 16'b0011111111111111 : 16'b0111111111111111;
														assign node16 = (inp[2]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node19 = (inp[12]) ? node23 : node20;
														assign node20 = (inp[5]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node23 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node26 = (inp[2]) ? node34 : node27;
													assign node27 = (inp[5]) ? node31 : node28;
														assign node28 = (inp[10]) ? 16'b0001111111111111 : 16'b0111111111111111;
														assign node31 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node34 = (inp[5]) ? node38 : node35;
														assign node35 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node38 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node41 = (inp[2]) ? node57 : node42;
												assign node42 = (inp[12]) ? node50 : node43;
													assign node43 = (inp[3]) ? node47 : node44;
														assign node44 = (inp[11]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node47 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node50 = (inp[3]) ? node54 : node51;
														assign node51 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node54 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node57 = (inp[10]) ? node65 : node58;
													assign node58 = (inp[12]) ? node62 : node59;
														assign node59 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node62 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node65 = (inp[11]) ? node69 : node66;
														assign node66 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node69 = (inp[5]) ? 16'b0000000111111111 : 16'b0000011111111111;
										assign node72 = (inp[10]) ? node102 : node73;
											assign node73 = (inp[3]) ? node87 : node74;
												assign node74 = (inp[0]) ? node80 : node75;
													assign node75 = (inp[12]) ? 16'b0000111111111111 : node76;
														assign node76 = (inp[11]) ? 16'b0001111111111111 : 16'b0011111111111111;
													assign node80 = (inp[5]) ? node84 : node81;
														assign node81 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node84 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node87 = (inp[11]) ? node95 : node88;
													assign node88 = (inp[5]) ? node92 : node89;
														assign node89 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node92 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node95 = (inp[12]) ? node99 : node96;
														assign node96 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node99 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node102 = (inp[2]) ? node118 : node103;
												assign node103 = (inp[3]) ? node111 : node104;
													assign node104 = (inp[12]) ? node108 : node105;
														assign node105 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node108 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node111 = (inp[5]) ? node115 : node112;
														assign node112 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node115 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node118 = (inp[0]) ? node126 : node119;
													assign node119 = (inp[3]) ? node123 : node120;
														assign node120 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node123 = (inp[11]) ? 16'b0000001111111111 : 16'b0000001111111111;
													assign node126 = (inp[12]) ? node130 : node127;
														assign node127 = (inp[3]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node130 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
									assign node133 = (inp[0]) ? node195 : node134;
										assign node134 = (inp[12]) ? node166 : node135;
											assign node135 = (inp[3]) ? node151 : node136;
												assign node136 = (inp[10]) ? node144 : node137;
													assign node137 = (inp[5]) ? node141 : node138;
														assign node138 = (inp[11]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node141 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node144 = (inp[5]) ? node148 : node145;
														assign node145 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node148 = (inp[11]) ? 16'b0000111111111111 : 16'b0000111111111111;
												assign node151 = (inp[10]) ? node159 : node152;
													assign node152 = (inp[7]) ? node156 : node153;
														assign node153 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node156 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node159 = (inp[11]) ? node163 : node160;
														assign node160 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node163 = (inp[2]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node166 = (inp[7]) ? node182 : node167;
												assign node167 = (inp[3]) ? node175 : node168;
													assign node168 = (inp[2]) ? node172 : node169;
														assign node169 = (inp[10]) ? 16'b0000111111111111 : 16'b0000111111111111;
														assign node172 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node175 = (inp[11]) ? node179 : node176;
														assign node176 = (inp[2]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node179 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node182 = (inp[10]) ? node188 : node183;
													assign node183 = (inp[5]) ? node185 : 16'b0000011111111111;
														assign node185 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node188 = (inp[2]) ? node192 : node189;
														assign node189 = (inp[11]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node192 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
										assign node195 = (inp[7]) ? node227 : node196;
											assign node196 = (inp[3]) ? node212 : node197;
												assign node197 = (inp[5]) ? node205 : node198;
													assign node198 = (inp[11]) ? node202 : node199;
														assign node199 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node202 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node205 = (inp[2]) ? node209 : node206;
														assign node206 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node209 = (inp[11]) ? 16'b0000001111111111 : 16'b0000001111111111;
												assign node212 = (inp[10]) ? node220 : node213;
													assign node213 = (inp[2]) ? node217 : node214;
														assign node214 = (inp[12]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node217 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node220 = (inp[11]) ? node224 : node221;
														assign node221 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node224 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node227 = (inp[5]) ? node243 : node228;
												assign node228 = (inp[10]) ? node236 : node229;
													assign node229 = (inp[12]) ? node233 : node230;
														assign node230 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node233 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node236 = (inp[11]) ? node240 : node237;
														assign node237 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node240 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node243 = (inp[11]) ? node249 : node244;
													assign node244 = (inp[3]) ? node246 : 16'b0000001111111111;
														assign node246 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node249 = (inp[2]) ? node253 : node250;
														assign node250 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node253 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
								assign node256 = (inp[5]) ? node372 : node257;
									assign node257 = (inp[2]) ? node313 : node258;
										assign node258 = (inp[11]) ? node288 : node259;
											assign node259 = (inp[10]) ? node275 : node260;
												assign node260 = (inp[7]) ? node268 : node261;
													assign node261 = (inp[0]) ? node265 : node262;
														assign node262 = (inp[3]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node265 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node268 = (inp[12]) ? node272 : node269;
														assign node269 = (inp[3]) ? 16'b0000111111111111 : 16'b0011111111111111;
														assign node272 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node275 = (inp[0]) ? node283 : node276;
													assign node276 = (inp[14]) ? node280 : node277;
														assign node277 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node280 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node283 = (inp[14]) ? node285 : 16'b0000111111111111;
														assign node285 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node288 = (inp[12]) ? node302 : node289;
												assign node289 = (inp[14]) ? node297 : node290;
													assign node290 = (inp[0]) ? node294 : node291;
														assign node291 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node294 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node297 = (inp[7]) ? 16'b0000011111111111 : node298;
														assign node298 = (inp[3]) ? 16'b0000011111111111 : 16'b0000011111111111;
												assign node302 = (inp[0]) ? node308 : node303;
													assign node303 = (inp[10]) ? node305 : 16'b0000011111111111;
														assign node305 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node308 = (inp[14]) ? 16'b0000001111111111 : node309;
														assign node309 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node313 = (inp[7]) ? node341 : node314;
											assign node314 = (inp[11]) ? node330 : node315;
												assign node315 = (inp[3]) ? node323 : node316;
													assign node316 = (inp[0]) ? node320 : node317;
														assign node317 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node320 = (inp[12]) ? 16'b0000011111111111 : 16'b0000011111111111;
													assign node323 = (inp[12]) ? node327 : node324;
														assign node324 = (inp[10]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node327 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node330 = (inp[14]) ? node336 : node331;
													assign node331 = (inp[0]) ? node333 : 16'b0000111111111111;
														assign node333 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node336 = (inp[10]) ? node338 : 16'b0000011111111111;
														assign node338 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node341 = (inp[0]) ? node357 : node342;
												assign node342 = (inp[10]) ? node350 : node343;
													assign node343 = (inp[3]) ? node347 : node344;
														assign node344 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node347 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node350 = (inp[12]) ? node354 : node351;
														assign node351 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node354 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node357 = (inp[3]) ? node365 : node358;
													assign node358 = (inp[14]) ? node362 : node359;
														assign node359 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node362 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node365 = (inp[12]) ? node369 : node366;
														assign node366 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node369 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
									assign node372 = (inp[2]) ? node426 : node373;
										assign node373 = (inp[7]) ? node401 : node374;
											assign node374 = (inp[3]) ? node388 : node375;
												assign node375 = (inp[11]) ? node381 : node376;
													assign node376 = (inp[12]) ? 16'b0000111111111111 : node377;
														assign node377 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node381 = (inp[12]) ? node385 : node382;
														assign node382 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node385 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node388 = (inp[12]) ? node396 : node389;
													assign node389 = (inp[14]) ? node393 : node390;
														assign node390 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node393 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node396 = (inp[14]) ? 16'b0000001111111111 : node397;
														assign node397 = (inp[11]) ? 16'b0000001111111111 : 16'b0000001111111111;
											assign node401 = (inp[11]) ? node411 : node402;
												assign node402 = (inp[14]) ? node406 : node403;
													assign node403 = (inp[3]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node406 = (inp[3]) ? 16'b0000001111111111 : node407;
														assign node407 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node411 = (inp[14]) ? node419 : node412;
													assign node412 = (inp[3]) ? node416 : node413;
														assign node413 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node416 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node419 = (inp[3]) ? node423 : node420;
														assign node420 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node423 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node426 = (inp[12]) ? node458 : node427;
											assign node427 = (inp[0]) ? node443 : node428;
												assign node428 = (inp[10]) ? node436 : node429;
													assign node429 = (inp[7]) ? node433 : node430;
														assign node430 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node433 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node436 = (inp[3]) ? node440 : node437;
														assign node437 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node440 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node443 = (inp[14]) ? node451 : node444;
													assign node444 = (inp[10]) ? node448 : node445;
														assign node445 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node448 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node451 = (inp[3]) ? node455 : node452;
														assign node452 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node455 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node458 = (inp[14]) ? node468 : node459;
												assign node459 = (inp[0]) ? node461 : 16'b0000001111111111;
													assign node461 = (inp[10]) ? node465 : node462;
														assign node462 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node465 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node468 = (inp[7]) ? node474 : node469;
													assign node469 = (inp[10]) ? node471 : 16'b0000001111111111;
														assign node471 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node474 = (inp[10]) ? node478 : node475;
														assign node475 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node478 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
							assign node481 = (inp[11]) ? node727 : node482;
								assign node482 = (inp[10]) ? node600 : node483;
									assign node483 = (inp[3]) ? node539 : node484;
										assign node484 = (inp[2]) ? node514 : node485;
											assign node485 = (inp[12]) ? node499 : node486;
												assign node486 = (inp[8]) ? node494 : node487;
													assign node487 = (inp[5]) ? node491 : node488;
														assign node488 = (inp[14]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node491 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node494 = (inp[0]) ? 16'b0000001111111111 : node495;
														assign node495 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
												assign node499 = (inp[0]) ? node507 : node500;
													assign node500 = (inp[7]) ? node504 : node501;
														assign node501 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node504 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node507 = (inp[5]) ? node511 : node508;
														assign node508 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node511 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node514 = (inp[7]) ? node526 : node515;
												assign node515 = (inp[5]) ? node521 : node516;
													assign node516 = (inp[0]) ? 16'b0000111111111111 : node517;
														assign node517 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node521 = (inp[12]) ? 16'b0000001111111111 : node522;
														assign node522 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node526 = (inp[0]) ? node534 : node527;
													assign node527 = (inp[12]) ? node531 : node528;
														assign node528 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node531 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node534 = (inp[12]) ? 16'b0000000111111111 : node535;
														assign node535 = (inp[8]) ? 16'b0000000111111111 : 16'b0000011111111111;
										assign node539 = (inp[12]) ? node571 : node540;
											assign node540 = (inp[7]) ? node556 : node541;
												assign node541 = (inp[0]) ? node549 : node542;
													assign node542 = (inp[14]) ? node546 : node543;
														assign node543 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node546 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node549 = (inp[8]) ? node553 : node550;
														assign node550 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node553 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node556 = (inp[14]) ? node564 : node557;
													assign node557 = (inp[5]) ? node561 : node558;
														assign node558 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node561 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node564 = (inp[8]) ? node568 : node565;
														assign node565 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node568 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node571 = (inp[0]) ? node585 : node572;
												assign node572 = (inp[14]) ? node580 : node573;
													assign node573 = (inp[2]) ? node577 : node574;
														assign node574 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node577 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node580 = (inp[2]) ? 16'b0000001111111111 : node581;
														assign node581 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node585 = (inp[14]) ? node593 : node586;
													assign node586 = (inp[5]) ? node590 : node587;
														assign node587 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node590 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node593 = (inp[5]) ? node597 : node594;
														assign node594 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node597 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node600 = (inp[7]) ? node664 : node601;
										assign node601 = (inp[0]) ? node633 : node602;
											assign node602 = (inp[14]) ? node618 : node603;
												assign node603 = (inp[8]) ? node611 : node604;
													assign node604 = (inp[5]) ? node608 : node605;
														assign node605 = (inp[12]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node608 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node611 = (inp[12]) ? node615 : node612;
														assign node612 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node615 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node618 = (inp[8]) ? node626 : node619;
													assign node619 = (inp[3]) ? node623 : node620;
														assign node620 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node623 = (inp[2]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node626 = (inp[12]) ? node630 : node627;
														assign node627 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node630 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node633 = (inp[8]) ? node649 : node634;
												assign node634 = (inp[2]) ? node642 : node635;
													assign node635 = (inp[5]) ? node639 : node636;
														assign node636 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node639 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node642 = (inp[5]) ? node646 : node643;
														assign node643 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node646 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node649 = (inp[14]) ? node657 : node650;
													assign node650 = (inp[3]) ? node654 : node651;
														assign node651 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node654 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node657 = (inp[12]) ? node661 : node658;
														assign node658 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node661 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node664 = (inp[3]) ? node696 : node665;
											assign node665 = (inp[2]) ? node681 : node666;
												assign node666 = (inp[8]) ? node674 : node667;
													assign node667 = (inp[14]) ? node671 : node668;
														assign node668 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node671 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node674 = (inp[5]) ? node678 : node675;
														assign node675 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node678 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node681 = (inp[14]) ? node689 : node682;
													assign node682 = (inp[12]) ? node686 : node683;
														assign node683 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node686 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node689 = (inp[12]) ? node693 : node690;
														assign node690 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node693 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node696 = (inp[5]) ? node712 : node697;
												assign node697 = (inp[8]) ? node705 : node698;
													assign node698 = (inp[2]) ? node702 : node699;
														assign node699 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node702 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node705 = (inp[0]) ? node709 : node706;
														assign node706 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node709 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node712 = (inp[8]) ? node720 : node713;
													assign node713 = (inp[14]) ? node717 : node714;
														assign node714 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node717 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node720 = (inp[14]) ? node724 : node721;
														assign node721 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node724 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
								assign node727 = (inp[2]) ? node849 : node728;
									assign node728 = (inp[7]) ? node790 : node729;
										assign node729 = (inp[12]) ? node761 : node730;
											assign node730 = (inp[5]) ? node746 : node731;
												assign node731 = (inp[10]) ? node739 : node732;
													assign node732 = (inp[14]) ? node736 : node733;
														assign node733 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node736 = (inp[3]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node739 = (inp[3]) ? node743 : node740;
														assign node740 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node743 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node746 = (inp[8]) ? node754 : node747;
													assign node747 = (inp[14]) ? node751 : node748;
														assign node748 = (inp[0]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node751 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node754 = (inp[0]) ? node758 : node755;
														assign node755 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node758 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node761 = (inp[8]) ? node777 : node762;
												assign node762 = (inp[0]) ? node770 : node763;
													assign node763 = (inp[3]) ? node767 : node764;
														assign node764 = (inp[5]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node767 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node770 = (inp[5]) ? node774 : node771;
														assign node771 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node774 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node777 = (inp[3]) ? node785 : node778;
													assign node778 = (inp[14]) ? node782 : node779;
														assign node779 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node782 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node785 = (inp[5]) ? node787 : 16'b0000000111111111;
														assign node787 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node790 = (inp[3]) ? node820 : node791;
											assign node791 = (inp[10]) ? node805 : node792;
												assign node792 = (inp[0]) ? node800 : node793;
													assign node793 = (inp[5]) ? node797 : node794;
														assign node794 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node797 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node800 = (inp[12]) ? 16'b0000000111111111 : node801;
														assign node801 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node805 = (inp[14]) ? node813 : node806;
													assign node806 = (inp[12]) ? node810 : node807;
														assign node807 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node810 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node813 = (inp[0]) ? node817 : node814;
														assign node814 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node817 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node820 = (inp[5]) ? node834 : node821;
												assign node821 = (inp[14]) ? node827 : node822;
													assign node822 = (inp[12]) ? 16'b0000001111111111 : node823;
														assign node823 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node827 = (inp[12]) ? node831 : node828;
														assign node828 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node831 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node834 = (inp[0]) ? node842 : node835;
													assign node835 = (inp[14]) ? node839 : node836;
														assign node836 = (inp[12]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node839 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node842 = (inp[12]) ? node846 : node843;
														assign node843 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node846 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node849 = (inp[8]) ? node911 : node850;
										assign node850 = (inp[3]) ? node882 : node851;
											assign node851 = (inp[5]) ? node867 : node852;
												assign node852 = (inp[0]) ? node860 : node853;
													assign node853 = (inp[7]) ? node857 : node854;
														assign node854 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node857 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node860 = (inp[12]) ? node864 : node861;
														assign node861 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node864 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000111111111;
												assign node867 = (inp[7]) ? node875 : node868;
													assign node868 = (inp[12]) ? node872 : node869;
														assign node869 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node872 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node875 = (inp[14]) ? node879 : node876;
														assign node876 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node879 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node882 = (inp[10]) ? node896 : node883;
												assign node883 = (inp[14]) ? node891 : node884;
													assign node884 = (inp[0]) ? node888 : node885;
														assign node885 = (inp[7]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node888 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node891 = (inp[7]) ? 16'b0000000111111111 : node892;
														assign node892 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node896 = (inp[7]) ? node904 : node897;
													assign node897 = (inp[12]) ? node901 : node898;
														assign node898 = (inp[0]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node901 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node904 = (inp[5]) ? node908 : node905;
														assign node905 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node908 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
										assign node911 = (inp[10]) ? node941 : node912;
											assign node912 = (inp[7]) ? node928 : node913;
												assign node913 = (inp[12]) ? node921 : node914;
													assign node914 = (inp[3]) ? node918 : node915;
														assign node915 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node918 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node921 = (inp[5]) ? node925 : node922;
														assign node922 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node925 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node928 = (inp[0]) ? node936 : node929;
													assign node929 = (inp[5]) ? node933 : node930;
														assign node930 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node933 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node936 = (inp[3]) ? node938 : 16'b0000000011111111;
														assign node938 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node941 = (inp[0]) ? node957 : node942;
												assign node942 = (inp[14]) ? node950 : node943;
													assign node943 = (inp[5]) ? node947 : node944;
														assign node944 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node947 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node950 = (inp[7]) ? node954 : node951;
														assign node951 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node954 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node957 = (inp[12]) ? node965 : node958;
													assign node958 = (inp[5]) ? node962 : node959;
														assign node959 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node962 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node965 = (inp[3]) ? node969 : node966;
														assign node966 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node969 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
						assign node972 = (inp[11]) ? node1470 : node973;
							assign node973 = (inp[5]) ? node1223 : node974;
								assign node974 = (inp[15]) ? node1102 : node975;
									assign node975 = (inp[14]) ? node1039 : node976;
										assign node976 = (inp[12]) ? node1008 : node977;
											assign node977 = (inp[7]) ? node993 : node978;
												assign node978 = (inp[0]) ? node986 : node979;
													assign node979 = (inp[3]) ? node983 : node980;
														assign node980 = (inp[8]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node983 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node986 = (inp[10]) ? node990 : node987;
														assign node987 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node990 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node993 = (inp[8]) ? node1001 : node994;
													assign node994 = (inp[0]) ? node998 : node995;
														assign node995 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node998 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1001 = (inp[2]) ? node1005 : node1002;
														assign node1002 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1005 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1008 = (inp[10]) ? node1024 : node1009;
												assign node1009 = (inp[3]) ? node1017 : node1010;
													assign node1010 = (inp[7]) ? node1014 : node1011;
														assign node1011 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1014 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1017 = (inp[7]) ? node1021 : node1018;
														assign node1018 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1021 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1024 = (inp[3]) ? node1032 : node1025;
													assign node1025 = (inp[7]) ? node1029 : node1026;
														assign node1026 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1029 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1032 = (inp[8]) ? node1036 : node1033;
														assign node1033 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1036 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node1039 = (inp[7]) ? node1071 : node1040;
											assign node1040 = (inp[10]) ? node1056 : node1041;
												assign node1041 = (inp[8]) ? node1049 : node1042;
													assign node1042 = (inp[12]) ? node1046 : node1043;
														assign node1043 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1046 = (inp[0]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node1049 = (inp[3]) ? node1053 : node1050;
														assign node1050 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1053 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1056 = (inp[2]) ? node1064 : node1057;
													assign node1057 = (inp[12]) ? node1061 : node1058;
														assign node1058 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1061 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1064 = (inp[8]) ? node1068 : node1065;
														assign node1065 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1068 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1071 = (inp[2]) ? node1087 : node1072;
												assign node1072 = (inp[3]) ? node1080 : node1073;
													assign node1073 = (inp[10]) ? node1077 : node1074;
														assign node1074 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1077 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1080 = (inp[8]) ? node1084 : node1081;
														assign node1081 = (inp[12]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node1084 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1087 = (inp[8]) ? node1095 : node1088;
													assign node1088 = (inp[3]) ? node1092 : node1089;
														assign node1089 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1092 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node1095 = (inp[0]) ? node1099 : node1096;
														assign node1096 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1099 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
									assign node1102 = (inp[12]) ? node1164 : node1103;
										assign node1103 = (inp[8]) ? node1133 : node1104;
											assign node1104 = (inp[14]) ? node1118 : node1105;
												assign node1105 = (inp[3]) ? node1113 : node1106;
													assign node1106 = (inp[0]) ? node1110 : node1107;
														assign node1107 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1110 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1113 = (inp[2]) ? 16'b0000011111111111 : node1114;
														assign node1114 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1118 = (inp[7]) ? node1126 : node1119;
													assign node1119 = (inp[0]) ? node1123 : node1120;
														assign node1120 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1123 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1126 = (inp[10]) ? node1130 : node1127;
														assign node1127 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1130 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
											assign node1133 = (inp[14]) ? node1149 : node1134;
												assign node1134 = (inp[10]) ? node1142 : node1135;
													assign node1135 = (inp[3]) ? node1139 : node1136;
														assign node1136 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1139 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1142 = (inp[2]) ? node1146 : node1143;
														assign node1143 = (inp[3]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node1146 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1149 = (inp[2]) ? node1157 : node1150;
													assign node1150 = (inp[3]) ? node1154 : node1151;
														assign node1151 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1154 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1157 = (inp[0]) ? node1161 : node1158;
														assign node1158 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node1161 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node1164 = (inp[7]) ? node1192 : node1165;
											assign node1165 = (inp[14]) ? node1181 : node1166;
												assign node1166 = (inp[3]) ? node1174 : node1167;
													assign node1167 = (inp[10]) ? node1171 : node1168;
														assign node1168 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1171 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1174 = (inp[2]) ? node1178 : node1175;
														assign node1175 = (inp[10]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node1178 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node1181 = (inp[0]) ? node1187 : node1182;
													assign node1182 = (inp[8]) ? node1184 : 16'b0000001111111111;
														assign node1184 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1187 = (inp[3]) ? 16'b0000000111111111 : node1188;
														assign node1188 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1192 = (inp[3]) ? node1208 : node1193;
												assign node1193 = (inp[2]) ? node1201 : node1194;
													assign node1194 = (inp[8]) ? node1198 : node1195;
														assign node1195 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1198 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1201 = (inp[0]) ? node1205 : node1202;
														assign node1202 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node1205 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node1208 = (inp[0]) ? node1216 : node1209;
													assign node1209 = (inp[2]) ? node1213 : node1210;
														assign node1210 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node1213 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1216 = (inp[8]) ? node1220 : node1217;
														assign node1217 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1220 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node1223 = (inp[12]) ? node1351 : node1224;
									assign node1224 = (inp[7]) ? node1288 : node1225;
										assign node1225 = (inp[2]) ? node1257 : node1226;
											assign node1226 = (inp[15]) ? node1242 : node1227;
												assign node1227 = (inp[14]) ? node1235 : node1228;
													assign node1228 = (inp[0]) ? node1232 : node1229;
														assign node1229 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1232 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1235 = (inp[0]) ? node1239 : node1236;
														assign node1236 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1239 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1242 = (inp[0]) ? node1250 : node1243;
													assign node1243 = (inp[8]) ? node1247 : node1244;
														assign node1244 = (inp[3]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node1247 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1250 = (inp[10]) ? node1254 : node1251;
														assign node1251 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1254 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1257 = (inp[14]) ? node1273 : node1258;
												assign node1258 = (inp[8]) ? node1266 : node1259;
													assign node1259 = (inp[3]) ? node1263 : node1260;
														assign node1260 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1263 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1266 = (inp[0]) ? node1270 : node1267;
														assign node1267 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1270 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1273 = (inp[3]) ? node1281 : node1274;
													assign node1274 = (inp[15]) ? node1278 : node1275;
														assign node1275 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1278 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1281 = (inp[10]) ? node1285 : node1282;
														assign node1282 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1285 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1288 = (inp[0]) ? node1320 : node1289;
											assign node1289 = (inp[10]) ? node1305 : node1290;
												assign node1290 = (inp[3]) ? node1298 : node1291;
													assign node1291 = (inp[2]) ? node1295 : node1292;
														assign node1292 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1295 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1298 = (inp[8]) ? node1302 : node1299;
														assign node1299 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1302 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1305 = (inp[8]) ? node1313 : node1306;
													assign node1306 = (inp[2]) ? node1310 : node1307;
														assign node1307 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1310 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1313 = (inp[2]) ? node1317 : node1314;
														assign node1314 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1317 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1320 = (inp[3]) ? node1336 : node1321;
												assign node1321 = (inp[10]) ? node1329 : node1322;
													assign node1322 = (inp[14]) ? node1326 : node1323;
														assign node1323 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1326 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1329 = (inp[14]) ? node1333 : node1330;
														assign node1330 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1333 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1336 = (inp[8]) ? node1344 : node1337;
													assign node1337 = (inp[14]) ? node1341 : node1338;
														assign node1338 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1341 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1344 = (inp[2]) ? node1348 : node1345;
														assign node1345 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1348 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
									assign node1351 = (inp[2]) ? node1411 : node1352;
										assign node1352 = (inp[8]) ? node1382 : node1353;
											assign node1353 = (inp[3]) ? node1367 : node1354;
												assign node1354 = (inp[0]) ? node1360 : node1355;
													assign node1355 = (inp[7]) ? node1357 : 16'b0000111111111111;
														assign node1357 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1360 = (inp[14]) ? node1364 : node1361;
														assign node1361 = (inp[10]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node1364 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1367 = (inp[15]) ? node1375 : node1368;
													assign node1368 = (inp[10]) ? node1372 : node1369;
														assign node1369 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1372 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1375 = (inp[7]) ? node1379 : node1376;
														assign node1376 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1379 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node1382 = (inp[15]) ? node1396 : node1383;
												assign node1383 = (inp[3]) ? node1389 : node1384;
													assign node1384 = (inp[14]) ? node1386 : 16'b0000011111111111;
														assign node1386 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1389 = (inp[0]) ? node1393 : node1390;
														assign node1390 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1393 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1396 = (inp[10]) ? node1404 : node1397;
													assign node1397 = (inp[0]) ? node1401 : node1398;
														assign node1398 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1401 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1404 = (inp[14]) ? node1408 : node1405;
														assign node1405 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1408 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1411 = (inp[8]) ? node1441 : node1412;
											assign node1412 = (inp[7]) ? node1428 : node1413;
												assign node1413 = (inp[14]) ? node1421 : node1414;
													assign node1414 = (inp[3]) ? node1418 : node1415;
														assign node1415 = (inp[15]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node1418 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1421 = (inp[3]) ? node1425 : node1422;
														assign node1422 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1425 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1428 = (inp[0]) ? node1434 : node1429;
													assign node1429 = (inp[10]) ? node1431 : 16'b0000001111111111;
														assign node1431 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1434 = (inp[15]) ? node1438 : node1435;
														assign node1435 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node1438 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1441 = (inp[15]) ? node1457 : node1442;
												assign node1442 = (inp[3]) ? node1450 : node1443;
													assign node1443 = (inp[14]) ? node1447 : node1444;
														assign node1444 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node1447 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node1450 = (inp[7]) ? node1454 : node1451;
														assign node1451 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node1454 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node1457 = (inp[7]) ? node1463 : node1458;
													assign node1458 = (inp[10]) ? node1460 : 16'b0000000011111111;
														assign node1460 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1463 = (inp[3]) ? node1467 : node1464;
														assign node1464 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node1467 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node1470 = (inp[0]) ? node1710 : node1471;
								assign node1471 = (inp[8]) ? node1593 : node1472;
									assign node1472 = (inp[7]) ? node1530 : node1473;
										assign node1473 = (inp[15]) ? node1503 : node1474;
											assign node1474 = (inp[12]) ? node1490 : node1475;
												assign node1475 = (inp[3]) ? node1483 : node1476;
													assign node1476 = (inp[5]) ? node1480 : node1477;
														assign node1477 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1480 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1483 = (inp[10]) ? node1487 : node1484;
														assign node1484 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1487 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1490 = (inp[2]) ? node1498 : node1491;
													assign node1491 = (inp[10]) ? node1495 : node1492;
														assign node1492 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1495 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1498 = (inp[5]) ? 16'b0000001111111111 : node1499;
														assign node1499 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1503 = (inp[3]) ? node1517 : node1504;
												assign node1504 = (inp[14]) ? node1510 : node1505;
													assign node1505 = (inp[12]) ? 16'b0000011111111111 : node1506;
														assign node1506 = (inp[2]) ? 16'b0000011111111111 : 16'b0000011111111111;
													assign node1510 = (inp[12]) ? node1514 : node1511;
														assign node1511 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1514 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1517 = (inp[10]) ? node1523 : node1518;
													assign node1518 = (inp[5]) ? 16'b0000000111111111 : node1519;
														assign node1519 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1523 = (inp[2]) ? node1527 : node1524;
														assign node1524 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1527 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node1530 = (inp[3]) ? node1562 : node1531;
											assign node1531 = (inp[15]) ? node1547 : node1532;
												assign node1532 = (inp[10]) ? node1540 : node1533;
													assign node1533 = (inp[2]) ? node1537 : node1534;
														assign node1534 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1537 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1540 = (inp[12]) ? node1544 : node1541;
														assign node1541 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1544 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1547 = (inp[14]) ? node1555 : node1548;
													assign node1548 = (inp[2]) ? node1552 : node1549;
														assign node1549 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1552 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1555 = (inp[10]) ? node1559 : node1556;
														assign node1556 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1559 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node1562 = (inp[5]) ? node1578 : node1563;
												assign node1563 = (inp[12]) ? node1571 : node1564;
													assign node1564 = (inp[10]) ? node1568 : node1565;
														assign node1565 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1568 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1571 = (inp[15]) ? node1575 : node1572;
														assign node1572 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node1575 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1578 = (inp[2]) ? node1586 : node1579;
													assign node1579 = (inp[14]) ? node1583 : node1580;
														assign node1580 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node1583 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1586 = (inp[12]) ? node1590 : node1587;
														assign node1587 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1590 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node1593 = (inp[5]) ? node1651 : node1594;
										assign node1594 = (inp[15]) ? node1626 : node1595;
											assign node1595 = (inp[2]) ? node1611 : node1596;
												assign node1596 = (inp[7]) ? node1604 : node1597;
													assign node1597 = (inp[12]) ? node1601 : node1598;
														assign node1598 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1601 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1604 = (inp[10]) ? node1608 : node1605;
														assign node1605 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1608 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node1611 = (inp[12]) ? node1619 : node1612;
													assign node1612 = (inp[7]) ? node1616 : node1613;
														assign node1613 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node1616 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1619 = (inp[14]) ? node1623 : node1620;
														assign node1620 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1623 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node1626 = (inp[14]) ? node1642 : node1627;
												assign node1627 = (inp[2]) ? node1635 : node1628;
													assign node1628 = (inp[7]) ? node1632 : node1629;
														assign node1629 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1632 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1635 = (inp[12]) ? node1639 : node1636;
														assign node1636 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1639 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node1642 = (inp[2]) ? node1648 : node1643;
													assign node1643 = (inp[10]) ? node1645 : 16'b0000000111111111;
														assign node1645 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1648 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node1651 = (inp[7]) ? node1681 : node1652;
											assign node1652 = (inp[15]) ? node1668 : node1653;
												assign node1653 = (inp[12]) ? node1661 : node1654;
													assign node1654 = (inp[2]) ? node1658 : node1655;
														assign node1655 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1658 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1661 = (inp[10]) ? node1665 : node1662;
														assign node1662 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1665 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1668 = (inp[12]) ? node1676 : node1669;
													assign node1669 = (inp[3]) ? node1673 : node1670;
														assign node1670 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1673 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node1676 = (inp[14]) ? 16'b0000000001111111 : node1677;
														assign node1677 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node1681 = (inp[10]) ? node1695 : node1682;
												assign node1682 = (inp[3]) ? node1688 : node1683;
													assign node1683 = (inp[2]) ? node1685 : 16'b0000000111111111;
														assign node1685 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node1688 = (inp[15]) ? node1692 : node1689;
														assign node1689 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node1692 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node1695 = (inp[15]) ? node1703 : node1696;
													assign node1696 = (inp[3]) ? node1700 : node1697;
														assign node1697 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node1700 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1703 = (inp[12]) ? node1707 : node1704;
														assign node1704 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node1707 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
								assign node1710 = (inp[14]) ? node1824 : node1711;
									assign node1711 = (inp[15]) ? node1761 : node1712;
										assign node1712 = (inp[2]) ? node1732 : node1713;
											assign node1713 = (inp[12]) ? node1725 : node1714;
												assign node1714 = (inp[8]) ? node1720 : node1715;
													assign node1715 = (inp[7]) ? node1717 : 16'b0000111111111111;
														assign node1717 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node1720 = (inp[3]) ? 16'b0000001111111111 : node1721;
														assign node1721 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1725 = (inp[3]) ? node1727 : 16'b0000001111111111;
													assign node1727 = (inp[10]) ? 16'b0000000111111111 : node1728;
														assign node1728 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node1732 = (inp[5]) ? node1746 : node1733;
												assign node1733 = (inp[10]) ? node1739 : node1734;
													assign node1734 = (inp[7]) ? node1736 : 16'b0000011111111111;
														assign node1736 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1739 = (inp[12]) ? node1743 : node1740;
														assign node1740 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1743 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node1746 = (inp[8]) ? node1754 : node1747;
													assign node1747 = (inp[12]) ? node1751 : node1748;
														assign node1748 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1751 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1754 = (inp[7]) ? node1758 : node1755;
														assign node1755 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node1758 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1761 = (inp[5]) ? node1793 : node1762;
											assign node1762 = (inp[12]) ? node1778 : node1763;
												assign node1763 = (inp[3]) ? node1771 : node1764;
													assign node1764 = (inp[7]) ? node1768 : node1765;
														assign node1765 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1768 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1771 = (inp[7]) ? node1775 : node1772;
														assign node1772 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1775 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node1778 = (inp[7]) ? node1786 : node1779;
													assign node1779 = (inp[10]) ? node1783 : node1780;
														assign node1780 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node1783 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1786 = (inp[8]) ? node1790 : node1787;
														assign node1787 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1790 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node1793 = (inp[12]) ? node1809 : node1794;
												assign node1794 = (inp[10]) ? node1802 : node1795;
													assign node1795 = (inp[3]) ? node1799 : node1796;
														assign node1796 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1799 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node1802 = (inp[3]) ? node1806 : node1803;
														assign node1803 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1806 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node1809 = (inp[2]) ? node1817 : node1810;
													assign node1810 = (inp[7]) ? node1814 : node1811;
														assign node1811 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1814 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1817 = (inp[10]) ? node1821 : node1818;
														assign node1818 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node1821 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
									assign node1824 = (inp[3]) ? node1884 : node1825;
										assign node1825 = (inp[10]) ? node1855 : node1826;
											assign node1826 = (inp[2]) ? node1842 : node1827;
												assign node1827 = (inp[12]) ? node1835 : node1828;
													assign node1828 = (inp[5]) ? node1832 : node1829;
														assign node1829 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node1832 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node1835 = (inp[15]) ? node1839 : node1836;
														assign node1836 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1839 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node1842 = (inp[8]) ? node1850 : node1843;
													assign node1843 = (inp[15]) ? node1847 : node1844;
														assign node1844 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1847 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node1850 = (inp[7]) ? node1852 : 16'b0000000011111111;
														assign node1852 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node1855 = (inp[2]) ? node1871 : node1856;
												assign node1856 = (inp[12]) ? node1864 : node1857;
													assign node1857 = (inp[7]) ? node1861 : node1858;
														assign node1858 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node1861 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node1864 = (inp[15]) ? node1868 : node1865;
														assign node1865 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node1868 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node1871 = (inp[8]) ? node1877 : node1872;
													assign node1872 = (inp[12]) ? node1874 : 16'b0000000011111111;
														assign node1874 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1877 = (inp[5]) ? node1881 : node1878;
														assign node1878 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node1881 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node1884 = (inp[15]) ? node1914 : node1885;
											assign node1885 = (inp[10]) ? node1899 : node1886;
												assign node1886 = (inp[7]) ? node1892 : node1887;
													assign node1887 = (inp[5]) ? node1889 : 16'b0000000111111111;
														assign node1889 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node1892 = (inp[5]) ? node1896 : node1893;
														assign node1893 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1896 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node1899 = (inp[12]) ? node1907 : node1900;
													assign node1900 = (inp[2]) ? node1904 : node1901;
														assign node1901 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1904 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1907 = (inp[8]) ? node1911 : node1908;
														assign node1908 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node1911 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node1914 = (inp[7]) ? node1930 : node1915;
												assign node1915 = (inp[5]) ? node1923 : node1916;
													assign node1916 = (inp[8]) ? node1920 : node1917;
														assign node1917 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node1920 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node1923 = (inp[12]) ? node1927 : node1924;
														assign node1924 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node1927 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node1930 = (inp[12]) ? node1938 : node1931;
													assign node1931 = (inp[8]) ? node1935 : node1932;
														assign node1932 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node1935 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node1938 = (inp[5]) ? node1942 : node1939;
														assign node1939 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node1942 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000011111;
					assign node1945 = (inp[12]) ? node2911 : node1946;
						assign node1946 = (inp[14]) ? node2440 : node1947;
							assign node1947 = (inp[7]) ? node2195 : node1948;
								assign node1948 = (inp[15]) ? node2070 : node1949;
									assign node1949 = (inp[2]) ? node2013 : node1950;
										assign node1950 = (inp[3]) ? node1982 : node1951;
											assign node1951 = (inp[4]) ? node1967 : node1952;
												assign node1952 = (inp[11]) ? node1960 : node1953;
													assign node1953 = (inp[5]) ? node1957 : node1954;
														assign node1954 = (inp[10]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node1957 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node1960 = (inp[10]) ? node1964 : node1961;
														assign node1961 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1964 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node1967 = (inp[8]) ? node1975 : node1968;
													assign node1968 = (inp[5]) ? node1972 : node1969;
														assign node1969 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1972 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node1975 = (inp[11]) ? node1979 : node1976;
														assign node1976 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1979 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node1982 = (inp[11]) ? node1998 : node1983;
												assign node1983 = (inp[8]) ? node1991 : node1984;
													assign node1984 = (inp[10]) ? node1988 : node1985;
														assign node1985 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node1988 = (inp[0]) ? 16'b0000001111111111 : 16'b0000111111111111;
													assign node1991 = (inp[10]) ? node1995 : node1992;
														assign node1992 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node1995 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node1998 = (inp[8]) ? node2006 : node1999;
													assign node1999 = (inp[5]) ? node2003 : node2000;
														assign node2000 = (inp[10]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node2003 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2006 = (inp[0]) ? node2010 : node2007;
														assign node2007 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2010 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2013 = (inp[5]) ? node2041 : node2014;
											assign node2014 = (inp[4]) ? node2028 : node2015;
												assign node2015 = (inp[8]) ? node2023 : node2016;
													assign node2016 = (inp[3]) ? node2020 : node2017;
														assign node2017 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node2020 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2023 = (inp[11]) ? 16'b0000011111111111 : node2024;
														assign node2024 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node2028 = (inp[11]) ? node2034 : node2029;
													assign node2029 = (inp[3]) ? node2031 : 16'b0000111111111111;
														assign node2031 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2034 = (inp[3]) ? node2038 : node2035;
														assign node2035 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2038 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node2041 = (inp[11]) ? node2057 : node2042;
												assign node2042 = (inp[0]) ? node2050 : node2043;
													assign node2043 = (inp[4]) ? node2047 : node2044;
														assign node2044 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2047 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2050 = (inp[8]) ? node2054 : node2051;
														assign node2051 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2054 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2057 = (inp[8]) ? node2063 : node2058;
													assign node2058 = (inp[4]) ? 16'b0000001111111111 : node2059;
														assign node2059 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2063 = (inp[4]) ? node2067 : node2064;
														assign node2064 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2067 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
									assign node2070 = (inp[10]) ? node2134 : node2071;
										assign node2071 = (inp[5]) ? node2103 : node2072;
											assign node2072 = (inp[8]) ? node2088 : node2073;
												assign node2073 = (inp[2]) ? node2081 : node2074;
													assign node2074 = (inp[0]) ? node2078 : node2075;
														assign node2075 = (inp[4]) ? 16'b0000111111111111 : 16'b0000111111111111;
														assign node2078 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2081 = (inp[0]) ? node2085 : node2082;
														assign node2082 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2085 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2088 = (inp[11]) ? node2096 : node2089;
													assign node2089 = (inp[2]) ? node2093 : node2090;
														assign node2090 = (inp[0]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node2093 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2096 = (inp[0]) ? node2100 : node2097;
														assign node2097 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2100 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2103 = (inp[3]) ? node2119 : node2104;
												assign node2104 = (inp[11]) ? node2112 : node2105;
													assign node2105 = (inp[4]) ? node2109 : node2106;
														assign node2106 = (inp[2]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node2109 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2112 = (inp[0]) ? node2116 : node2113;
														assign node2113 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2116 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node2119 = (inp[2]) ? node2127 : node2120;
													assign node2120 = (inp[0]) ? node2124 : node2121;
														assign node2121 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2124 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2127 = (inp[4]) ? node2131 : node2128;
														assign node2128 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node2131 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2134 = (inp[8]) ? node2164 : node2135;
											assign node2135 = (inp[3]) ? node2151 : node2136;
												assign node2136 = (inp[5]) ? node2144 : node2137;
													assign node2137 = (inp[0]) ? node2141 : node2138;
														assign node2138 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2141 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2144 = (inp[4]) ? node2148 : node2145;
														assign node2145 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2148 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node2151 = (inp[2]) ? node2157 : node2152;
													assign node2152 = (inp[5]) ? 16'b0000001111111111 : node2153;
														assign node2153 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2157 = (inp[0]) ? node2161 : node2158;
														assign node2158 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2161 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node2164 = (inp[2]) ? node2180 : node2165;
												assign node2165 = (inp[11]) ? node2173 : node2166;
													assign node2166 = (inp[5]) ? node2170 : node2167;
														assign node2167 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2170 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2173 = (inp[3]) ? node2177 : node2174;
														assign node2174 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2177 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2180 = (inp[11]) ? node2188 : node2181;
													assign node2181 = (inp[0]) ? node2185 : node2182;
														assign node2182 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2185 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2188 = (inp[5]) ? node2192 : node2189;
														assign node2189 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2192 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
								assign node2195 = (inp[4]) ? node2319 : node2196;
									assign node2196 = (inp[0]) ? node2256 : node2197;
										assign node2197 = (inp[3]) ? node2229 : node2198;
											assign node2198 = (inp[15]) ? node2214 : node2199;
												assign node2199 = (inp[8]) ? node2207 : node2200;
													assign node2200 = (inp[10]) ? node2204 : node2201;
														assign node2201 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node2204 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2207 = (inp[10]) ? node2211 : node2208;
														assign node2208 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2211 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2214 = (inp[2]) ? node2222 : node2215;
													assign node2215 = (inp[5]) ? node2219 : node2216;
														assign node2216 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2219 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2222 = (inp[8]) ? node2226 : node2223;
														assign node2223 = (inp[10]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node2226 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node2229 = (inp[5]) ? node2245 : node2230;
												assign node2230 = (inp[8]) ? node2238 : node2231;
													assign node2231 = (inp[10]) ? node2235 : node2232;
														assign node2232 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2235 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2238 = (inp[15]) ? node2242 : node2239;
														assign node2239 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2242 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2245 = (inp[11]) ? node2251 : node2246;
													assign node2246 = (inp[8]) ? 16'b0000001111111111 : node2247;
														assign node2247 = (inp[10]) ? 16'b0000001111111111 : 16'b0000001111111111;
													assign node2251 = (inp[15]) ? 16'b0000000111111111 : node2252;
														assign node2252 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2256 = (inp[3]) ? node2288 : node2257;
											assign node2257 = (inp[10]) ? node2273 : node2258;
												assign node2258 = (inp[11]) ? node2266 : node2259;
													assign node2259 = (inp[8]) ? node2263 : node2260;
														assign node2260 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2263 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2266 = (inp[8]) ? node2270 : node2267;
														assign node2267 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2270 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2273 = (inp[2]) ? node2281 : node2274;
													assign node2274 = (inp[11]) ? node2278 : node2275;
														assign node2275 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2278 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2281 = (inp[8]) ? node2285 : node2282;
														assign node2282 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node2285 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2288 = (inp[10]) ? node2304 : node2289;
												assign node2289 = (inp[5]) ? node2297 : node2290;
													assign node2290 = (inp[11]) ? node2294 : node2291;
														assign node2291 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2294 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2297 = (inp[2]) ? node2301 : node2298;
														assign node2298 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2301 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2304 = (inp[15]) ? node2312 : node2305;
													assign node2305 = (inp[5]) ? node2309 : node2306;
														assign node2306 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2309 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2312 = (inp[8]) ? node2316 : node2313;
														assign node2313 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2316 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node2319 = (inp[11]) ? node2379 : node2320;
										assign node2320 = (inp[2]) ? node2352 : node2321;
											assign node2321 = (inp[10]) ? node2337 : node2322;
												assign node2322 = (inp[15]) ? node2330 : node2323;
													assign node2323 = (inp[0]) ? node2327 : node2324;
														assign node2324 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2327 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2330 = (inp[8]) ? node2334 : node2331;
														assign node2331 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2334 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2337 = (inp[15]) ? node2345 : node2338;
													assign node2338 = (inp[5]) ? node2342 : node2339;
														assign node2339 = (inp[3]) ? 16'b0000011111111111 : 16'b0000001111111111;
														assign node2342 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2345 = (inp[5]) ? node2349 : node2346;
														assign node2346 = (inp[3]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node2349 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2352 = (inp[8]) ? node2366 : node2353;
												assign node2353 = (inp[15]) ? node2361 : node2354;
													assign node2354 = (inp[3]) ? node2358 : node2355;
														assign node2355 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2358 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2361 = (inp[3]) ? 16'b0000000111111111 : node2362;
														assign node2362 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2366 = (inp[5]) ? node2372 : node2367;
													assign node2367 = (inp[0]) ? 16'b0000000111111111 : node2368;
														assign node2368 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2372 = (inp[10]) ? node2376 : node2373;
														assign node2373 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2376 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node2379 = (inp[2]) ? node2411 : node2380;
											assign node2380 = (inp[0]) ? node2396 : node2381;
												assign node2381 = (inp[5]) ? node2389 : node2382;
													assign node2382 = (inp[3]) ? node2386 : node2383;
														assign node2383 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2386 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2389 = (inp[15]) ? node2393 : node2390;
														assign node2390 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node2393 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2396 = (inp[5]) ? node2404 : node2397;
													assign node2397 = (inp[15]) ? node2401 : node2398;
														assign node2398 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node2401 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2404 = (inp[15]) ? node2408 : node2405;
														assign node2405 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2408 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node2411 = (inp[3]) ? node2427 : node2412;
												assign node2412 = (inp[5]) ? node2420 : node2413;
													assign node2413 = (inp[15]) ? node2417 : node2414;
														assign node2414 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2417 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2420 = (inp[10]) ? node2424 : node2421;
														assign node2421 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2424 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node2427 = (inp[5]) ? node2433 : node2428;
													assign node2428 = (inp[10]) ? node2430 : 16'b0000000011111111;
														assign node2430 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node2433 = (inp[8]) ? node2437 : node2434;
														assign node2434 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node2437 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
							assign node2440 = (inp[2]) ? node2672 : node2441;
								assign node2441 = (inp[11]) ? node2555 : node2442;
									assign node2442 = (inp[0]) ? node2500 : node2443;
										assign node2443 = (inp[4]) ? node2471 : node2444;
											assign node2444 = (inp[7]) ? node2458 : node2445;
												assign node2445 = (inp[15]) ? node2451 : node2446;
													assign node2446 = (inp[3]) ? 16'b0000111111111111 : node2447;
														assign node2447 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node2451 = (inp[10]) ? node2455 : node2452;
														assign node2452 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2455 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2458 = (inp[10]) ? node2466 : node2459;
													assign node2459 = (inp[8]) ? node2463 : node2460;
														assign node2460 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2463 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2466 = (inp[5]) ? 16'b0000001111111111 : node2467;
														assign node2467 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2471 = (inp[3]) ? node2487 : node2472;
												assign node2472 = (inp[8]) ? node2480 : node2473;
													assign node2473 = (inp[7]) ? node2477 : node2474;
														assign node2474 = (inp[15]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node2477 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2480 = (inp[10]) ? node2484 : node2481;
														assign node2481 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2484 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2487 = (inp[8]) ? node2495 : node2488;
													assign node2488 = (inp[7]) ? node2492 : node2489;
														assign node2489 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2492 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node2495 = (inp[5]) ? 16'b0000000111111111 : node2496;
														assign node2496 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node2500 = (inp[15]) ? node2530 : node2501;
											assign node2501 = (inp[3]) ? node2515 : node2502;
												assign node2502 = (inp[4]) ? node2510 : node2503;
													assign node2503 = (inp[7]) ? node2507 : node2504;
														assign node2504 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2507 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2510 = (inp[10]) ? 16'b0000001111111111 : node2511;
														assign node2511 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node2515 = (inp[10]) ? node2523 : node2516;
													assign node2516 = (inp[8]) ? node2520 : node2517;
														assign node2517 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2520 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2523 = (inp[7]) ? node2527 : node2524;
														assign node2524 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2527 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2530 = (inp[5]) ? node2542 : node2531;
												assign node2531 = (inp[4]) ? node2537 : node2532;
													assign node2532 = (inp[8]) ? 16'b0000001111111111 : node2533;
														assign node2533 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2537 = (inp[7]) ? 16'b0000000111111111 : node2538;
														assign node2538 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2542 = (inp[10]) ? node2550 : node2543;
													assign node2543 = (inp[4]) ? node2547 : node2544;
														assign node2544 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2547 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2550 = (inp[7]) ? node2552 : 16'b0000000111111111;
														assign node2552 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000001111111;
									assign node2555 = (inp[4]) ? node2613 : node2556;
										assign node2556 = (inp[0]) ? node2588 : node2557;
											assign node2557 = (inp[10]) ? node2573 : node2558;
												assign node2558 = (inp[15]) ? node2566 : node2559;
													assign node2559 = (inp[7]) ? node2563 : node2560;
														assign node2560 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2563 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2566 = (inp[5]) ? node2570 : node2567;
														assign node2567 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2570 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2573 = (inp[3]) ? node2581 : node2574;
													assign node2574 = (inp[8]) ? node2578 : node2575;
														assign node2575 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2578 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2581 = (inp[5]) ? node2585 : node2582;
														assign node2582 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2585 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node2588 = (inp[10]) ? node2604 : node2589;
												assign node2589 = (inp[7]) ? node2597 : node2590;
													assign node2590 = (inp[15]) ? node2594 : node2591;
														assign node2591 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2594 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2597 = (inp[3]) ? node2601 : node2598;
														assign node2598 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2601 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node2604 = (inp[5]) ? 16'b0000000011111111 : node2605;
													assign node2605 = (inp[3]) ? node2609 : node2606;
														assign node2606 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2609 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node2613 = (inp[7]) ? node2643 : node2614;
											assign node2614 = (inp[10]) ? node2628 : node2615;
												assign node2615 = (inp[15]) ? node2623 : node2616;
													assign node2616 = (inp[0]) ? node2620 : node2617;
														assign node2617 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2620 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node2623 = (inp[8]) ? 16'b0000000111111111 : node2624;
														assign node2624 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2628 = (inp[0]) ? node2636 : node2629;
													assign node2629 = (inp[3]) ? node2633 : node2630;
														assign node2630 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2633 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2636 = (inp[8]) ? node2640 : node2637;
														assign node2637 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2640 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2643 = (inp[3]) ? node2659 : node2644;
												assign node2644 = (inp[10]) ? node2652 : node2645;
													assign node2645 = (inp[8]) ? node2649 : node2646;
														assign node2646 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node2649 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2652 = (inp[5]) ? node2656 : node2653;
														assign node2653 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node2656 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2659 = (inp[15]) ? node2667 : node2660;
													assign node2660 = (inp[0]) ? node2664 : node2661;
														assign node2661 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2664 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2667 = (inp[8]) ? node2669 : 16'b0000000011111111;
														assign node2669 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node2672 = (inp[7]) ? node2796 : node2673;
									assign node2673 = (inp[0]) ? node2737 : node2674;
										assign node2674 = (inp[15]) ? node2706 : node2675;
											assign node2675 = (inp[8]) ? node2691 : node2676;
												assign node2676 = (inp[3]) ? node2684 : node2677;
													assign node2677 = (inp[11]) ? node2681 : node2678;
														assign node2678 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2681 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2684 = (inp[5]) ? node2688 : node2685;
														assign node2685 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2688 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2691 = (inp[4]) ? node2699 : node2692;
													assign node2692 = (inp[10]) ? node2696 : node2693;
														assign node2693 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2696 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
													assign node2699 = (inp[3]) ? node2703 : node2700;
														assign node2700 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2703 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node2706 = (inp[11]) ? node2722 : node2707;
												assign node2707 = (inp[5]) ? node2715 : node2708;
													assign node2708 = (inp[10]) ? node2712 : node2709;
														assign node2709 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2712 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2715 = (inp[4]) ? node2719 : node2716;
														assign node2716 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2719 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2722 = (inp[3]) ? node2730 : node2723;
													assign node2723 = (inp[5]) ? node2727 : node2724;
														assign node2724 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2727 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2730 = (inp[10]) ? node2734 : node2731;
														assign node2731 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2734 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node2737 = (inp[5]) ? node2767 : node2738;
											assign node2738 = (inp[10]) ? node2752 : node2739;
												assign node2739 = (inp[15]) ? node2747 : node2740;
													assign node2740 = (inp[3]) ? node2744 : node2741;
														assign node2741 = (inp[11]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node2744 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2747 = (inp[4]) ? 16'b0000000111111111 : node2748;
														assign node2748 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2752 = (inp[3]) ? node2760 : node2753;
													assign node2753 = (inp[11]) ? node2757 : node2754;
														assign node2754 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node2757 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2760 = (inp[4]) ? node2764 : node2761;
														assign node2761 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2764 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2767 = (inp[15]) ? node2781 : node2768;
												assign node2768 = (inp[10]) ? node2776 : node2769;
													assign node2769 = (inp[4]) ? node2773 : node2770;
														assign node2770 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2773 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2776 = (inp[3]) ? 16'b0000000011111111 : node2777;
														assign node2777 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node2781 = (inp[4]) ? node2789 : node2782;
													assign node2782 = (inp[8]) ? node2786 : node2783;
														assign node2783 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node2786 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2789 = (inp[3]) ? node2793 : node2790;
														assign node2790 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node2793 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
									assign node2796 = (inp[5]) ? node2856 : node2797;
										assign node2797 = (inp[0]) ? node2825 : node2798;
											assign node2798 = (inp[3]) ? node2810 : node2799;
												assign node2799 = (inp[8]) ? node2807 : node2800;
													assign node2800 = (inp[11]) ? node2804 : node2801;
														assign node2801 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2804 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2807 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node2810 = (inp[11]) ? node2818 : node2811;
													assign node2811 = (inp[15]) ? node2815 : node2812;
														assign node2812 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2815 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2818 = (inp[10]) ? node2822 : node2819;
														assign node2819 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2822 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2825 = (inp[15]) ? node2841 : node2826;
												assign node2826 = (inp[4]) ? node2834 : node2827;
													assign node2827 = (inp[3]) ? node2831 : node2828;
														assign node2828 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2831 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2834 = (inp[10]) ? node2838 : node2835;
														assign node2835 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2838 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2841 = (inp[3]) ? node2849 : node2842;
													assign node2842 = (inp[8]) ? node2846 : node2843;
														assign node2843 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node2846 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2849 = (inp[4]) ? node2853 : node2850;
														assign node2850 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node2853 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node2856 = (inp[11]) ? node2882 : node2857;
											assign node2857 = (inp[15]) ? node2873 : node2858;
												assign node2858 = (inp[3]) ? node2866 : node2859;
													assign node2859 = (inp[10]) ? node2863 : node2860;
														assign node2860 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2863 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node2866 = (inp[0]) ? node2870 : node2867;
														assign node2867 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2870 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node2873 = (inp[10]) ? 16'b0000000001111111 : node2874;
													assign node2874 = (inp[4]) ? node2878 : node2875;
														assign node2875 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2878 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node2882 = (inp[4]) ? node2898 : node2883;
												assign node2883 = (inp[3]) ? node2891 : node2884;
													assign node2884 = (inp[15]) ? node2888 : node2885;
														assign node2885 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node2888 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node2891 = (inp[10]) ? node2895 : node2892;
														assign node2892 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node2895 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node2898 = (inp[15]) ? node2904 : node2899;
													assign node2899 = (inp[8]) ? node2901 : 16'b0000000001111111;
														assign node2901 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node2904 = (inp[10]) ? node2908 : node2905;
														assign node2905 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node2908 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node2911 = (inp[14]) ? node3403 : node2912;
							assign node2912 = (inp[10]) ? node3154 : node2913;
								assign node2913 = (inp[2]) ? node3033 : node2914;
									assign node2914 = (inp[11]) ? node2970 : node2915;
										assign node2915 = (inp[5]) ? node2941 : node2916;
											assign node2916 = (inp[3]) ? node2930 : node2917;
												assign node2917 = (inp[7]) ? node2925 : node2918;
													assign node2918 = (inp[0]) ? node2922 : node2919;
														assign node2919 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node2922 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2925 = (inp[15]) ? node2927 : 16'b0000111111111111;
														assign node2927 = (inp[4]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node2930 = (inp[0]) ? node2936 : node2931;
													assign node2931 = (inp[8]) ? 16'b0000001111111111 : node2932;
														assign node2932 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node2936 = (inp[15]) ? 16'b0000001111111111 : node2937;
														assign node2937 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node2941 = (inp[4]) ? node2957 : node2942;
												assign node2942 = (inp[8]) ? node2950 : node2943;
													assign node2943 = (inp[0]) ? node2947 : node2944;
														assign node2944 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2947 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2950 = (inp[0]) ? node2954 : node2951;
														assign node2951 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node2954 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2957 = (inp[3]) ? node2963 : node2958;
													assign node2958 = (inp[15]) ? node2960 : 16'b0000001111111111;
														assign node2960 = (inp[0]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node2963 = (inp[15]) ? node2967 : node2964;
														assign node2964 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2967 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
										assign node2970 = (inp[5]) ? node3002 : node2971;
											assign node2971 = (inp[7]) ? node2987 : node2972;
												assign node2972 = (inp[15]) ? node2980 : node2973;
													assign node2973 = (inp[4]) ? node2977 : node2974;
														assign node2974 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node2977 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node2980 = (inp[0]) ? node2984 : node2981;
														assign node2981 = (inp[8]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node2984 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node2987 = (inp[3]) ? node2995 : node2988;
													assign node2988 = (inp[4]) ? node2992 : node2989;
														assign node2989 = (inp[15]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node2992 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node2995 = (inp[0]) ? node2999 : node2996;
														assign node2996 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node2999 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3002 = (inp[7]) ? node3018 : node3003;
												assign node3003 = (inp[8]) ? node3011 : node3004;
													assign node3004 = (inp[15]) ? node3008 : node3005;
														assign node3005 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3008 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3011 = (inp[15]) ? node3015 : node3012;
														assign node3012 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node3015 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3018 = (inp[3]) ? node3026 : node3019;
													assign node3019 = (inp[0]) ? node3023 : node3020;
														assign node3020 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node3023 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3026 = (inp[8]) ? node3030 : node3027;
														assign node3027 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3030 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node3033 = (inp[8]) ? node3095 : node3034;
										assign node3034 = (inp[3]) ? node3066 : node3035;
											assign node3035 = (inp[7]) ? node3051 : node3036;
												assign node3036 = (inp[5]) ? node3044 : node3037;
													assign node3037 = (inp[0]) ? node3041 : node3038;
														assign node3038 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3041 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3044 = (inp[11]) ? node3048 : node3045;
														assign node3045 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3048 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3051 = (inp[4]) ? node3059 : node3052;
													assign node3052 = (inp[5]) ? node3056 : node3053;
														assign node3053 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3056 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3059 = (inp[0]) ? node3063 : node3060;
														assign node3060 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3063 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node3066 = (inp[11]) ? node3082 : node3067;
												assign node3067 = (inp[5]) ? node3075 : node3068;
													assign node3068 = (inp[7]) ? node3072 : node3069;
														assign node3069 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3072 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3075 = (inp[15]) ? node3079 : node3076;
														assign node3076 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3079 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3082 = (inp[15]) ? node3090 : node3083;
													assign node3083 = (inp[4]) ? node3087 : node3084;
														assign node3084 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3087 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node3090 = (inp[5]) ? 16'b0000000011111111 : node3091;
														assign node3091 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3095 = (inp[11]) ? node3127 : node3096;
											assign node3096 = (inp[0]) ? node3112 : node3097;
												assign node3097 = (inp[4]) ? node3105 : node3098;
													assign node3098 = (inp[7]) ? node3102 : node3099;
														assign node3099 = (inp[3]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node3102 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3105 = (inp[3]) ? node3109 : node3106;
														assign node3106 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3109 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3112 = (inp[15]) ? node3120 : node3113;
													assign node3113 = (inp[5]) ? node3117 : node3114;
														assign node3114 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3117 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3120 = (inp[4]) ? node3124 : node3121;
														assign node3121 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3124 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node3127 = (inp[5]) ? node3139 : node3128;
												assign node3128 = (inp[7]) ? node3134 : node3129;
													assign node3129 = (inp[0]) ? node3131 : 16'b0000000111111111;
														assign node3131 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3134 = (inp[3]) ? node3136 : 16'b0000000011111111;
														assign node3136 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3139 = (inp[3]) ? node3147 : node3140;
													assign node3140 = (inp[0]) ? node3144 : node3141;
														assign node3141 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node3144 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3147 = (inp[15]) ? node3151 : node3148;
														assign node3148 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3151 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node3154 = (inp[0]) ? node3280 : node3155;
									assign node3155 = (inp[8]) ? node3217 : node3156;
										assign node3156 = (inp[7]) ? node3188 : node3157;
											assign node3157 = (inp[4]) ? node3173 : node3158;
												assign node3158 = (inp[15]) ? node3166 : node3159;
													assign node3159 = (inp[11]) ? node3163 : node3160;
														assign node3160 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3163 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3166 = (inp[11]) ? node3170 : node3167;
														assign node3167 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3170 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node3173 = (inp[2]) ? node3181 : node3174;
													assign node3174 = (inp[5]) ? node3178 : node3175;
														assign node3175 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3178 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3181 = (inp[11]) ? node3185 : node3182;
														assign node3182 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3185 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node3188 = (inp[15]) ? node3204 : node3189;
												assign node3189 = (inp[4]) ? node3197 : node3190;
													assign node3190 = (inp[5]) ? node3194 : node3191;
														assign node3191 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3194 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3197 = (inp[3]) ? node3201 : node3198;
														assign node3198 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3201 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3204 = (inp[5]) ? node3212 : node3205;
													assign node3205 = (inp[3]) ? node3209 : node3206;
														assign node3206 = (inp[2]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node3209 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3212 = (inp[3]) ? node3214 : 16'b0000000011111111;
														assign node3214 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3217 = (inp[3]) ? node3249 : node3218;
											assign node3218 = (inp[2]) ? node3234 : node3219;
												assign node3219 = (inp[4]) ? node3227 : node3220;
													assign node3220 = (inp[11]) ? node3224 : node3221;
														assign node3221 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3224 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3227 = (inp[5]) ? node3231 : node3228;
														assign node3228 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3231 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node3234 = (inp[11]) ? node3242 : node3235;
													assign node3235 = (inp[7]) ? node3239 : node3236;
														assign node3236 = (inp[5]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node3239 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3242 = (inp[7]) ? node3246 : node3243;
														assign node3243 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node3246 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3249 = (inp[11]) ? node3265 : node3250;
												assign node3250 = (inp[2]) ? node3258 : node3251;
													assign node3251 = (inp[5]) ? node3255 : node3252;
														assign node3252 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3255 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3258 = (inp[4]) ? node3262 : node3259;
														assign node3259 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3262 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node3265 = (inp[15]) ? node3273 : node3266;
													assign node3266 = (inp[4]) ? node3270 : node3267;
														assign node3267 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node3270 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3273 = (inp[2]) ? node3277 : node3274;
														assign node3274 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3277 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node3280 = (inp[2]) ? node3344 : node3281;
										assign node3281 = (inp[15]) ? node3313 : node3282;
											assign node3282 = (inp[11]) ? node3298 : node3283;
												assign node3283 = (inp[3]) ? node3291 : node3284;
													assign node3284 = (inp[5]) ? node3288 : node3285;
														assign node3285 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3288 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3291 = (inp[4]) ? node3295 : node3292;
														assign node3292 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3295 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3298 = (inp[3]) ? node3306 : node3299;
													assign node3299 = (inp[5]) ? node3303 : node3300;
														assign node3300 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3303 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3306 = (inp[7]) ? node3310 : node3307;
														assign node3307 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3310 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node3313 = (inp[4]) ? node3329 : node3314;
												assign node3314 = (inp[7]) ? node3322 : node3315;
													assign node3315 = (inp[11]) ? node3319 : node3316;
														assign node3316 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3319 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3322 = (inp[5]) ? node3326 : node3323;
														assign node3323 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3326 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node3329 = (inp[3]) ? node3337 : node3330;
													assign node3330 = (inp[8]) ? node3334 : node3331;
														assign node3331 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3334 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3337 = (inp[7]) ? node3341 : node3338;
														assign node3338 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3341 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3344 = (inp[3]) ? node3372 : node3345;
											assign node3345 = (inp[11]) ? node3361 : node3346;
												assign node3346 = (inp[4]) ? node3354 : node3347;
													assign node3347 = (inp[5]) ? node3351 : node3348;
														assign node3348 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3351 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3354 = (inp[5]) ? node3358 : node3355;
														assign node3355 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3358 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3361 = (inp[4]) ? node3367 : node3362;
													assign node3362 = (inp[5]) ? node3364 : 16'b0000000011111111;
														assign node3364 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3367 = (inp[8]) ? 16'b0000000000111111 : node3368;
														assign node3368 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node3372 = (inp[15]) ? node3388 : node3373;
												assign node3373 = (inp[8]) ? node3381 : node3374;
													assign node3374 = (inp[5]) ? node3378 : node3375;
														assign node3375 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3378 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3381 = (inp[7]) ? node3385 : node3382;
														assign node3382 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3385 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3388 = (inp[11]) ? node3396 : node3389;
													assign node3389 = (inp[7]) ? node3393 : node3390;
														assign node3390 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node3393 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node3396 = (inp[7]) ? node3400 : node3397;
														assign node3397 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node3400 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node3403 = (inp[15]) ? node3645 : node3404;
								assign node3404 = (inp[10]) ? node3526 : node3405;
									assign node3405 = (inp[7]) ? node3465 : node3406;
										assign node3406 = (inp[5]) ? node3436 : node3407;
											assign node3407 = (inp[11]) ? node3423 : node3408;
												assign node3408 = (inp[2]) ? node3416 : node3409;
													assign node3409 = (inp[3]) ? node3413 : node3410;
														assign node3410 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3413 = (inp[0]) ? 16'b0000011111111111 : 16'b0000011111111111;
													assign node3416 = (inp[0]) ? node3420 : node3417;
														assign node3417 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3420 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
												assign node3423 = (inp[2]) ? node3431 : node3424;
													assign node3424 = (inp[0]) ? node3428 : node3425;
														assign node3425 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3428 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3431 = (inp[4]) ? 16'b0000000011111111 : node3432;
														assign node3432 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3436 = (inp[3]) ? node3450 : node3437;
												assign node3437 = (inp[11]) ? node3445 : node3438;
													assign node3438 = (inp[4]) ? node3442 : node3439;
														assign node3439 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3442 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3445 = (inp[0]) ? 16'b0000000111111111 : node3446;
														assign node3446 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3450 = (inp[11]) ? node3458 : node3451;
													assign node3451 = (inp[0]) ? node3455 : node3452;
														assign node3452 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3455 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3458 = (inp[2]) ? node3462 : node3459;
														assign node3459 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3462 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node3465 = (inp[3]) ? node3497 : node3466;
											assign node3466 = (inp[0]) ? node3482 : node3467;
												assign node3467 = (inp[8]) ? node3475 : node3468;
													assign node3468 = (inp[5]) ? node3472 : node3469;
														assign node3469 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3472 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3475 = (inp[11]) ? node3479 : node3476;
														assign node3476 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node3479 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3482 = (inp[2]) ? node3490 : node3483;
													assign node3483 = (inp[4]) ? node3487 : node3484;
														assign node3484 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3487 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3490 = (inp[8]) ? node3494 : node3491;
														assign node3491 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3494 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3497 = (inp[11]) ? node3513 : node3498;
												assign node3498 = (inp[4]) ? node3506 : node3499;
													assign node3499 = (inp[2]) ? node3503 : node3500;
														assign node3500 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3503 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3506 = (inp[8]) ? node3510 : node3507;
														assign node3507 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node3510 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3513 = (inp[4]) ? node3519 : node3514;
													assign node3514 = (inp[2]) ? 16'b0000000111111111 : node3515;
														assign node3515 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node3519 = (inp[0]) ? node3523 : node3520;
														assign node3520 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3523 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
									assign node3526 = (inp[4]) ? node3588 : node3527;
										assign node3527 = (inp[2]) ? node3559 : node3528;
											assign node3528 = (inp[7]) ? node3544 : node3529;
												assign node3529 = (inp[3]) ? node3537 : node3530;
													assign node3530 = (inp[11]) ? node3534 : node3531;
														assign node3531 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3534 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3537 = (inp[5]) ? node3541 : node3538;
														assign node3538 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3541 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node3544 = (inp[5]) ? node3552 : node3545;
													assign node3545 = (inp[11]) ? node3549 : node3546;
														assign node3546 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node3549 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3552 = (inp[0]) ? node3556 : node3553;
														assign node3553 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node3556 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node3559 = (inp[11]) ? node3575 : node3560;
												assign node3560 = (inp[8]) ? node3568 : node3561;
													assign node3561 = (inp[3]) ? node3565 : node3562;
														assign node3562 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node3565 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3568 = (inp[7]) ? node3572 : node3569;
														assign node3569 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3572 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3575 = (inp[3]) ? node3581 : node3576;
													assign node3576 = (inp[7]) ? node3578 : 16'b0000000011111111;
														assign node3578 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3581 = (inp[8]) ? node3585 : node3582;
														assign node3582 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node3585 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3588 = (inp[8]) ? node3616 : node3589;
											assign node3589 = (inp[2]) ? node3605 : node3590;
												assign node3590 = (inp[0]) ? node3598 : node3591;
													assign node3591 = (inp[7]) ? node3595 : node3592;
														assign node3592 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node3595 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node3598 = (inp[11]) ? node3602 : node3599;
														assign node3599 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3602 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3605 = (inp[0]) ? node3613 : node3606;
													assign node3606 = (inp[5]) ? node3610 : node3607;
														assign node3607 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node3610 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3613 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3616 = (inp[3]) ? node3632 : node3617;
												assign node3617 = (inp[0]) ? node3625 : node3618;
													assign node3618 = (inp[11]) ? node3622 : node3619;
														assign node3619 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node3622 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3625 = (inp[5]) ? node3629 : node3626;
														assign node3626 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3629 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3632 = (inp[7]) ? node3638 : node3633;
													assign node3633 = (inp[0]) ? node3635 : 16'b0000000001111111;
														assign node3635 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node3638 = (inp[0]) ? node3642 : node3639;
														assign node3639 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node3642 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node3645 = (inp[7]) ? node3771 : node3646;
									assign node3646 = (inp[8]) ? node3708 : node3647;
										assign node3647 = (inp[0]) ? node3677 : node3648;
											assign node3648 = (inp[11]) ? node3662 : node3649;
												assign node3649 = (inp[2]) ? node3657 : node3650;
													assign node3650 = (inp[4]) ? node3654 : node3651;
														assign node3651 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3654 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node3657 = (inp[5]) ? 16'b0000000111111111 : node3658;
														assign node3658 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node3662 = (inp[2]) ? node3670 : node3663;
													assign node3663 = (inp[3]) ? node3667 : node3664;
														assign node3664 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3667 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node3670 = (inp[4]) ? node3674 : node3671;
														assign node3671 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node3674 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node3677 = (inp[3]) ? node3693 : node3678;
												assign node3678 = (inp[10]) ? node3686 : node3679;
													assign node3679 = (inp[5]) ? node3683 : node3680;
														assign node3680 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node3683 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node3686 = (inp[4]) ? node3690 : node3687;
														assign node3687 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3690 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3693 = (inp[11]) ? node3701 : node3694;
													assign node3694 = (inp[10]) ? node3698 : node3695;
														assign node3695 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node3698 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3701 = (inp[10]) ? node3705 : node3702;
														assign node3702 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3705 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node3708 = (inp[11]) ? node3740 : node3709;
											assign node3709 = (inp[10]) ? node3725 : node3710;
												assign node3710 = (inp[0]) ? node3718 : node3711;
													assign node3711 = (inp[4]) ? node3715 : node3712;
														assign node3712 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node3715 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node3718 = (inp[2]) ? node3722 : node3719;
														assign node3719 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3722 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3725 = (inp[2]) ? node3733 : node3726;
													assign node3726 = (inp[4]) ? node3730 : node3727;
														assign node3727 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node3730 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3733 = (inp[3]) ? node3737 : node3734;
														assign node3734 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node3737 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3740 = (inp[5]) ? node3756 : node3741;
												assign node3741 = (inp[3]) ? node3749 : node3742;
													assign node3742 = (inp[4]) ? node3746 : node3743;
														assign node3743 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3746 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node3749 = (inp[0]) ? node3753 : node3750;
														assign node3750 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3753 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3756 = (inp[3]) ? node3764 : node3757;
													assign node3757 = (inp[4]) ? node3761 : node3758;
														assign node3758 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node3761 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node3764 = (inp[2]) ? node3768 : node3765;
														assign node3765 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node3768 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node3771 = (inp[0]) ? node3831 : node3772;
										assign node3772 = (inp[11]) ? node3800 : node3773;
											assign node3773 = (inp[8]) ? node3787 : node3774;
												assign node3774 = (inp[10]) ? node3780 : node3775;
													assign node3775 = (inp[2]) ? 16'b0000000111111111 : node3776;
														assign node3776 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node3780 = (inp[3]) ? node3784 : node3781;
														assign node3781 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3784 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node3787 = (inp[3]) ? node3795 : node3788;
													assign node3788 = (inp[10]) ? node3792 : node3789;
														assign node3789 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node3792 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node3795 = (inp[10]) ? 16'b0000000000011111 : node3796;
														assign node3796 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node3800 = (inp[5]) ? node3816 : node3801;
												assign node3801 = (inp[10]) ? node3809 : node3802;
													assign node3802 = (inp[4]) ? node3806 : node3803;
														assign node3803 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node3806 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node3809 = (inp[4]) ? node3813 : node3810;
														assign node3810 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3813 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3816 = (inp[10]) ? node3824 : node3817;
													assign node3817 = (inp[8]) ? node3821 : node3818;
														assign node3818 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node3821 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node3824 = (inp[8]) ? node3828 : node3825;
														assign node3825 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node3828 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000011111;
										assign node3831 = (inp[8]) ? node3859 : node3832;
											assign node3832 = (inp[2]) ? node3844 : node3833;
												assign node3833 = (inp[10]) ? node3839 : node3834;
													assign node3834 = (inp[4]) ? node3836 : 16'b0000000111111111;
														assign node3836 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node3839 = (inp[5]) ? node3841 : 16'b0000000001111111;
														assign node3841 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node3844 = (inp[10]) ? node3852 : node3845;
													assign node3845 = (inp[5]) ? node3849 : node3846;
														assign node3846 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node3849 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node3852 = (inp[4]) ? node3856 : node3853;
														assign node3853 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node3856 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node3859 = (inp[4]) ? node3873 : node3860;
												assign node3860 = (inp[2]) ? node3866 : node3861;
													assign node3861 = (inp[3]) ? node3863 : 16'b0000000011111111;
														assign node3863 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node3866 = (inp[5]) ? node3870 : node3867;
														assign node3867 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node3870 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node3873 = (inp[3]) ? node3881 : node3874;
													assign node3874 = (inp[11]) ? node3878 : node3875;
														assign node3875 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node3878 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node3881 = (inp[10]) ? node3885 : node3882;
														assign node3882 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node3885 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
				assign node3888 = (inp[13]) ? node5846 : node3889;
					assign node3889 = (inp[14]) ? node4877 : node3890;
						assign node3890 = (inp[12]) ? node4386 : node3891;
							assign node3891 = (inp[7]) ? node4137 : node3892;
								assign node3892 = (inp[8]) ? node4014 : node3893;
									assign node3893 = (inp[3]) ? node3953 : node3894;
										assign node3894 = (inp[15]) ? node3926 : node3895;
											assign node3895 = (inp[5]) ? node3911 : node3896;
												assign node3896 = (inp[0]) ? node3904 : node3897;
													assign node3897 = (inp[10]) ? node3901 : node3898;
														assign node3898 = (inp[11]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node3901 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node3904 = (inp[4]) ? node3908 : node3905;
														assign node3905 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node3908 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3911 = (inp[11]) ? node3919 : node3912;
													assign node3912 = (inp[4]) ? node3916 : node3913;
														assign node3913 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node3916 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3919 = (inp[10]) ? node3923 : node3920;
														assign node3920 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3923 = (inp[0]) ? 16'b0000000111111111 : 16'b0000011111111111;
											assign node3926 = (inp[11]) ? node3940 : node3927;
												assign node3927 = (inp[5]) ? node3935 : node3928;
													assign node3928 = (inp[2]) ? node3932 : node3929;
														assign node3929 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node3932 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node3935 = (inp[2]) ? 16'b0000011111111111 : node3936;
														assign node3936 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node3940 = (inp[4]) ? node3946 : node3941;
													assign node3941 = (inp[10]) ? node3943 : 16'b0000111111111111;
														assign node3943 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3946 = (inp[10]) ? node3950 : node3947;
														assign node3947 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3950 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node3953 = (inp[5]) ? node3985 : node3954;
											assign node3954 = (inp[0]) ? node3970 : node3955;
												assign node3955 = (inp[4]) ? node3963 : node3956;
													assign node3956 = (inp[15]) ? node3960 : node3957;
														assign node3957 = (inp[10]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node3960 = (inp[2]) ? 16'b0000111111111111 : 16'b0000111111111111;
													assign node3963 = (inp[10]) ? node3967 : node3964;
														assign node3964 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3967 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node3970 = (inp[2]) ? node3978 : node3971;
													assign node3971 = (inp[15]) ? node3975 : node3972;
														assign node3972 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3975 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3978 = (inp[15]) ? node3982 : node3979;
														assign node3979 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3982 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node3985 = (inp[0]) ? node4001 : node3986;
												assign node3986 = (inp[2]) ? node3994 : node3987;
													assign node3987 = (inp[11]) ? node3991 : node3988;
														assign node3988 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node3991 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node3994 = (inp[10]) ? node3998 : node3995;
														assign node3995 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node3998 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node4001 = (inp[10]) ? node4009 : node4002;
													assign node4002 = (inp[15]) ? node4006 : node4003;
														assign node4003 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4006 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4009 = (inp[2]) ? 16'b0000000111111111 : node4010;
														assign node4010 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
									assign node4014 = (inp[4]) ? node4076 : node4015;
										assign node4015 = (inp[15]) ? node4047 : node4016;
											assign node4016 = (inp[5]) ? node4032 : node4017;
												assign node4017 = (inp[10]) ? node4025 : node4018;
													assign node4018 = (inp[11]) ? node4022 : node4019;
														assign node4019 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node4022 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4025 = (inp[2]) ? node4029 : node4026;
														assign node4026 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4029 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4032 = (inp[3]) ? node4040 : node4033;
													assign node4033 = (inp[0]) ? node4037 : node4034;
														assign node4034 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4037 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4040 = (inp[11]) ? node4044 : node4041;
														assign node4041 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4044 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4047 = (inp[2]) ? node4061 : node4048;
												assign node4048 = (inp[3]) ? node4054 : node4049;
													assign node4049 = (inp[5]) ? 16'b0000011111111111 : node4050;
														assign node4050 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4054 = (inp[5]) ? node4058 : node4055;
														assign node4055 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4058 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4061 = (inp[11]) ? node4069 : node4062;
													assign node4062 = (inp[5]) ? node4066 : node4063;
														assign node4063 = (inp[3]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node4066 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4069 = (inp[0]) ? node4073 : node4070;
														assign node4070 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4073 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4076 = (inp[3]) ? node4108 : node4077;
											assign node4077 = (inp[2]) ? node4093 : node4078;
												assign node4078 = (inp[11]) ? node4086 : node4079;
													assign node4079 = (inp[5]) ? node4083 : node4080;
														assign node4080 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4083 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4086 = (inp[15]) ? node4090 : node4087;
														assign node4087 = (inp[0]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node4090 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4093 = (inp[5]) ? node4101 : node4094;
													assign node4094 = (inp[0]) ? node4098 : node4095;
														assign node4095 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4098 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4101 = (inp[0]) ? node4105 : node4102;
														assign node4102 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4105 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4108 = (inp[15]) ? node4122 : node4109;
												assign node4109 = (inp[10]) ? node4115 : node4110;
													assign node4110 = (inp[11]) ? 16'b0000001111111111 : node4111;
														assign node4111 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4115 = (inp[2]) ? node4119 : node4116;
														assign node4116 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4119 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4122 = (inp[2]) ? node4130 : node4123;
													assign node4123 = (inp[5]) ? node4127 : node4124;
														assign node4124 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node4127 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node4130 = (inp[10]) ? node4134 : node4131;
														assign node4131 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4134 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000001111111;
								assign node4137 = (inp[4]) ? node4263 : node4138;
									assign node4138 = (inp[3]) ? node4202 : node4139;
										assign node4139 = (inp[0]) ? node4171 : node4140;
											assign node4140 = (inp[11]) ? node4156 : node4141;
												assign node4141 = (inp[8]) ? node4149 : node4142;
													assign node4142 = (inp[15]) ? node4146 : node4143;
														assign node4143 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node4146 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4149 = (inp[2]) ? node4153 : node4150;
														assign node4150 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4153 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4156 = (inp[10]) ? node4164 : node4157;
													assign node4157 = (inp[8]) ? node4161 : node4158;
														assign node4158 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4161 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4164 = (inp[5]) ? node4168 : node4165;
														assign node4165 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4168 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4171 = (inp[5]) ? node4187 : node4172;
												assign node4172 = (inp[15]) ? node4180 : node4173;
													assign node4173 = (inp[8]) ? node4177 : node4174;
														assign node4174 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4177 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4180 = (inp[8]) ? node4184 : node4181;
														assign node4181 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4184 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4187 = (inp[11]) ? node4195 : node4188;
													assign node4188 = (inp[8]) ? node4192 : node4189;
														assign node4189 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4192 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4195 = (inp[10]) ? node4199 : node4196;
														assign node4196 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4199 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
										assign node4202 = (inp[10]) ? node4232 : node4203;
											assign node4203 = (inp[2]) ? node4217 : node4204;
												assign node4204 = (inp[11]) ? node4212 : node4205;
													assign node4205 = (inp[8]) ? node4209 : node4206;
														assign node4206 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4209 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4212 = (inp[0]) ? 16'b0000001111111111 : node4213;
														assign node4213 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4217 = (inp[11]) ? node4225 : node4218;
													assign node4218 = (inp[8]) ? node4222 : node4219;
														assign node4219 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4222 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4225 = (inp[5]) ? node4229 : node4226;
														assign node4226 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node4229 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4232 = (inp[5]) ? node4248 : node4233;
												assign node4233 = (inp[15]) ? node4241 : node4234;
													assign node4234 = (inp[11]) ? node4238 : node4235;
														assign node4235 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4238 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4241 = (inp[8]) ? node4245 : node4242;
														assign node4242 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4245 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node4248 = (inp[0]) ? node4256 : node4249;
													assign node4249 = (inp[2]) ? node4253 : node4250;
														assign node4250 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node4253 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4256 = (inp[15]) ? node4260 : node4257;
														assign node4257 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4260 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node4263 = (inp[2]) ? node4325 : node4264;
										assign node4264 = (inp[8]) ? node4296 : node4265;
											assign node4265 = (inp[10]) ? node4281 : node4266;
												assign node4266 = (inp[15]) ? node4274 : node4267;
													assign node4267 = (inp[0]) ? node4271 : node4268;
														assign node4268 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4271 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4274 = (inp[11]) ? node4278 : node4275;
														assign node4275 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4278 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node4281 = (inp[3]) ? node4289 : node4282;
													assign node4282 = (inp[11]) ? node4286 : node4283;
														assign node4283 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4286 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4289 = (inp[5]) ? node4293 : node4290;
														assign node4290 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4293 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4296 = (inp[5]) ? node4312 : node4297;
												assign node4297 = (inp[3]) ? node4305 : node4298;
													assign node4298 = (inp[11]) ? node4302 : node4299;
														assign node4299 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4302 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4305 = (inp[0]) ? node4309 : node4306;
														assign node4306 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4309 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node4312 = (inp[0]) ? node4318 : node4313;
													assign node4313 = (inp[10]) ? node4315 : 16'b0000000111111111;
														assign node4315 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4318 = (inp[15]) ? node4322 : node4319;
														assign node4319 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4322 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node4325 = (inp[5]) ? node4355 : node4326;
											assign node4326 = (inp[0]) ? node4340 : node4327;
												assign node4327 = (inp[10]) ? node4333 : node4328;
													assign node4328 = (inp[3]) ? node4330 : 16'b0000001111111111;
														assign node4330 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4333 = (inp[8]) ? node4337 : node4334;
														assign node4334 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4337 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4340 = (inp[11]) ? node4348 : node4341;
													assign node4341 = (inp[8]) ? node4345 : node4342;
														assign node4342 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4345 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4348 = (inp[15]) ? node4352 : node4349;
														assign node4349 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4352 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4355 = (inp[15]) ? node4371 : node4356;
												assign node4356 = (inp[3]) ? node4364 : node4357;
													assign node4357 = (inp[10]) ? node4361 : node4358;
														assign node4358 = (inp[0]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node4361 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4364 = (inp[10]) ? node4368 : node4365;
														assign node4365 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4368 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4371 = (inp[10]) ? node4379 : node4372;
													assign node4372 = (inp[0]) ? node4376 : node4373;
														assign node4373 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4376 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node4379 = (inp[8]) ? node4383 : node4380;
														assign node4380 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4383 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node4386 = (inp[8]) ? node4634 : node4387;
								assign node4387 = (inp[15]) ? node4509 : node4388;
									assign node4388 = (inp[10]) ? node4450 : node4389;
										assign node4389 = (inp[3]) ? node4421 : node4390;
											assign node4390 = (inp[11]) ? node4406 : node4391;
												assign node4391 = (inp[5]) ? node4399 : node4392;
													assign node4392 = (inp[0]) ? node4396 : node4393;
														assign node4393 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node4396 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4399 = (inp[2]) ? node4403 : node4400;
														assign node4400 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4403 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4406 = (inp[2]) ? node4414 : node4407;
													assign node4407 = (inp[5]) ? node4411 : node4408;
														assign node4408 = (inp[0]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node4411 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4414 = (inp[5]) ? node4418 : node4415;
														assign node4415 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4418 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4421 = (inp[4]) ? node4437 : node4422;
												assign node4422 = (inp[5]) ? node4430 : node4423;
													assign node4423 = (inp[7]) ? node4427 : node4424;
														assign node4424 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4427 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4430 = (inp[2]) ? node4434 : node4431;
														assign node4431 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4434 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
												assign node4437 = (inp[0]) ? node4443 : node4438;
													assign node4438 = (inp[5]) ? node4440 : 16'b0000001111111111;
														assign node4440 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4443 = (inp[2]) ? node4447 : node4444;
														assign node4444 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4447 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node4450 = (inp[11]) ? node4478 : node4451;
											assign node4451 = (inp[7]) ? node4463 : node4452;
												assign node4452 = (inp[3]) ? node4458 : node4453;
													assign node4453 = (inp[2]) ? 16'b0000011111111111 : node4454;
														assign node4454 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node4458 = (inp[2]) ? 16'b0000001111111111 : node4459;
														assign node4459 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4463 = (inp[2]) ? node4471 : node4464;
													assign node4464 = (inp[4]) ? node4468 : node4465;
														assign node4465 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4468 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4471 = (inp[3]) ? node4475 : node4472;
														assign node4472 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4475 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4478 = (inp[4]) ? node4494 : node4479;
												assign node4479 = (inp[0]) ? node4487 : node4480;
													assign node4480 = (inp[5]) ? node4484 : node4481;
														assign node4481 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4484 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4487 = (inp[5]) ? node4491 : node4488;
														assign node4488 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4491 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4494 = (inp[3]) ? node4502 : node4495;
													assign node4495 = (inp[5]) ? node4499 : node4496;
														assign node4496 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4499 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4502 = (inp[0]) ? node4506 : node4503;
														assign node4503 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4506 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node4509 = (inp[7]) ? node4573 : node4510;
										assign node4510 = (inp[5]) ? node4542 : node4511;
											assign node4511 = (inp[2]) ? node4527 : node4512;
												assign node4512 = (inp[11]) ? node4520 : node4513;
													assign node4513 = (inp[4]) ? node4517 : node4514;
														assign node4514 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4517 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4520 = (inp[0]) ? node4524 : node4521;
														assign node4521 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4524 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4527 = (inp[0]) ? node4535 : node4528;
													assign node4528 = (inp[10]) ? node4532 : node4529;
														assign node4529 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4532 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4535 = (inp[4]) ? node4539 : node4536;
														assign node4536 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node4539 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4542 = (inp[3]) ? node4558 : node4543;
												assign node4543 = (inp[0]) ? node4551 : node4544;
													assign node4544 = (inp[10]) ? node4548 : node4545;
														assign node4545 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4548 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node4551 = (inp[2]) ? node4555 : node4552;
														assign node4552 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4555 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4558 = (inp[11]) ? node4566 : node4559;
													assign node4559 = (inp[10]) ? node4563 : node4560;
														assign node4560 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node4563 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4566 = (inp[2]) ? node4570 : node4567;
														assign node4567 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4570 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4573 = (inp[2]) ? node4603 : node4574;
											assign node4574 = (inp[3]) ? node4588 : node4575;
												assign node4575 = (inp[4]) ? node4583 : node4576;
													assign node4576 = (inp[0]) ? node4580 : node4577;
														assign node4577 = (inp[5]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node4580 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4583 = (inp[5]) ? 16'b0000000111111111 : node4584;
														assign node4584 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4588 = (inp[4]) ? node4596 : node4589;
													assign node4589 = (inp[11]) ? node4593 : node4590;
														assign node4590 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4593 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node4596 = (inp[10]) ? node4600 : node4597;
														assign node4597 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4600 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4603 = (inp[5]) ? node4619 : node4604;
												assign node4604 = (inp[11]) ? node4612 : node4605;
													assign node4605 = (inp[0]) ? node4609 : node4606;
														assign node4606 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4609 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4612 = (inp[3]) ? node4616 : node4613;
														assign node4613 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4616 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node4619 = (inp[4]) ? node4627 : node4620;
													assign node4620 = (inp[3]) ? node4624 : node4621;
														assign node4621 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node4624 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4627 = (inp[11]) ? node4631 : node4628;
														assign node4628 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node4631 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
								assign node4634 = (inp[15]) ? node4754 : node4635;
									assign node4635 = (inp[5]) ? node4695 : node4636;
										assign node4636 = (inp[2]) ? node4664 : node4637;
											assign node4637 = (inp[0]) ? node4649 : node4638;
												assign node4638 = (inp[3]) ? node4644 : node4639;
													assign node4639 = (inp[4]) ? node4641 : 16'b0000111111111111;
														assign node4641 = (inp[11]) ? 16'b0000011111111111 : 16'b0000011111111111;
													assign node4644 = (inp[11]) ? 16'b0000001111111111 : node4645;
														assign node4645 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4649 = (inp[4]) ? node4657 : node4650;
													assign node4650 = (inp[11]) ? node4654 : node4651;
														assign node4651 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4654 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4657 = (inp[3]) ? node4661 : node4658;
														assign node4658 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4661 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4664 = (inp[4]) ? node4680 : node4665;
												assign node4665 = (inp[3]) ? node4673 : node4666;
													assign node4666 = (inp[10]) ? node4670 : node4667;
														assign node4667 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4670 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4673 = (inp[11]) ? node4677 : node4674;
														assign node4674 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4677 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node4680 = (inp[11]) ? node4688 : node4681;
													assign node4681 = (inp[7]) ? node4685 : node4682;
														assign node4682 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4685 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4688 = (inp[10]) ? node4692 : node4689;
														assign node4689 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4692 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node4695 = (inp[0]) ? node4723 : node4696;
											assign node4696 = (inp[10]) ? node4710 : node4697;
												assign node4697 = (inp[2]) ? node4705 : node4698;
													assign node4698 = (inp[4]) ? node4702 : node4699;
														assign node4699 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4702 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4705 = (inp[4]) ? 16'b0000000111111111 : node4706;
														assign node4706 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4710 = (inp[3]) ? node4716 : node4711;
													assign node4711 = (inp[7]) ? node4713 : 16'b0000001111111111;
														assign node4713 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4716 = (inp[2]) ? node4720 : node4717;
														assign node4717 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4720 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4723 = (inp[7]) ? node4739 : node4724;
												assign node4724 = (inp[11]) ? node4732 : node4725;
													assign node4725 = (inp[10]) ? node4729 : node4726;
														assign node4726 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node4729 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4732 = (inp[2]) ? node4736 : node4733;
														assign node4733 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4736 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4739 = (inp[4]) ? node4747 : node4740;
													assign node4740 = (inp[2]) ? node4744 : node4741;
														assign node4741 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4744 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4747 = (inp[3]) ? node4751 : node4748;
														assign node4748 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4751 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node4754 = (inp[10]) ? node4818 : node4755;
										assign node4755 = (inp[5]) ? node4787 : node4756;
											assign node4756 = (inp[2]) ? node4772 : node4757;
												assign node4757 = (inp[7]) ? node4765 : node4758;
													assign node4758 = (inp[0]) ? node4762 : node4759;
														assign node4759 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4762 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4765 = (inp[4]) ? node4769 : node4766;
														assign node4766 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4769 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4772 = (inp[0]) ? node4780 : node4773;
													assign node4773 = (inp[3]) ? node4777 : node4774;
														assign node4774 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4777 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4780 = (inp[3]) ? node4784 : node4781;
														assign node4781 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4784 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node4787 = (inp[3]) ? node4803 : node4788;
												assign node4788 = (inp[4]) ? node4796 : node4789;
													assign node4789 = (inp[11]) ? node4793 : node4790;
														assign node4790 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4793 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4796 = (inp[2]) ? node4800 : node4797;
														assign node4797 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4800 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node4803 = (inp[11]) ? node4811 : node4804;
													assign node4804 = (inp[0]) ? node4808 : node4805;
														assign node4805 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4808 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4811 = (inp[7]) ? node4815 : node4812;
														assign node4812 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node4815 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node4818 = (inp[11]) ? node4846 : node4819;
											assign node4819 = (inp[2]) ? node4833 : node4820;
												assign node4820 = (inp[5]) ? node4826 : node4821;
													assign node4821 = (inp[4]) ? 16'b0000000111111111 : node4822;
														assign node4822 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4826 = (inp[4]) ? node4830 : node4827;
														assign node4827 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4830 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4833 = (inp[0]) ? node4841 : node4834;
													assign node4834 = (inp[4]) ? node4838 : node4835;
														assign node4835 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4838 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node4841 = (inp[7]) ? node4843 : 16'b0000000001111111;
														assign node4843 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node4846 = (inp[7]) ? node4862 : node4847;
												assign node4847 = (inp[3]) ? node4855 : node4848;
													assign node4848 = (inp[4]) ? node4852 : node4849;
														assign node4849 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node4852 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node4855 = (inp[4]) ? node4859 : node4856;
														assign node4856 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4859 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node4862 = (inp[0]) ? node4870 : node4863;
													assign node4863 = (inp[3]) ? node4867 : node4864;
														assign node4864 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node4867 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node4870 = (inp[3]) ? node4874 : node4871;
														assign node4871 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node4874 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node4877 = (inp[15]) ? node5359 : node4878;
							assign node4878 = (inp[12]) ? node5124 : node4879;
								assign node4879 = (inp[11]) ? node5001 : node4880;
									assign node4880 = (inp[10]) ? node4940 : node4881;
										assign node4881 = (inp[4]) ? node4911 : node4882;
											assign node4882 = (inp[5]) ? node4898 : node4883;
												assign node4883 = (inp[3]) ? node4891 : node4884;
													assign node4884 = (inp[0]) ? node4888 : node4885;
														assign node4885 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node4888 = (inp[2]) ? 16'b0000111111111111 : 16'b0000011111111111;
													assign node4891 = (inp[7]) ? node4895 : node4892;
														assign node4892 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4895 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node4898 = (inp[8]) ? node4904 : node4899;
													assign node4899 = (inp[7]) ? node4901 : 16'b0000011111111111;
														assign node4901 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4904 = (inp[7]) ? node4908 : node4905;
														assign node4905 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4908 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node4911 = (inp[8]) ? node4925 : node4912;
												assign node4912 = (inp[7]) ? node4918 : node4913;
													assign node4913 = (inp[3]) ? node4915 : 16'b0000011111111111;
														assign node4915 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node4918 = (inp[2]) ? node4922 : node4919;
														assign node4919 = (inp[5]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node4922 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node4925 = (inp[5]) ? node4933 : node4926;
													assign node4926 = (inp[2]) ? node4930 : node4927;
														assign node4927 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4930 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4933 = (inp[3]) ? node4937 : node4934;
														assign node4934 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4937 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node4940 = (inp[2]) ? node4970 : node4941;
											assign node4941 = (inp[0]) ? node4955 : node4942;
												assign node4942 = (inp[4]) ? node4950 : node4943;
													assign node4943 = (inp[7]) ? node4947 : node4944;
														assign node4944 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node4947 = (inp[8]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node4950 = (inp[8]) ? node4952 : 16'b0000001111111111;
														assign node4952 = (inp[3]) ? 16'b0000001111111111 : 16'b0000001111111111;
												assign node4955 = (inp[5]) ? node4963 : node4956;
													assign node4956 = (inp[4]) ? node4960 : node4957;
														assign node4957 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4960 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4963 = (inp[4]) ? node4967 : node4964;
														assign node4964 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4967 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node4970 = (inp[7]) ? node4986 : node4971;
												assign node4971 = (inp[8]) ? node4979 : node4972;
													assign node4972 = (inp[3]) ? node4976 : node4973;
														assign node4973 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node4976 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node4979 = (inp[5]) ? node4983 : node4980;
														assign node4980 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node4983 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node4986 = (inp[5]) ? node4994 : node4987;
													assign node4987 = (inp[0]) ? node4991 : node4988;
														assign node4988 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node4991 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node4994 = (inp[3]) ? node4998 : node4995;
														assign node4995 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node4998 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
									assign node5001 = (inp[3]) ? node5063 : node5002;
										assign node5002 = (inp[4]) ? node5034 : node5003;
											assign node5003 = (inp[10]) ? node5019 : node5004;
												assign node5004 = (inp[5]) ? node5012 : node5005;
													assign node5005 = (inp[8]) ? node5009 : node5006;
														assign node5006 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node5009 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5012 = (inp[7]) ? node5016 : node5013;
														assign node5013 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5016 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5019 = (inp[0]) ? node5027 : node5020;
													assign node5020 = (inp[5]) ? node5024 : node5021;
														assign node5021 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5024 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5027 = (inp[2]) ? node5031 : node5028;
														assign node5028 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5031 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5034 = (inp[5]) ? node5050 : node5035;
												assign node5035 = (inp[2]) ? node5043 : node5036;
													assign node5036 = (inp[8]) ? node5040 : node5037;
														assign node5037 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5040 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5043 = (inp[0]) ? node5047 : node5044;
														assign node5044 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5047 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5050 = (inp[0]) ? node5056 : node5051;
													assign node5051 = (inp[10]) ? node5053 : 16'b0000000111111111;
														assign node5053 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5056 = (inp[8]) ? node5060 : node5057;
														assign node5057 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5060 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node5063 = (inp[4]) ? node5095 : node5064;
											assign node5064 = (inp[5]) ? node5080 : node5065;
												assign node5065 = (inp[10]) ? node5073 : node5066;
													assign node5066 = (inp[7]) ? node5070 : node5067;
														assign node5067 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5070 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5073 = (inp[8]) ? node5077 : node5074;
														assign node5074 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5077 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5080 = (inp[0]) ? node5088 : node5081;
													assign node5081 = (inp[2]) ? node5085 : node5082;
														assign node5082 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5085 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5088 = (inp[7]) ? node5092 : node5089;
														assign node5089 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5092 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node5095 = (inp[7]) ? node5109 : node5096;
												assign node5096 = (inp[10]) ? node5102 : node5097;
													assign node5097 = (inp[5]) ? node5099 : 16'b0000001111111111;
														assign node5099 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5102 = (inp[5]) ? node5106 : node5103;
														assign node5103 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5106 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node5109 = (inp[2]) ? node5117 : node5110;
													assign node5110 = (inp[10]) ? node5114 : node5111;
														assign node5111 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node5114 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5117 = (inp[0]) ? node5121 : node5118;
														assign node5118 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node5121 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node5124 = (inp[4]) ? node5246 : node5125;
									assign node5125 = (inp[3]) ? node5187 : node5126;
										assign node5126 = (inp[8]) ? node5156 : node5127;
											assign node5127 = (inp[2]) ? node5143 : node5128;
												assign node5128 = (inp[5]) ? node5136 : node5129;
													assign node5129 = (inp[7]) ? node5133 : node5130;
														assign node5130 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node5133 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5136 = (inp[0]) ? node5140 : node5137;
														assign node5137 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5140 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5143 = (inp[11]) ? node5151 : node5144;
													assign node5144 = (inp[7]) ? node5148 : node5145;
														assign node5145 = (inp[5]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node5148 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5151 = (inp[5]) ? 16'b0000000011111111 : node5152;
														assign node5152 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5156 = (inp[0]) ? node5172 : node5157;
												assign node5157 = (inp[7]) ? node5165 : node5158;
													assign node5158 = (inp[5]) ? node5162 : node5159;
														assign node5159 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5162 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5165 = (inp[10]) ? node5169 : node5166;
														assign node5166 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node5169 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5172 = (inp[11]) ? node5180 : node5173;
													assign node5173 = (inp[10]) ? node5177 : node5174;
														assign node5174 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5177 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5180 = (inp[2]) ? node5184 : node5181;
														assign node5181 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5184 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000001111111;
										assign node5187 = (inp[7]) ? node5219 : node5188;
											assign node5188 = (inp[11]) ? node5204 : node5189;
												assign node5189 = (inp[0]) ? node5197 : node5190;
													assign node5190 = (inp[2]) ? node5194 : node5191;
														assign node5191 = (inp[10]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node5194 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5197 = (inp[2]) ? node5201 : node5198;
														assign node5198 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5201 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5204 = (inp[8]) ? node5212 : node5205;
													assign node5205 = (inp[10]) ? node5209 : node5206;
														assign node5206 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5209 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5212 = (inp[0]) ? node5216 : node5213;
														assign node5213 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5216 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5219 = (inp[11]) ? node5233 : node5220;
												assign node5220 = (inp[0]) ? node5226 : node5221;
													assign node5221 = (inp[2]) ? node5223 : 16'b0000001111111111;
														assign node5223 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5226 = (inp[10]) ? node5230 : node5227;
														assign node5227 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5230 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5233 = (inp[5]) ? node5241 : node5234;
													assign node5234 = (inp[8]) ? node5238 : node5235;
														assign node5235 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node5238 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5241 = (inp[2]) ? 16'b0000000000111111 : node5242;
														assign node5242 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node5246 = (inp[0]) ? node5306 : node5247;
										assign node5247 = (inp[8]) ? node5275 : node5248;
											assign node5248 = (inp[2]) ? node5262 : node5249;
												assign node5249 = (inp[7]) ? node5255 : node5250;
													assign node5250 = (inp[10]) ? 16'b0000001111111111 : node5251;
														assign node5251 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5255 = (inp[10]) ? node5259 : node5256;
														assign node5256 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5259 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node5262 = (inp[3]) ? node5270 : node5263;
													assign node5263 = (inp[11]) ? node5267 : node5264;
														assign node5264 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5267 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node5270 = (inp[11]) ? 16'b0000000011111111 : node5271;
														assign node5271 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5275 = (inp[10]) ? node5291 : node5276;
												assign node5276 = (inp[7]) ? node5284 : node5277;
													assign node5277 = (inp[5]) ? node5281 : node5278;
														assign node5278 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5281 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5284 = (inp[2]) ? node5288 : node5285;
														assign node5285 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5288 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5291 = (inp[3]) ? node5299 : node5292;
													assign node5292 = (inp[11]) ? node5296 : node5293;
														assign node5293 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node5296 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5299 = (inp[2]) ? node5303 : node5300;
														assign node5300 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node5303 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node5306 = (inp[2]) ? node5336 : node5307;
											assign node5307 = (inp[7]) ? node5321 : node5308;
												assign node5308 = (inp[11]) ? node5314 : node5309;
													assign node5309 = (inp[5]) ? node5311 : 16'b0000000111111111;
														assign node5311 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5314 = (inp[8]) ? node5318 : node5315;
														assign node5315 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5318 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5321 = (inp[10]) ? node5329 : node5322;
													assign node5322 = (inp[5]) ? node5326 : node5323;
														assign node5323 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node5326 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5329 = (inp[8]) ? node5333 : node5330;
														assign node5330 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5333 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5336 = (inp[5]) ? node5344 : node5337;
												assign node5337 = (inp[3]) ? node5339 : 16'b0000000011111111;
													assign node5339 = (inp[11]) ? node5341 : 16'b0000000011111111;
														assign node5341 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5344 = (inp[11]) ? node5352 : node5345;
													assign node5345 = (inp[7]) ? node5349 : node5346;
														assign node5346 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5349 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node5352 = (inp[10]) ? node5356 : node5353;
														assign node5353 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5356 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
							assign node5359 = (inp[12]) ? node5601 : node5360;
								assign node5360 = (inp[7]) ? node5478 : node5361;
									assign node5361 = (inp[2]) ? node5415 : node5362;
										assign node5362 = (inp[3]) ? node5390 : node5363;
											assign node5363 = (inp[5]) ? node5379 : node5364;
												assign node5364 = (inp[10]) ? node5372 : node5365;
													assign node5365 = (inp[8]) ? node5369 : node5366;
														assign node5366 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node5369 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5372 = (inp[8]) ? node5376 : node5373;
														assign node5373 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5376 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5379 = (inp[8]) ? node5387 : node5380;
													assign node5380 = (inp[11]) ? node5384 : node5381;
														assign node5381 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5384 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5387 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5390 = (inp[11]) ? node5402 : node5391;
												assign node5391 = (inp[0]) ? node5399 : node5392;
													assign node5392 = (inp[4]) ? node5396 : node5393;
														assign node5393 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5396 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5399 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5402 = (inp[5]) ? node5410 : node5403;
													assign node5403 = (inp[0]) ? node5407 : node5404;
														assign node5404 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5407 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5410 = (inp[8]) ? node5412 : 16'b0000000011111111;
														assign node5412 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
										assign node5415 = (inp[0]) ? node5447 : node5416;
											assign node5416 = (inp[4]) ? node5432 : node5417;
												assign node5417 = (inp[10]) ? node5425 : node5418;
													assign node5418 = (inp[5]) ? node5422 : node5419;
														assign node5419 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5422 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5425 = (inp[3]) ? node5429 : node5426;
														assign node5426 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5429 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5432 = (inp[3]) ? node5440 : node5433;
													assign node5433 = (inp[11]) ? node5437 : node5434;
														assign node5434 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5437 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5440 = (inp[8]) ? node5444 : node5441;
														assign node5441 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node5444 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5447 = (inp[5]) ? node5463 : node5448;
												assign node5448 = (inp[10]) ? node5456 : node5449;
													assign node5449 = (inp[8]) ? node5453 : node5450;
														assign node5450 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5453 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node5456 = (inp[11]) ? node5460 : node5457;
														assign node5457 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5460 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5463 = (inp[8]) ? node5471 : node5464;
													assign node5464 = (inp[10]) ? node5468 : node5465;
														assign node5465 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5468 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5471 = (inp[10]) ? node5475 : node5472;
														assign node5472 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node5475 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5478 = (inp[4]) ? node5540 : node5479;
										assign node5479 = (inp[10]) ? node5511 : node5480;
											assign node5480 = (inp[8]) ? node5496 : node5481;
												assign node5481 = (inp[0]) ? node5489 : node5482;
													assign node5482 = (inp[2]) ? node5486 : node5483;
														assign node5483 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5486 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5489 = (inp[2]) ? node5493 : node5490;
														assign node5490 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5493 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5496 = (inp[3]) ? node5504 : node5497;
													assign node5497 = (inp[5]) ? node5501 : node5498;
														assign node5498 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5501 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5504 = (inp[11]) ? node5508 : node5505;
														assign node5505 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5508 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5511 = (inp[5]) ? node5527 : node5512;
												assign node5512 = (inp[3]) ? node5520 : node5513;
													assign node5513 = (inp[8]) ? node5517 : node5514;
														assign node5514 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5517 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5520 = (inp[11]) ? node5524 : node5521;
														assign node5521 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5524 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5527 = (inp[3]) ? node5533 : node5528;
													assign node5528 = (inp[11]) ? node5530 : 16'b0000000011111111;
														assign node5530 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5533 = (inp[2]) ? node5537 : node5534;
														assign node5534 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5537 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
										assign node5540 = (inp[5]) ? node5572 : node5541;
											assign node5541 = (inp[10]) ? node5557 : node5542;
												assign node5542 = (inp[3]) ? node5550 : node5543;
													assign node5543 = (inp[2]) ? node5547 : node5544;
														assign node5544 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node5547 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5550 = (inp[0]) ? node5554 : node5551;
														assign node5551 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5554 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5557 = (inp[0]) ? node5565 : node5558;
													assign node5558 = (inp[8]) ? node5562 : node5559;
														assign node5559 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node5562 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5565 = (inp[2]) ? node5569 : node5566;
														assign node5566 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node5569 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node5572 = (inp[3]) ? node5586 : node5573;
												assign node5573 = (inp[0]) ? node5579 : node5574;
													assign node5574 = (inp[8]) ? node5576 : 16'b0000000011111111;
														assign node5576 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5579 = (inp[2]) ? node5583 : node5580;
														assign node5580 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5583 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5586 = (inp[0]) ? node5594 : node5587;
													assign node5587 = (inp[2]) ? node5591 : node5588;
														assign node5588 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node5591 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5594 = (inp[2]) ? node5598 : node5595;
														assign node5595 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node5598 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000011111;
								assign node5601 = (inp[0]) ? node5723 : node5602;
									assign node5602 = (inp[8]) ? node5662 : node5603;
										assign node5603 = (inp[3]) ? node5631 : node5604;
											assign node5604 = (inp[11]) ? node5618 : node5605;
												assign node5605 = (inp[7]) ? node5611 : node5606;
													assign node5606 = (inp[5]) ? node5608 : 16'b0000001111111111;
														assign node5608 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5611 = (inp[2]) ? node5615 : node5612;
														assign node5612 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5615 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node5618 = (inp[2]) ? node5626 : node5619;
													assign node5619 = (inp[5]) ? node5623 : node5620;
														assign node5620 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node5623 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5626 = (inp[5]) ? node5628 : 16'b0000000111111111;
														assign node5628 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node5631 = (inp[10]) ? node5647 : node5632;
												assign node5632 = (inp[2]) ? node5640 : node5633;
													assign node5633 = (inp[11]) ? node5637 : node5634;
														assign node5634 = (inp[4]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node5637 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5640 = (inp[4]) ? node5644 : node5641;
														assign node5641 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5644 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node5647 = (inp[4]) ? node5655 : node5648;
													assign node5648 = (inp[7]) ? node5652 : node5649;
														assign node5649 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5652 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5655 = (inp[5]) ? node5659 : node5656;
														assign node5656 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5659 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
										assign node5662 = (inp[4]) ? node5692 : node5663;
											assign node5663 = (inp[11]) ? node5679 : node5664;
												assign node5664 = (inp[2]) ? node5672 : node5665;
													assign node5665 = (inp[5]) ? node5669 : node5666;
														assign node5666 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5669 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5672 = (inp[3]) ? node5676 : node5673;
														assign node5673 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node5676 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5679 = (inp[5]) ? node5685 : node5680;
													assign node5680 = (inp[7]) ? node5682 : 16'b0000000111111111;
														assign node5682 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5685 = (inp[7]) ? node5689 : node5686;
														assign node5686 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5689 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node5692 = (inp[11]) ? node5708 : node5693;
												assign node5693 = (inp[7]) ? node5701 : node5694;
													assign node5694 = (inp[2]) ? node5698 : node5695;
														assign node5695 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node5698 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5701 = (inp[3]) ? node5705 : node5702;
														assign node5702 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5705 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5708 = (inp[7]) ? node5716 : node5709;
													assign node5709 = (inp[3]) ? node5713 : node5710;
														assign node5710 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node5713 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5716 = (inp[10]) ? node5720 : node5717;
														assign node5717 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5720 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node5723 = (inp[4]) ? node5783 : node5724;
										assign node5724 = (inp[8]) ? node5754 : node5725;
											assign node5725 = (inp[11]) ? node5739 : node5726;
												assign node5726 = (inp[3]) ? node5732 : node5727;
													assign node5727 = (inp[7]) ? node5729 : 16'b0000001111111111;
														assign node5729 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5732 = (inp[5]) ? node5736 : node5733;
														assign node5733 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5736 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node5739 = (inp[2]) ? node5747 : node5740;
													assign node5740 = (inp[3]) ? node5744 : node5741;
														assign node5741 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5744 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node5747 = (inp[10]) ? node5751 : node5748;
														assign node5748 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5751 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node5754 = (inp[10]) ? node5768 : node5755;
												assign node5755 = (inp[7]) ? node5761 : node5756;
													assign node5756 = (inp[2]) ? 16'b0000000011111111 : node5757;
														assign node5757 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node5761 = (inp[2]) ? node5765 : node5762;
														assign node5762 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5765 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node5768 = (inp[3]) ? node5776 : node5769;
													assign node5769 = (inp[5]) ? node5773 : node5770;
														assign node5770 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5773 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5776 = (inp[7]) ? node5780 : node5777;
														assign node5777 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5780 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node5783 = (inp[7]) ? node5815 : node5784;
											assign node5784 = (inp[2]) ? node5800 : node5785;
												assign node5785 = (inp[8]) ? node5793 : node5786;
													assign node5786 = (inp[5]) ? node5790 : node5787;
														assign node5787 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node5790 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node5793 = (inp[11]) ? node5797 : node5794;
														assign node5794 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node5797 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node5800 = (inp[11]) ? node5808 : node5801;
													assign node5801 = (inp[3]) ? node5805 : node5802;
														assign node5802 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node5805 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5808 = (inp[5]) ? node5812 : node5809;
														assign node5809 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5812 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node5815 = (inp[2]) ? node5831 : node5816;
												assign node5816 = (inp[8]) ? node5824 : node5817;
													assign node5817 = (inp[3]) ? node5821 : node5818;
														assign node5818 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node5821 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node5824 = (inp[3]) ? node5828 : node5825;
														assign node5825 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5828 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node5831 = (inp[3]) ? node5839 : node5832;
													assign node5832 = (inp[5]) ? node5836 : node5833;
														assign node5833 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node5836 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node5839 = (inp[11]) ? node5843 : node5840;
														assign node5840 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node5843 = (inp[10]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node5846 = (inp[0]) ? node6824 : node5847;
						assign node5847 = (inp[3]) ? node6329 : node5848;
							assign node5848 = (inp[7]) ? node6086 : node5849;
								assign node5849 = (inp[14]) ? node5969 : node5850;
									assign node5850 = (inp[12]) ? node5910 : node5851;
										assign node5851 = (inp[15]) ? node5883 : node5852;
											assign node5852 = (inp[11]) ? node5868 : node5853;
												assign node5853 = (inp[2]) ? node5861 : node5854;
													assign node5854 = (inp[4]) ? node5858 : node5855;
														assign node5855 = (inp[10]) ? 16'b0001111111111111 : 16'b0001111111111111;
														assign node5858 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5861 = (inp[8]) ? node5865 : node5862;
														assign node5862 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node5865 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5868 = (inp[4]) ? node5876 : node5869;
													assign node5869 = (inp[10]) ? node5873 : node5870;
														assign node5870 = (inp[8]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node5873 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5876 = (inp[10]) ? node5880 : node5877;
														assign node5877 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5880 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node5883 = (inp[8]) ? node5897 : node5884;
												assign node5884 = (inp[11]) ? node5892 : node5885;
													assign node5885 = (inp[10]) ? node5889 : node5886;
														assign node5886 = (inp[5]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node5889 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5892 = (inp[2]) ? 16'b0000001111111111 : node5893;
														assign node5893 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5897 = (inp[10]) ? node5905 : node5898;
													assign node5898 = (inp[2]) ? node5902 : node5899;
														assign node5899 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5902 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5905 = (inp[11]) ? 16'b0000000111111111 : node5906;
														assign node5906 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node5910 = (inp[10]) ? node5940 : node5911;
											assign node5911 = (inp[8]) ? node5925 : node5912;
												assign node5912 = (inp[2]) ? node5918 : node5913;
													assign node5913 = (inp[11]) ? 16'b0000011111111111 : node5914;
														assign node5914 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node5918 = (inp[4]) ? node5922 : node5919;
														assign node5919 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5922 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node5925 = (inp[15]) ? node5933 : node5926;
													assign node5926 = (inp[11]) ? node5930 : node5927;
														assign node5927 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5930 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node5933 = (inp[11]) ? node5937 : node5934;
														assign node5934 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5937 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node5940 = (inp[5]) ? node5954 : node5941;
												assign node5941 = (inp[11]) ? node5947 : node5942;
													assign node5942 = (inp[15]) ? 16'b0000001111111111 : node5943;
														assign node5943 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5947 = (inp[8]) ? node5951 : node5948;
														assign node5948 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node5951 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node5954 = (inp[2]) ? node5962 : node5955;
													assign node5955 = (inp[15]) ? node5959 : node5956;
														assign node5956 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node5959 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node5962 = (inp[15]) ? node5966 : node5963;
														assign node5963 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node5966 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node5969 = (inp[4]) ? node6027 : node5970;
										assign node5970 = (inp[2]) ? node6000 : node5971;
											assign node5971 = (inp[8]) ? node5985 : node5972;
												assign node5972 = (inp[11]) ? node5980 : node5973;
													assign node5973 = (inp[12]) ? node5977 : node5974;
														assign node5974 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node5977 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node5980 = (inp[10]) ? 16'b0000001111111111 : node5981;
														assign node5981 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node5985 = (inp[5]) ? node5993 : node5986;
													assign node5986 = (inp[11]) ? node5990 : node5987;
														assign node5987 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node5990 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node5993 = (inp[12]) ? node5997 : node5994;
														assign node5994 = (inp[10]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node5997 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6000 = (inp[15]) ? node6014 : node6001;
												assign node6001 = (inp[11]) ? node6009 : node6002;
													assign node6002 = (inp[8]) ? node6006 : node6003;
														assign node6003 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6006 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6009 = (inp[8]) ? node6011 : 16'b0000000111111111;
														assign node6011 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6014 = (inp[8]) ? node6020 : node6015;
													assign node6015 = (inp[10]) ? 16'b0000000111111111 : node6016;
														assign node6016 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node6020 = (inp[10]) ? node6024 : node6021;
														assign node6021 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6024 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6027 = (inp[12]) ? node6057 : node6028;
											assign node6028 = (inp[11]) ? node6044 : node6029;
												assign node6029 = (inp[10]) ? node6037 : node6030;
													assign node6030 = (inp[5]) ? node6034 : node6031;
														assign node6031 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6034 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6037 = (inp[5]) ? node6041 : node6038;
														assign node6038 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6041 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6044 = (inp[2]) ? node6052 : node6045;
													assign node6045 = (inp[8]) ? node6049 : node6046;
														assign node6046 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6049 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6052 = (inp[8]) ? 16'b0000000011111111 : node6053;
														assign node6053 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6057 = (inp[15]) ? node6073 : node6058;
												assign node6058 = (inp[2]) ? node6066 : node6059;
													assign node6059 = (inp[8]) ? node6063 : node6060;
														assign node6060 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6063 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6066 = (inp[11]) ? node6070 : node6067;
														assign node6067 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node6070 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node6073 = (inp[5]) ? node6081 : node6074;
													assign node6074 = (inp[11]) ? node6078 : node6075;
														assign node6075 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6078 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6081 = (inp[8]) ? 16'b0000000001111111 : node6082;
														assign node6082 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000001111111;
								assign node6086 = (inp[5]) ? node6208 : node6087;
									assign node6087 = (inp[10]) ? node6147 : node6088;
										assign node6088 = (inp[8]) ? node6118 : node6089;
											assign node6089 = (inp[12]) ? node6103 : node6090;
												assign node6090 = (inp[11]) ? node6098 : node6091;
													assign node6091 = (inp[14]) ? node6095 : node6092;
														assign node6092 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6095 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6098 = (inp[15]) ? 16'b0000000111111111 : node6099;
														assign node6099 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node6103 = (inp[14]) ? node6111 : node6104;
													assign node6104 = (inp[2]) ? node6108 : node6105;
														assign node6105 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6108 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6111 = (inp[15]) ? node6115 : node6112;
														assign node6112 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6115 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node6118 = (inp[2]) ? node6132 : node6119;
												assign node6119 = (inp[11]) ? node6125 : node6120;
													assign node6120 = (inp[12]) ? 16'b0000001111111111 : node6121;
														assign node6121 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6125 = (inp[14]) ? node6129 : node6126;
														assign node6126 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6129 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node6132 = (inp[14]) ? node6140 : node6133;
													assign node6133 = (inp[4]) ? node6137 : node6134;
														assign node6134 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6137 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6140 = (inp[15]) ? node6144 : node6141;
														assign node6141 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6144 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6147 = (inp[15]) ? node6177 : node6148;
											assign node6148 = (inp[12]) ? node6162 : node6149;
												assign node6149 = (inp[2]) ? node6157 : node6150;
													assign node6150 = (inp[8]) ? node6154 : node6151;
														assign node6151 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6154 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6157 = (inp[14]) ? 16'b0000000011111111 : node6158;
														assign node6158 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6162 = (inp[2]) ? node6170 : node6163;
													assign node6163 = (inp[4]) ? node6167 : node6164;
														assign node6164 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node6167 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6170 = (inp[8]) ? node6174 : node6171;
														assign node6171 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6174 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6177 = (inp[14]) ? node6193 : node6178;
												assign node6178 = (inp[4]) ? node6186 : node6179;
													assign node6179 = (inp[11]) ? node6183 : node6180;
														assign node6180 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6183 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6186 = (inp[11]) ? node6190 : node6187;
														assign node6187 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6190 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node6193 = (inp[12]) ? node6201 : node6194;
													assign node6194 = (inp[8]) ? node6198 : node6195;
														assign node6195 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node6198 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6201 = (inp[4]) ? node6205 : node6202;
														assign node6202 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node6205 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
									assign node6208 = (inp[2]) ? node6270 : node6209;
										assign node6209 = (inp[4]) ? node6239 : node6210;
											assign node6210 = (inp[11]) ? node6226 : node6211;
												assign node6211 = (inp[14]) ? node6219 : node6212;
													assign node6212 = (inp[10]) ? node6216 : node6213;
														assign node6213 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6216 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6219 = (inp[15]) ? node6223 : node6220;
														assign node6220 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6223 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6226 = (inp[8]) ? node6232 : node6227;
													assign node6227 = (inp[15]) ? node6229 : 16'b0000001111111111;
														assign node6229 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6232 = (inp[12]) ? node6236 : node6233;
														assign node6233 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6236 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node6239 = (inp[10]) ? node6255 : node6240;
												assign node6240 = (inp[8]) ? node6248 : node6241;
													assign node6241 = (inp[12]) ? node6245 : node6242;
														assign node6242 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6245 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6248 = (inp[14]) ? node6252 : node6249;
														assign node6249 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6252 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6255 = (inp[15]) ? node6263 : node6256;
													assign node6256 = (inp[11]) ? node6260 : node6257;
														assign node6257 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6260 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6263 = (inp[8]) ? node6267 : node6264;
														assign node6264 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6267 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node6270 = (inp[12]) ? node6300 : node6271;
											assign node6271 = (inp[14]) ? node6287 : node6272;
												assign node6272 = (inp[15]) ? node6280 : node6273;
													assign node6273 = (inp[11]) ? node6277 : node6274;
														assign node6274 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6277 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6280 = (inp[4]) ? node6284 : node6281;
														assign node6281 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6284 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6287 = (inp[4]) ? node6293 : node6288;
													assign node6288 = (inp[10]) ? node6290 : 16'b0000001111111111;
														assign node6290 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6293 = (inp[15]) ? node6297 : node6294;
														assign node6294 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node6297 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6300 = (inp[11]) ? node6314 : node6301;
												assign node6301 = (inp[15]) ? node6309 : node6302;
													assign node6302 = (inp[8]) ? node6306 : node6303;
														assign node6303 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6306 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6309 = (inp[4]) ? node6311 : 16'b0000000001111111;
														assign node6311 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6314 = (inp[10]) ? node6322 : node6315;
													assign node6315 = (inp[4]) ? node6319 : node6316;
														assign node6316 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node6319 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6322 = (inp[14]) ? node6326 : node6323;
														assign node6323 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node6326 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node6329 = (inp[8]) ? node6579 : node6330;
								assign node6330 = (inp[14]) ? node6454 : node6331;
									assign node6331 = (inp[15]) ? node6393 : node6332;
										assign node6332 = (inp[11]) ? node6364 : node6333;
											assign node6333 = (inp[4]) ? node6349 : node6334;
												assign node6334 = (inp[12]) ? node6342 : node6335;
													assign node6335 = (inp[2]) ? node6339 : node6336;
														assign node6336 = (inp[10]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6339 = (inp[5]) ? 16'b0000001111111111 : 16'b0000001111111111;
													assign node6342 = (inp[7]) ? node6346 : node6343;
														assign node6343 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6346 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6349 = (inp[2]) ? node6357 : node6350;
													assign node6350 = (inp[12]) ? node6354 : node6351;
														assign node6351 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6354 = (inp[10]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6357 = (inp[12]) ? node6361 : node6358;
														assign node6358 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6361 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node6364 = (inp[7]) ? node6380 : node6365;
												assign node6365 = (inp[4]) ? node6373 : node6366;
													assign node6366 = (inp[5]) ? node6370 : node6367;
														assign node6367 = (inp[10]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6370 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6373 = (inp[12]) ? node6377 : node6374;
														assign node6374 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node6377 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6380 = (inp[4]) ? node6388 : node6381;
													assign node6381 = (inp[2]) ? node6385 : node6382;
														assign node6382 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6385 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6388 = (inp[5]) ? 16'b0000000011111111 : node6389;
														assign node6389 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
										assign node6393 = (inp[5]) ? node6425 : node6394;
											assign node6394 = (inp[4]) ? node6410 : node6395;
												assign node6395 = (inp[10]) ? node6403 : node6396;
													assign node6396 = (inp[2]) ? node6400 : node6397;
														assign node6397 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6400 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6403 = (inp[2]) ? node6407 : node6404;
														assign node6404 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6407 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6410 = (inp[11]) ? node6418 : node6411;
													assign node6411 = (inp[10]) ? node6415 : node6412;
														assign node6412 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6415 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6418 = (inp[2]) ? node6422 : node6419;
														assign node6419 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6422 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node6425 = (inp[7]) ? node6439 : node6426;
												assign node6426 = (inp[11]) ? node6432 : node6427;
													assign node6427 = (inp[10]) ? 16'b0000000111111111 : node6428;
														assign node6428 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6432 = (inp[10]) ? node6436 : node6433;
														assign node6433 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6436 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6439 = (inp[12]) ? node6447 : node6440;
													assign node6440 = (inp[4]) ? node6444 : node6441;
														assign node6441 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6444 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node6447 = (inp[10]) ? node6451 : node6448;
														assign node6448 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6451 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node6454 = (inp[7]) ? node6518 : node6455;
										assign node6455 = (inp[12]) ? node6487 : node6456;
											assign node6456 = (inp[11]) ? node6472 : node6457;
												assign node6457 = (inp[10]) ? node6465 : node6458;
													assign node6458 = (inp[2]) ? node6462 : node6459;
														assign node6459 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6462 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6465 = (inp[4]) ? node6469 : node6466;
														assign node6466 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6469 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6472 = (inp[2]) ? node6480 : node6473;
													assign node6473 = (inp[10]) ? node6477 : node6474;
														assign node6474 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6477 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6480 = (inp[4]) ? node6484 : node6481;
														assign node6481 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6484 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6487 = (inp[11]) ? node6503 : node6488;
												assign node6488 = (inp[2]) ? node6496 : node6489;
													assign node6489 = (inp[4]) ? node6493 : node6490;
														assign node6490 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6493 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node6496 = (inp[5]) ? node6500 : node6497;
														assign node6497 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6500 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6503 = (inp[10]) ? node6511 : node6504;
													assign node6504 = (inp[2]) ? node6508 : node6505;
														assign node6505 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6508 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node6511 = (inp[5]) ? node6515 : node6512;
														assign node6512 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node6515 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6518 = (inp[10]) ? node6548 : node6519;
											assign node6519 = (inp[11]) ? node6535 : node6520;
												assign node6520 = (inp[2]) ? node6528 : node6521;
													assign node6521 = (inp[12]) ? node6525 : node6522;
														assign node6522 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6525 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6528 = (inp[5]) ? node6532 : node6529;
														assign node6529 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6532 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6535 = (inp[15]) ? node6541 : node6536;
													assign node6536 = (inp[4]) ? node6538 : 16'b0000000111111111;
														assign node6538 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6541 = (inp[2]) ? node6545 : node6542;
														assign node6542 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6545 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node6548 = (inp[4]) ? node6564 : node6549;
												assign node6549 = (inp[5]) ? node6557 : node6550;
													assign node6550 = (inp[2]) ? node6554 : node6551;
														assign node6551 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6554 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6557 = (inp[2]) ? node6561 : node6558;
														assign node6558 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6561 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node6564 = (inp[2]) ? node6572 : node6565;
													assign node6565 = (inp[15]) ? node6569 : node6566;
														assign node6566 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6569 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6572 = (inp[12]) ? node6576 : node6573;
														assign node6573 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node6576 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node6579 = (inp[4]) ? node6701 : node6580;
									assign node6580 = (inp[5]) ? node6640 : node6581;
										assign node6581 = (inp[11]) ? node6613 : node6582;
											assign node6582 = (inp[2]) ? node6598 : node6583;
												assign node6583 = (inp[10]) ? node6591 : node6584;
													assign node6584 = (inp[14]) ? node6588 : node6585;
														assign node6585 = (inp[7]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node6588 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6591 = (inp[12]) ? node6595 : node6592;
														assign node6592 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node6595 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node6598 = (inp[12]) ? node6606 : node6599;
													assign node6599 = (inp[7]) ? node6603 : node6600;
														assign node6600 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node6603 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6606 = (inp[10]) ? node6610 : node6607;
														assign node6607 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6610 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6613 = (inp[7]) ? node6627 : node6614;
												assign node6614 = (inp[15]) ? node6622 : node6615;
													assign node6615 = (inp[10]) ? node6619 : node6616;
														assign node6616 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6619 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node6622 = (inp[10]) ? 16'b0000000011111111 : node6623;
														assign node6623 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node6627 = (inp[14]) ? node6635 : node6628;
													assign node6628 = (inp[2]) ? node6632 : node6629;
														assign node6629 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6632 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node6635 = (inp[12]) ? 16'b0000000001111111 : node6636;
														assign node6636 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6640 = (inp[10]) ? node6672 : node6641;
											assign node6641 = (inp[15]) ? node6657 : node6642;
												assign node6642 = (inp[14]) ? node6650 : node6643;
													assign node6643 = (inp[11]) ? node6647 : node6644;
														assign node6644 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6647 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6650 = (inp[12]) ? node6654 : node6651;
														assign node6651 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node6654 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6657 = (inp[7]) ? node6665 : node6658;
													assign node6658 = (inp[12]) ? node6662 : node6659;
														assign node6659 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6662 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6665 = (inp[2]) ? node6669 : node6666;
														assign node6666 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6669 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node6672 = (inp[15]) ? node6686 : node6673;
												assign node6673 = (inp[14]) ? node6679 : node6674;
													assign node6674 = (inp[11]) ? 16'b0000000011111111 : node6675;
														assign node6675 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6679 = (inp[11]) ? node6683 : node6680;
														assign node6680 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6683 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6686 = (inp[7]) ? node6694 : node6687;
													assign node6687 = (inp[2]) ? node6691 : node6688;
														assign node6688 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node6691 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6694 = (inp[12]) ? node6698 : node6695;
														assign node6695 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node6698 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node6701 = (inp[15]) ? node6763 : node6702;
										assign node6702 = (inp[10]) ? node6732 : node6703;
											assign node6703 = (inp[2]) ? node6719 : node6704;
												assign node6704 = (inp[7]) ? node6712 : node6705;
													assign node6705 = (inp[5]) ? node6709 : node6706;
														assign node6706 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6709 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6712 = (inp[11]) ? node6716 : node6713;
														assign node6713 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node6716 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6719 = (inp[14]) ? node6725 : node6720;
													assign node6720 = (inp[7]) ? node6722 : 16'b0000000011111111;
														assign node6722 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6725 = (inp[12]) ? node6729 : node6726;
														assign node6726 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node6729 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node6732 = (inp[5]) ? node6748 : node6733;
												assign node6733 = (inp[7]) ? node6741 : node6734;
													assign node6734 = (inp[14]) ? node6738 : node6735;
														assign node6735 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6738 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node6741 = (inp[11]) ? node6745 : node6742;
														assign node6742 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node6745 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6748 = (inp[12]) ? node6756 : node6749;
													assign node6749 = (inp[7]) ? node6753 : node6750;
														assign node6750 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node6753 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node6756 = (inp[2]) ? node6760 : node6757;
														assign node6757 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node6760 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node6763 = (inp[12]) ? node6795 : node6764;
											assign node6764 = (inp[7]) ? node6780 : node6765;
												assign node6765 = (inp[11]) ? node6773 : node6766;
													assign node6766 = (inp[14]) ? node6770 : node6767;
														assign node6767 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6770 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6773 = (inp[2]) ? node6777 : node6774;
														assign node6774 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node6777 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node6780 = (inp[5]) ? node6788 : node6781;
													assign node6781 = (inp[11]) ? node6785 : node6782;
														assign node6782 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node6785 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node6788 = (inp[14]) ? node6792 : node6789;
														assign node6789 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node6792 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node6795 = (inp[2]) ? node6809 : node6796;
												assign node6796 = (inp[7]) ? node6804 : node6797;
													assign node6797 = (inp[5]) ? node6801 : node6798;
														assign node6798 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node6801 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node6804 = (inp[11]) ? 16'b0000000000011111 : node6805;
														assign node6805 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node6809 = (inp[10]) ? node6817 : node6810;
													assign node6810 = (inp[5]) ? node6814 : node6811;
														assign node6811 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node6814 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node6817 = (inp[14]) ? node6821 : node6818;
														assign node6818 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node6821 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node6824 = (inp[2]) ? node7308 : node6825;
							assign node6825 = (inp[12]) ? node7065 : node6826;
								assign node6826 = (inp[7]) ? node6944 : node6827;
									assign node6827 = (inp[8]) ? node6885 : node6828;
										assign node6828 = (inp[3]) ? node6856 : node6829;
											assign node6829 = (inp[11]) ? node6845 : node6830;
												assign node6830 = (inp[4]) ? node6838 : node6831;
													assign node6831 = (inp[14]) ? node6835 : node6832;
														assign node6832 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node6835 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6838 = (inp[15]) ? node6842 : node6839;
														assign node6839 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6842 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node6845 = (inp[15]) ? node6851 : node6846;
													assign node6846 = (inp[5]) ? node6848 : 16'b0000011111111111;
														assign node6848 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6851 = (inp[5]) ? 16'b0000000001111111 : node6852;
														assign node6852 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node6856 = (inp[15]) ? node6870 : node6857;
												assign node6857 = (inp[4]) ? node6863 : node6858;
													assign node6858 = (inp[10]) ? 16'b0000001111111111 : node6859;
														assign node6859 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node6863 = (inp[5]) ? node6867 : node6864;
														assign node6864 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node6867 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6870 = (inp[10]) ? node6878 : node6871;
													assign node6871 = (inp[11]) ? node6875 : node6872;
														assign node6872 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6875 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6878 = (inp[5]) ? node6882 : node6879;
														assign node6879 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6882 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node6885 = (inp[10]) ? node6913 : node6886;
											assign node6886 = (inp[3]) ? node6900 : node6887;
												assign node6887 = (inp[4]) ? node6893 : node6888;
													assign node6888 = (inp[11]) ? 16'b0000001111111111 : node6889;
														assign node6889 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node6893 = (inp[11]) ? node6897 : node6894;
														assign node6894 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node6897 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6900 = (inp[11]) ? node6908 : node6901;
													assign node6901 = (inp[14]) ? node6905 : node6902;
														assign node6902 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6905 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6908 = (inp[14]) ? 16'b0000000011111111 : node6909;
														assign node6909 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node6913 = (inp[15]) ? node6929 : node6914;
												assign node6914 = (inp[14]) ? node6922 : node6915;
													assign node6915 = (inp[5]) ? node6919 : node6916;
														assign node6916 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6919 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6922 = (inp[4]) ? node6926 : node6923;
														assign node6923 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6926 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node6929 = (inp[14]) ? node6937 : node6930;
													assign node6930 = (inp[3]) ? node6934 : node6931;
														assign node6931 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node6934 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6937 = (inp[4]) ? node6941 : node6938;
														assign node6938 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node6941 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node6944 = (inp[11]) ? node7004 : node6945;
										assign node6945 = (inp[3]) ? node6973 : node6946;
											assign node6946 = (inp[15]) ? node6960 : node6947;
												assign node6947 = (inp[10]) ? node6955 : node6948;
													assign node6948 = (inp[5]) ? node6952 : node6949;
														assign node6949 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node6952 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node6955 = (inp[5]) ? node6957 : 16'b0000000111111111;
														assign node6957 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node6960 = (inp[4]) ? node6966 : node6961;
													assign node6961 = (inp[14]) ? node6963 : 16'b0000000111111111;
														assign node6963 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6966 = (inp[8]) ? node6970 : node6967;
														assign node6967 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6970 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node6973 = (inp[5]) ? node6989 : node6974;
												assign node6974 = (inp[10]) ? node6982 : node6975;
													assign node6975 = (inp[4]) ? node6979 : node6976;
														assign node6976 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node6979 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node6982 = (inp[4]) ? node6986 : node6983;
														assign node6983 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6986 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node6989 = (inp[4]) ? node6997 : node6990;
													assign node6990 = (inp[10]) ? node6994 : node6991;
														assign node6991 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node6994 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node6997 = (inp[15]) ? node7001 : node6998;
														assign node6998 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7001 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node7004 = (inp[14]) ? node7034 : node7005;
											assign node7005 = (inp[10]) ? node7021 : node7006;
												assign node7006 = (inp[8]) ? node7014 : node7007;
													assign node7007 = (inp[15]) ? node7011 : node7008;
														assign node7008 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7011 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7014 = (inp[4]) ? node7018 : node7015;
														assign node7015 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7018 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7021 = (inp[5]) ? node7029 : node7022;
													assign node7022 = (inp[8]) ? node7026 : node7023;
														assign node7023 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7026 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node7029 = (inp[8]) ? node7031 : 16'b0000000001111111;
														assign node7031 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7034 = (inp[4]) ? node7050 : node7035;
												assign node7035 = (inp[3]) ? node7043 : node7036;
													assign node7036 = (inp[15]) ? node7040 : node7037;
														assign node7037 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7040 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7043 = (inp[8]) ? node7047 : node7044;
														assign node7044 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7047 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7050 = (inp[5]) ? node7058 : node7051;
													assign node7051 = (inp[15]) ? node7055 : node7052;
														assign node7052 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node7055 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7058 = (inp[15]) ? node7062 : node7059;
														assign node7059 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7062 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node7065 = (inp[3]) ? node7187 : node7066;
									assign node7066 = (inp[4]) ? node7124 : node7067;
										assign node7067 = (inp[10]) ? node7095 : node7068;
											assign node7068 = (inp[7]) ? node7084 : node7069;
												assign node7069 = (inp[5]) ? node7077 : node7070;
													assign node7070 = (inp[11]) ? node7074 : node7071;
														assign node7071 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7074 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7077 = (inp[14]) ? node7081 : node7078;
														assign node7078 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7081 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node7084 = (inp[11]) ? node7090 : node7085;
													assign node7085 = (inp[8]) ? 16'b0000000111111111 : node7086;
														assign node7086 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7090 = (inp[8]) ? 16'b0000000011111111 : node7091;
														assign node7091 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node7095 = (inp[5]) ? node7111 : node7096;
												assign node7096 = (inp[7]) ? node7104 : node7097;
													assign node7097 = (inp[15]) ? node7101 : node7098;
														assign node7098 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7101 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7104 = (inp[8]) ? node7108 : node7105;
														assign node7105 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7108 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7111 = (inp[7]) ? node7119 : node7112;
													assign node7112 = (inp[15]) ? node7116 : node7113;
														assign node7113 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7116 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node7119 = (inp[8]) ? node7121 : 16'b0000000001111111;
														assign node7121 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7124 = (inp[11]) ? node7156 : node7125;
											assign node7125 = (inp[5]) ? node7141 : node7126;
												assign node7126 = (inp[15]) ? node7134 : node7127;
													assign node7127 = (inp[14]) ? node7131 : node7128;
														assign node7128 = (inp[10]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node7131 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7134 = (inp[7]) ? node7138 : node7135;
														assign node7135 = (inp[10]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7138 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7141 = (inp[8]) ? node7149 : node7142;
													assign node7142 = (inp[10]) ? node7146 : node7143;
														assign node7143 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7146 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000001111111;
													assign node7149 = (inp[7]) ? node7153 : node7150;
														assign node7150 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7153 = (inp[10]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node7156 = (inp[7]) ? node7172 : node7157;
												assign node7157 = (inp[10]) ? node7165 : node7158;
													assign node7158 = (inp[15]) ? node7162 : node7159;
														assign node7159 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7162 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7165 = (inp[8]) ? node7169 : node7166;
														assign node7166 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7169 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7172 = (inp[10]) ? node7180 : node7173;
													assign node7173 = (inp[5]) ? node7177 : node7174;
														assign node7174 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7177 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7180 = (inp[15]) ? node7184 : node7181;
														assign node7181 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7184 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7187 = (inp[8]) ? node7247 : node7188;
										assign node7188 = (inp[11]) ? node7216 : node7189;
											assign node7189 = (inp[10]) ? node7203 : node7190;
												assign node7190 = (inp[7]) ? node7196 : node7191;
													assign node7191 = (inp[14]) ? 16'b0000000111111111 : node7192;
														assign node7192 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7196 = (inp[5]) ? node7200 : node7197;
														assign node7197 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7200 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7203 = (inp[4]) ? node7211 : node7204;
													assign node7204 = (inp[5]) ? node7208 : node7205;
														assign node7205 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7208 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7211 = (inp[15]) ? node7213 : 16'b0000000011111111;
														assign node7213 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node7216 = (inp[5]) ? node7232 : node7217;
												assign node7217 = (inp[14]) ? node7225 : node7218;
													assign node7218 = (inp[15]) ? node7222 : node7219;
														assign node7219 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7222 = (inp[10]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node7225 = (inp[4]) ? node7229 : node7226;
														assign node7226 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7229 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7232 = (inp[7]) ? node7240 : node7233;
													assign node7233 = (inp[15]) ? node7237 : node7234;
														assign node7234 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7237 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node7240 = (inp[4]) ? node7244 : node7241;
														assign node7241 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node7244 = (inp[10]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7247 = (inp[4]) ? node7277 : node7248;
											assign node7248 = (inp[14]) ? node7262 : node7249;
												assign node7249 = (inp[10]) ? node7255 : node7250;
													assign node7250 = (inp[5]) ? 16'b0000000011111111 : node7251;
														assign node7251 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7255 = (inp[15]) ? node7259 : node7256;
														assign node7256 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7259 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7262 = (inp[5]) ? node7270 : node7263;
													assign node7263 = (inp[11]) ? node7267 : node7264;
														assign node7264 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node7267 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node7270 = (inp[10]) ? node7274 : node7271;
														assign node7271 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7274 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7277 = (inp[7]) ? node7293 : node7278;
												assign node7278 = (inp[5]) ? node7286 : node7279;
													assign node7279 = (inp[15]) ? node7283 : node7280;
														assign node7280 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7283 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7286 = (inp[15]) ? node7290 : node7287;
														assign node7287 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node7290 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7293 = (inp[5]) ? node7301 : node7294;
													assign node7294 = (inp[11]) ? node7298 : node7295;
														assign node7295 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node7298 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node7301 = (inp[10]) ? node7305 : node7302;
														assign node7302 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node7305 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node7308 = (inp[10]) ? node7548 : node7309;
								assign node7309 = (inp[3]) ? node7429 : node7310;
									assign node7310 = (inp[7]) ? node7368 : node7311;
										assign node7311 = (inp[12]) ? node7341 : node7312;
											assign node7312 = (inp[5]) ? node7328 : node7313;
												assign node7313 = (inp[15]) ? node7321 : node7314;
													assign node7314 = (inp[4]) ? node7318 : node7315;
														assign node7315 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7318 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7321 = (inp[14]) ? node7325 : node7322;
														assign node7322 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7325 = (inp[8]) ? 16'b0000000001111111 : 16'b0000001111111111;
												assign node7328 = (inp[4]) ? node7336 : node7329;
													assign node7329 = (inp[15]) ? node7333 : node7330;
														assign node7330 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7333 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7336 = (inp[14]) ? 16'b0000000001111111 : node7337;
														assign node7337 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node7341 = (inp[11]) ? node7355 : node7342;
												assign node7342 = (inp[8]) ? node7348 : node7343;
													assign node7343 = (inp[4]) ? node7345 : 16'b0000001111111111;
														assign node7345 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7348 = (inp[5]) ? node7352 : node7349;
														assign node7349 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7352 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7355 = (inp[4]) ? node7361 : node7356;
													assign node7356 = (inp[5]) ? 16'b0000000001111111 : node7357;
														assign node7357 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node7361 = (inp[8]) ? node7365 : node7362;
														assign node7362 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7365 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7368 = (inp[12]) ? node7400 : node7369;
											assign node7369 = (inp[11]) ? node7385 : node7370;
												assign node7370 = (inp[4]) ? node7378 : node7371;
													assign node7371 = (inp[5]) ? node7375 : node7372;
														assign node7372 = (inp[15]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node7375 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7378 = (inp[15]) ? node7382 : node7379;
														assign node7379 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7382 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7385 = (inp[5]) ? node7393 : node7386;
													assign node7386 = (inp[14]) ? node7390 : node7387;
														assign node7387 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7390 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node7393 = (inp[8]) ? node7397 : node7394;
														assign node7394 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7397 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7400 = (inp[8]) ? node7414 : node7401;
												assign node7401 = (inp[11]) ? node7407 : node7402;
													assign node7402 = (inp[5]) ? 16'b0000000011111111 : node7403;
														assign node7403 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7407 = (inp[14]) ? node7411 : node7408;
														assign node7408 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7411 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node7414 = (inp[4]) ? node7422 : node7415;
													assign node7415 = (inp[11]) ? node7419 : node7416;
														assign node7416 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node7419 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7422 = (inp[5]) ? node7426 : node7423;
														assign node7423 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7426 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node7429 = (inp[4]) ? node7487 : node7430;
										assign node7430 = (inp[7]) ? node7458 : node7431;
											assign node7431 = (inp[8]) ? node7445 : node7432;
												assign node7432 = (inp[11]) ? node7438 : node7433;
													assign node7433 = (inp[12]) ? node7435 : 16'b0000000111111111;
														assign node7435 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7438 = (inp[15]) ? node7442 : node7439;
														assign node7439 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7442 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7445 = (inp[11]) ? node7453 : node7446;
													assign node7446 = (inp[5]) ? node7450 : node7447;
														assign node7447 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7450 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7453 = (inp[15]) ? node7455 : 16'b0000000001111111;
														assign node7455 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7458 = (inp[15]) ? node7474 : node7459;
												assign node7459 = (inp[11]) ? node7467 : node7460;
													assign node7460 = (inp[12]) ? node7464 : node7461;
														assign node7461 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7464 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7467 = (inp[14]) ? node7471 : node7468;
														assign node7468 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7471 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7474 = (inp[5]) ? node7482 : node7475;
													assign node7475 = (inp[8]) ? node7479 : node7476;
														assign node7476 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7479 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7482 = (inp[12]) ? node7484 : 16'b0000000000111111;
														assign node7484 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node7487 = (inp[12]) ? node7519 : node7488;
											assign node7488 = (inp[8]) ? node7504 : node7489;
												assign node7489 = (inp[14]) ? node7497 : node7490;
													assign node7490 = (inp[15]) ? node7494 : node7491;
														assign node7491 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7494 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7497 = (inp[11]) ? node7501 : node7498;
														assign node7498 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7501 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node7504 = (inp[15]) ? node7512 : node7505;
													assign node7505 = (inp[5]) ? node7509 : node7506;
														assign node7506 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node7509 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7512 = (inp[14]) ? node7516 : node7513;
														assign node7513 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7516 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node7519 = (inp[8]) ? node7535 : node7520;
												assign node7520 = (inp[11]) ? node7528 : node7521;
													assign node7521 = (inp[5]) ? node7525 : node7522;
														assign node7522 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node7525 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7528 = (inp[5]) ? node7532 : node7529;
														assign node7529 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node7532 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node7535 = (inp[14]) ? node7543 : node7536;
													assign node7536 = (inp[15]) ? node7540 : node7537;
														assign node7537 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7540 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node7543 = (inp[5]) ? node7545 : 16'b0000000000011111;
														assign node7545 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node7548 = (inp[5]) ? node7668 : node7549;
									assign node7549 = (inp[14]) ? node7613 : node7550;
										assign node7550 = (inp[4]) ? node7582 : node7551;
											assign node7551 = (inp[15]) ? node7567 : node7552;
												assign node7552 = (inp[12]) ? node7560 : node7553;
													assign node7553 = (inp[11]) ? node7557 : node7554;
														assign node7554 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7557 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7560 = (inp[3]) ? node7564 : node7561;
														assign node7561 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7564 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node7567 = (inp[7]) ? node7575 : node7568;
													assign node7568 = (inp[8]) ? node7572 : node7569;
														assign node7569 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7572 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7575 = (inp[11]) ? node7579 : node7576;
														assign node7576 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node7579 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node7582 = (inp[7]) ? node7598 : node7583;
												assign node7583 = (inp[3]) ? node7591 : node7584;
													assign node7584 = (inp[12]) ? node7588 : node7585;
														assign node7585 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node7588 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node7591 = (inp[11]) ? node7595 : node7592;
														assign node7592 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node7595 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node7598 = (inp[12]) ? node7606 : node7599;
													assign node7599 = (inp[15]) ? node7603 : node7600;
														assign node7600 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7603 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node7606 = (inp[8]) ? node7610 : node7607;
														assign node7607 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node7610 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node7613 = (inp[12]) ? node7645 : node7614;
											assign node7614 = (inp[11]) ? node7630 : node7615;
												assign node7615 = (inp[3]) ? node7623 : node7616;
													assign node7616 = (inp[15]) ? node7620 : node7617;
														assign node7617 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node7620 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node7623 = (inp[7]) ? node7627 : node7624;
														assign node7624 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7627 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node7630 = (inp[15]) ? node7638 : node7631;
													assign node7631 = (inp[3]) ? node7635 : node7632;
														assign node7632 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7635 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7638 = (inp[4]) ? node7642 : node7639;
														assign node7639 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7642 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node7645 = (inp[4]) ? node7659 : node7646;
												assign node7646 = (inp[7]) ? node7652 : node7647;
													assign node7647 = (inp[11]) ? node7649 : 16'b0000000001111111;
														assign node7649 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7652 = (inp[11]) ? node7656 : node7653;
														assign node7653 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7656 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7659 = (inp[8]) ? node7665 : node7660;
													assign node7660 = (inp[15]) ? node7662 : 16'b0000000000111111;
														assign node7662 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
													assign node7665 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node7668 = (inp[11]) ? node7726 : node7669;
										assign node7669 = (inp[7]) ? node7697 : node7670;
											assign node7670 = (inp[4]) ? node7682 : node7671;
												assign node7671 = (inp[15]) ? node7675 : node7672;
													assign node7672 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node7675 = (inp[3]) ? node7679 : node7676;
														assign node7676 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7679 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node7682 = (inp[12]) ? node7690 : node7683;
													assign node7683 = (inp[15]) ? node7687 : node7684;
														assign node7684 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node7687 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7690 = (inp[8]) ? node7694 : node7691;
														assign node7691 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7694 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node7697 = (inp[4]) ? node7713 : node7698;
												assign node7698 = (inp[15]) ? node7706 : node7699;
													assign node7699 = (inp[14]) ? node7703 : node7700;
														assign node7700 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7703 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node7706 = (inp[3]) ? node7710 : node7707;
														assign node7707 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node7710 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node7713 = (inp[12]) ? node7719 : node7714;
													assign node7714 = (inp[3]) ? node7716 : 16'b0000000000111111;
														assign node7716 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node7719 = (inp[8]) ? node7723 : node7720;
														assign node7720 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node7723 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node7726 = (inp[7]) ? node7756 : node7727;
											assign node7727 = (inp[12]) ? node7743 : node7728;
												assign node7728 = (inp[15]) ? node7736 : node7729;
													assign node7729 = (inp[4]) ? node7733 : node7730;
														assign node7730 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node7733 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node7736 = (inp[14]) ? node7740 : node7737;
														assign node7737 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node7740 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node7743 = (inp[3]) ? node7751 : node7744;
													assign node7744 = (inp[4]) ? node7748 : node7745;
														assign node7745 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7748 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node7751 = (inp[15]) ? node7753 : 16'b0000000000011111;
														assign node7753 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node7756 = (inp[3]) ? node7772 : node7757;
												assign node7757 = (inp[4]) ? node7765 : node7758;
													assign node7758 = (inp[8]) ? node7762 : node7759;
														assign node7759 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node7762 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node7765 = (inp[8]) ? node7769 : node7766;
														assign node7766 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node7769 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node7772 = (inp[15]) ? node7778 : node7773;
													assign node7773 = (inp[14]) ? node7775 : 16'b0000000000111111;
														assign node7775 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node7778 = (inp[12]) ? node7782 : node7779;
														assign node7779 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node7782 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
			assign node7785 = (inp[10]) ? node11665 : node7786;
				assign node7786 = (inp[2]) ? node9724 : node7787;
					assign node7787 = (inp[15]) ? node8757 : node7788;
						assign node7788 = (inp[4]) ? node8272 : node7789;
							assign node7789 = (inp[13]) ? node8033 : node7790;
								assign node7790 = (inp[11]) ? node7918 : node7791;
									assign node7791 = (inp[3]) ? node7855 : node7792;
										assign node7792 = (inp[5]) ? node7824 : node7793;
											assign node7793 = (inp[14]) ? node7809 : node7794;
												assign node7794 = (inp[12]) ? node7802 : node7795;
													assign node7795 = (inp[9]) ? node7799 : node7796;
														assign node7796 = (inp[8]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node7799 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node7802 = (inp[7]) ? node7806 : node7803;
														assign node7803 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node7806 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node7809 = (inp[8]) ? node7817 : node7810;
													assign node7810 = (inp[9]) ? node7814 : node7811;
														assign node7811 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node7814 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7817 = (inp[7]) ? node7821 : node7818;
														assign node7818 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node7821 = (inp[0]) ? 16'b0000011111111111 : 16'b0000001111111111;
											assign node7824 = (inp[7]) ? node7840 : node7825;
												assign node7825 = (inp[9]) ? node7833 : node7826;
													assign node7826 = (inp[8]) ? node7830 : node7827;
														assign node7827 = (inp[12]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node7830 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7833 = (inp[0]) ? node7837 : node7834;
														assign node7834 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node7837 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7840 = (inp[0]) ? node7848 : node7841;
													assign node7841 = (inp[8]) ? node7845 : node7842;
														assign node7842 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node7845 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7848 = (inp[8]) ? node7852 : node7849;
														assign node7849 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7852 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node7855 = (inp[5]) ? node7887 : node7856;
											assign node7856 = (inp[0]) ? node7872 : node7857;
												assign node7857 = (inp[8]) ? node7865 : node7858;
													assign node7858 = (inp[14]) ? node7862 : node7859;
														assign node7859 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node7862 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7865 = (inp[14]) ? node7869 : node7866;
														assign node7866 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node7869 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7872 = (inp[12]) ? node7880 : node7873;
													assign node7873 = (inp[9]) ? node7877 : node7874;
														assign node7874 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node7877 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7880 = (inp[7]) ? node7884 : node7881;
														assign node7881 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7884 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7887 = (inp[9]) ? node7903 : node7888;
												assign node7888 = (inp[14]) ? node7896 : node7889;
													assign node7889 = (inp[8]) ? node7893 : node7890;
														assign node7890 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node7893 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7896 = (inp[7]) ? node7900 : node7897;
														assign node7897 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7900 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node7903 = (inp[7]) ? node7911 : node7904;
													assign node7904 = (inp[0]) ? node7908 : node7905;
														assign node7905 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7908 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7911 = (inp[14]) ? node7915 : node7912;
														assign node7912 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node7915 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node7918 = (inp[0]) ? node7976 : node7919;
										assign node7919 = (inp[12]) ? node7949 : node7920;
											assign node7920 = (inp[14]) ? node7936 : node7921;
												assign node7921 = (inp[9]) ? node7929 : node7922;
													assign node7922 = (inp[8]) ? node7926 : node7923;
														assign node7923 = (inp[5]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node7926 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7929 = (inp[5]) ? node7933 : node7930;
														assign node7930 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node7933 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7936 = (inp[3]) ? node7942 : node7937;
													assign node7937 = (inp[7]) ? 16'b0000011111111111 : node7938;
														assign node7938 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node7942 = (inp[9]) ? node7946 : node7943;
														assign node7943 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7946 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node7949 = (inp[5]) ? node7963 : node7950;
												assign node7950 = (inp[7]) ? node7956 : node7951;
													assign node7951 = (inp[14]) ? node7953 : 16'b0001111111111111;
														assign node7953 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node7956 = (inp[9]) ? node7960 : node7957;
														assign node7957 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7960 = (inp[14]) ? 16'b0000001111111111 : 16'b0000001111111111;
												assign node7963 = (inp[7]) ? node7971 : node7964;
													assign node7964 = (inp[3]) ? node7968 : node7965;
														assign node7965 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node7968 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7971 = (inp[14]) ? 16'b0000000111111111 : node7972;
														assign node7972 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node7976 = (inp[5]) ? node8006 : node7977;
											assign node7977 = (inp[9]) ? node7991 : node7978;
												assign node7978 = (inp[7]) ? node7986 : node7979;
													assign node7979 = (inp[14]) ? node7983 : node7980;
														assign node7980 = (inp[3]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node7983 = (inp[3]) ? 16'b0000011111111111 : 16'b0000001111111111;
													assign node7986 = (inp[14]) ? 16'b0000001111111111 : node7987;
														assign node7987 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node7991 = (inp[7]) ? node7999 : node7992;
													assign node7992 = (inp[14]) ? node7996 : node7993;
														assign node7993 = (inp[8]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node7996 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node7999 = (inp[14]) ? node8003 : node8000;
														assign node8000 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node8003 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8006 = (inp[8]) ? node8020 : node8007;
												assign node8007 = (inp[12]) ? node8015 : node8008;
													assign node8008 = (inp[14]) ? node8012 : node8009;
														assign node8009 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8012 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8015 = (inp[9]) ? node8017 : 16'b0000000111111111;
														assign node8017 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8020 = (inp[14]) ? node8026 : node8021;
													assign node8021 = (inp[3]) ? node8023 : 16'b0000001111111111;
														assign node8023 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8026 = (inp[12]) ? node8030 : node8027;
														assign node8027 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node8030 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
								assign node8033 = (inp[7]) ? node8153 : node8034;
									assign node8034 = (inp[9]) ? node8096 : node8035;
										assign node8035 = (inp[12]) ? node8067 : node8036;
											assign node8036 = (inp[3]) ? node8052 : node8037;
												assign node8037 = (inp[8]) ? node8045 : node8038;
													assign node8038 = (inp[5]) ? node8042 : node8039;
														assign node8039 = (inp[14]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node8042 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8045 = (inp[14]) ? node8049 : node8046;
														assign node8046 = (inp[11]) ? 16'b0000111111111111 : 16'b0000111111111111;
														assign node8049 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8052 = (inp[5]) ? node8060 : node8053;
													assign node8053 = (inp[14]) ? node8057 : node8054;
														assign node8054 = (inp[8]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node8057 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8060 = (inp[14]) ? node8064 : node8061;
														assign node8061 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8064 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node8067 = (inp[14]) ? node8081 : node8068;
												assign node8068 = (inp[8]) ? node8076 : node8069;
													assign node8069 = (inp[3]) ? node8073 : node8070;
														assign node8070 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8073 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8076 = (inp[3]) ? 16'b0000000111111111 : node8077;
														assign node8077 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8081 = (inp[0]) ? node8089 : node8082;
													assign node8082 = (inp[5]) ? node8086 : node8083;
														assign node8083 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8086 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node8089 = (inp[3]) ? node8093 : node8090;
														assign node8090 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8093 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node8096 = (inp[5]) ? node8126 : node8097;
											assign node8097 = (inp[14]) ? node8113 : node8098;
												assign node8098 = (inp[3]) ? node8106 : node8099;
													assign node8099 = (inp[11]) ? node8103 : node8100;
														assign node8100 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8103 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8106 = (inp[8]) ? node8110 : node8107;
														assign node8107 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8110 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8113 = (inp[0]) ? node8121 : node8114;
													assign node8114 = (inp[3]) ? node8118 : node8115;
														assign node8115 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8118 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node8121 = (inp[12]) ? node8123 : 16'b0000000111111111;
														assign node8123 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8126 = (inp[14]) ? node8140 : node8127;
												assign node8127 = (inp[0]) ? node8133 : node8128;
													assign node8128 = (inp[3]) ? 16'b0000001111111111 : node8129;
														assign node8129 = (inp[11]) ? 16'b0000001111111111 : 16'b0000001111111111;
													assign node8133 = (inp[12]) ? node8137 : node8134;
														assign node8134 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8137 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8140 = (inp[3]) ? node8146 : node8141;
													assign node8141 = (inp[11]) ? 16'b0000000011111111 : node8142;
														assign node8142 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8146 = (inp[12]) ? node8150 : node8147;
														assign node8147 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8150 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
									assign node8153 = (inp[8]) ? node8209 : node8154;
										assign node8154 = (inp[5]) ? node8184 : node8155;
											assign node8155 = (inp[0]) ? node8169 : node8156;
												assign node8156 = (inp[14]) ? node8162 : node8157;
													assign node8157 = (inp[3]) ? node8159 : 16'b0000011111111111;
														assign node8159 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8162 = (inp[3]) ? node8166 : node8163;
														assign node8163 = (inp[9]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node8166 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8169 = (inp[9]) ? node8177 : node8170;
													assign node8170 = (inp[12]) ? node8174 : node8171;
														assign node8171 = (inp[14]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node8174 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8177 = (inp[11]) ? node8181 : node8178;
														assign node8178 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8181 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8184 = (inp[3]) ? node8200 : node8185;
												assign node8185 = (inp[12]) ? node8193 : node8186;
													assign node8186 = (inp[0]) ? node8190 : node8187;
														assign node8187 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8190 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8193 = (inp[14]) ? node8197 : node8194;
														assign node8194 = (inp[9]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node8197 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8200 = (inp[11]) ? node8204 : node8201;
													assign node8201 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8204 = (inp[0]) ? node8206 : 16'b0000000111111111;
														assign node8206 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8209 = (inp[14]) ? node8241 : node8210;
											assign node8210 = (inp[11]) ? node8226 : node8211;
												assign node8211 = (inp[9]) ? node8219 : node8212;
													assign node8212 = (inp[0]) ? node8216 : node8213;
														assign node8213 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8216 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8219 = (inp[3]) ? node8223 : node8220;
														assign node8220 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node8223 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8226 = (inp[5]) ? node8234 : node8227;
													assign node8227 = (inp[3]) ? node8231 : node8228;
														assign node8228 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8231 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node8234 = (inp[3]) ? node8238 : node8235;
														assign node8235 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8238 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8241 = (inp[9]) ? node8257 : node8242;
												assign node8242 = (inp[3]) ? node8250 : node8243;
													assign node8243 = (inp[12]) ? node8247 : node8244;
														assign node8244 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8247 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8250 = (inp[5]) ? node8254 : node8251;
														assign node8251 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8254 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8257 = (inp[5]) ? node8265 : node8258;
													assign node8258 = (inp[3]) ? node8262 : node8259;
														assign node8259 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node8262 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8265 = (inp[3]) ? node8269 : node8266;
														assign node8266 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8269 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node8272 = (inp[0]) ? node8518 : node8273;
								assign node8273 = (inp[12]) ? node8399 : node8274;
									assign node8274 = (inp[9]) ? node8336 : node8275;
										assign node8275 = (inp[13]) ? node8305 : node8276;
											assign node8276 = (inp[5]) ? node8292 : node8277;
												assign node8277 = (inp[11]) ? node8285 : node8278;
													assign node8278 = (inp[7]) ? node8282 : node8279;
														assign node8279 = (inp[8]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node8282 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8285 = (inp[3]) ? node8289 : node8286;
														assign node8286 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8289 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8292 = (inp[14]) ? node8298 : node8293;
													assign node8293 = (inp[7]) ? node8295 : 16'b0000111111111111;
														assign node8295 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8298 = (inp[3]) ? node8302 : node8299;
														assign node8299 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8302 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node8305 = (inp[8]) ? node8321 : node8306;
												assign node8306 = (inp[5]) ? node8314 : node8307;
													assign node8307 = (inp[3]) ? node8311 : node8308;
														assign node8308 = (inp[14]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node8311 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8314 = (inp[11]) ? node8318 : node8315;
														assign node8315 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node8318 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8321 = (inp[5]) ? node8329 : node8322;
													assign node8322 = (inp[11]) ? node8326 : node8323;
														assign node8323 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8326 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8329 = (inp[11]) ? node8333 : node8330;
														assign node8330 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8333 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
										assign node8336 = (inp[7]) ? node8368 : node8337;
											assign node8337 = (inp[14]) ? node8353 : node8338;
												assign node8338 = (inp[3]) ? node8346 : node8339;
													assign node8339 = (inp[5]) ? node8343 : node8340;
														assign node8340 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8343 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8346 = (inp[8]) ? node8350 : node8347;
														assign node8347 = (inp[5]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node8350 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8353 = (inp[13]) ? node8361 : node8354;
													assign node8354 = (inp[5]) ? node8358 : node8355;
														assign node8355 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8358 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8361 = (inp[11]) ? node8365 : node8362;
														assign node8362 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8365 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8368 = (inp[14]) ? node8384 : node8369;
												assign node8369 = (inp[11]) ? node8377 : node8370;
													assign node8370 = (inp[13]) ? node8374 : node8371;
														assign node8371 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8374 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8377 = (inp[8]) ? node8381 : node8378;
														assign node8378 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8381 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node8384 = (inp[3]) ? node8392 : node8385;
													assign node8385 = (inp[8]) ? node8389 : node8386;
														assign node8386 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8389 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node8392 = (inp[13]) ? node8396 : node8393;
														assign node8393 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8396 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node8399 = (inp[3]) ? node8457 : node8400;
										assign node8400 = (inp[7]) ? node8428 : node8401;
											assign node8401 = (inp[14]) ? node8415 : node8402;
												assign node8402 = (inp[13]) ? node8408 : node8403;
													assign node8403 = (inp[8]) ? node8405 : 16'b0000011111111111;
														assign node8405 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8408 = (inp[11]) ? node8412 : node8409;
														assign node8409 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8412 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8415 = (inp[8]) ? node8423 : node8416;
													assign node8416 = (inp[5]) ? node8420 : node8417;
														assign node8417 = (inp[11]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node8420 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8423 = (inp[11]) ? 16'b0000000111111111 : node8424;
														assign node8424 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node8428 = (inp[13]) ? node8442 : node8429;
												assign node8429 = (inp[9]) ? node8437 : node8430;
													assign node8430 = (inp[14]) ? node8434 : node8431;
														assign node8431 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8434 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8437 = (inp[5]) ? node8439 : 16'b0000001111111111;
														assign node8439 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node8442 = (inp[11]) ? node8450 : node8443;
													assign node8443 = (inp[14]) ? node8447 : node8444;
														assign node8444 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node8447 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8450 = (inp[9]) ? node8454 : node8451;
														assign node8451 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8454 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node8457 = (inp[13]) ? node8489 : node8458;
											assign node8458 = (inp[8]) ? node8474 : node8459;
												assign node8459 = (inp[9]) ? node8467 : node8460;
													assign node8460 = (inp[11]) ? node8464 : node8461;
														assign node8461 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8464 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8467 = (inp[7]) ? node8471 : node8468;
														assign node8468 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8471 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8474 = (inp[11]) ? node8482 : node8475;
													assign node8475 = (inp[5]) ? node8479 : node8476;
														assign node8476 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8479 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8482 = (inp[9]) ? node8486 : node8483;
														assign node8483 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8486 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node8489 = (inp[14]) ? node8505 : node8490;
												assign node8490 = (inp[11]) ? node8498 : node8491;
													assign node8491 = (inp[8]) ? node8495 : node8492;
														assign node8492 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8495 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node8498 = (inp[7]) ? node8502 : node8499;
														assign node8499 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node8502 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node8505 = (inp[7]) ? node8511 : node8506;
													assign node8506 = (inp[5]) ? node8508 : 16'b0000000011111111;
														assign node8508 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8511 = (inp[9]) ? node8515 : node8512;
														assign node8512 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8515 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node8518 = (inp[7]) ? node8642 : node8519;
									assign node8519 = (inp[3]) ? node8583 : node8520;
										assign node8520 = (inp[5]) ? node8552 : node8521;
											assign node8521 = (inp[9]) ? node8537 : node8522;
												assign node8522 = (inp[8]) ? node8530 : node8523;
													assign node8523 = (inp[13]) ? node8527 : node8524;
														assign node8524 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8527 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8530 = (inp[14]) ? node8534 : node8531;
														assign node8531 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8534 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8537 = (inp[14]) ? node8545 : node8538;
													assign node8538 = (inp[11]) ? node8542 : node8539;
														assign node8539 = (inp[8]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node8542 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8545 = (inp[13]) ? node8549 : node8546;
														assign node8546 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8549 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8552 = (inp[11]) ? node8568 : node8553;
												assign node8553 = (inp[9]) ? node8561 : node8554;
													assign node8554 = (inp[14]) ? node8558 : node8555;
														assign node8555 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8558 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8561 = (inp[8]) ? node8565 : node8562;
														assign node8562 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8565 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8568 = (inp[13]) ? node8576 : node8569;
													assign node8569 = (inp[9]) ? node8573 : node8570;
														assign node8570 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node8573 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8576 = (inp[12]) ? node8580 : node8577;
														assign node8577 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8580 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8583 = (inp[8]) ? node8611 : node8584;
											assign node8584 = (inp[12]) ? node8598 : node8585;
												assign node8585 = (inp[13]) ? node8591 : node8586;
													assign node8586 = (inp[5]) ? node8588 : 16'b0000011111111111;
														assign node8588 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8591 = (inp[5]) ? node8595 : node8592;
														assign node8592 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8595 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8598 = (inp[5]) ? node8606 : node8599;
													assign node8599 = (inp[11]) ? node8603 : node8600;
														assign node8600 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8603 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8606 = (inp[11]) ? 16'b0000000001111111 : node8607;
														assign node8607 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node8611 = (inp[11]) ? node8627 : node8612;
												assign node8612 = (inp[13]) ? node8620 : node8613;
													assign node8613 = (inp[9]) ? node8617 : node8614;
														assign node8614 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8617 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8620 = (inp[14]) ? node8624 : node8621;
														assign node8621 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8624 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8627 = (inp[5]) ? node8635 : node8628;
													assign node8628 = (inp[14]) ? node8632 : node8629;
														assign node8629 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8632 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8635 = (inp[13]) ? node8639 : node8636;
														assign node8636 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8639 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node8642 = (inp[13]) ? node8704 : node8643;
										assign node8643 = (inp[9]) ? node8673 : node8644;
											assign node8644 = (inp[5]) ? node8660 : node8645;
												assign node8645 = (inp[3]) ? node8653 : node8646;
													assign node8646 = (inp[12]) ? node8650 : node8647;
														assign node8647 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8650 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node8653 = (inp[8]) ? node8657 : node8654;
														assign node8654 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8657 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8660 = (inp[14]) ? node8666 : node8661;
													assign node8661 = (inp[11]) ? 16'b0000000011111111 : node8662;
														assign node8662 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node8666 = (inp[3]) ? node8670 : node8667;
														assign node8667 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8670 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node8673 = (inp[3]) ? node8689 : node8674;
												assign node8674 = (inp[14]) ? node8682 : node8675;
													assign node8675 = (inp[12]) ? node8679 : node8676;
														assign node8676 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8679 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8682 = (inp[5]) ? node8686 : node8683;
														assign node8683 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8686 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8689 = (inp[12]) ? node8697 : node8690;
													assign node8690 = (inp[8]) ? node8694 : node8691;
														assign node8691 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node8694 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node8697 = (inp[14]) ? node8701 : node8698;
														assign node8698 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8701 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
										assign node8704 = (inp[11]) ? node8726 : node8705;
											assign node8705 = (inp[3]) ? node8719 : node8706;
												assign node8706 = (inp[8]) ? node8712 : node8707;
													assign node8707 = (inp[5]) ? node8709 : 16'b0000000111111111;
														assign node8709 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8712 = (inp[14]) ? node8716 : node8713;
														assign node8713 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node8716 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node8719 = (inp[8]) ? 16'b0000000001111111 : node8720;
													assign node8720 = (inp[14]) ? node8722 : 16'b0000000011111111;
														assign node8722 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node8726 = (inp[12]) ? node8742 : node8727;
												assign node8727 = (inp[8]) ? node8735 : node8728;
													assign node8728 = (inp[3]) ? node8732 : node8729;
														assign node8729 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node8732 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8735 = (inp[9]) ? node8739 : node8736;
														assign node8736 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8739 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node8742 = (inp[5]) ? node8750 : node8743;
													assign node8743 = (inp[3]) ? node8747 : node8744;
														assign node8744 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node8747 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node8750 = (inp[14]) ? node8754 : node8751;
														assign node8751 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node8754 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
						assign node8757 = (inp[7]) ? node9241 : node8758;
							assign node8758 = (inp[11]) ? node8998 : node8759;
								assign node8759 = (inp[9]) ? node8877 : node8760;
									assign node8760 = (inp[12]) ? node8820 : node8761;
										assign node8761 = (inp[4]) ? node8789 : node8762;
											assign node8762 = (inp[13]) ? node8776 : node8763;
												assign node8763 = (inp[14]) ? node8771 : node8764;
													assign node8764 = (inp[0]) ? node8768 : node8765;
														assign node8765 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node8768 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8771 = (inp[0]) ? 16'b0000011111111111 : node8772;
														assign node8772 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node8776 = (inp[8]) ? node8782 : node8777;
													assign node8777 = (inp[0]) ? 16'b0000001111111111 : node8778;
														assign node8778 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node8782 = (inp[3]) ? node8786 : node8783;
														assign node8783 = (inp[14]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node8786 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node8789 = (inp[14]) ? node8805 : node8790;
												assign node8790 = (inp[8]) ? node8798 : node8791;
													assign node8791 = (inp[0]) ? node8795 : node8792;
														assign node8792 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8795 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8798 = (inp[3]) ? node8802 : node8799;
														assign node8799 = (inp[13]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node8802 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8805 = (inp[0]) ? node8813 : node8806;
													assign node8806 = (inp[3]) ? node8810 : node8807;
														assign node8807 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8810 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node8813 = (inp[13]) ? node8817 : node8814;
														assign node8814 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8817 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node8820 = (inp[3]) ? node8848 : node8821;
											assign node8821 = (inp[8]) ? node8835 : node8822;
												assign node8822 = (inp[13]) ? node8830 : node8823;
													assign node8823 = (inp[14]) ? node8827 : node8824;
														assign node8824 = (inp[0]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node8827 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8830 = (inp[5]) ? 16'b0000001111111111 : node8831;
														assign node8831 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node8835 = (inp[0]) ? node8843 : node8836;
													assign node8836 = (inp[14]) ? node8840 : node8837;
														assign node8837 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8840 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8843 = (inp[13]) ? 16'b0000000011111111 : node8844;
														assign node8844 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
											assign node8848 = (inp[5]) ? node8864 : node8849;
												assign node8849 = (inp[13]) ? node8857 : node8850;
													assign node8850 = (inp[4]) ? node8854 : node8851;
														assign node8851 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8854 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8857 = (inp[0]) ? node8861 : node8858;
														assign node8858 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8861 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8864 = (inp[14]) ? node8870 : node8865;
													assign node8865 = (inp[8]) ? node8867 : 16'b0000001111111111;
														assign node8867 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8870 = (inp[0]) ? node8874 : node8871;
														assign node8871 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node8874 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node8877 = (inp[12]) ? node8939 : node8878;
										assign node8878 = (inp[0]) ? node8910 : node8879;
											assign node8879 = (inp[14]) ? node8895 : node8880;
												assign node8880 = (inp[13]) ? node8888 : node8881;
													assign node8881 = (inp[5]) ? node8885 : node8882;
														assign node8882 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node8885 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node8888 = (inp[8]) ? node8892 : node8889;
														assign node8889 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8892 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node8895 = (inp[3]) ? node8903 : node8896;
													assign node8896 = (inp[5]) ? node8900 : node8897;
														assign node8897 = (inp[8]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node8900 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8903 = (inp[13]) ? node8907 : node8904;
														assign node8904 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8907 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node8910 = (inp[3]) ? node8926 : node8911;
												assign node8911 = (inp[5]) ? node8919 : node8912;
													assign node8912 = (inp[14]) ? node8916 : node8913;
														assign node8913 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8916 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8919 = (inp[4]) ? node8923 : node8920;
														assign node8920 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8923 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8926 = (inp[13]) ? node8932 : node8927;
													assign node8927 = (inp[14]) ? node8929 : 16'b0000000111111111;
														assign node8929 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8932 = (inp[8]) ? node8936 : node8933;
														assign node8933 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node8936 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node8939 = (inp[14]) ? node8971 : node8940;
											assign node8940 = (inp[5]) ? node8956 : node8941;
												assign node8941 = (inp[4]) ? node8949 : node8942;
													assign node8942 = (inp[0]) ? node8946 : node8943;
														assign node8943 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node8946 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node8949 = (inp[3]) ? node8953 : node8950;
														assign node8950 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8953 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8956 = (inp[8]) ? node8964 : node8957;
													assign node8957 = (inp[13]) ? node8961 : node8958;
														assign node8958 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8961 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node8964 = (inp[0]) ? node8968 : node8965;
														assign node8965 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node8968 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node8971 = (inp[4]) ? node8985 : node8972;
												assign node8972 = (inp[13]) ? node8980 : node8973;
													assign node8973 = (inp[3]) ? node8977 : node8974;
														assign node8974 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node8977 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node8980 = (inp[8]) ? 16'b0000000011111111 : node8981;
														assign node8981 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node8985 = (inp[8]) ? node8991 : node8986;
													assign node8986 = (inp[13]) ? node8988 : 16'b0000000011111111;
														assign node8988 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node8991 = (inp[13]) ? node8995 : node8992;
														assign node8992 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node8995 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
								assign node8998 = (inp[13]) ? node9120 : node8999;
									assign node8999 = (inp[9]) ? node9059 : node9000;
										assign node9000 = (inp[14]) ? node9030 : node9001;
											assign node9001 = (inp[8]) ? node9017 : node9002;
												assign node9002 = (inp[4]) ? node9010 : node9003;
													assign node9003 = (inp[5]) ? node9007 : node9004;
														assign node9004 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9007 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9010 = (inp[3]) ? node9014 : node9011;
														assign node9011 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9014 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9017 = (inp[0]) ? node9023 : node9018;
													assign node9018 = (inp[5]) ? 16'b0000000111111111 : node9019;
														assign node9019 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9023 = (inp[4]) ? node9027 : node9024;
														assign node9024 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node9027 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node9030 = (inp[0]) ? node9044 : node9031;
												assign node9031 = (inp[4]) ? node9039 : node9032;
													assign node9032 = (inp[3]) ? node9036 : node9033;
														assign node9033 = (inp[5]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node9036 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node9039 = (inp[8]) ? node9041 : 16'b0000000111111111;
														assign node9041 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9044 = (inp[8]) ? node9052 : node9045;
													assign node9045 = (inp[3]) ? node9049 : node9046;
														assign node9046 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9049 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
													assign node9052 = (inp[3]) ? node9056 : node9053;
														assign node9053 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9056 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9059 = (inp[3]) ? node9091 : node9060;
											assign node9060 = (inp[5]) ? node9076 : node9061;
												assign node9061 = (inp[8]) ? node9069 : node9062;
													assign node9062 = (inp[4]) ? node9066 : node9063;
														assign node9063 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9066 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9069 = (inp[4]) ? node9073 : node9070;
														assign node9070 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node9073 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node9076 = (inp[0]) ? node9084 : node9077;
													assign node9077 = (inp[8]) ? node9081 : node9078;
														assign node9078 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node9081 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node9084 = (inp[12]) ? node9088 : node9085;
														assign node9085 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9088 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9091 = (inp[0]) ? node9105 : node9092;
												assign node9092 = (inp[4]) ? node9098 : node9093;
													assign node9093 = (inp[5]) ? 16'b0000000111111111 : node9094;
														assign node9094 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9098 = (inp[12]) ? node9102 : node9099;
														assign node9099 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9102 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node9105 = (inp[4]) ? node9113 : node9106;
													assign node9106 = (inp[14]) ? node9110 : node9107;
														assign node9107 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9110 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9113 = (inp[8]) ? node9117 : node9114;
														assign node9114 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9117 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node9120 = (inp[8]) ? node9182 : node9121;
										assign node9121 = (inp[14]) ? node9153 : node9122;
											assign node9122 = (inp[3]) ? node9138 : node9123;
												assign node9123 = (inp[12]) ? node9131 : node9124;
													assign node9124 = (inp[4]) ? node9128 : node9125;
														assign node9125 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9128 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9131 = (inp[4]) ? node9135 : node9132;
														assign node9132 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9135 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9138 = (inp[5]) ? node9146 : node9139;
													assign node9139 = (inp[0]) ? node9143 : node9140;
														assign node9140 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9143 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9146 = (inp[0]) ? node9150 : node9147;
														assign node9147 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9150 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9153 = (inp[0]) ? node9167 : node9154;
												assign node9154 = (inp[9]) ? node9160 : node9155;
													assign node9155 = (inp[5]) ? node9157 : 16'b0000001111111111;
														assign node9157 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9160 = (inp[12]) ? node9164 : node9161;
														assign node9161 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9164 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9167 = (inp[12]) ? node9175 : node9168;
													assign node9168 = (inp[3]) ? node9172 : node9169;
														assign node9169 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9172 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9175 = (inp[5]) ? node9179 : node9176;
														assign node9176 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9179 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node9182 = (inp[5]) ? node9212 : node9183;
											assign node9183 = (inp[0]) ? node9197 : node9184;
												assign node9184 = (inp[3]) ? node9190 : node9185;
													assign node9185 = (inp[12]) ? node9187 : 16'b0000000111111111;
														assign node9187 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9190 = (inp[4]) ? node9194 : node9191;
														assign node9191 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9194 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9197 = (inp[9]) ? node9205 : node9198;
													assign node9198 = (inp[12]) ? node9202 : node9199;
														assign node9199 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9202 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9205 = (inp[12]) ? node9209 : node9206;
														assign node9206 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9209 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9212 = (inp[3]) ? node9226 : node9213;
												assign node9213 = (inp[9]) ? node9221 : node9214;
													assign node9214 = (inp[0]) ? node9218 : node9215;
														assign node9215 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node9218 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9221 = (inp[0]) ? node9223 : 16'b0000000001111111;
														assign node9223 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node9226 = (inp[4]) ? node9234 : node9227;
													assign node9227 = (inp[0]) ? node9231 : node9228;
														assign node9228 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9231 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9234 = (inp[12]) ? node9238 : node9235;
														assign node9235 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node9238 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node9241 = (inp[3]) ? node9483 : node9242;
								assign node9242 = (inp[9]) ? node9362 : node9243;
									assign node9243 = (inp[0]) ? node9301 : node9244;
										assign node9244 = (inp[8]) ? node9270 : node9245;
											assign node9245 = (inp[13]) ? node9261 : node9246;
												assign node9246 = (inp[12]) ? node9254 : node9247;
													assign node9247 = (inp[11]) ? node9251 : node9248;
														assign node9248 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9251 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9254 = (inp[5]) ? node9258 : node9255;
														assign node9255 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node9258 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9261 = (inp[11]) ? 16'b0000000111111111 : node9262;
													assign node9262 = (inp[4]) ? node9266 : node9263;
														assign node9263 = (inp[12]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node9266 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9270 = (inp[4]) ? node9286 : node9271;
												assign node9271 = (inp[12]) ? node9279 : node9272;
													assign node9272 = (inp[11]) ? node9276 : node9273;
														assign node9273 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9276 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9279 = (inp[14]) ? node9283 : node9280;
														assign node9280 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9283 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9286 = (inp[13]) ? node9294 : node9287;
													assign node9287 = (inp[14]) ? node9291 : node9288;
														assign node9288 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9291 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9294 = (inp[14]) ? node9298 : node9295;
														assign node9295 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9298 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9301 = (inp[14]) ? node9331 : node9302;
											assign node9302 = (inp[5]) ? node9318 : node9303;
												assign node9303 = (inp[11]) ? node9311 : node9304;
													assign node9304 = (inp[13]) ? node9308 : node9305;
														assign node9305 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9308 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9311 = (inp[13]) ? node9315 : node9312;
														assign node9312 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9315 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node9318 = (inp[13]) ? node9326 : node9319;
													assign node9319 = (inp[12]) ? node9323 : node9320;
														assign node9320 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9323 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9326 = (inp[11]) ? 16'b0000000011111111 : node9327;
														assign node9327 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9331 = (inp[13]) ? node9347 : node9332;
												assign node9332 = (inp[12]) ? node9340 : node9333;
													assign node9333 = (inp[11]) ? node9337 : node9334;
														assign node9334 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9337 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node9340 = (inp[5]) ? node9344 : node9341;
														assign node9341 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9344 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9347 = (inp[5]) ? node9355 : node9348;
													assign node9348 = (inp[12]) ? node9352 : node9349;
														assign node9349 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9352 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node9355 = (inp[4]) ? node9359 : node9356;
														assign node9356 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9359 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node9362 = (inp[8]) ? node9420 : node9363;
										assign node9363 = (inp[12]) ? node9389 : node9364;
											assign node9364 = (inp[14]) ? node9376 : node9365;
												assign node9365 = (inp[13]) ? node9371 : node9366;
													assign node9366 = (inp[4]) ? 16'b0000001111111111 : node9367;
														assign node9367 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9371 = (inp[4]) ? node9373 : 16'b0000001111111111;
														assign node9373 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9376 = (inp[11]) ? node9384 : node9377;
													assign node9377 = (inp[13]) ? node9381 : node9378;
														assign node9378 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9381 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9384 = (inp[13]) ? 16'b0000000011111111 : node9385;
														assign node9385 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9389 = (inp[13]) ? node9405 : node9390;
												assign node9390 = (inp[14]) ? node9398 : node9391;
													assign node9391 = (inp[5]) ? node9395 : node9392;
														assign node9392 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9395 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9398 = (inp[0]) ? node9402 : node9399;
														assign node9399 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9402 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node9405 = (inp[11]) ? node9413 : node9406;
													assign node9406 = (inp[14]) ? node9410 : node9407;
														assign node9407 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9410 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9413 = (inp[4]) ? node9417 : node9414;
														assign node9414 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9417 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node9420 = (inp[5]) ? node9452 : node9421;
											assign node9421 = (inp[12]) ? node9437 : node9422;
												assign node9422 = (inp[4]) ? node9430 : node9423;
													assign node9423 = (inp[0]) ? node9427 : node9424;
														assign node9424 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9427 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9430 = (inp[11]) ? node9434 : node9431;
														assign node9431 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9434 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9437 = (inp[0]) ? node9445 : node9438;
													assign node9438 = (inp[4]) ? node9442 : node9439;
														assign node9439 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9442 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9445 = (inp[11]) ? node9449 : node9446;
														assign node9446 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9449 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9452 = (inp[4]) ? node9468 : node9453;
												assign node9453 = (inp[13]) ? node9461 : node9454;
													assign node9454 = (inp[11]) ? node9458 : node9455;
														assign node9455 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9458 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9461 = (inp[12]) ? node9465 : node9462;
														assign node9462 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9465 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9468 = (inp[11]) ? node9476 : node9469;
													assign node9469 = (inp[13]) ? node9473 : node9470;
														assign node9470 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9473 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9476 = (inp[0]) ? node9480 : node9477;
														assign node9477 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node9480 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000011111;
								assign node9483 = (inp[0]) ? node9605 : node9484;
									assign node9484 = (inp[13]) ? node9546 : node9485;
										assign node9485 = (inp[8]) ? node9515 : node9486;
											assign node9486 = (inp[5]) ? node9500 : node9487;
												assign node9487 = (inp[12]) ? node9495 : node9488;
													assign node9488 = (inp[14]) ? node9492 : node9489;
														assign node9489 = (inp[9]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node9492 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9495 = (inp[4]) ? node9497 : 16'b0000011111111111;
														assign node9497 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9500 = (inp[4]) ? node9508 : node9501;
													assign node9501 = (inp[12]) ? node9505 : node9502;
														assign node9502 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9505 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9508 = (inp[9]) ? node9512 : node9509;
														assign node9509 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9512 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9515 = (inp[12]) ? node9531 : node9516;
												assign node9516 = (inp[4]) ? node9524 : node9517;
													assign node9517 = (inp[14]) ? node9521 : node9518;
														assign node9518 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9521 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9524 = (inp[11]) ? node9528 : node9525;
														assign node9525 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9528 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9531 = (inp[14]) ? node9539 : node9532;
													assign node9532 = (inp[11]) ? node9536 : node9533;
														assign node9533 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9536 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9539 = (inp[9]) ? node9543 : node9540;
														assign node9540 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9543 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node9546 = (inp[5]) ? node9576 : node9547;
											assign node9547 = (inp[9]) ? node9561 : node9548;
												assign node9548 = (inp[12]) ? node9554 : node9549;
													assign node9549 = (inp[11]) ? node9551 : 16'b0000000111111111;
														assign node9551 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9554 = (inp[4]) ? node9558 : node9555;
														assign node9555 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9558 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9561 = (inp[11]) ? node9569 : node9562;
													assign node9562 = (inp[4]) ? node9566 : node9563;
														assign node9563 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9566 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9569 = (inp[8]) ? node9573 : node9570;
														assign node9570 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9573 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9576 = (inp[9]) ? node9592 : node9577;
												assign node9577 = (inp[14]) ? node9585 : node9578;
													assign node9578 = (inp[12]) ? node9582 : node9579;
														assign node9579 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9582 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9585 = (inp[8]) ? node9589 : node9586;
														assign node9586 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9589 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9592 = (inp[14]) ? node9598 : node9593;
													assign node9593 = (inp[11]) ? node9595 : 16'b0000000011111111;
														assign node9595 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9598 = (inp[12]) ? node9602 : node9599;
														assign node9599 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node9602 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node9605 = (inp[8]) ? node9665 : node9606;
										assign node9606 = (inp[13]) ? node9636 : node9607;
											assign node9607 = (inp[11]) ? node9621 : node9608;
												assign node9608 = (inp[4]) ? node9616 : node9609;
													assign node9609 = (inp[9]) ? node9613 : node9610;
														assign node9610 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node9613 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9616 = (inp[14]) ? 16'b0000000011111111 : node9617;
														assign node9617 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9621 = (inp[12]) ? node9629 : node9622;
													assign node9622 = (inp[4]) ? node9626 : node9623;
														assign node9623 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9626 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9629 = (inp[4]) ? node9633 : node9630;
														assign node9630 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9633 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9636 = (inp[11]) ? node9650 : node9637;
												assign node9637 = (inp[4]) ? node9645 : node9638;
													assign node9638 = (inp[9]) ? node9642 : node9639;
														assign node9639 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9642 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9645 = (inp[5]) ? node9647 : 16'b0000000011111111;
														assign node9647 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node9650 = (inp[5]) ? node9658 : node9651;
													assign node9651 = (inp[12]) ? node9655 : node9652;
														assign node9652 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9655 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9658 = (inp[14]) ? node9662 : node9659;
														assign node9659 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node9662 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node9665 = (inp[9]) ? node9695 : node9666;
											assign node9666 = (inp[5]) ? node9682 : node9667;
												assign node9667 = (inp[12]) ? node9675 : node9668;
													assign node9668 = (inp[11]) ? node9672 : node9669;
														assign node9669 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node9672 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node9675 = (inp[4]) ? node9679 : node9676;
														assign node9676 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node9679 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node9682 = (inp[11]) ? node9690 : node9683;
													assign node9683 = (inp[4]) ? node9687 : node9684;
														assign node9684 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node9687 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9690 = (inp[4]) ? 16'b0000000000111111 : node9691;
														assign node9691 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node9695 = (inp[12]) ? node9711 : node9696;
												assign node9696 = (inp[4]) ? node9704 : node9697;
													assign node9697 = (inp[13]) ? node9701 : node9698;
														assign node9698 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node9701 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node9704 = (inp[14]) ? node9708 : node9705;
														assign node9705 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node9708 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node9711 = (inp[11]) ? node9719 : node9712;
													assign node9712 = (inp[5]) ? node9716 : node9713;
														assign node9713 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node9716 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node9719 = (inp[4]) ? node9721 : 16'b0000000000011111;
														assign node9721 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node9724 = (inp[5]) ? node10698 : node9725;
						assign node9725 = (inp[7]) ? node10215 : node9726;
							assign node9726 = (inp[9]) ? node9968 : node9727;
								assign node9727 = (inp[11]) ? node9849 : node9728;
									assign node9728 = (inp[4]) ? node9788 : node9729;
										assign node9729 = (inp[14]) ? node9761 : node9730;
											assign node9730 = (inp[8]) ? node9746 : node9731;
												assign node9731 = (inp[0]) ? node9739 : node9732;
													assign node9732 = (inp[13]) ? node9736 : node9733;
														assign node9733 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node9736 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node9739 = (inp[3]) ? node9743 : node9740;
														assign node9740 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9743 = (inp[13]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node9746 = (inp[0]) ? node9754 : node9747;
													assign node9747 = (inp[15]) ? node9751 : node9748;
														assign node9748 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9751 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9754 = (inp[12]) ? node9758 : node9755;
														assign node9755 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9758 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node9761 = (inp[12]) ? node9777 : node9762;
												assign node9762 = (inp[3]) ? node9770 : node9763;
													assign node9763 = (inp[15]) ? node9767 : node9764;
														assign node9764 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9767 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9770 = (inp[13]) ? node9774 : node9771;
														assign node9771 = (inp[8]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node9774 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9777 = (inp[13]) ? node9783 : node9778;
													assign node9778 = (inp[0]) ? 16'b0000001111111111 : node9779;
														assign node9779 = (inp[8]) ? 16'b0000001111111111 : 16'b0000001111111111;
													assign node9783 = (inp[8]) ? 16'b0000000011111111 : node9784;
														assign node9784 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node9788 = (inp[13]) ? node9818 : node9789;
											assign node9789 = (inp[3]) ? node9803 : node9790;
												assign node9790 = (inp[15]) ? node9796 : node9791;
													assign node9791 = (inp[12]) ? 16'b0000011111111111 : node9792;
														assign node9792 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node9796 = (inp[8]) ? node9800 : node9797;
														assign node9797 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9800 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9803 = (inp[15]) ? node9811 : node9804;
													assign node9804 = (inp[14]) ? node9808 : node9805;
														assign node9805 = (inp[8]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node9808 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9811 = (inp[8]) ? node9815 : node9812;
														assign node9812 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node9815 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9818 = (inp[3]) ? node9834 : node9819;
												assign node9819 = (inp[14]) ? node9827 : node9820;
													assign node9820 = (inp[8]) ? node9824 : node9821;
														assign node9821 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9824 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9827 = (inp[0]) ? node9831 : node9828;
														assign node9828 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9831 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9834 = (inp[15]) ? node9842 : node9835;
													assign node9835 = (inp[12]) ? node9839 : node9836;
														assign node9836 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9839 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node9842 = (inp[0]) ? node9846 : node9843;
														assign node9843 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9846 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node9849 = (inp[0]) ? node9907 : node9850;
										assign node9850 = (inp[4]) ? node9880 : node9851;
											assign node9851 = (inp[13]) ? node9867 : node9852;
												assign node9852 = (inp[8]) ? node9860 : node9853;
													assign node9853 = (inp[12]) ? node9857 : node9854;
														assign node9854 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9857 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9860 = (inp[3]) ? node9864 : node9861;
														assign node9861 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9864 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node9867 = (inp[15]) ? node9873 : node9868;
													assign node9868 = (inp[12]) ? 16'b0000001111111111 : node9869;
														assign node9869 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9873 = (inp[3]) ? node9877 : node9874;
														assign node9874 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9877 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node9880 = (inp[14]) ? node9894 : node9881;
												assign node9881 = (inp[15]) ? node9887 : node9882;
													assign node9882 = (inp[13]) ? 16'b0000001111111111 : node9883;
														assign node9883 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9887 = (inp[12]) ? node9891 : node9888;
														assign node9888 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node9891 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node9894 = (inp[8]) ? node9902 : node9895;
													assign node9895 = (inp[3]) ? node9899 : node9896;
														assign node9896 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9899 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9902 = (inp[15]) ? node9904 : 16'b0000000011111111;
														assign node9904 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node9907 = (inp[15]) ? node9939 : node9908;
											assign node9908 = (inp[3]) ? node9924 : node9909;
												assign node9909 = (inp[8]) ? node9917 : node9910;
													assign node9910 = (inp[13]) ? node9914 : node9911;
														assign node9911 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9914 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9917 = (inp[14]) ? node9921 : node9918;
														assign node9918 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9921 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node9924 = (inp[12]) ? node9932 : node9925;
													assign node9925 = (inp[8]) ? node9929 : node9926;
														assign node9926 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9929 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node9932 = (inp[14]) ? node9936 : node9933;
														assign node9933 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node9936 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node9939 = (inp[8]) ? node9955 : node9940;
												assign node9940 = (inp[13]) ? node9948 : node9941;
													assign node9941 = (inp[14]) ? node9945 : node9942;
														assign node9942 = (inp[12]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node9945 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node9948 = (inp[12]) ? node9952 : node9949;
														assign node9949 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node9952 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node9955 = (inp[4]) ? node9963 : node9956;
													assign node9956 = (inp[12]) ? node9960 : node9957;
														assign node9957 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node9960 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node9963 = (inp[3]) ? 16'b0000000001111111 : node9964;
														assign node9964 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node9968 = (inp[8]) ? node10090 : node9969;
									assign node9969 = (inp[15]) ? node10031 : node9970;
										assign node9970 = (inp[0]) ? node10002 : node9971;
											assign node9971 = (inp[3]) ? node9987 : node9972;
												assign node9972 = (inp[12]) ? node9980 : node9973;
													assign node9973 = (inp[14]) ? node9977 : node9974;
														assign node9974 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node9977 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node9980 = (inp[11]) ? node9984 : node9981;
														assign node9981 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9984 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node9987 = (inp[4]) ? node9995 : node9988;
													assign node9988 = (inp[14]) ? node9992 : node9989;
														assign node9989 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node9992 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node9995 = (inp[11]) ? node9999 : node9996;
														assign node9996 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node9999 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10002 = (inp[12]) ? node10018 : node10003;
												assign node10003 = (inp[3]) ? node10011 : node10004;
													assign node10004 = (inp[14]) ? node10008 : node10005;
														assign node10005 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10008 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10011 = (inp[14]) ? node10015 : node10012;
														assign node10012 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10015 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10018 = (inp[14]) ? node10026 : node10019;
													assign node10019 = (inp[4]) ? node10023 : node10020;
														assign node10020 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node10023 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10026 = (inp[13]) ? node10028 : 16'b0000000011111111;
														assign node10028 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10031 = (inp[11]) ? node10061 : node10032;
											assign node10032 = (inp[14]) ? node10046 : node10033;
												assign node10033 = (inp[12]) ? node10039 : node10034;
													assign node10034 = (inp[4]) ? 16'b0000001111111111 : node10035;
														assign node10035 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10039 = (inp[3]) ? node10043 : node10040;
														assign node10040 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10043 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node10046 = (inp[12]) ? node10054 : node10047;
													assign node10047 = (inp[3]) ? node10051 : node10048;
														assign node10048 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10051 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10054 = (inp[13]) ? node10058 : node10055;
														assign node10055 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10058 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10061 = (inp[0]) ? node10077 : node10062;
												assign node10062 = (inp[12]) ? node10070 : node10063;
													assign node10063 = (inp[4]) ? node10067 : node10064;
														assign node10064 = (inp[13]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node10067 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node10070 = (inp[4]) ? node10074 : node10071;
														assign node10071 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10074 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10077 = (inp[3]) ? node10083 : node10078;
													assign node10078 = (inp[13]) ? node10080 : 16'b0000000011111111;
														assign node10080 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10083 = (inp[12]) ? node10087 : node10084;
														assign node10084 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node10087 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
									assign node10090 = (inp[4]) ? node10154 : node10091;
										assign node10091 = (inp[15]) ? node10123 : node10092;
											assign node10092 = (inp[3]) ? node10108 : node10093;
												assign node10093 = (inp[0]) ? node10101 : node10094;
													assign node10094 = (inp[11]) ? node10098 : node10095;
														assign node10095 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10098 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10101 = (inp[11]) ? node10105 : node10102;
														assign node10102 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node10105 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10108 = (inp[11]) ? node10116 : node10109;
													assign node10109 = (inp[13]) ? node10113 : node10110;
														assign node10110 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10113 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10116 = (inp[0]) ? node10120 : node10117;
														assign node10117 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10120 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10123 = (inp[12]) ? node10139 : node10124;
												assign node10124 = (inp[0]) ? node10132 : node10125;
													assign node10125 = (inp[3]) ? node10129 : node10126;
														assign node10126 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10129 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10132 = (inp[14]) ? node10136 : node10133;
														assign node10133 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10136 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10139 = (inp[0]) ? node10147 : node10140;
													assign node10140 = (inp[14]) ? node10144 : node10141;
														assign node10141 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10144 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node10147 = (inp[11]) ? node10151 : node10148;
														assign node10148 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10151 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node10154 = (inp[3]) ? node10184 : node10155;
											assign node10155 = (inp[11]) ? node10169 : node10156;
												assign node10156 = (inp[14]) ? node10162 : node10157;
													assign node10157 = (inp[12]) ? node10159 : 16'b0000001111111111;
														assign node10159 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node10162 = (inp[12]) ? node10166 : node10163;
														assign node10163 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10166 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10169 = (inp[12]) ? node10177 : node10170;
													assign node10170 = (inp[13]) ? node10174 : node10171;
														assign node10171 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10174 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10177 = (inp[13]) ? node10181 : node10178;
														assign node10178 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10181 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node10184 = (inp[15]) ? node10200 : node10185;
												assign node10185 = (inp[12]) ? node10193 : node10186;
													assign node10186 = (inp[11]) ? node10190 : node10187;
														assign node10187 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10190 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10193 = (inp[0]) ? node10197 : node10194;
														assign node10194 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10197 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10200 = (inp[14]) ? node10208 : node10201;
													assign node10201 = (inp[11]) ? node10205 : node10202;
														assign node10202 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node10205 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10208 = (inp[11]) ? node10212 : node10209;
														assign node10209 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node10212 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000011111;
							assign node10215 = (inp[11]) ? node10451 : node10216;
								assign node10216 = (inp[9]) ? node10332 : node10217;
									assign node10217 = (inp[0]) ? node10281 : node10218;
										assign node10218 = (inp[13]) ? node10250 : node10219;
											assign node10219 = (inp[8]) ? node10235 : node10220;
												assign node10220 = (inp[14]) ? node10228 : node10221;
													assign node10221 = (inp[4]) ? node10225 : node10222;
														assign node10222 = (inp[3]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node10225 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10228 = (inp[4]) ? node10232 : node10229;
														assign node10229 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10232 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10235 = (inp[3]) ? node10243 : node10236;
													assign node10236 = (inp[14]) ? node10240 : node10237;
														assign node10237 = (inp[12]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node10240 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10243 = (inp[12]) ? node10247 : node10244;
														assign node10244 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10247 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10250 = (inp[4]) ? node10266 : node10251;
												assign node10251 = (inp[3]) ? node10259 : node10252;
													assign node10252 = (inp[15]) ? node10256 : node10253;
														assign node10253 = (inp[12]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node10256 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10259 = (inp[15]) ? node10263 : node10260;
														assign node10260 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10263 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10266 = (inp[3]) ? node10274 : node10267;
													assign node10267 = (inp[15]) ? node10271 : node10268;
														assign node10268 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10271 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10274 = (inp[14]) ? node10278 : node10275;
														assign node10275 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10278 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
										assign node10281 = (inp[8]) ? node10309 : node10282;
											assign node10282 = (inp[13]) ? node10294 : node10283;
												assign node10283 = (inp[4]) ? node10291 : node10284;
													assign node10284 = (inp[12]) ? node10288 : node10285;
														assign node10285 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10288 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10291 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
												assign node10294 = (inp[14]) ? node10302 : node10295;
													assign node10295 = (inp[12]) ? node10299 : node10296;
														assign node10296 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10299 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10302 = (inp[15]) ? node10306 : node10303;
														assign node10303 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node10306 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10309 = (inp[4]) ? node10323 : node10310;
												assign node10310 = (inp[14]) ? node10316 : node10311;
													assign node10311 = (inp[13]) ? node10313 : 16'b0000001111111111;
														assign node10313 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10316 = (inp[13]) ? node10320 : node10317;
														assign node10317 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10320 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10323 = (inp[15]) ? 16'b0000000001111111 : node10324;
													assign node10324 = (inp[3]) ? node10328 : node10325;
														assign node10325 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10328 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
									assign node10332 = (inp[4]) ? node10392 : node10333;
										assign node10333 = (inp[12]) ? node10363 : node10334;
											assign node10334 = (inp[13]) ? node10350 : node10335;
												assign node10335 = (inp[15]) ? node10343 : node10336;
													assign node10336 = (inp[3]) ? node10340 : node10337;
														assign node10337 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10340 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node10343 = (inp[8]) ? node10347 : node10344;
														assign node10344 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node10347 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10350 = (inp[3]) ? node10356 : node10351;
													assign node10351 = (inp[14]) ? node10353 : 16'b0000001111111111;
														assign node10353 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10356 = (inp[0]) ? node10360 : node10357;
														assign node10357 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10360 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10363 = (inp[14]) ? node10377 : node10364;
												assign node10364 = (inp[15]) ? node10372 : node10365;
													assign node10365 = (inp[0]) ? node10369 : node10366;
														assign node10366 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node10369 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10372 = (inp[8]) ? 16'b0000000001111111 : node10373;
														assign node10373 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node10377 = (inp[15]) ? node10385 : node10378;
													assign node10378 = (inp[8]) ? node10382 : node10379;
														assign node10379 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10382 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node10385 = (inp[13]) ? node10389 : node10386;
														assign node10386 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10389 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node10392 = (inp[15]) ? node10422 : node10393;
											assign node10393 = (inp[8]) ? node10407 : node10394;
												assign node10394 = (inp[12]) ? node10400 : node10395;
													assign node10395 = (inp[13]) ? node10397 : 16'b0000001111111111;
														assign node10397 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10400 = (inp[14]) ? node10404 : node10401;
														assign node10401 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10404 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10407 = (inp[12]) ? node10415 : node10408;
													assign node10408 = (inp[13]) ? node10412 : node10409;
														assign node10409 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10412 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10415 = (inp[14]) ? node10419 : node10416;
														assign node10416 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node10419 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10422 = (inp[13]) ? node10436 : node10423;
												assign node10423 = (inp[3]) ? node10429 : node10424;
													assign node10424 = (inp[0]) ? 16'b0000000001111111 : node10425;
														assign node10425 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10429 = (inp[14]) ? node10433 : node10430;
														assign node10430 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10433 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10436 = (inp[8]) ? node10444 : node10437;
													assign node10437 = (inp[12]) ? node10441 : node10438;
														assign node10438 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node10441 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10444 = (inp[3]) ? node10448 : node10445;
														assign node10445 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10448 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node10451 = (inp[3]) ? node10575 : node10452;
									assign node10452 = (inp[12]) ? node10516 : node10453;
										assign node10453 = (inp[15]) ? node10485 : node10454;
											assign node10454 = (inp[14]) ? node10470 : node10455;
												assign node10455 = (inp[0]) ? node10463 : node10456;
													assign node10456 = (inp[8]) ? node10460 : node10457;
														assign node10457 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10460 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10463 = (inp[13]) ? node10467 : node10464;
														assign node10464 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10467 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10470 = (inp[4]) ? node10478 : node10471;
													assign node10471 = (inp[0]) ? node10475 : node10472;
														assign node10472 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10475 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node10478 = (inp[13]) ? node10482 : node10479;
														assign node10479 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node10482 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10485 = (inp[14]) ? node10501 : node10486;
												assign node10486 = (inp[13]) ? node10494 : node10487;
													assign node10487 = (inp[4]) ? node10491 : node10488;
														assign node10488 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10491 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10494 = (inp[9]) ? node10498 : node10495;
														assign node10495 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10498 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10501 = (inp[4]) ? node10509 : node10502;
													assign node10502 = (inp[9]) ? node10506 : node10503;
														assign node10503 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10506 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10509 = (inp[0]) ? node10513 : node10510;
														assign node10510 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10513 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10516 = (inp[13]) ? node10544 : node10517;
											assign node10517 = (inp[9]) ? node10531 : node10518;
												assign node10518 = (inp[15]) ? node10524 : node10519;
													assign node10519 = (inp[0]) ? 16'b0000000011111111 : node10520;
														assign node10520 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10524 = (inp[14]) ? node10528 : node10525;
														assign node10525 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10528 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10531 = (inp[0]) ? node10537 : node10532;
													assign node10532 = (inp[8]) ? node10534 : 16'b0000000011111111;
														assign node10534 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node10537 = (inp[14]) ? node10541 : node10538;
														assign node10538 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node10541 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node10544 = (inp[8]) ? node10560 : node10545;
												assign node10545 = (inp[0]) ? node10553 : node10546;
													assign node10546 = (inp[14]) ? node10550 : node10547;
														assign node10547 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10550 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10553 = (inp[9]) ? node10557 : node10554;
														assign node10554 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node10557 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10560 = (inp[9]) ? node10568 : node10561;
													assign node10561 = (inp[4]) ? node10565 : node10562;
														assign node10562 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10565 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node10568 = (inp[4]) ? node10572 : node10569;
														assign node10569 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10572 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node10575 = (inp[9]) ? node10639 : node10576;
										assign node10576 = (inp[15]) ? node10608 : node10577;
											assign node10577 = (inp[13]) ? node10593 : node10578;
												assign node10578 = (inp[4]) ? node10586 : node10579;
													assign node10579 = (inp[8]) ? node10583 : node10580;
														assign node10580 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node10583 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10586 = (inp[0]) ? node10590 : node10587;
														assign node10587 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node10590 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10593 = (inp[0]) ? node10601 : node10594;
													assign node10594 = (inp[12]) ? node10598 : node10595;
														assign node10595 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10598 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10601 = (inp[4]) ? node10605 : node10602;
														assign node10602 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10605 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10608 = (inp[12]) ? node10624 : node10609;
												assign node10609 = (inp[4]) ? node10617 : node10610;
													assign node10610 = (inp[14]) ? node10614 : node10611;
														assign node10611 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10614 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10617 = (inp[13]) ? node10621 : node10618;
														assign node10618 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node10621 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10624 = (inp[0]) ? node10632 : node10625;
													assign node10625 = (inp[14]) ? node10629 : node10626;
														assign node10626 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10629 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node10632 = (inp[14]) ? node10636 : node10633;
														assign node10633 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node10636 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node10639 = (inp[15]) ? node10669 : node10640;
											assign node10640 = (inp[8]) ? node10656 : node10641;
												assign node10641 = (inp[0]) ? node10649 : node10642;
													assign node10642 = (inp[14]) ? node10646 : node10643;
														assign node10643 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node10646 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10649 = (inp[12]) ? node10653 : node10650;
														assign node10650 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10653 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10656 = (inp[0]) ? node10664 : node10657;
													assign node10657 = (inp[4]) ? node10661 : node10658;
														assign node10658 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10661 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10664 = (inp[4]) ? node10666 : 16'b0000000000111111;
														assign node10666 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node10669 = (inp[13]) ? node10683 : node10670;
												assign node10670 = (inp[14]) ? node10676 : node10671;
													assign node10671 = (inp[0]) ? node10673 : 16'b0000000001111111;
														assign node10673 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10676 = (inp[4]) ? node10680 : node10677;
														assign node10677 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10680 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node10683 = (inp[12]) ? node10691 : node10684;
													assign node10684 = (inp[4]) ? node10688 : node10685;
														assign node10685 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node10688 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node10691 = (inp[14]) ? node10695 : node10692;
														assign node10692 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node10695 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node10698 = (inp[4]) ? node11184 : node10699;
							assign node10699 = (inp[14]) ? node10945 : node10700;
								assign node10700 = (inp[12]) ? node10822 : node10701;
									assign node10701 = (inp[7]) ? node10763 : node10702;
										assign node10702 = (inp[15]) ? node10734 : node10703;
											assign node10703 = (inp[0]) ? node10719 : node10704;
												assign node10704 = (inp[8]) ? node10712 : node10705;
													assign node10705 = (inp[11]) ? node10709 : node10706;
														assign node10706 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node10709 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10712 = (inp[9]) ? node10716 : node10713;
														assign node10713 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10716 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10719 = (inp[11]) ? node10727 : node10720;
													assign node10720 = (inp[9]) ? node10724 : node10721;
														assign node10721 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10724 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10727 = (inp[13]) ? node10731 : node10728;
														assign node10728 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10731 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node10734 = (inp[11]) ? node10750 : node10735;
												assign node10735 = (inp[13]) ? node10743 : node10736;
													assign node10736 = (inp[0]) ? node10740 : node10737;
														assign node10737 = (inp[9]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node10740 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node10743 = (inp[3]) ? node10747 : node10744;
														assign node10744 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10747 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10750 = (inp[0]) ? node10758 : node10751;
													assign node10751 = (inp[3]) ? node10755 : node10752;
														assign node10752 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10755 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node10758 = (inp[8]) ? 16'b0000000001111111 : node10759;
														assign node10759 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node10763 = (inp[11]) ? node10793 : node10764;
											assign node10764 = (inp[8]) ? node10778 : node10765;
												assign node10765 = (inp[15]) ? node10773 : node10766;
													assign node10766 = (inp[3]) ? node10770 : node10767;
														assign node10767 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10770 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node10773 = (inp[0]) ? 16'b0000000111111111 : node10774;
														assign node10774 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node10778 = (inp[13]) ? node10786 : node10779;
													assign node10779 = (inp[15]) ? node10783 : node10780;
														assign node10780 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10783 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node10786 = (inp[9]) ? node10790 : node10787;
														assign node10787 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10790 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10793 = (inp[13]) ? node10809 : node10794;
												assign node10794 = (inp[0]) ? node10802 : node10795;
													assign node10795 = (inp[9]) ? node10799 : node10796;
														assign node10796 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10799 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10802 = (inp[8]) ? node10806 : node10803;
														assign node10803 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node10806 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node10809 = (inp[9]) ? node10815 : node10810;
													assign node10810 = (inp[3]) ? node10812 : 16'b0000000011111111;
														assign node10812 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10815 = (inp[8]) ? node10819 : node10816;
														assign node10816 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node10819 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node10822 = (inp[0]) ? node10884 : node10823;
										assign node10823 = (inp[9]) ? node10853 : node10824;
											assign node10824 = (inp[11]) ? node10838 : node10825;
												assign node10825 = (inp[8]) ? node10831 : node10826;
													assign node10826 = (inp[13]) ? 16'b0000001111111111 : node10827;
														assign node10827 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node10831 = (inp[15]) ? node10835 : node10832;
														assign node10832 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10835 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node10838 = (inp[3]) ? node10846 : node10839;
													assign node10839 = (inp[13]) ? node10843 : node10840;
														assign node10840 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10843 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10846 = (inp[8]) ? node10850 : node10847;
														assign node10847 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10850 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10853 = (inp[13]) ? node10869 : node10854;
												assign node10854 = (inp[15]) ? node10862 : node10855;
													assign node10855 = (inp[8]) ? node10859 : node10856;
														assign node10856 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10859 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10862 = (inp[11]) ? node10866 : node10863;
														assign node10863 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10866 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node10869 = (inp[7]) ? node10877 : node10870;
													assign node10870 = (inp[3]) ? node10874 : node10871;
														assign node10871 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10874 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10877 = (inp[15]) ? node10881 : node10878;
														assign node10878 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10881 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node10884 = (inp[3]) ? node10914 : node10885;
											assign node10885 = (inp[11]) ? node10899 : node10886;
												assign node10886 = (inp[13]) ? node10894 : node10887;
													assign node10887 = (inp[9]) ? node10891 : node10888;
														assign node10888 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10891 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10894 = (inp[15]) ? 16'b0000000011111111 : node10895;
														assign node10895 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node10899 = (inp[8]) ? node10907 : node10900;
													assign node10900 = (inp[7]) ? node10904 : node10901;
														assign node10901 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10904 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10907 = (inp[15]) ? node10911 : node10908;
														assign node10908 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10911 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node10914 = (inp[13]) ? node10930 : node10915;
												assign node10915 = (inp[11]) ? node10923 : node10916;
													assign node10916 = (inp[15]) ? node10920 : node10917;
														assign node10917 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node10920 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node10923 = (inp[8]) ? node10927 : node10924;
														assign node10924 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10927 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node10930 = (inp[15]) ? node10938 : node10931;
													assign node10931 = (inp[11]) ? node10935 : node10932;
														assign node10932 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node10935 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node10938 = (inp[11]) ? node10942 : node10939;
														assign node10939 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node10942 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node10945 = (inp[7]) ? node11071 : node10946;
									assign node10946 = (inp[3]) ? node11008 : node10947;
										assign node10947 = (inp[0]) ? node10979 : node10948;
											assign node10948 = (inp[12]) ? node10964 : node10949;
												assign node10949 = (inp[11]) ? node10957 : node10950;
													assign node10950 = (inp[15]) ? node10954 : node10951;
														assign node10951 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node10954 = (inp[8]) ? 16'b0000001111111111 : 16'b0000001111111111;
													assign node10957 = (inp[15]) ? node10961 : node10958;
														assign node10958 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node10961 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node10964 = (inp[13]) ? node10972 : node10965;
													assign node10965 = (inp[8]) ? node10969 : node10966;
														assign node10966 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node10969 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10972 = (inp[15]) ? node10976 : node10973;
														assign node10973 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node10976 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node10979 = (inp[9]) ? node10995 : node10980;
												assign node10980 = (inp[13]) ? node10988 : node10981;
													assign node10981 = (inp[8]) ? node10985 : node10982;
														assign node10982 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node10985 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node10988 = (inp[11]) ? node10992 : node10989;
														assign node10989 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node10992 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node10995 = (inp[12]) ? node11001 : node10996;
													assign node10996 = (inp[15]) ? 16'b0000000011111111 : node10997;
														assign node10997 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11001 = (inp[15]) ? node11005 : node11002;
														assign node11002 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11005 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11008 = (inp[0]) ? node11040 : node11009;
											assign node11009 = (inp[8]) ? node11025 : node11010;
												assign node11010 = (inp[11]) ? node11018 : node11011;
													assign node11011 = (inp[12]) ? node11015 : node11012;
														assign node11012 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11015 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11018 = (inp[12]) ? node11022 : node11019;
														assign node11019 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11022 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11025 = (inp[11]) ? node11033 : node11026;
													assign node11026 = (inp[13]) ? node11030 : node11027;
														assign node11027 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node11030 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11033 = (inp[12]) ? node11037 : node11034;
														assign node11034 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11037 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11040 = (inp[9]) ? node11056 : node11041;
												assign node11041 = (inp[12]) ? node11049 : node11042;
													assign node11042 = (inp[11]) ? node11046 : node11043;
														assign node11043 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11046 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11049 = (inp[8]) ? node11053 : node11050;
														assign node11050 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11053 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11056 = (inp[15]) ? node11064 : node11057;
													assign node11057 = (inp[12]) ? node11061 : node11058;
														assign node11058 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11061 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11064 = (inp[11]) ? node11068 : node11065;
														assign node11065 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node11068 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node11071 = (inp[0]) ? node11129 : node11072;
										assign node11072 = (inp[8]) ? node11102 : node11073;
											assign node11073 = (inp[15]) ? node11087 : node11074;
												assign node11074 = (inp[9]) ? node11082 : node11075;
													assign node11075 = (inp[11]) ? node11079 : node11076;
														assign node11076 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11079 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11082 = (inp[11]) ? 16'b0000000011111111 : node11083;
														assign node11083 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11087 = (inp[13]) ? node11095 : node11088;
													assign node11088 = (inp[11]) ? node11092 : node11089;
														assign node11089 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11092 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11095 = (inp[12]) ? node11099 : node11096;
														assign node11096 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11099 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node11102 = (inp[9]) ? node11118 : node11103;
												assign node11103 = (inp[13]) ? node11111 : node11104;
													assign node11104 = (inp[12]) ? node11108 : node11105;
														assign node11105 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11108 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11111 = (inp[15]) ? node11115 : node11112;
														assign node11112 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11115 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node11118 = (inp[15]) ? node11126 : node11119;
													assign node11119 = (inp[11]) ? node11123 : node11120;
														assign node11120 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11123 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11126 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node11129 = (inp[11]) ? node11155 : node11130;
											assign node11130 = (inp[15]) ? node11142 : node11131;
												assign node11131 = (inp[9]) ? node11135 : node11132;
													assign node11132 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11135 = (inp[13]) ? node11139 : node11136;
														assign node11136 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11139 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node11142 = (inp[12]) ? node11150 : node11143;
													assign node11143 = (inp[13]) ? node11147 : node11144;
														assign node11144 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11147 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node11150 = (inp[3]) ? node11152 : 16'b0000000000111111;
														assign node11152 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node11155 = (inp[15]) ? node11171 : node11156;
												assign node11156 = (inp[3]) ? node11164 : node11157;
													assign node11157 = (inp[8]) ? node11161 : node11158;
														assign node11158 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node11161 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node11164 = (inp[13]) ? node11168 : node11165;
														assign node11165 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node11168 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11171 = (inp[8]) ? node11179 : node11172;
													assign node11172 = (inp[13]) ? node11176 : node11173;
														assign node11173 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node11176 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11179 = (inp[13]) ? node11181 : 16'b0000000000011111;
														assign node11181 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000011111;
							assign node11184 = (inp[15]) ? node11424 : node11185;
								assign node11185 = (inp[3]) ? node11305 : node11186;
									assign node11186 = (inp[9]) ? node11248 : node11187;
										assign node11187 = (inp[0]) ? node11217 : node11188;
											assign node11188 = (inp[12]) ? node11202 : node11189;
												assign node11189 = (inp[8]) ? node11197 : node11190;
													assign node11190 = (inp[7]) ? node11194 : node11191;
														assign node11191 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11194 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node11197 = (inp[14]) ? 16'b0000000111111111 : node11198;
														assign node11198 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11202 = (inp[7]) ? node11210 : node11203;
													assign node11203 = (inp[8]) ? node11207 : node11204;
														assign node11204 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11207 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11210 = (inp[14]) ? node11214 : node11211;
														assign node11211 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11214 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node11217 = (inp[8]) ? node11233 : node11218;
												assign node11218 = (inp[14]) ? node11226 : node11219;
													assign node11219 = (inp[13]) ? node11223 : node11220;
														assign node11220 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11223 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11226 = (inp[7]) ? node11230 : node11227;
														assign node11227 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11230 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11233 = (inp[11]) ? node11241 : node11234;
													assign node11234 = (inp[7]) ? node11238 : node11235;
														assign node11235 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node11238 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11241 = (inp[12]) ? node11245 : node11242;
														assign node11242 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11245 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11248 = (inp[13]) ? node11278 : node11249;
											assign node11249 = (inp[8]) ? node11265 : node11250;
												assign node11250 = (inp[0]) ? node11258 : node11251;
													assign node11251 = (inp[7]) ? node11255 : node11252;
														assign node11252 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11255 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11258 = (inp[11]) ? node11262 : node11259;
														assign node11259 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11262 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11265 = (inp[11]) ? node11273 : node11266;
													assign node11266 = (inp[7]) ? node11270 : node11267;
														assign node11267 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node11270 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11273 = (inp[7]) ? node11275 : 16'b0000000001111111;
														assign node11275 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node11278 = (inp[0]) ? node11292 : node11279;
												assign node11279 = (inp[11]) ? node11285 : node11280;
													assign node11280 = (inp[7]) ? node11282 : 16'b0000000011111111;
														assign node11282 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11285 = (inp[12]) ? node11289 : node11286;
														assign node11286 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11289 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11292 = (inp[14]) ? node11298 : node11293;
													assign node11293 = (inp[11]) ? node11295 : 16'b0000000001111111;
														assign node11295 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11298 = (inp[8]) ? node11302 : node11299;
														assign node11299 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11302 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node11305 = (inp[13]) ? node11363 : node11306;
										assign node11306 = (inp[14]) ? node11334 : node11307;
											assign node11307 = (inp[9]) ? node11323 : node11308;
												assign node11308 = (inp[11]) ? node11316 : node11309;
													assign node11309 = (inp[12]) ? node11313 : node11310;
														assign node11310 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11313 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11316 = (inp[7]) ? node11320 : node11317;
														assign node11317 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11320 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node11323 = (inp[0]) ? node11327 : node11324;
													assign node11324 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11327 = (inp[8]) ? node11331 : node11328;
														assign node11328 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node11331 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node11334 = (inp[12]) ? node11350 : node11335;
												assign node11335 = (inp[0]) ? node11343 : node11336;
													assign node11336 = (inp[9]) ? node11340 : node11337;
														assign node11337 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11340 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11343 = (inp[11]) ? node11347 : node11344;
														assign node11344 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11347 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node11350 = (inp[9]) ? node11358 : node11351;
													assign node11351 = (inp[7]) ? node11355 : node11352;
														assign node11352 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11355 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11358 = (inp[11]) ? 16'b0000000000111111 : node11359;
														assign node11359 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11363 = (inp[0]) ? node11395 : node11364;
											assign node11364 = (inp[12]) ? node11380 : node11365;
												assign node11365 = (inp[7]) ? node11373 : node11366;
													assign node11366 = (inp[8]) ? node11370 : node11367;
														assign node11367 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11370 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11373 = (inp[9]) ? node11377 : node11374;
														assign node11374 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11377 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11380 = (inp[9]) ? node11388 : node11381;
													assign node11381 = (inp[7]) ? node11385 : node11382;
														assign node11382 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node11385 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node11388 = (inp[14]) ? node11392 : node11389;
														assign node11389 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node11392 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node11395 = (inp[11]) ? node11409 : node11396;
												assign node11396 = (inp[8]) ? node11404 : node11397;
													assign node11397 = (inp[12]) ? node11401 : node11398;
														assign node11398 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11401 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11404 = (inp[7]) ? 16'b0000000000111111 : node11405;
														assign node11405 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11409 = (inp[14]) ? node11417 : node11410;
													assign node11410 = (inp[12]) ? node11414 : node11411;
														assign node11411 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node11414 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11417 = (inp[8]) ? node11421 : node11418;
														assign node11418 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node11421 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node11424 = (inp[14]) ? node11542 : node11425;
									assign node11425 = (inp[3]) ? node11481 : node11426;
										assign node11426 = (inp[12]) ? node11456 : node11427;
											assign node11427 = (inp[7]) ? node11441 : node11428;
												assign node11428 = (inp[0]) ? node11434 : node11429;
													assign node11429 = (inp[8]) ? 16'b0000000111111111 : node11430;
														assign node11430 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11434 = (inp[8]) ? node11438 : node11435;
														assign node11435 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node11438 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11441 = (inp[8]) ? node11449 : node11442;
													assign node11442 = (inp[13]) ? node11446 : node11443;
														assign node11443 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11446 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node11449 = (inp[0]) ? node11453 : node11450;
														assign node11450 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11453 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node11456 = (inp[0]) ? node11472 : node11457;
												assign node11457 = (inp[9]) ? node11465 : node11458;
													assign node11458 = (inp[8]) ? node11462 : node11459;
														assign node11459 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node11462 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11465 = (inp[7]) ? node11469 : node11466;
														assign node11466 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11469 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11472 = (inp[13]) ? node11476 : node11473;
													assign node11473 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11476 = (inp[9]) ? 16'b0000000000111111 : node11477;
														assign node11477 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node11481 = (inp[13]) ? node11513 : node11482;
											assign node11482 = (inp[0]) ? node11498 : node11483;
												assign node11483 = (inp[11]) ? node11491 : node11484;
													assign node11484 = (inp[8]) ? node11488 : node11485;
														assign node11485 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11488 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11491 = (inp[7]) ? node11495 : node11492;
														assign node11492 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11495 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node11498 = (inp[9]) ? node11506 : node11499;
													assign node11499 = (inp[12]) ? node11503 : node11500;
														assign node11500 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11503 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11506 = (inp[7]) ? node11510 : node11507;
														assign node11507 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11510 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node11513 = (inp[8]) ? node11527 : node11514;
												assign node11514 = (inp[0]) ? node11522 : node11515;
													assign node11515 = (inp[7]) ? node11519 : node11516;
														assign node11516 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11519 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11522 = (inp[9]) ? node11524 : 16'b0000000011111111;
														assign node11524 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11527 = (inp[7]) ? node11535 : node11528;
													assign node11528 = (inp[9]) ? node11532 : node11529;
														assign node11529 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11532 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node11535 = (inp[0]) ? node11539 : node11536;
														assign node11536 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node11539 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000001111;
									assign node11542 = (inp[9]) ? node11602 : node11543;
										assign node11543 = (inp[8]) ? node11575 : node11544;
											assign node11544 = (inp[13]) ? node11560 : node11545;
												assign node11545 = (inp[3]) ? node11553 : node11546;
													assign node11546 = (inp[0]) ? node11550 : node11547;
														assign node11547 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11550 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node11553 = (inp[11]) ? node11557 : node11554;
														assign node11554 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11557 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11560 = (inp[12]) ? node11568 : node11561;
													assign node11561 = (inp[3]) ? node11565 : node11562;
														assign node11562 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11565 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node11568 = (inp[0]) ? node11572 : node11569;
														assign node11569 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11572 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node11575 = (inp[7]) ? node11587 : node11576;
												assign node11576 = (inp[3]) ? node11582 : node11577;
													assign node11577 = (inp[0]) ? 16'b0000000001111111 : node11578;
														assign node11578 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node11582 = (inp[12]) ? 16'b0000000000011111 : node11583;
														assign node11583 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node11587 = (inp[13]) ? node11595 : node11588;
													assign node11588 = (inp[11]) ? node11592 : node11589;
														assign node11589 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11592 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11595 = (inp[3]) ? node11599 : node11596;
														assign node11596 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node11599 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node11602 = (inp[7]) ? node11634 : node11603;
											assign node11603 = (inp[8]) ? node11619 : node11604;
												assign node11604 = (inp[12]) ? node11612 : node11605;
													assign node11605 = (inp[3]) ? node11609 : node11606;
														assign node11606 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11609 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node11612 = (inp[13]) ? node11616 : node11613;
														assign node11613 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node11616 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node11619 = (inp[3]) ? node11627 : node11620;
													assign node11620 = (inp[0]) ? node11624 : node11621;
														assign node11621 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node11624 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11627 = (inp[11]) ? node11631 : node11628;
														assign node11628 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node11631 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node11634 = (inp[13]) ? node11650 : node11635;
												assign node11635 = (inp[12]) ? node11643 : node11636;
													assign node11636 = (inp[0]) ? node11640 : node11637;
														assign node11637 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node11640 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node11643 = (inp[3]) ? node11647 : node11644;
														assign node11644 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node11647 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node11650 = (inp[12]) ? node11658 : node11651;
													assign node11651 = (inp[8]) ? node11655 : node11652;
														assign node11652 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node11655 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node11658 = (inp[0]) ? node11662 : node11659;
														assign node11659 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node11662 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
				assign node11665 = (inp[5]) ? node13595 : node11666;
					assign node11666 = (inp[4]) ? node12630 : node11667;
						assign node11667 = (inp[11]) ? node12157 : node11668;
							assign node11668 = (inp[2]) ? node11918 : node11669;
								assign node11669 = (inp[0]) ? node11793 : node11670;
									assign node11670 = (inp[9]) ? node11732 : node11671;
										assign node11671 = (inp[13]) ? node11701 : node11672;
											assign node11672 = (inp[8]) ? node11686 : node11673;
												assign node11673 = (inp[14]) ? node11679 : node11674;
													assign node11674 = (inp[12]) ? 16'b0000111111111111 : node11675;
														assign node11675 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node11679 = (inp[7]) ? node11683 : node11680;
														assign node11680 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node11683 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node11686 = (inp[14]) ? node11694 : node11687;
													assign node11687 = (inp[15]) ? node11691 : node11688;
														assign node11688 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node11691 = (inp[3]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node11694 = (inp[7]) ? node11698 : node11695;
														assign node11695 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11698 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node11701 = (inp[12]) ? node11717 : node11702;
												assign node11702 = (inp[15]) ? node11710 : node11703;
													assign node11703 = (inp[7]) ? node11707 : node11704;
														assign node11704 = (inp[14]) ? 16'b0000011111111111 : 16'b0001111111111111;
														assign node11707 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node11710 = (inp[7]) ? node11714 : node11711;
														assign node11711 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11714 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11717 = (inp[8]) ? node11725 : node11718;
													assign node11718 = (inp[3]) ? node11722 : node11719;
														assign node11719 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11722 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11725 = (inp[14]) ? node11729 : node11726;
														assign node11726 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node11729 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000011111111;
										assign node11732 = (inp[14]) ? node11762 : node11733;
											assign node11733 = (inp[13]) ? node11749 : node11734;
												assign node11734 = (inp[15]) ? node11742 : node11735;
													assign node11735 = (inp[12]) ? node11739 : node11736;
														assign node11736 = (inp[7]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node11739 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node11742 = (inp[7]) ? node11746 : node11743;
														assign node11743 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11746 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node11749 = (inp[15]) ? node11755 : node11750;
													assign node11750 = (inp[3]) ? node11752 : 16'b0000001111111111;
														assign node11752 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11755 = (inp[12]) ? node11759 : node11756;
														assign node11756 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11759 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11762 = (inp[15]) ? node11778 : node11763;
												assign node11763 = (inp[3]) ? node11771 : node11764;
													assign node11764 = (inp[7]) ? node11768 : node11765;
														assign node11765 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11768 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11771 = (inp[13]) ? node11775 : node11772;
														assign node11772 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11775 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node11778 = (inp[3]) ? node11786 : node11779;
													assign node11779 = (inp[7]) ? node11783 : node11780;
														assign node11780 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11783 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11786 = (inp[13]) ? node11790 : node11787;
														assign node11787 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11790 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node11793 = (inp[3]) ? node11857 : node11794;
										assign node11794 = (inp[9]) ? node11826 : node11795;
											assign node11795 = (inp[14]) ? node11811 : node11796;
												assign node11796 = (inp[8]) ? node11804 : node11797;
													assign node11797 = (inp[7]) ? node11801 : node11798;
														assign node11798 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node11801 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node11804 = (inp[7]) ? node11808 : node11805;
														assign node11805 = (inp[12]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node11808 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node11811 = (inp[13]) ? node11819 : node11812;
													assign node11812 = (inp[7]) ? node11816 : node11813;
														assign node11813 = (inp[12]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node11816 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11819 = (inp[7]) ? node11823 : node11820;
														assign node11820 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node11823 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
											assign node11826 = (inp[12]) ? node11842 : node11827;
												assign node11827 = (inp[15]) ? node11835 : node11828;
													assign node11828 = (inp[7]) ? node11832 : node11829;
														assign node11829 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11832 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node11835 = (inp[14]) ? node11839 : node11836;
														assign node11836 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11839 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11842 = (inp[15]) ? node11850 : node11843;
													assign node11843 = (inp[14]) ? node11847 : node11844;
														assign node11844 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11847 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11850 = (inp[14]) ? node11854 : node11851;
														assign node11851 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node11854 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node11857 = (inp[12]) ? node11887 : node11858;
											assign node11858 = (inp[8]) ? node11874 : node11859;
												assign node11859 = (inp[14]) ? node11867 : node11860;
													assign node11860 = (inp[9]) ? node11864 : node11861;
														assign node11861 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11864 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11867 = (inp[9]) ? node11871 : node11868;
														assign node11868 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node11871 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11874 = (inp[7]) ? node11880 : node11875;
													assign node11875 = (inp[14]) ? 16'b0000000111111111 : node11876;
														assign node11876 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11880 = (inp[14]) ? node11884 : node11881;
														assign node11881 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node11884 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node11887 = (inp[13]) ? node11903 : node11888;
												assign node11888 = (inp[9]) ? node11896 : node11889;
													assign node11889 = (inp[15]) ? node11893 : node11890;
														assign node11890 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node11893 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11896 = (inp[7]) ? node11900 : node11897;
														assign node11897 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node11900 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node11903 = (inp[9]) ? node11911 : node11904;
													assign node11904 = (inp[14]) ? node11908 : node11905;
														assign node11905 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node11908 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node11911 = (inp[15]) ? node11915 : node11912;
														assign node11912 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node11915 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node11918 = (inp[12]) ? node12038 : node11919;
									assign node11919 = (inp[0]) ? node11979 : node11920;
										assign node11920 = (inp[8]) ? node11948 : node11921;
											assign node11921 = (inp[15]) ? node11935 : node11922;
												assign node11922 = (inp[9]) ? node11930 : node11923;
													assign node11923 = (inp[3]) ? node11927 : node11924;
														assign node11924 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node11927 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node11930 = (inp[13]) ? 16'b0000000111111111 : node11931;
														assign node11931 = (inp[14]) ? 16'b0000011111111111 : 16'b0000001111111111;
												assign node11935 = (inp[14]) ? node11941 : node11936;
													assign node11936 = (inp[7]) ? node11938 : 16'b0000011111111111;
														assign node11938 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11941 = (inp[13]) ? node11945 : node11942;
														assign node11942 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11945 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node11948 = (inp[3]) ? node11964 : node11949;
												assign node11949 = (inp[9]) ? node11957 : node11950;
													assign node11950 = (inp[14]) ? node11954 : node11951;
														assign node11951 = (inp[15]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node11954 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11957 = (inp[7]) ? node11961 : node11958;
														assign node11958 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11961 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11964 = (inp[14]) ? node11972 : node11965;
													assign node11965 = (inp[9]) ? node11969 : node11966;
														assign node11966 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node11969 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node11972 = (inp[7]) ? node11976 : node11973;
														assign node11973 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node11976 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node11979 = (inp[8]) ? node12011 : node11980;
											assign node11980 = (inp[13]) ? node11996 : node11981;
												assign node11981 = (inp[3]) ? node11989 : node11982;
													assign node11982 = (inp[14]) ? node11986 : node11983;
														assign node11983 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node11986 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node11989 = (inp[9]) ? node11993 : node11990;
														assign node11990 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node11993 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node11996 = (inp[15]) ? node12004 : node11997;
													assign node11997 = (inp[14]) ? node12001 : node11998;
														assign node11998 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12001 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12004 = (inp[7]) ? node12008 : node12005;
														assign node12005 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12008 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node12011 = (inp[15]) ? node12027 : node12012;
												assign node12012 = (inp[7]) ? node12020 : node12013;
													assign node12013 = (inp[9]) ? node12017 : node12014;
														assign node12014 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12017 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12020 = (inp[13]) ? node12024 : node12021;
														assign node12021 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12024 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node12027 = (inp[7]) ? node12033 : node12028;
													assign node12028 = (inp[14]) ? node12030 : 16'b0000000111111111;
														assign node12030 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12033 = (inp[9]) ? node12035 : 16'b0000000001111111;
														assign node12035 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
									assign node12038 = (inp[7]) ? node12098 : node12039;
										assign node12039 = (inp[9]) ? node12067 : node12040;
											assign node12040 = (inp[3]) ? node12052 : node12041;
												assign node12041 = (inp[8]) ? node12049 : node12042;
													assign node12042 = (inp[14]) ? node12046 : node12043;
														assign node12043 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12046 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12049 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12052 = (inp[15]) ? node12060 : node12053;
													assign node12053 = (inp[13]) ? node12057 : node12054;
														assign node12054 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12057 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12060 = (inp[8]) ? node12064 : node12061;
														assign node12061 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12064 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node12067 = (inp[14]) ? node12083 : node12068;
												assign node12068 = (inp[13]) ? node12076 : node12069;
													assign node12069 = (inp[3]) ? node12073 : node12070;
														assign node12070 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12073 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12076 = (inp[0]) ? node12080 : node12077;
														assign node12077 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12080 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12083 = (inp[13]) ? node12091 : node12084;
													assign node12084 = (inp[3]) ? node12088 : node12085;
														assign node12085 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12088 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12091 = (inp[8]) ? node12095 : node12092;
														assign node12092 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12095 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node12098 = (inp[15]) ? node12126 : node12099;
											assign node12099 = (inp[8]) ? node12113 : node12100;
												assign node12100 = (inp[0]) ? node12106 : node12101;
													assign node12101 = (inp[3]) ? node12103 : 16'b0000001111111111;
														assign node12103 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node12106 = (inp[13]) ? node12110 : node12107;
														assign node12107 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12110 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12113 = (inp[0]) ? node12121 : node12114;
													assign node12114 = (inp[13]) ? node12118 : node12115;
														assign node12115 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12118 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node12121 = (inp[3]) ? node12123 : 16'b0000000011111111;
														assign node12123 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node12126 = (inp[3]) ? node12142 : node12127;
												assign node12127 = (inp[14]) ? node12135 : node12128;
													assign node12128 = (inp[9]) ? node12132 : node12129;
														assign node12129 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12132 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12135 = (inp[9]) ? node12139 : node12136;
														assign node12136 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node12139 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12142 = (inp[9]) ? node12150 : node12143;
													assign node12143 = (inp[13]) ? node12147 : node12144;
														assign node12144 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12147 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12150 = (inp[8]) ? node12154 : node12151;
														assign node12151 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12154 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node12157 = (inp[15]) ? node12393 : node12158;
								assign node12158 = (inp[13]) ? node12278 : node12159;
									assign node12159 = (inp[7]) ? node12219 : node12160;
										assign node12160 = (inp[8]) ? node12192 : node12161;
											assign node12161 = (inp[0]) ? node12177 : node12162;
												assign node12162 = (inp[9]) ? node12170 : node12163;
													assign node12163 = (inp[14]) ? node12167 : node12164;
														assign node12164 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node12167 = (inp[12]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node12170 = (inp[2]) ? node12174 : node12171;
														assign node12171 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12174 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12177 = (inp[2]) ? node12185 : node12178;
													assign node12178 = (inp[3]) ? node12182 : node12179;
														assign node12179 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12182 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node12185 = (inp[12]) ? node12189 : node12186;
														assign node12186 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12189 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node12192 = (inp[3]) ? node12206 : node12193;
												assign node12193 = (inp[14]) ? node12201 : node12194;
													assign node12194 = (inp[0]) ? node12198 : node12195;
														assign node12195 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12198 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12201 = (inp[12]) ? 16'b0000000111111111 : node12202;
														assign node12202 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12206 = (inp[0]) ? node12212 : node12207;
													assign node12207 = (inp[9]) ? 16'b0000000111111111 : node12208;
														assign node12208 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12212 = (inp[12]) ? node12216 : node12213;
														assign node12213 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node12216 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
										assign node12219 = (inp[14]) ? node12249 : node12220;
											assign node12220 = (inp[12]) ? node12234 : node12221;
												assign node12221 = (inp[9]) ? node12227 : node12222;
													assign node12222 = (inp[0]) ? node12224 : 16'b0000011111111111;
														assign node12224 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12227 = (inp[2]) ? node12231 : node12228;
														assign node12228 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12231 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12234 = (inp[9]) ? node12242 : node12235;
													assign node12235 = (inp[3]) ? node12239 : node12236;
														assign node12236 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12239 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12242 = (inp[8]) ? node12246 : node12243;
														assign node12243 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node12246 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node12249 = (inp[3]) ? node12263 : node12250;
												assign node12250 = (inp[9]) ? node12258 : node12251;
													assign node12251 = (inp[2]) ? node12255 : node12252;
														assign node12252 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12255 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12258 = (inp[8]) ? 16'b0000000011111111 : node12259;
														assign node12259 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node12263 = (inp[0]) ? node12271 : node12264;
													assign node12264 = (inp[8]) ? node12268 : node12265;
														assign node12265 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12268 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12271 = (inp[9]) ? node12275 : node12272;
														assign node12272 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12275 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node12278 = (inp[3]) ? node12334 : node12279;
										assign node12279 = (inp[8]) ? node12305 : node12280;
											assign node12280 = (inp[0]) ? node12290 : node12281;
												assign node12281 = (inp[7]) ? 16'b0000000111111111 : node12282;
													assign node12282 = (inp[2]) ? node12286 : node12283;
														assign node12283 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12286 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12290 = (inp[12]) ? node12298 : node12291;
													assign node12291 = (inp[2]) ? node12295 : node12292;
														assign node12292 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12295 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12298 = (inp[2]) ? node12302 : node12299;
														assign node12299 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12302 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node12305 = (inp[12]) ? node12321 : node12306;
												assign node12306 = (inp[14]) ? node12314 : node12307;
													assign node12307 = (inp[7]) ? node12311 : node12308;
														assign node12308 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12311 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12314 = (inp[9]) ? node12318 : node12315;
														assign node12315 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12318 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12321 = (inp[2]) ? node12329 : node12322;
													assign node12322 = (inp[7]) ? node12326 : node12323;
														assign node12323 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12326 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12329 = (inp[0]) ? node12331 : 16'b0000000001111111;
														assign node12331 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node12334 = (inp[14]) ? node12366 : node12335;
											assign node12335 = (inp[8]) ? node12351 : node12336;
												assign node12336 = (inp[12]) ? node12344 : node12337;
													assign node12337 = (inp[9]) ? node12341 : node12338;
														assign node12338 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12341 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12344 = (inp[0]) ? node12348 : node12345;
														assign node12345 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12348 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12351 = (inp[2]) ? node12359 : node12352;
													assign node12352 = (inp[7]) ? node12356 : node12353;
														assign node12353 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12356 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12359 = (inp[0]) ? node12363 : node12360;
														assign node12360 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12363 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node12366 = (inp[8]) ? node12380 : node12367;
												assign node12367 = (inp[9]) ? node12375 : node12368;
													assign node12368 = (inp[2]) ? node12372 : node12369;
														assign node12369 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12372 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node12375 = (inp[2]) ? node12377 : 16'b0000000001111111;
														assign node12377 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12380 = (inp[2]) ? node12388 : node12381;
													assign node12381 = (inp[9]) ? node12385 : node12382;
														assign node12382 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12385 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12388 = (inp[9]) ? node12390 : 16'b0000000000111111;
														assign node12390 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node12393 = (inp[0]) ? node12509 : node12394;
									assign node12394 = (inp[14]) ? node12450 : node12395;
										assign node12395 = (inp[12]) ? node12425 : node12396;
											assign node12396 = (inp[13]) ? node12410 : node12397;
												assign node12397 = (inp[9]) ? node12403 : node12398;
													assign node12398 = (inp[8]) ? node12400 : 16'b0000011111111111;
														assign node12400 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12403 = (inp[8]) ? node12407 : node12404;
														assign node12404 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12407 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12410 = (inp[9]) ? node12418 : node12411;
													assign node12411 = (inp[8]) ? node12415 : node12412;
														assign node12412 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12415 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node12418 = (inp[7]) ? node12422 : node12419;
														assign node12419 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12422 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node12425 = (inp[3]) ? node12439 : node12426;
												assign node12426 = (inp[9]) ? node12434 : node12427;
													assign node12427 = (inp[13]) ? node12431 : node12428;
														assign node12428 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12431 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node12434 = (inp[2]) ? 16'b0000000001111111 : node12435;
														assign node12435 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12439 = (inp[8]) ? node12445 : node12440;
													assign node12440 = (inp[9]) ? node12442 : 16'b0000000011111111;
														assign node12442 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12445 = (inp[2]) ? 16'b0000000001111111 : node12446;
														assign node12446 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node12450 = (inp[13]) ? node12480 : node12451;
											assign node12451 = (inp[7]) ? node12465 : node12452;
												assign node12452 = (inp[2]) ? node12458 : node12453;
													assign node12453 = (inp[9]) ? 16'b0000000111111111 : node12454;
														assign node12454 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12458 = (inp[8]) ? node12462 : node12459;
														assign node12459 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12462 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12465 = (inp[8]) ? node12473 : node12466;
													assign node12466 = (inp[9]) ? node12470 : node12467;
														assign node12467 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12470 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node12473 = (inp[3]) ? node12477 : node12474;
														assign node12474 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12477 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node12480 = (inp[2]) ? node12496 : node12481;
												assign node12481 = (inp[7]) ? node12489 : node12482;
													assign node12482 = (inp[8]) ? node12486 : node12483;
														assign node12483 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12486 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12489 = (inp[3]) ? node12493 : node12490;
														assign node12490 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12493 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12496 = (inp[9]) ? node12502 : node12497;
													assign node12497 = (inp[7]) ? node12499 : 16'b0000000001111111;
														assign node12499 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12502 = (inp[7]) ? node12506 : node12503;
														assign node12503 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12506 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node12509 = (inp[2]) ? node12571 : node12510;
										assign node12510 = (inp[13]) ? node12542 : node12511;
											assign node12511 = (inp[12]) ? node12527 : node12512;
												assign node12512 = (inp[3]) ? node12520 : node12513;
													assign node12513 = (inp[9]) ? node12517 : node12514;
														assign node12514 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12517 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12520 = (inp[7]) ? node12524 : node12521;
														assign node12521 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12524 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12527 = (inp[8]) ? node12535 : node12528;
													assign node12528 = (inp[3]) ? node12532 : node12529;
														assign node12529 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node12532 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12535 = (inp[14]) ? node12539 : node12536;
														assign node12536 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12539 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node12542 = (inp[9]) ? node12556 : node12543;
												assign node12543 = (inp[3]) ? node12549 : node12544;
													assign node12544 = (inp[8]) ? node12546 : 16'b0000000011111111;
														assign node12546 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12549 = (inp[7]) ? node12553 : node12550;
														assign node12550 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node12553 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12556 = (inp[8]) ? node12564 : node12557;
													assign node12557 = (inp[14]) ? node12561 : node12558;
														assign node12558 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12561 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12564 = (inp[12]) ? node12568 : node12565;
														assign node12565 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node12568 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node12571 = (inp[14]) ? node12603 : node12572;
											assign node12572 = (inp[8]) ? node12588 : node12573;
												assign node12573 = (inp[13]) ? node12581 : node12574;
													assign node12574 = (inp[9]) ? node12578 : node12575;
														assign node12575 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12578 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12581 = (inp[7]) ? node12585 : node12582;
														assign node12582 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12585 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node12588 = (inp[3]) ? node12596 : node12589;
													assign node12589 = (inp[13]) ? node12593 : node12590;
														assign node12590 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12593 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12596 = (inp[12]) ? node12600 : node12597;
														assign node12597 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12600 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node12603 = (inp[12]) ? node12617 : node12604;
												assign node12604 = (inp[3]) ? node12610 : node12605;
													assign node12605 = (inp[13]) ? 16'b0000000001111111 : node12606;
														assign node12606 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12610 = (inp[13]) ? node12614 : node12611;
														assign node12611 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12614 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node12617 = (inp[9]) ? node12623 : node12618;
													assign node12618 = (inp[8]) ? 16'b0000000000111111 : node12619;
														assign node12619 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node12623 = (inp[7]) ? node12627 : node12624;
														assign node12624 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node12627 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node12630 = (inp[15]) ? node13132 : node12631;
							assign node12631 = (inp[0]) ? node12883 : node12632;
								assign node12632 = (inp[7]) ? node12756 : node12633;
									assign node12633 = (inp[2]) ? node12697 : node12634;
										assign node12634 = (inp[11]) ? node12666 : node12635;
											assign node12635 = (inp[13]) ? node12651 : node12636;
												assign node12636 = (inp[8]) ? node12644 : node12637;
													assign node12637 = (inp[3]) ? node12641 : node12638;
														assign node12638 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node12641 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node12644 = (inp[3]) ? node12648 : node12645;
														assign node12645 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12648 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node12651 = (inp[14]) ? node12659 : node12652;
													assign node12652 = (inp[8]) ? node12656 : node12653;
														assign node12653 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12656 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12659 = (inp[9]) ? node12663 : node12660;
														assign node12660 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12663 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node12666 = (inp[14]) ? node12682 : node12667;
												assign node12667 = (inp[3]) ? node12675 : node12668;
													assign node12668 = (inp[13]) ? node12672 : node12669;
														assign node12669 = (inp[12]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node12672 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12675 = (inp[12]) ? node12679 : node12676;
														assign node12676 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12679 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12682 = (inp[9]) ? node12690 : node12683;
													assign node12683 = (inp[12]) ? node12687 : node12684;
														assign node12684 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12687 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12690 = (inp[13]) ? node12694 : node12691;
														assign node12691 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12694 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node12697 = (inp[12]) ? node12727 : node12698;
											assign node12698 = (inp[13]) ? node12712 : node12699;
												assign node12699 = (inp[14]) ? node12707 : node12700;
													assign node12700 = (inp[11]) ? node12704 : node12701;
														assign node12701 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12704 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12707 = (inp[9]) ? 16'b0000000011111111 : node12708;
														assign node12708 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node12712 = (inp[14]) ? node12720 : node12713;
													assign node12713 = (inp[3]) ? node12717 : node12714;
														assign node12714 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12717 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12720 = (inp[11]) ? node12724 : node12721;
														assign node12721 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12724 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node12727 = (inp[9]) ? node12743 : node12728;
												assign node12728 = (inp[3]) ? node12736 : node12729;
													assign node12729 = (inp[8]) ? node12733 : node12730;
														assign node12730 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12733 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12736 = (inp[14]) ? node12740 : node12737;
														assign node12737 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12740 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node12743 = (inp[8]) ? node12749 : node12744;
													assign node12744 = (inp[14]) ? node12746 : 16'b0000000111111111;
														assign node12746 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12749 = (inp[13]) ? node12753 : node12750;
														assign node12750 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12753 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node12756 = (inp[3]) ? node12820 : node12757;
										assign node12757 = (inp[12]) ? node12789 : node12758;
											assign node12758 = (inp[9]) ? node12774 : node12759;
												assign node12759 = (inp[8]) ? node12767 : node12760;
													assign node12760 = (inp[11]) ? node12764 : node12761;
														assign node12761 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12764 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12767 = (inp[14]) ? node12771 : node12768;
														assign node12768 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node12771 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12774 = (inp[13]) ? node12782 : node12775;
													assign node12775 = (inp[11]) ? node12779 : node12776;
														assign node12776 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12779 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12782 = (inp[14]) ? node12786 : node12783;
														assign node12783 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node12786 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
											assign node12789 = (inp[2]) ? node12805 : node12790;
												assign node12790 = (inp[9]) ? node12798 : node12791;
													assign node12791 = (inp[8]) ? node12795 : node12792;
														assign node12792 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12795 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12798 = (inp[8]) ? node12802 : node12799;
														assign node12799 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12802 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12805 = (inp[11]) ? node12813 : node12806;
													assign node12806 = (inp[14]) ? node12810 : node12807;
														assign node12807 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12810 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12813 = (inp[9]) ? node12817 : node12814;
														assign node12814 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12817 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
										assign node12820 = (inp[14]) ? node12852 : node12821;
											assign node12821 = (inp[13]) ? node12837 : node12822;
												assign node12822 = (inp[12]) ? node12830 : node12823;
													assign node12823 = (inp[9]) ? node12827 : node12824;
														assign node12824 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12827 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12830 = (inp[9]) ? node12834 : node12831;
														assign node12831 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12834 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12837 = (inp[8]) ? node12845 : node12838;
													assign node12838 = (inp[2]) ? node12842 : node12839;
														assign node12839 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node12842 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12845 = (inp[2]) ? node12849 : node12846;
														assign node12846 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node12849 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node12852 = (inp[11]) ? node12868 : node12853;
												assign node12853 = (inp[8]) ? node12861 : node12854;
													assign node12854 = (inp[9]) ? node12858 : node12855;
														assign node12855 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node12858 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12861 = (inp[12]) ? node12865 : node12862;
														assign node12862 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node12865 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node12868 = (inp[2]) ? node12876 : node12869;
													assign node12869 = (inp[13]) ? node12873 : node12870;
														assign node12870 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12873 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node12876 = (inp[12]) ? node12880 : node12877;
														assign node12877 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node12880 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node12883 = (inp[8]) ? node13009 : node12884;
									assign node12884 = (inp[14]) ? node12946 : node12885;
										assign node12885 = (inp[3]) ? node12917 : node12886;
											assign node12886 = (inp[11]) ? node12902 : node12887;
												assign node12887 = (inp[13]) ? node12895 : node12888;
													assign node12888 = (inp[2]) ? node12892 : node12889;
														assign node12889 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node12892 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node12895 = (inp[9]) ? node12899 : node12896;
														assign node12896 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12899 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node12902 = (inp[7]) ? node12910 : node12903;
													assign node12903 = (inp[2]) ? node12907 : node12904;
														assign node12904 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12907 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12910 = (inp[13]) ? node12914 : node12911;
														assign node12911 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12914 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node12917 = (inp[12]) ? node12933 : node12918;
												assign node12918 = (inp[11]) ? node12926 : node12919;
													assign node12919 = (inp[13]) ? node12923 : node12920;
														assign node12920 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12923 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12926 = (inp[13]) ? node12930 : node12927;
														assign node12927 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12930 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12933 = (inp[2]) ? node12939 : node12934;
													assign node12934 = (inp[9]) ? 16'b0000000011111111 : node12935;
														assign node12935 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node12939 = (inp[13]) ? node12943 : node12940;
														assign node12940 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node12943 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node12946 = (inp[7]) ? node12978 : node12947;
											assign node12947 = (inp[12]) ? node12963 : node12948;
												assign node12948 = (inp[2]) ? node12956 : node12949;
													assign node12949 = (inp[11]) ? node12953 : node12950;
														assign node12950 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node12953 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node12956 = (inp[13]) ? node12960 : node12957;
														assign node12957 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12960 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node12963 = (inp[11]) ? node12971 : node12964;
													assign node12964 = (inp[9]) ? node12968 : node12965;
														assign node12965 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node12968 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12971 = (inp[9]) ? node12975 : node12972;
														assign node12972 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12975 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node12978 = (inp[13]) ? node12994 : node12979;
												assign node12979 = (inp[11]) ? node12987 : node12980;
													assign node12980 = (inp[2]) ? node12984 : node12981;
														assign node12981 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node12984 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node12987 = (inp[9]) ? node12991 : node12988;
														assign node12988 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12991 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node12994 = (inp[9]) ? node13002 : node12995;
													assign node12995 = (inp[2]) ? node12999 : node12996;
														assign node12996 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node12999 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13002 = (inp[2]) ? node13006 : node13003;
														assign node13003 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13006 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node13009 = (inp[3]) ? node13073 : node13010;
										assign node13010 = (inp[7]) ? node13042 : node13011;
											assign node13011 = (inp[14]) ? node13027 : node13012;
												assign node13012 = (inp[13]) ? node13020 : node13013;
													assign node13013 = (inp[11]) ? node13017 : node13014;
														assign node13014 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13017 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13020 = (inp[12]) ? node13024 : node13021;
														assign node13021 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13024 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13027 = (inp[11]) ? node13035 : node13028;
													assign node13028 = (inp[2]) ? node13032 : node13029;
														assign node13029 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node13032 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13035 = (inp[9]) ? node13039 : node13036;
														assign node13036 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13039 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13042 = (inp[11]) ? node13058 : node13043;
												assign node13043 = (inp[14]) ? node13051 : node13044;
													assign node13044 = (inp[2]) ? node13048 : node13045;
														assign node13045 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13048 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13051 = (inp[9]) ? node13055 : node13052;
														assign node13052 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13055 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node13058 = (inp[13]) ? node13066 : node13059;
													assign node13059 = (inp[9]) ? node13063 : node13060;
														assign node13060 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13063 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node13066 = (inp[12]) ? node13070 : node13067;
														assign node13067 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node13070 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node13073 = (inp[11]) ? node13101 : node13074;
											assign node13074 = (inp[7]) ? node13088 : node13075;
												assign node13075 = (inp[9]) ? node13081 : node13076;
													assign node13076 = (inp[14]) ? 16'b0000000011111111 : node13077;
														assign node13077 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13081 = (inp[14]) ? node13085 : node13082;
														assign node13082 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13085 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node13088 = (inp[13]) ? node13094 : node13089;
													assign node13089 = (inp[2]) ? node13091 : 16'b0000000001111111;
														assign node13091 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13094 = (inp[12]) ? node13098 : node13095;
														assign node13095 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13098 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node13101 = (inp[9]) ? node13117 : node13102;
												assign node13102 = (inp[12]) ? node13110 : node13103;
													assign node13103 = (inp[13]) ? node13107 : node13104;
														assign node13104 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13107 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13110 = (inp[2]) ? node13114 : node13111;
														assign node13111 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13114 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node13117 = (inp[14]) ? node13125 : node13118;
													assign node13118 = (inp[12]) ? node13122 : node13119;
														assign node13119 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13122 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node13125 = (inp[7]) ? node13129 : node13126;
														assign node13126 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node13129 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node13132 = (inp[13]) ? node13374 : node13133;
								assign node13133 = (inp[12]) ? node13253 : node13134;
									assign node13134 = (inp[0]) ? node13194 : node13135;
										assign node13135 = (inp[8]) ? node13165 : node13136;
											assign node13136 = (inp[7]) ? node13150 : node13137;
												assign node13137 = (inp[2]) ? node13145 : node13138;
													assign node13138 = (inp[11]) ? node13142 : node13139;
														assign node13139 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13142 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13145 = (inp[11]) ? 16'b0000000111111111 : node13146;
														assign node13146 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node13150 = (inp[2]) ? node13158 : node13151;
													assign node13151 = (inp[14]) ? node13155 : node13152;
														assign node13152 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13155 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13158 = (inp[3]) ? node13162 : node13159;
														assign node13159 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13162 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node13165 = (inp[7]) ? node13181 : node13166;
												assign node13166 = (inp[9]) ? node13174 : node13167;
													assign node13167 = (inp[14]) ? node13171 : node13168;
														assign node13168 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13171 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13174 = (inp[3]) ? node13178 : node13175;
														assign node13175 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13178 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13181 = (inp[3]) ? node13187 : node13182;
													assign node13182 = (inp[2]) ? 16'b0000000001111111 : node13183;
														assign node13183 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13187 = (inp[14]) ? node13191 : node13188;
														assign node13188 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13191 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node13194 = (inp[8]) ? node13224 : node13195;
											assign node13195 = (inp[14]) ? node13211 : node13196;
												assign node13196 = (inp[3]) ? node13204 : node13197;
													assign node13197 = (inp[7]) ? node13201 : node13198;
														assign node13198 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13201 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node13204 = (inp[7]) ? node13208 : node13205;
														assign node13205 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node13208 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13211 = (inp[3]) ? node13219 : node13212;
													assign node13212 = (inp[7]) ? node13216 : node13213;
														assign node13213 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13216 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node13219 = (inp[7]) ? node13221 : 16'b0000000001111111;
														assign node13221 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13224 = (inp[2]) ? node13238 : node13225;
												assign node13225 = (inp[11]) ? node13231 : node13226;
													assign node13226 = (inp[14]) ? node13228 : 16'b0000000111111111;
														assign node13228 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13231 = (inp[14]) ? node13235 : node13232;
														assign node13232 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13235 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13238 = (inp[3]) ? node13246 : node13239;
													assign node13239 = (inp[11]) ? node13243 : node13240;
														assign node13240 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13243 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13246 = (inp[9]) ? node13250 : node13247;
														assign node13247 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13250 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node13253 = (inp[7]) ? node13313 : node13254;
										assign node13254 = (inp[9]) ? node13282 : node13255;
											assign node13255 = (inp[2]) ? node13267 : node13256;
												assign node13256 = (inp[11]) ? node13262 : node13257;
													assign node13257 = (inp[8]) ? node13259 : 16'b0000001111111111;
														assign node13259 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node13262 = (inp[8]) ? node13264 : 16'b0000000011111111;
														assign node13264 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13267 = (inp[8]) ? node13275 : node13268;
													assign node13268 = (inp[11]) ? node13272 : node13269;
														assign node13269 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13272 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node13275 = (inp[11]) ? node13279 : node13276;
														assign node13276 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13279 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node13282 = (inp[14]) ? node13298 : node13283;
												assign node13283 = (inp[2]) ? node13291 : node13284;
													assign node13284 = (inp[3]) ? node13288 : node13285;
														assign node13285 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node13288 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node13291 = (inp[0]) ? node13295 : node13292;
														assign node13292 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13295 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node13298 = (inp[11]) ? node13306 : node13299;
													assign node13299 = (inp[8]) ? node13303 : node13300;
														assign node13300 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13303 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13306 = (inp[3]) ? node13310 : node13307;
														assign node13307 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13310 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node13313 = (inp[14]) ? node13343 : node13314;
											assign node13314 = (inp[3]) ? node13328 : node13315;
												assign node13315 = (inp[0]) ? node13323 : node13316;
													assign node13316 = (inp[8]) ? node13320 : node13317;
														assign node13317 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13320 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13323 = (inp[8]) ? 16'b0000000000111111 : node13324;
														assign node13324 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node13328 = (inp[9]) ? node13336 : node13329;
													assign node13329 = (inp[11]) ? node13333 : node13330;
														assign node13330 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13333 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13336 = (inp[2]) ? node13340 : node13337;
														assign node13337 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13340 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node13343 = (inp[3]) ? node13359 : node13344;
												assign node13344 = (inp[11]) ? node13352 : node13345;
													assign node13345 = (inp[9]) ? node13349 : node13346;
														assign node13346 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13349 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node13352 = (inp[9]) ? node13356 : node13353;
														assign node13353 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node13356 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node13359 = (inp[2]) ? node13367 : node13360;
													assign node13360 = (inp[8]) ? node13364 : node13361;
														assign node13361 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13364 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node13367 = (inp[0]) ? node13371 : node13368;
														assign node13368 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node13371 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node13374 = (inp[9]) ? node13478 : node13375;
									assign node13375 = (inp[2]) ? node13431 : node13376;
										assign node13376 = (inp[14]) ? node13400 : node13377;
											assign node13377 = (inp[3]) ? node13391 : node13378;
												assign node13378 = (inp[0]) ? node13384 : node13379;
													assign node13379 = (inp[12]) ? node13381 : 16'b0000000111111111;
														assign node13381 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13384 = (inp[8]) ? node13388 : node13385;
														assign node13385 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13388 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13391 = (inp[11]) ? node13393 : 16'b0000000011111111;
													assign node13393 = (inp[12]) ? node13397 : node13394;
														assign node13394 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13397 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node13400 = (inp[12]) ? node13416 : node13401;
												assign node13401 = (inp[11]) ? node13409 : node13402;
													assign node13402 = (inp[8]) ? node13406 : node13403;
														assign node13403 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node13406 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13409 = (inp[0]) ? node13413 : node13410;
														assign node13410 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13413 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13416 = (inp[3]) ? node13424 : node13417;
													assign node13417 = (inp[11]) ? node13421 : node13418;
														assign node13418 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13421 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13424 = (inp[0]) ? node13428 : node13425;
														assign node13425 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node13428 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node13431 = (inp[0]) ? node13457 : node13432;
											assign node13432 = (inp[3]) ? node13444 : node13433;
												assign node13433 = (inp[11]) ? node13439 : node13434;
													assign node13434 = (inp[12]) ? node13436 : 16'b0000000011111111;
														assign node13436 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13439 = (inp[14]) ? 16'b0000000001111111 : node13440;
														assign node13440 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13444 = (inp[11]) ? node13450 : node13445;
													assign node13445 = (inp[8]) ? 16'b0000000001111111 : node13446;
														assign node13446 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13450 = (inp[12]) ? node13454 : node13451;
														assign node13451 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node13454 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node13457 = (inp[7]) ? node13465 : node13458;
												assign node13458 = (inp[14]) ? 16'b0000000000111111 : node13459;
													assign node13459 = (inp[8]) ? node13461 : 16'b0000000001111111;
														assign node13461 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13465 = (inp[12]) ? node13473 : node13466;
													assign node13466 = (inp[8]) ? node13470 : node13467;
														assign node13467 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13470 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node13473 = (inp[14]) ? 16'b0000000000001111 : node13474;
														assign node13474 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node13478 = (inp[8]) ? node13532 : node13479;
										assign node13479 = (inp[14]) ? node13509 : node13480;
											assign node13480 = (inp[12]) ? node13494 : node13481;
												assign node13481 = (inp[0]) ? node13489 : node13482;
													assign node13482 = (inp[3]) ? node13486 : node13483;
														assign node13483 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13486 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13489 = (inp[7]) ? 16'b0000000000111111 : node13490;
														assign node13490 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node13494 = (inp[2]) ? node13502 : node13495;
													assign node13495 = (inp[3]) ? node13499 : node13496;
														assign node13496 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13499 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13502 = (inp[7]) ? node13506 : node13503;
														assign node13503 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node13506 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node13509 = (inp[7]) ? node13523 : node13510;
												assign node13510 = (inp[11]) ? node13518 : node13511;
													assign node13511 = (inp[0]) ? node13515 : node13512;
														assign node13512 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13515 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13518 = (inp[2]) ? node13520 : 16'b0000000000111111;
														assign node13520 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node13523 = (inp[12]) ? node13527 : node13524;
													assign node13524 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node13527 = (inp[3]) ? node13529 : 16'b0000000000011111;
														assign node13529 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node13532 = (inp[12]) ? node13564 : node13533;
											assign node13533 = (inp[11]) ? node13549 : node13534;
												assign node13534 = (inp[14]) ? node13542 : node13535;
													assign node13535 = (inp[3]) ? node13539 : node13536;
														assign node13536 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13539 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13542 = (inp[3]) ? node13546 : node13543;
														assign node13543 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node13546 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node13549 = (inp[7]) ? node13557 : node13550;
													assign node13550 = (inp[0]) ? node13554 : node13551;
														assign node13551 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13554 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node13557 = (inp[14]) ? node13561 : node13558;
														assign node13558 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node13561 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000001111;
											assign node13564 = (inp[14]) ? node13580 : node13565;
												assign node13565 = (inp[7]) ? node13573 : node13566;
													assign node13566 = (inp[2]) ? node13570 : node13567;
														assign node13567 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13570 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node13573 = (inp[11]) ? node13577 : node13574;
														assign node13574 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node13577 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node13580 = (inp[2]) ? node13588 : node13581;
													assign node13581 = (inp[0]) ? node13585 : node13582;
														assign node13582 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node13585 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node13588 = (inp[7]) ? node13592 : node13589;
														assign node13589 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node13592 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000000111;
					assign node13595 = (inp[12]) ? node14575 : node13596;
						assign node13596 = (inp[0]) ? node14084 : node13597;
							assign node13597 = (inp[8]) ? node13845 : node13598;
								assign node13598 = (inp[3]) ? node13720 : node13599;
									assign node13599 = (inp[14]) ? node13659 : node13600;
										assign node13600 = (inp[11]) ? node13630 : node13601;
											assign node13601 = (inp[2]) ? node13615 : node13602;
												assign node13602 = (inp[9]) ? node13610 : node13603;
													assign node13603 = (inp[7]) ? node13607 : node13604;
														assign node13604 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node13607 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13610 = (inp[4]) ? 16'b0000001111111111 : node13611;
														assign node13611 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node13615 = (inp[13]) ? node13623 : node13616;
													assign node13616 = (inp[4]) ? node13620 : node13617;
														assign node13617 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13620 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13623 = (inp[15]) ? node13627 : node13624;
														assign node13624 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13627 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node13630 = (inp[2]) ? node13646 : node13631;
												assign node13631 = (inp[7]) ? node13639 : node13632;
													assign node13632 = (inp[13]) ? node13636 : node13633;
														assign node13633 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13636 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13639 = (inp[4]) ? node13643 : node13640;
														assign node13640 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13643 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13646 = (inp[15]) ? node13652 : node13647;
													assign node13647 = (inp[9]) ? 16'b0000000111111111 : node13648;
														assign node13648 = (inp[13]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node13652 = (inp[7]) ? node13656 : node13653;
														assign node13653 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13656 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node13659 = (inp[9]) ? node13691 : node13660;
											assign node13660 = (inp[11]) ? node13676 : node13661;
												assign node13661 = (inp[13]) ? node13669 : node13662;
													assign node13662 = (inp[15]) ? node13666 : node13663;
														assign node13663 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13666 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13669 = (inp[4]) ? node13673 : node13670;
														assign node13670 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node13673 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13676 = (inp[4]) ? node13684 : node13677;
													assign node13677 = (inp[7]) ? node13681 : node13678;
														assign node13678 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13681 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node13684 = (inp[15]) ? node13688 : node13685;
														assign node13685 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13688 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node13691 = (inp[15]) ? node13705 : node13692;
												assign node13692 = (inp[4]) ? node13700 : node13693;
													assign node13693 = (inp[2]) ? node13697 : node13694;
														assign node13694 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node13697 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node13700 = (inp[13]) ? node13702 : 16'b0000000011111111;
														assign node13702 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13705 = (inp[7]) ? node13713 : node13706;
													assign node13706 = (inp[2]) ? node13710 : node13707;
														assign node13707 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13710 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13713 = (inp[2]) ? node13717 : node13714;
														assign node13714 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13717 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node13720 = (inp[15]) ? node13784 : node13721;
										assign node13721 = (inp[14]) ? node13753 : node13722;
											assign node13722 = (inp[7]) ? node13738 : node13723;
												assign node13723 = (inp[11]) ? node13731 : node13724;
													assign node13724 = (inp[4]) ? node13728 : node13725;
														assign node13725 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node13728 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node13731 = (inp[9]) ? node13735 : node13732;
														assign node13732 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13735 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13738 = (inp[2]) ? node13746 : node13739;
													assign node13739 = (inp[4]) ? node13743 : node13740;
														assign node13740 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13743 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13746 = (inp[11]) ? node13750 : node13747;
														assign node13747 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13750 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node13753 = (inp[7]) ? node13769 : node13754;
												assign node13754 = (inp[2]) ? node13762 : node13755;
													assign node13755 = (inp[9]) ? node13759 : node13756;
														assign node13756 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13759 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node13762 = (inp[11]) ? node13766 : node13763;
														assign node13763 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13766 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node13769 = (inp[9]) ? node13777 : node13770;
													assign node13770 = (inp[4]) ? node13774 : node13771;
														assign node13771 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13774 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node13777 = (inp[2]) ? node13781 : node13778;
														assign node13778 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13781 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node13784 = (inp[13]) ? node13816 : node13785;
											assign node13785 = (inp[9]) ? node13801 : node13786;
												assign node13786 = (inp[7]) ? node13794 : node13787;
													assign node13787 = (inp[4]) ? node13791 : node13788;
														assign node13788 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13791 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13794 = (inp[11]) ? node13798 : node13795;
														assign node13795 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13798 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node13801 = (inp[4]) ? node13809 : node13802;
													assign node13802 = (inp[11]) ? node13806 : node13803;
														assign node13803 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node13806 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node13809 = (inp[14]) ? node13813 : node13810;
														assign node13810 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13813 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13816 = (inp[11]) ? node13830 : node13817;
												assign node13817 = (inp[14]) ? node13823 : node13818;
													assign node13818 = (inp[9]) ? node13820 : 16'b0000000011111111;
														assign node13820 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13823 = (inp[2]) ? node13827 : node13824;
														assign node13824 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13827 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13830 = (inp[2]) ? node13838 : node13831;
													assign node13831 = (inp[4]) ? node13835 : node13832;
														assign node13832 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13835 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13838 = (inp[14]) ? node13842 : node13839;
														assign node13839 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node13842 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node13845 = (inp[11]) ? node13965 : node13846;
									assign node13846 = (inp[2]) ? node13902 : node13847;
										assign node13847 = (inp[3]) ? node13875 : node13848;
											assign node13848 = (inp[13]) ? node13862 : node13849;
												assign node13849 = (inp[7]) ? node13855 : node13850;
													assign node13850 = (inp[4]) ? 16'b0000001111111111 : node13851;
														assign node13851 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node13855 = (inp[9]) ? node13859 : node13856;
														assign node13856 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13859 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node13862 = (inp[7]) ? node13870 : node13863;
													assign node13863 = (inp[4]) ? node13867 : node13864;
														assign node13864 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node13867 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13870 = (inp[14]) ? 16'b0000000011111111 : node13871;
														assign node13871 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node13875 = (inp[9]) ? node13889 : node13876;
												assign node13876 = (inp[7]) ? node13884 : node13877;
													assign node13877 = (inp[15]) ? node13881 : node13878;
														assign node13878 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node13881 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13884 = (inp[15]) ? 16'b0000000001111111 : node13885;
														assign node13885 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node13889 = (inp[4]) ? node13897 : node13890;
													assign node13890 = (inp[14]) ? node13894 : node13891;
														assign node13891 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13894 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13897 = (inp[13]) ? node13899 : 16'b0000000001111111;
														assign node13899 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node13902 = (inp[14]) ? node13934 : node13903;
											assign node13903 = (inp[15]) ? node13919 : node13904;
												assign node13904 = (inp[3]) ? node13912 : node13905;
													assign node13905 = (inp[7]) ? node13909 : node13906;
														assign node13906 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node13909 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13912 = (inp[9]) ? node13916 : node13913;
														assign node13913 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node13916 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13919 = (inp[4]) ? node13927 : node13920;
													assign node13920 = (inp[7]) ? node13924 : node13921;
														assign node13921 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13924 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13927 = (inp[13]) ? node13931 : node13928;
														assign node13928 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node13931 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node13934 = (inp[7]) ? node13950 : node13935;
												assign node13935 = (inp[15]) ? node13943 : node13936;
													assign node13936 = (inp[3]) ? node13940 : node13937;
														assign node13937 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13940 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13943 = (inp[4]) ? node13947 : node13944;
														assign node13944 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13947 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node13950 = (inp[3]) ? node13958 : node13951;
													assign node13951 = (inp[4]) ? node13955 : node13952;
														assign node13952 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node13955 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node13958 = (inp[13]) ? node13962 : node13959;
														assign node13959 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node13962 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node13965 = (inp[9]) ? node14023 : node13966;
										assign node13966 = (inp[2]) ? node13996 : node13967;
											assign node13967 = (inp[13]) ? node13983 : node13968;
												assign node13968 = (inp[14]) ? node13976 : node13969;
													assign node13969 = (inp[4]) ? node13973 : node13970;
														assign node13970 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node13973 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node13976 = (inp[15]) ? node13980 : node13977;
														assign node13977 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node13980 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node13983 = (inp[15]) ? node13991 : node13984;
													assign node13984 = (inp[3]) ? node13988 : node13985;
														assign node13985 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node13988 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node13991 = (inp[3]) ? 16'b0000000000111111 : node13992;
														assign node13992 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node13996 = (inp[14]) ? node14012 : node13997;
												assign node13997 = (inp[7]) ? node14005 : node13998;
													assign node13998 = (inp[13]) ? node14002 : node13999;
														assign node13999 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14002 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14005 = (inp[3]) ? node14009 : node14006;
														assign node14006 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14009 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14012 = (inp[3]) ? node14016 : node14013;
													assign node14013 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node14016 = (inp[15]) ? node14020 : node14017;
														assign node14017 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14020 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node14023 = (inp[13]) ? node14055 : node14024;
											assign node14024 = (inp[3]) ? node14040 : node14025;
												assign node14025 = (inp[15]) ? node14033 : node14026;
													assign node14026 = (inp[14]) ? node14030 : node14027;
														assign node14027 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14030 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14033 = (inp[2]) ? node14037 : node14034;
														assign node14034 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14037 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14040 = (inp[14]) ? node14048 : node14041;
													assign node14041 = (inp[7]) ? node14045 : node14042;
														assign node14042 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14045 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node14048 = (inp[7]) ? node14052 : node14049;
														assign node14049 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node14052 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node14055 = (inp[15]) ? node14069 : node14056;
												assign node14056 = (inp[2]) ? node14064 : node14057;
													assign node14057 = (inp[14]) ? node14061 : node14058;
														assign node14058 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node14061 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14064 = (inp[7]) ? node14066 : 16'b0000000000111111;
														assign node14066 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14069 = (inp[7]) ? node14077 : node14070;
													assign node14070 = (inp[4]) ? node14074 : node14071;
														assign node14071 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node14074 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node14077 = (inp[14]) ? node14081 : node14078;
														assign node14078 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node14081 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node14084 = (inp[14]) ? node14330 : node14085;
								assign node14085 = (inp[15]) ? node14207 : node14086;
									assign node14086 = (inp[11]) ? node14146 : node14087;
										assign node14087 = (inp[13]) ? node14115 : node14088;
											assign node14088 = (inp[2]) ? node14102 : node14089;
												assign node14089 = (inp[8]) ? node14097 : node14090;
													assign node14090 = (inp[9]) ? node14094 : node14091;
														assign node14091 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node14094 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node14097 = (inp[3]) ? 16'b0000000111111111 : node14098;
														assign node14098 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000111111111;
												assign node14102 = (inp[3]) ? node14110 : node14103;
													assign node14103 = (inp[4]) ? node14107 : node14104;
														assign node14104 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14107 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node14110 = (inp[7]) ? 16'b0000000001111111 : node14111;
														assign node14111 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node14115 = (inp[8]) ? node14131 : node14116;
												assign node14116 = (inp[3]) ? node14124 : node14117;
													assign node14117 = (inp[4]) ? node14121 : node14118;
														assign node14118 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14121 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14124 = (inp[9]) ? node14128 : node14125;
														assign node14125 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14128 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14131 = (inp[3]) ? node14139 : node14132;
													assign node14132 = (inp[4]) ? node14136 : node14133;
														assign node14133 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14136 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14139 = (inp[9]) ? node14143 : node14140;
														assign node14140 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14143 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14146 = (inp[9]) ? node14176 : node14147;
											assign node14147 = (inp[8]) ? node14163 : node14148;
												assign node14148 = (inp[7]) ? node14156 : node14149;
													assign node14149 = (inp[13]) ? node14153 : node14150;
														assign node14150 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14153 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14156 = (inp[4]) ? node14160 : node14157;
														assign node14157 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14160 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14163 = (inp[2]) ? node14171 : node14164;
													assign node14164 = (inp[3]) ? node14168 : node14165;
														assign node14165 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node14168 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node14171 = (inp[7]) ? 16'b0000000001111111 : node14172;
														assign node14172 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14176 = (inp[7]) ? node14192 : node14177;
												assign node14177 = (inp[2]) ? node14185 : node14178;
													assign node14178 = (inp[13]) ? node14182 : node14179;
														assign node14179 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14182 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14185 = (inp[8]) ? node14189 : node14186;
														assign node14186 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14189 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node14192 = (inp[13]) ? node14200 : node14193;
													assign node14193 = (inp[2]) ? node14197 : node14194;
														assign node14194 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14197 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14200 = (inp[2]) ? node14204 : node14201;
														assign node14201 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node14204 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
									assign node14207 = (inp[8]) ? node14271 : node14208;
										assign node14208 = (inp[7]) ? node14240 : node14209;
											assign node14209 = (inp[11]) ? node14225 : node14210;
												assign node14210 = (inp[13]) ? node14218 : node14211;
													assign node14211 = (inp[3]) ? node14215 : node14212;
														assign node14212 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14215 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node14218 = (inp[3]) ? node14222 : node14219;
														assign node14219 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14222 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node14225 = (inp[2]) ? node14233 : node14226;
													assign node14226 = (inp[13]) ? node14230 : node14227;
														assign node14227 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14230 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node14233 = (inp[4]) ? node14237 : node14234;
														assign node14234 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14237 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node14240 = (inp[9]) ? node14256 : node14241;
												assign node14241 = (inp[13]) ? node14249 : node14242;
													assign node14242 = (inp[2]) ? node14246 : node14243;
														assign node14243 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14246 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14249 = (inp[3]) ? node14253 : node14250;
														assign node14250 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14253 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14256 = (inp[2]) ? node14264 : node14257;
													assign node14257 = (inp[3]) ? node14261 : node14258;
														assign node14258 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14261 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14264 = (inp[13]) ? node14268 : node14265;
														assign node14265 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14268 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node14271 = (inp[11]) ? node14301 : node14272;
											assign node14272 = (inp[7]) ? node14288 : node14273;
												assign node14273 = (inp[13]) ? node14281 : node14274;
													assign node14274 = (inp[9]) ? node14278 : node14275;
														assign node14275 = (inp[2]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node14278 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14281 = (inp[2]) ? node14285 : node14282;
														assign node14282 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14285 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node14288 = (inp[9]) ? node14296 : node14289;
													assign node14289 = (inp[13]) ? node14293 : node14290;
														assign node14290 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14293 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14296 = (inp[4]) ? node14298 : 16'b0000000000111111;
														assign node14298 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node14301 = (inp[13]) ? node14315 : node14302;
												assign node14302 = (inp[2]) ? node14308 : node14303;
													assign node14303 = (inp[9]) ? node14305 : 16'b0000000001111111;
														assign node14305 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14308 = (inp[7]) ? node14312 : node14309;
														assign node14309 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node14312 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14315 = (inp[9]) ? node14323 : node14316;
													assign node14316 = (inp[7]) ? node14320 : node14317;
														assign node14317 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14320 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14323 = (inp[2]) ? node14327 : node14324;
														assign node14324 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node14327 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node14330 = (inp[3]) ? node14454 : node14331;
									assign node14331 = (inp[9]) ? node14393 : node14332;
										assign node14332 = (inp[2]) ? node14364 : node14333;
											assign node14333 = (inp[11]) ? node14349 : node14334;
												assign node14334 = (inp[7]) ? node14342 : node14335;
													assign node14335 = (inp[4]) ? node14339 : node14336;
														assign node14336 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14339 = (inp[13]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node14342 = (inp[8]) ? node14346 : node14343;
														assign node14343 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14346 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14349 = (inp[8]) ? node14357 : node14350;
													assign node14350 = (inp[7]) ? node14354 : node14351;
														assign node14351 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14354 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14357 = (inp[4]) ? node14361 : node14358;
														assign node14358 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14361 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node14364 = (inp[13]) ? node14380 : node14365;
												assign node14365 = (inp[4]) ? node14373 : node14366;
													assign node14366 = (inp[7]) ? node14370 : node14367;
														assign node14367 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14370 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14373 = (inp[15]) ? node14377 : node14374;
														assign node14374 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14377 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14380 = (inp[11]) ? node14386 : node14381;
													assign node14381 = (inp[15]) ? node14383 : 16'b0000000011111111;
														assign node14383 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14386 = (inp[15]) ? node14390 : node14387;
														assign node14387 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node14390 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node14393 = (inp[2]) ? node14425 : node14394;
											assign node14394 = (inp[4]) ? node14410 : node14395;
												assign node14395 = (inp[15]) ? node14403 : node14396;
													assign node14396 = (inp[13]) ? node14400 : node14397;
														assign node14397 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14400 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14403 = (inp[13]) ? node14407 : node14404;
														assign node14404 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14407 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14410 = (inp[11]) ? node14418 : node14411;
													assign node14411 = (inp[7]) ? node14415 : node14412;
														assign node14412 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node14415 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14418 = (inp[8]) ? node14422 : node14419;
														assign node14419 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node14422 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14425 = (inp[11]) ? node14441 : node14426;
												assign node14426 = (inp[4]) ? node14434 : node14427;
													assign node14427 = (inp[15]) ? node14431 : node14428;
														assign node14428 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14431 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14434 = (inp[13]) ? node14438 : node14435;
														assign node14435 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14438 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14441 = (inp[4]) ? node14447 : node14442;
													assign node14442 = (inp[13]) ? node14444 : 16'b0000000000111111;
														assign node14444 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14447 = (inp[7]) ? node14451 : node14448;
														assign node14448 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node14451 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node14454 = (inp[13]) ? node14514 : node14455;
										assign node14455 = (inp[2]) ? node14483 : node14456;
											assign node14456 = (inp[4]) ? node14470 : node14457;
												assign node14457 = (inp[15]) ? node14465 : node14458;
													assign node14458 = (inp[8]) ? node14462 : node14459;
														assign node14459 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node14462 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14465 = (inp[8]) ? 16'b0000000001111111 : node14466;
														assign node14466 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14470 = (inp[7]) ? node14476 : node14471;
													assign node14471 = (inp[15]) ? node14473 : 16'b0000000011111111;
														assign node14473 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14476 = (inp[11]) ? node14480 : node14477;
														assign node14477 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14480 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14483 = (inp[9]) ? node14499 : node14484;
												assign node14484 = (inp[11]) ? node14492 : node14485;
													assign node14485 = (inp[8]) ? node14489 : node14486;
														assign node14486 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14489 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14492 = (inp[4]) ? node14496 : node14493;
														assign node14493 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14496 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14499 = (inp[7]) ? node14507 : node14500;
													assign node14500 = (inp[8]) ? node14504 : node14501;
														assign node14501 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14504 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14507 = (inp[11]) ? node14511 : node14508;
														assign node14508 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node14511 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node14514 = (inp[8]) ? node14546 : node14515;
											assign node14515 = (inp[11]) ? node14531 : node14516;
												assign node14516 = (inp[9]) ? node14524 : node14517;
													assign node14517 = (inp[2]) ? node14521 : node14518;
														assign node14518 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14521 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14524 = (inp[4]) ? node14528 : node14525;
														assign node14525 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14528 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14531 = (inp[15]) ? node14539 : node14532;
													assign node14532 = (inp[2]) ? node14536 : node14533;
														assign node14533 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node14536 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node14539 = (inp[9]) ? node14543 : node14540;
														assign node14540 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node14543 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000001111;
											assign node14546 = (inp[9]) ? node14560 : node14547;
												assign node14547 = (inp[4]) ? node14553 : node14548;
													assign node14548 = (inp[11]) ? 16'b0000000000111111 : node14549;
														assign node14549 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14553 = (inp[2]) ? node14557 : node14554;
														assign node14554 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node14557 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node14560 = (inp[11]) ? node14568 : node14561;
													assign node14561 = (inp[15]) ? node14565 : node14562;
														assign node14562 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node14565 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node14568 = (inp[7]) ? node14572 : node14569;
														assign node14569 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000011111;
														assign node14572 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node14575 = (inp[4]) ? node15069 : node14576;
							assign node14576 = (inp[13]) ? node14824 : node14577;
								assign node14577 = (inp[15]) ? node14699 : node14578;
									assign node14578 = (inp[8]) ? node14638 : node14579;
										assign node14579 = (inp[7]) ? node14609 : node14580;
											assign node14580 = (inp[0]) ? node14594 : node14581;
												assign node14581 = (inp[2]) ? node14587 : node14582;
													assign node14582 = (inp[14]) ? 16'b0000001111111111 : node14583;
														assign node14583 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node14587 = (inp[9]) ? node14591 : node14588;
														assign node14588 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14591 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node14594 = (inp[14]) ? node14602 : node14595;
													assign node14595 = (inp[11]) ? node14599 : node14596;
														assign node14596 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14599 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14602 = (inp[3]) ? node14606 : node14603;
														assign node14603 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14606 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node14609 = (inp[0]) ? node14625 : node14610;
												assign node14610 = (inp[2]) ? node14618 : node14611;
													assign node14611 = (inp[9]) ? node14615 : node14612;
														assign node14612 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14615 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14618 = (inp[11]) ? node14622 : node14619;
														assign node14619 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14622 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node14625 = (inp[11]) ? node14633 : node14626;
													assign node14626 = (inp[3]) ? node14630 : node14627;
														assign node14627 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node14630 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14633 = (inp[2]) ? node14635 : 16'b0000000001111111;
														assign node14635 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node14638 = (inp[0]) ? node14668 : node14639;
											assign node14639 = (inp[3]) ? node14655 : node14640;
												assign node14640 = (inp[9]) ? node14648 : node14641;
													assign node14641 = (inp[2]) ? node14645 : node14642;
														assign node14642 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node14645 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14648 = (inp[14]) ? node14652 : node14649;
														assign node14649 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node14652 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node14655 = (inp[11]) ? node14661 : node14656;
													assign node14656 = (inp[9]) ? 16'b0000000001111111 : node14657;
														assign node14657 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14661 = (inp[9]) ? node14665 : node14662;
														assign node14662 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node14665 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node14668 = (inp[14]) ? node14684 : node14669;
												assign node14669 = (inp[9]) ? node14677 : node14670;
													assign node14670 = (inp[3]) ? node14674 : node14671;
														assign node14671 = (inp[11]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node14674 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14677 = (inp[3]) ? node14681 : node14678;
														assign node14678 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14681 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14684 = (inp[11]) ? node14692 : node14685;
													assign node14685 = (inp[3]) ? node14689 : node14686;
														assign node14686 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node14689 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14692 = (inp[2]) ? node14696 : node14693;
														assign node14693 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14696 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node14699 = (inp[0]) ? node14761 : node14700;
										assign node14700 = (inp[7]) ? node14732 : node14701;
											assign node14701 = (inp[2]) ? node14717 : node14702;
												assign node14702 = (inp[11]) ? node14710 : node14703;
													assign node14703 = (inp[8]) ? node14707 : node14704;
														assign node14704 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14707 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14710 = (inp[8]) ? node14714 : node14711;
														assign node14711 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14714 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14717 = (inp[14]) ? node14725 : node14718;
													assign node14718 = (inp[9]) ? node14722 : node14719;
														assign node14719 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14722 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14725 = (inp[11]) ? node14729 : node14726;
														assign node14726 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14729 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node14732 = (inp[3]) ? node14748 : node14733;
												assign node14733 = (inp[14]) ? node14741 : node14734;
													assign node14734 = (inp[11]) ? node14738 : node14735;
														assign node14735 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14738 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14741 = (inp[9]) ? node14745 : node14742;
														assign node14742 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14745 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14748 = (inp[2]) ? node14754 : node14749;
													assign node14749 = (inp[8]) ? node14751 : 16'b0000000001111111;
														assign node14751 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14754 = (inp[14]) ? node14758 : node14755;
														assign node14755 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node14758 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node14761 = (inp[9]) ? node14793 : node14762;
											assign node14762 = (inp[7]) ? node14778 : node14763;
												assign node14763 = (inp[3]) ? node14771 : node14764;
													assign node14764 = (inp[8]) ? node14768 : node14765;
														assign node14765 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14768 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14771 = (inp[2]) ? node14775 : node14772;
														assign node14772 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14775 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14778 = (inp[11]) ? node14786 : node14779;
													assign node14779 = (inp[3]) ? node14783 : node14780;
														assign node14780 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14783 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14786 = (inp[3]) ? node14790 : node14787;
														assign node14787 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node14790 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node14793 = (inp[11]) ? node14809 : node14794;
												assign node14794 = (inp[7]) ? node14802 : node14795;
													assign node14795 = (inp[3]) ? node14799 : node14796;
														assign node14796 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14799 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14802 = (inp[14]) ? node14806 : node14803;
														assign node14803 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node14806 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node14809 = (inp[2]) ? node14817 : node14810;
													assign node14810 = (inp[8]) ? node14814 : node14811;
														assign node14811 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14814 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14817 = (inp[14]) ? node14821 : node14818;
														assign node14818 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node14821 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node14824 = (inp[8]) ? node14946 : node14825;
									assign node14825 = (inp[2]) ? node14885 : node14826;
										assign node14826 = (inp[11]) ? node14856 : node14827;
											assign node14827 = (inp[15]) ? node14841 : node14828;
												assign node14828 = (inp[14]) ? node14836 : node14829;
													assign node14829 = (inp[0]) ? node14833 : node14830;
														assign node14830 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node14833 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node14836 = (inp[7]) ? 16'b0000000001111111 : node14837;
														assign node14837 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node14841 = (inp[9]) ? node14849 : node14842;
													assign node14842 = (inp[3]) ? node14846 : node14843;
														assign node14843 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14846 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14849 = (inp[7]) ? node14853 : node14850;
														assign node14850 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14853 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node14856 = (inp[0]) ? node14872 : node14857;
												assign node14857 = (inp[9]) ? node14865 : node14858;
													assign node14858 = (inp[3]) ? node14862 : node14859;
														assign node14859 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node14862 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14865 = (inp[14]) ? node14869 : node14866;
														assign node14866 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14869 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14872 = (inp[9]) ? node14880 : node14873;
													assign node14873 = (inp[7]) ? node14877 : node14874;
														assign node14874 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14877 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node14880 = (inp[14]) ? node14882 : 16'b0000000000111111;
														assign node14882 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node14885 = (inp[7]) ? node14917 : node14886;
											assign node14886 = (inp[0]) ? node14902 : node14887;
												assign node14887 = (inp[11]) ? node14895 : node14888;
													assign node14888 = (inp[15]) ? node14892 : node14889;
														assign node14889 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node14892 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14895 = (inp[14]) ? node14899 : node14896;
														assign node14896 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14899 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14902 = (inp[15]) ? node14910 : node14903;
													assign node14903 = (inp[14]) ? node14907 : node14904;
														assign node14904 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14907 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14910 = (inp[9]) ? node14914 : node14911;
														assign node14911 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node14914 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node14917 = (inp[14]) ? node14931 : node14918;
												assign node14918 = (inp[9]) ? node14924 : node14919;
													assign node14919 = (inp[0]) ? node14921 : 16'b0000000001111111;
														assign node14921 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14924 = (inp[11]) ? node14928 : node14925;
														assign node14925 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14928 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node14931 = (inp[9]) ? node14939 : node14932;
													assign node14932 = (inp[15]) ? node14936 : node14933;
														assign node14933 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14936 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node14939 = (inp[15]) ? node14943 : node14940;
														assign node14940 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node14943 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node14946 = (inp[7]) ? node15008 : node14947;
										assign node14947 = (inp[0]) ? node14977 : node14948;
											assign node14948 = (inp[14]) ? node14964 : node14949;
												assign node14949 = (inp[15]) ? node14957 : node14950;
													assign node14950 = (inp[11]) ? node14954 : node14951;
														assign node14951 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node14954 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node14957 = (inp[9]) ? node14961 : node14958;
														assign node14958 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node14961 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node14964 = (inp[11]) ? node14972 : node14965;
													assign node14965 = (inp[3]) ? node14969 : node14966;
														assign node14966 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14969 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node14972 = (inp[15]) ? 16'b0000000000011111 : node14973;
														assign node14973 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node14977 = (inp[3]) ? node14993 : node14978;
												assign node14978 = (inp[9]) ? node14986 : node14979;
													assign node14979 = (inp[2]) ? node14983 : node14980;
														assign node14980 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node14983 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node14986 = (inp[15]) ? node14990 : node14987;
														assign node14987 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14990 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node14993 = (inp[14]) ? node15001 : node14994;
													assign node14994 = (inp[2]) ? node14998 : node14995;
														assign node14995 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node14998 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15001 = (inp[9]) ? node15005 : node15002;
														assign node15002 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15005 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node15008 = (inp[15]) ? node15040 : node15009;
											assign node15009 = (inp[11]) ? node15025 : node15010;
												assign node15010 = (inp[14]) ? node15018 : node15011;
													assign node15011 = (inp[3]) ? node15015 : node15012;
														assign node15012 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15015 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15018 = (inp[2]) ? node15022 : node15019;
														assign node15019 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15022 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15025 = (inp[2]) ? node15033 : node15026;
													assign node15026 = (inp[14]) ? node15030 : node15027;
														assign node15027 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15030 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15033 = (inp[0]) ? node15037 : node15034;
														assign node15034 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15037 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node15040 = (inp[2]) ? node15056 : node15041;
												assign node15041 = (inp[0]) ? node15049 : node15042;
													assign node15042 = (inp[11]) ? node15046 : node15043;
														assign node15043 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15046 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node15049 = (inp[14]) ? node15053 : node15050;
														assign node15050 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15053 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000001111;
												assign node15056 = (inp[11]) ? node15062 : node15057;
													assign node15057 = (inp[3]) ? node15059 : 16'b0000000000011111;
														assign node15059 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node15062 = (inp[3]) ? node15066 : node15063;
														assign node15063 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node15066 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node15069 = (inp[14]) ? node15313 : node15070;
								assign node15070 = (inp[0]) ? node15192 : node15071;
									assign node15071 = (inp[9]) ? node15133 : node15072;
										assign node15072 = (inp[3]) ? node15104 : node15073;
											assign node15073 = (inp[8]) ? node15089 : node15074;
												assign node15074 = (inp[11]) ? node15082 : node15075;
													assign node15075 = (inp[13]) ? node15079 : node15076;
														assign node15076 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15079 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15082 = (inp[2]) ? node15086 : node15083;
														assign node15083 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15086 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15089 = (inp[7]) ? node15097 : node15090;
													assign node15090 = (inp[13]) ? node15094 : node15091;
														assign node15091 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15094 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15097 = (inp[11]) ? node15101 : node15098;
														assign node15098 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15101 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node15104 = (inp[8]) ? node15118 : node15105;
												assign node15105 = (inp[11]) ? node15111 : node15106;
													assign node15106 = (inp[15]) ? node15108 : 16'b0000000111111111;
														assign node15108 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15111 = (inp[13]) ? node15115 : node15112;
														assign node15112 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15115 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15118 = (inp[13]) ? node15126 : node15119;
													assign node15119 = (inp[7]) ? node15123 : node15120;
														assign node15120 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node15123 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15126 = (inp[15]) ? node15130 : node15127;
														assign node15127 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node15130 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node15133 = (inp[11]) ? node15163 : node15134;
											assign node15134 = (inp[8]) ? node15150 : node15135;
												assign node15135 = (inp[13]) ? node15143 : node15136;
													assign node15136 = (inp[3]) ? node15140 : node15137;
														assign node15137 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15140 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15143 = (inp[7]) ? node15147 : node15144;
														assign node15144 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15147 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15150 = (inp[2]) ? node15156 : node15151;
													assign node15151 = (inp[3]) ? node15153 : 16'b0000000001111111;
														assign node15153 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15156 = (inp[15]) ? node15160 : node15157;
														assign node15157 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15160 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node15163 = (inp[2]) ? node15179 : node15164;
												assign node15164 = (inp[15]) ? node15172 : node15165;
													assign node15165 = (inp[7]) ? node15169 : node15166;
														assign node15166 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15169 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15172 = (inp[3]) ? node15176 : node15173;
														assign node15173 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15176 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15179 = (inp[7]) ? node15187 : node15180;
													assign node15180 = (inp[13]) ? node15184 : node15181;
														assign node15181 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15184 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15187 = (inp[15]) ? node15189 : 16'b0000000000011111;
														assign node15189 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node15192 = (inp[15]) ? node15254 : node15193;
										assign node15193 = (inp[7]) ? node15223 : node15194;
											assign node15194 = (inp[13]) ? node15208 : node15195;
												assign node15195 = (inp[9]) ? node15201 : node15196;
													assign node15196 = (inp[8]) ? node15198 : 16'b0000000111111111;
														assign node15198 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15201 = (inp[11]) ? node15205 : node15202;
														assign node15202 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15205 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15208 = (inp[8]) ? node15216 : node15209;
													assign node15209 = (inp[11]) ? node15213 : node15210;
														assign node15210 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15213 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15216 = (inp[3]) ? node15220 : node15217;
														assign node15217 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15220 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node15223 = (inp[2]) ? node15239 : node15224;
												assign node15224 = (inp[11]) ? node15232 : node15225;
													assign node15225 = (inp[8]) ? node15229 : node15226;
														assign node15226 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node15229 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node15232 = (inp[9]) ? node15236 : node15233;
														assign node15233 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15236 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15239 = (inp[3]) ? node15247 : node15240;
													assign node15240 = (inp[8]) ? node15244 : node15241;
														assign node15241 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15244 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15247 = (inp[9]) ? node15251 : node15248;
														assign node15248 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node15251 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node15254 = (inp[3]) ? node15284 : node15255;
											assign node15255 = (inp[13]) ? node15269 : node15256;
												assign node15256 = (inp[11]) ? node15262 : node15257;
													assign node15257 = (inp[2]) ? node15259 : 16'b0000000011111111;
														assign node15259 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15262 = (inp[2]) ? node15266 : node15263;
														assign node15263 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15266 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node15269 = (inp[7]) ? node15277 : node15270;
													assign node15270 = (inp[9]) ? node15274 : node15271;
														assign node15271 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15274 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15277 = (inp[9]) ? node15281 : node15278;
														assign node15278 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15281 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node15284 = (inp[2]) ? node15300 : node15285;
												assign node15285 = (inp[8]) ? node15293 : node15286;
													assign node15286 = (inp[13]) ? node15290 : node15287;
														assign node15287 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node15290 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node15293 = (inp[13]) ? node15297 : node15294;
														assign node15294 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15297 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node15300 = (inp[11]) ? node15306 : node15301;
													assign node15301 = (inp[9]) ? node15303 : 16'b0000000000011111;
														assign node15303 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node15306 = (inp[8]) ? node15310 : node15307;
														assign node15307 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node15310 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node15313 = (inp[3]) ? node15439 : node15314;
									assign node15314 = (inp[2]) ? node15378 : node15315;
										assign node15315 = (inp[7]) ? node15347 : node15316;
											assign node15316 = (inp[8]) ? node15332 : node15317;
												assign node15317 = (inp[9]) ? node15325 : node15318;
													assign node15318 = (inp[13]) ? node15322 : node15319;
														assign node15319 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node15322 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node15325 = (inp[11]) ? node15329 : node15326;
														assign node15326 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node15329 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node15332 = (inp[9]) ? node15340 : node15333;
													assign node15333 = (inp[15]) ? node15337 : node15334;
														assign node15334 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15337 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15340 = (inp[0]) ? node15344 : node15341;
														assign node15341 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15344 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node15347 = (inp[0]) ? node15363 : node15348;
												assign node15348 = (inp[15]) ? node15356 : node15349;
													assign node15349 = (inp[13]) ? node15353 : node15350;
														assign node15350 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node15353 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15356 = (inp[9]) ? node15360 : node15357;
														assign node15357 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15360 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15363 = (inp[15]) ? node15371 : node15364;
													assign node15364 = (inp[13]) ? node15368 : node15365;
														assign node15365 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15368 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15371 = (inp[9]) ? node15375 : node15372;
														assign node15372 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node15375 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node15378 = (inp[9]) ? node15408 : node15379;
											assign node15379 = (inp[7]) ? node15395 : node15380;
												assign node15380 = (inp[0]) ? node15388 : node15381;
													assign node15381 = (inp[13]) ? node15385 : node15382;
														assign node15382 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node15385 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15388 = (inp[13]) ? node15392 : node15389;
														assign node15389 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node15392 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15395 = (inp[15]) ? node15401 : node15396;
													assign node15396 = (inp[13]) ? node15398 : 16'b0000000000111111;
														assign node15398 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15401 = (inp[8]) ? node15405 : node15402;
														assign node15402 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15405 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node15408 = (inp[8]) ? node15424 : node15409;
												assign node15409 = (inp[11]) ? node15417 : node15410;
													assign node15410 = (inp[13]) ? node15414 : node15411;
														assign node15411 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15414 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15417 = (inp[7]) ? node15421 : node15418;
														assign node15418 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15421 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node15424 = (inp[11]) ? node15432 : node15425;
													assign node15425 = (inp[0]) ? node15429 : node15426;
														assign node15426 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15429 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node15432 = (inp[13]) ? node15436 : node15433;
														assign node15433 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node15436 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node15439 = (inp[8]) ? node15503 : node15440;
										assign node15440 = (inp[15]) ? node15472 : node15441;
											assign node15441 = (inp[2]) ? node15457 : node15442;
												assign node15442 = (inp[11]) ? node15450 : node15443;
													assign node15443 = (inp[9]) ? node15447 : node15444;
														assign node15444 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node15447 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node15450 = (inp[13]) ? node15454 : node15451;
														assign node15451 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15454 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node15457 = (inp[0]) ? node15465 : node15458;
													assign node15458 = (inp[11]) ? node15462 : node15459;
														assign node15459 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15462 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15465 = (inp[9]) ? node15469 : node15466;
														assign node15466 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15469 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node15472 = (inp[11]) ? node15488 : node15473;
												assign node15473 = (inp[0]) ? node15481 : node15474;
													assign node15474 = (inp[9]) ? node15478 : node15475;
														assign node15475 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node15478 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000011111;
													assign node15481 = (inp[13]) ? node15485 : node15482;
														assign node15482 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15485 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node15488 = (inp[13]) ? node15496 : node15489;
													assign node15489 = (inp[9]) ? node15493 : node15490;
														assign node15490 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15493 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node15496 = (inp[2]) ? node15500 : node15497;
														assign node15497 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node15500 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node15503 = (inp[7]) ? node15531 : node15504;
											assign node15504 = (inp[13]) ? node15518 : node15505;
												assign node15505 = (inp[9]) ? node15511 : node15506;
													assign node15506 = (inp[0]) ? node15508 : 16'b0000000000111111;
														assign node15508 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node15511 = (inp[15]) ? node15515 : node15512;
														assign node15512 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15515 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node15518 = (inp[11]) ? node15526 : node15519;
													assign node15519 = (inp[2]) ? node15523 : node15520;
														assign node15520 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node15523 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node15526 = (inp[15]) ? node15528 : 16'b0000000000001111;
														assign node15528 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000000111;
											assign node15531 = (inp[2]) ? node15545 : node15532;
												assign node15532 = (inp[0]) ? node15538 : node15533;
													assign node15533 = (inp[9]) ? node15535 : 16'b0000000000011111;
														assign node15535 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node15538 = (inp[9]) ? node15542 : node15539;
														assign node15539 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node15542 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node15545 = (inp[15]) ? node15553 : node15546;
													assign node15546 = (inp[9]) ? node15550 : node15547;
														assign node15547 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node15550 = (inp[13]) ? 16'b0000000000000011 : 16'b0000000000001111;
													assign node15553 = (inp[9]) ? node15555 : 16'b0000000000000111;
														assign node15555 = (inp[0]) ? 16'b0000000000000011 : 16'b0000000000000111;
		assign node15558 = (inp[10]) ? node23388 : node15559;
			assign node15559 = (inp[12]) ? node19479 : node15560;
				assign node15560 = (inp[13]) ? node17506 : node15561;
					assign node15561 = (inp[11]) ? node16537 : node15562;
						assign node15562 = (inp[8]) ? node16050 : node15563;
							assign node15563 = (inp[9]) ? node15803 : node15564;
								assign node15564 = (inp[5]) ? node15682 : node15565;
									assign node15565 = (inp[15]) ? node15623 : node15566;
										assign node15566 = (inp[2]) ? node15596 : node15567;
											assign node15567 = (inp[7]) ? node15583 : node15568;
												assign node15568 = (inp[14]) ? node15576 : node15569;
													assign node15569 = (inp[0]) ? node15573 : node15570;
														assign node15570 = (inp[1]) ? 16'b0001111111111111 : 16'b0011111111111111;
														assign node15573 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node15576 = (inp[3]) ? node15580 : node15577;
														assign node15577 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node15580 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
												assign node15583 = (inp[3]) ? node15591 : node15584;
													assign node15584 = (inp[4]) ? node15588 : node15585;
														assign node15585 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node15588 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node15591 = (inp[0]) ? 16'b0000011111111111 : node15592;
														assign node15592 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
											assign node15596 = (inp[0]) ? node15610 : node15597;
												assign node15597 = (inp[3]) ? node15603 : node15598;
													assign node15598 = (inp[7]) ? 16'b0000111111111111 : node15599;
														assign node15599 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node15603 = (inp[14]) ? node15607 : node15604;
														assign node15604 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15607 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node15610 = (inp[7]) ? node15618 : node15611;
													assign node15611 = (inp[1]) ? node15615 : node15612;
														assign node15612 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15615 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15618 = (inp[3]) ? 16'b0000000111111111 : node15619;
														assign node15619 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
										assign node15623 = (inp[14]) ? node15653 : node15624;
											assign node15624 = (inp[4]) ? node15638 : node15625;
												assign node15625 = (inp[2]) ? node15631 : node15626;
													assign node15626 = (inp[0]) ? 16'b0000111111111111 : node15627;
														assign node15627 = (inp[7]) ? 16'b0000111111111111 : 16'b0001111111111111;
													assign node15631 = (inp[0]) ? node15635 : node15632;
														assign node15632 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15635 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node15638 = (inp[0]) ? node15646 : node15639;
													assign node15639 = (inp[3]) ? node15643 : node15640;
														assign node15640 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15643 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15646 = (inp[1]) ? node15650 : node15647;
														assign node15647 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15650 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node15653 = (inp[3]) ? node15667 : node15654;
												assign node15654 = (inp[0]) ? node15660 : node15655;
													assign node15655 = (inp[4]) ? node15657 : 16'b0000111111111111;
														assign node15657 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15660 = (inp[4]) ? node15664 : node15661;
														assign node15661 = (inp[2]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node15664 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15667 = (inp[0]) ? node15675 : node15668;
													assign node15668 = (inp[1]) ? node15672 : node15669;
														assign node15669 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15672 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15675 = (inp[7]) ? node15679 : node15676;
														assign node15676 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15679 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
									assign node15682 = (inp[3]) ? node15742 : node15683;
										assign node15683 = (inp[7]) ? node15715 : node15684;
											assign node15684 = (inp[1]) ? node15700 : node15685;
												assign node15685 = (inp[15]) ? node15693 : node15686;
													assign node15686 = (inp[2]) ? node15690 : node15687;
														assign node15687 = (inp[4]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node15690 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node15693 = (inp[2]) ? node15697 : node15694;
														assign node15694 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15697 = (inp[0]) ? 16'b0000001111111111 : 16'b0000001111111111;
												assign node15700 = (inp[4]) ? node15708 : node15701;
													assign node15701 = (inp[14]) ? node15705 : node15702;
														assign node15702 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15705 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15708 = (inp[0]) ? node15712 : node15709;
														assign node15709 = (inp[14]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node15712 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node15715 = (inp[4]) ? node15729 : node15716;
												assign node15716 = (inp[0]) ? node15722 : node15717;
													assign node15717 = (inp[15]) ? 16'b0000001111111111 : node15718;
														assign node15718 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node15722 = (inp[1]) ? node15726 : node15723;
														assign node15723 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15726 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15729 = (inp[14]) ? node15735 : node15730;
													assign node15730 = (inp[15]) ? node15732 : 16'b0000001111111111;
														assign node15732 = (inp[1]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node15735 = (inp[15]) ? node15739 : node15736;
														assign node15736 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node15739 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node15742 = (inp[4]) ? node15774 : node15743;
											assign node15743 = (inp[2]) ? node15759 : node15744;
												assign node15744 = (inp[0]) ? node15752 : node15745;
													assign node15745 = (inp[7]) ? node15749 : node15746;
														assign node15746 = (inp[1]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node15749 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15752 = (inp[7]) ? node15756 : node15753;
														assign node15753 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15756 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15759 = (inp[15]) ? node15767 : node15760;
													assign node15760 = (inp[7]) ? node15764 : node15761;
														assign node15761 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15764 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15767 = (inp[14]) ? node15771 : node15768;
														assign node15768 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node15771 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node15774 = (inp[7]) ? node15790 : node15775;
												assign node15775 = (inp[0]) ? node15783 : node15776;
													assign node15776 = (inp[2]) ? node15780 : node15777;
														assign node15777 = (inp[14]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node15780 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15783 = (inp[15]) ? node15787 : node15784;
														assign node15784 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15787 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15790 = (inp[15]) ? node15798 : node15791;
													assign node15791 = (inp[14]) ? node15795 : node15792;
														assign node15792 = (inp[1]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node15795 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15798 = (inp[1]) ? node15800 : 16'b0000000011111111;
														assign node15800 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node15803 = (inp[1]) ? node15927 : node15804;
									assign node15804 = (inp[0]) ? node15864 : node15805;
										assign node15805 = (inp[3]) ? node15835 : node15806;
											assign node15806 = (inp[14]) ? node15820 : node15807;
												assign node15807 = (inp[5]) ? node15813 : node15808;
													assign node15808 = (inp[15]) ? node15810 : 16'b0001111111111111;
														assign node15810 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node15813 = (inp[15]) ? node15817 : node15814;
														assign node15814 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15817 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node15820 = (inp[7]) ? node15828 : node15821;
													assign node15821 = (inp[15]) ? node15825 : node15822;
														assign node15822 = (inp[4]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15825 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15828 = (inp[5]) ? node15832 : node15829;
														assign node15829 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15832 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node15835 = (inp[15]) ? node15851 : node15836;
												assign node15836 = (inp[14]) ? node15844 : node15837;
													assign node15837 = (inp[5]) ? node15841 : node15838;
														assign node15838 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15841 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15844 = (inp[2]) ? node15848 : node15845;
														assign node15845 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15848 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15851 = (inp[2]) ? node15859 : node15852;
													assign node15852 = (inp[14]) ? node15856 : node15853;
														assign node15853 = (inp[4]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node15856 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15859 = (inp[7]) ? 16'b0000000111111111 : node15860;
														assign node15860 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
										assign node15864 = (inp[3]) ? node15896 : node15865;
											assign node15865 = (inp[2]) ? node15881 : node15866;
												assign node15866 = (inp[4]) ? node15874 : node15867;
													assign node15867 = (inp[14]) ? node15871 : node15868;
														assign node15868 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15871 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node15874 = (inp[15]) ? node15878 : node15875;
														assign node15875 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15878 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15881 = (inp[5]) ? node15889 : node15882;
													assign node15882 = (inp[7]) ? node15886 : node15883;
														assign node15883 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15886 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15889 = (inp[14]) ? node15893 : node15890;
														assign node15890 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15893 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node15896 = (inp[4]) ? node15912 : node15897;
												assign node15897 = (inp[14]) ? node15905 : node15898;
													assign node15898 = (inp[2]) ? node15902 : node15899;
														assign node15899 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15902 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15905 = (inp[2]) ? node15909 : node15906;
														assign node15906 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15909 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15912 = (inp[5]) ? node15920 : node15913;
													assign node15913 = (inp[14]) ? node15917 : node15914;
														assign node15914 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node15917 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15920 = (inp[14]) ? node15924 : node15921;
														assign node15921 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node15924 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node15927 = (inp[2]) ? node15991 : node15928;
										assign node15928 = (inp[15]) ? node15960 : node15929;
											assign node15929 = (inp[7]) ? node15945 : node15930;
												assign node15930 = (inp[5]) ? node15938 : node15931;
													assign node15931 = (inp[3]) ? node15935 : node15932;
														assign node15932 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node15935 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node15938 = (inp[4]) ? node15942 : node15939;
														assign node15939 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15942 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node15945 = (inp[5]) ? node15953 : node15946;
													assign node15946 = (inp[0]) ? node15950 : node15947;
														assign node15947 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15950 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15953 = (inp[4]) ? node15957 : node15954;
														assign node15954 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15957 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node15960 = (inp[3]) ? node15976 : node15961;
												assign node15961 = (inp[5]) ? node15969 : node15962;
													assign node15962 = (inp[0]) ? node15966 : node15963;
														assign node15963 = (inp[4]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node15966 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node15969 = (inp[0]) ? node15973 : node15970;
														assign node15970 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node15973 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node15976 = (inp[5]) ? node15984 : node15977;
													assign node15977 = (inp[4]) ? node15981 : node15978;
														assign node15978 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node15981 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node15984 = (inp[4]) ? node15988 : node15985;
														assign node15985 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node15988 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node15991 = (inp[7]) ? node16019 : node15992;
											assign node15992 = (inp[5]) ? node16006 : node15993;
												assign node15993 = (inp[14]) ? node16001 : node15994;
													assign node15994 = (inp[0]) ? node15998 : node15995;
														assign node15995 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node15998 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16001 = (inp[15]) ? node16003 : 16'b0000001111111111;
														assign node16003 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16006 = (inp[4]) ? node16014 : node16007;
													assign node16007 = (inp[15]) ? node16011 : node16008;
														assign node16008 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16011 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16014 = (inp[14]) ? 16'b0000000011111111 : node16015;
														assign node16015 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16019 = (inp[0]) ? node16035 : node16020;
												assign node16020 = (inp[15]) ? node16028 : node16021;
													assign node16021 = (inp[4]) ? node16025 : node16022;
														assign node16022 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16025 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16028 = (inp[3]) ? node16032 : node16029;
														assign node16029 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16032 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16035 = (inp[4]) ? node16043 : node16036;
													assign node16036 = (inp[5]) ? node16040 : node16037;
														assign node16037 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16040 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16043 = (inp[14]) ? node16047 : node16044;
														assign node16044 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16047 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
							assign node16050 = (inp[1]) ? node16294 : node16051;
								assign node16051 = (inp[7]) ? node16175 : node16052;
									assign node16052 = (inp[15]) ? node16114 : node16053;
										assign node16053 = (inp[14]) ? node16083 : node16054;
											assign node16054 = (inp[4]) ? node16070 : node16055;
												assign node16055 = (inp[5]) ? node16063 : node16056;
													assign node16056 = (inp[3]) ? node16060 : node16057;
														assign node16057 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node16060 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node16063 = (inp[0]) ? node16067 : node16064;
														assign node16064 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16067 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16070 = (inp[9]) ? node16078 : node16071;
													assign node16071 = (inp[0]) ? node16075 : node16072;
														assign node16072 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16075 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16078 = (inp[0]) ? 16'b0000000111111111 : node16079;
														assign node16079 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node16083 = (inp[3]) ? node16099 : node16084;
												assign node16084 = (inp[4]) ? node16092 : node16085;
													assign node16085 = (inp[0]) ? node16089 : node16086;
														assign node16086 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16089 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16092 = (inp[9]) ? node16096 : node16093;
														assign node16093 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16096 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16099 = (inp[4]) ? node16107 : node16100;
													assign node16100 = (inp[0]) ? node16104 : node16101;
														assign node16101 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16104 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16107 = (inp[0]) ? node16111 : node16108;
														assign node16108 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16111 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node16114 = (inp[2]) ? node16146 : node16115;
											assign node16115 = (inp[14]) ? node16131 : node16116;
												assign node16116 = (inp[0]) ? node16124 : node16117;
													assign node16117 = (inp[5]) ? node16121 : node16118;
														assign node16118 = (inp[9]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16121 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16124 = (inp[9]) ? node16128 : node16125;
														assign node16125 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16128 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node16131 = (inp[3]) ? node16139 : node16132;
													assign node16132 = (inp[5]) ? node16136 : node16133;
														assign node16133 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16136 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16139 = (inp[5]) ? node16143 : node16140;
														assign node16140 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16143 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16146 = (inp[0]) ? node16162 : node16147;
												assign node16147 = (inp[3]) ? node16155 : node16148;
													assign node16148 = (inp[9]) ? node16152 : node16149;
														assign node16149 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16152 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16155 = (inp[4]) ? node16159 : node16156;
														assign node16156 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16159 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16162 = (inp[14]) ? node16168 : node16163;
													assign node16163 = (inp[9]) ? node16165 : 16'b0000000111111111;
														assign node16165 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16168 = (inp[3]) ? node16172 : node16169;
														assign node16169 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16172 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node16175 = (inp[3]) ? node16235 : node16176;
										assign node16176 = (inp[14]) ? node16206 : node16177;
											assign node16177 = (inp[0]) ? node16193 : node16178;
												assign node16178 = (inp[2]) ? node16186 : node16179;
													assign node16179 = (inp[4]) ? node16183 : node16180;
														assign node16180 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16183 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16186 = (inp[5]) ? node16190 : node16187;
														assign node16187 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16190 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16193 = (inp[15]) ? node16201 : node16194;
													assign node16194 = (inp[5]) ? node16198 : node16195;
														assign node16195 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16198 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16201 = (inp[5]) ? 16'b0000000011111111 : node16202;
														assign node16202 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node16206 = (inp[4]) ? node16222 : node16207;
												assign node16207 = (inp[5]) ? node16215 : node16208;
													assign node16208 = (inp[0]) ? node16212 : node16209;
														assign node16209 = (inp[15]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node16212 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16215 = (inp[2]) ? node16219 : node16216;
														assign node16216 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node16219 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16222 = (inp[0]) ? node16228 : node16223;
													assign node16223 = (inp[15]) ? 16'b0000000011111111 : node16224;
														assign node16224 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16228 = (inp[5]) ? node16232 : node16229;
														assign node16229 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16232 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node16235 = (inp[9]) ? node16267 : node16236;
											assign node16236 = (inp[14]) ? node16252 : node16237;
												assign node16237 = (inp[5]) ? node16245 : node16238;
													assign node16238 = (inp[0]) ? node16242 : node16239;
														assign node16239 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16242 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16245 = (inp[4]) ? node16249 : node16246;
														assign node16246 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16249 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16252 = (inp[4]) ? node16260 : node16253;
													assign node16253 = (inp[0]) ? node16257 : node16254;
														assign node16254 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node16257 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node16260 = (inp[5]) ? node16264 : node16261;
														assign node16261 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16264 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node16267 = (inp[2]) ? node16281 : node16268;
												assign node16268 = (inp[14]) ? node16276 : node16269;
													assign node16269 = (inp[4]) ? node16273 : node16270;
														assign node16270 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16273 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16276 = (inp[0]) ? 16'b0000000011111111 : node16277;
														assign node16277 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16281 = (inp[15]) ? node16287 : node16282;
													assign node16282 = (inp[4]) ? node16284 : 16'b0000000111111111;
														assign node16284 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16287 = (inp[4]) ? node16291 : node16288;
														assign node16288 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16291 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node16294 = (inp[0]) ? node16416 : node16295;
									assign node16295 = (inp[14]) ? node16355 : node16296;
										assign node16296 = (inp[15]) ? node16326 : node16297;
											assign node16297 = (inp[4]) ? node16311 : node16298;
												assign node16298 = (inp[5]) ? node16306 : node16299;
													assign node16299 = (inp[7]) ? node16303 : node16300;
														assign node16300 = (inp[9]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node16303 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16306 = (inp[2]) ? 16'b0000001111111111 : node16307;
														assign node16307 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16311 = (inp[5]) ? node16319 : node16312;
													assign node16312 = (inp[7]) ? node16316 : node16313;
														assign node16313 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16316 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16319 = (inp[9]) ? node16323 : node16320;
														assign node16320 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16323 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16326 = (inp[2]) ? node16340 : node16327;
												assign node16327 = (inp[7]) ? node16335 : node16328;
													assign node16328 = (inp[5]) ? node16332 : node16329;
														assign node16329 = (inp[4]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node16332 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16335 = (inp[4]) ? 16'b0000000011111111 : node16336;
														assign node16336 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16340 = (inp[3]) ? node16348 : node16341;
													assign node16341 = (inp[5]) ? node16345 : node16342;
														assign node16342 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16345 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16348 = (inp[7]) ? node16352 : node16349;
														assign node16349 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node16352 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node16355 = (inp[4]) ? node16385 : node16356;
											assign node16356 = (inp[9]) ? node16370 : node16357;
												assign node16357 = (inp[2]) ? node16365 : node16358;
													assign node16358 = (inp[5]) ? node16362 : node16359;
														assign node16359 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16362 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node16365 = (inp[15]) ? 16'b0000000111111111 : node16366;
														assign node16366 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16370 = (inp[2]) ? node16378 : node16371;
													assign node16371 = (inp[3]) ? node16375 : node16372;
														assign node16372 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16375 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16378 = (inp[15]) ? node16382 : node16379;
														assign node16379 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16382 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node16385 = (inp[3]) ? node16401 : node16386;
												assign node16386 = (inp[9]) ? node16394 : node16387;
													assign node16387 = (inp[7]) ? node16391 : node16388;
														assign node16388 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16391 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16394 = (inp[2]) ? node16398 : node16395;
														assign node16395 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16398 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node16401 = (inp[7]) ? node16409 : node16402;
													assign node16402 = (inp[9]) ? node16406 : node16403;
														assign node16403 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16406 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16409 = (inp[5]) ? node16413 : node16410;
														assign node16410 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16413 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node16416 = (inp[7]) ? node16478 : node16417;
										assign node16417 = (inp[9]) ? node16447 : node16418;
											assign node16418 = (inp[14]) ? node16434 : node16419;
												assign node16419 = (inp[15]) ? node16427 : node16420;
													assign node16420 = (inp[5]) ? node16424 : node16421;
														assign node16421 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16424 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16427 = (inp[2]) ? node16431 : node16428;
														assign node16428 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16431 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16434 = (inp[15]) ? node16442 : node16435;
													assign node16435 = (inp[4]) ? node16439 : node16436;
														assign node16436 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16439 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16442 = (inp[5]) ? 16'b0000000011111111 : node16443;
														assign node16443 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node16447 = (inp[15]) ? node16463 : node16448;
												assign node16448 = (inp[5]) ? node16456 : node16449;
													assign node16449 = (inp[4]) ? node16453 : node16450;
														assign node16450 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node16453 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16456 = (inp[14]) ? node16460 : node16457;
														assign node16457 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16460 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node16463 = (inp[2]) ? node16471 : node16464;
													assign node16464 = (inp[4]) ? node16468 : node16465;
														assign node16465 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node16468 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16471 = (inp[4]) ? node16475 : node16472;
														assign node16472 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node16475 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node16478 = (inp[5]) ? node16506 : node16479;
											assign node16479 = (inp[14]) ? node16491 : node16480;
												assign node16480 = (inp[2]) ? node16486 : node16481;
													assign node16481 = (inp[4]) ? 16'b0000000111111111 : node16482;
														assign node16482 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16486 = (inp[15]) ? 16'b0000000011111111 : node16487;
														assign node16487 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16491 = (inp[2]) ? node16499 : node16492;
													assign node16492 = (inp[9]) ? node16496 : node16493;
														assign node16493 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16496 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16499 = (inp[3]) ? node16503 : node16500;
														assign node16500 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16503 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node16506 = (inp[15]) ? node16522 : node16507;
												assign node16507 = (inp[3]) ? node16515 : node16508;
													assign node16508 = (inp[2]) ? node16512 : node16509;
														assign node16509 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node16512 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16515 = (inp[14]) ? node16519 : node16516;
														assign node16516 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16519 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node16522 = (inp[2]) ? node16530 : node16523;
													assign node16523 = (inp[14]) ? node16527 : node16524;
														assign node16524 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16527 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node16530 = (inp[4]) ? node16534 : node16531;
														assign node16531 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node16534 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
						assign node16537 = (inp[4]) ? node17025 : node16538;
							assign node16538 = (inp[5]) ? node16780 : node16539;
								assign node16539 = (inp[7]) ? node16661 : node16540;
									assign node16540 = (inp[3]) ? node16600 : node16541;
										assign node16541 = (inp[9]) ? node16571 : node16542;
											assign node16542 = (inp[14]) ? node16558 : node16543;
												assign node16543 = (inp[15]) ? node16551 : node16544;
													assign node16544 = (inp[2]) ? node16548 : node16545;
														assign node16545 = (inp[0]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node16548 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node16551 = (inp[1]) ? node16555 : node16552;
														assign node16552 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16555 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node16558 = (inp[15]) ? node16564 : node16559;
													assign node16559 = (inp[1]) ? 16'b0000011111111111 : node16560;
														assign node16560 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node16564 = (inp[2]) ? node16568 : node16565;
														assign node16565 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16568 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
											assign node16571 = (inp[0]) ? node16587 : node16572;
												assign node16572 = (inp[2]) ? node16580 : node16573;
													assign node16573 = (inp[8]) ? node16577 : node16574;
														assign node16574 = (inp[1]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node16577 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16580 = (inp[14]) ? node16584 : node16581;
														assign node16581 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16584 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16587 = (inp[2]) ? node16595 : node16588;
													assign node16588 = (inp[14]) ? node16592 : node16589;
														assign node16589 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16592 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16595 = (inp[8]) ? node16597 : 16'b0000000111111111;
														assign node16597 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node16600 = (inp[15]) ? node16632 : node16601;
											assign node16601 = (inp[14]) ? node16617 : node16602;
												assign node16602 = (inp[2]) ? node16610 : node16603;
													assign node16603 = (inp[1]) ? node16607 : node16604;
														assign node16604 = (inp[8]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node16607 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16610 = (inp[8]) ? node16614 : node16611;
														assign node16611 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16614 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16617 = (inp[1]) ? node16625 : node16618;
													assign node16618 = (inp[8]) ? node16622 : node16619;
														assign node16619 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16622 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16625 = (inp[2]) ? node16629 : node16626;
														assign node16626 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16629 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16632 = (inp[2]) ? node16648 : node16633;
												assign node16633 = (inp[8]) ? node16641 : node16634;
													assign node16634 = (inp[9]) ? node16638 : node16635;
														assign node16635 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16638 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16641 = (inp[1]) ? node16645 : node16642;
														assign node16642 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16645 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16648 = (inp[8]) ? node16656 : node16649;
													assign node16649 = (inp[1]) ? node16653 : node16650;
														assign node16650 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16653 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16656 = (inp[9]) ? 16'b0000000011111111 : node16657;
														assign node16657 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node16661 = (inp[14]) ? node16721 : node16662;
										assign node16662 = (inp[9]) ? node16692 : node16663;
											assign node16663 = (inp[1]) ? node16677 : node16664;
												assign node16664 = (inp[8]) ? node16670 : node16665;
													assign node16665 = (inp[15]) ? 16'b0000011111111111 : node16666;
														assign node16666 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node16670 = (inp[3]) ? node16674 : node16671;
														assign node16671 = (inp[0]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node16674 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16677 = (inp[15]) ? node16685 : node16678;
													assign node16678 = (inp[0]) ? node16682 : node16679;
														assign node16679 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16682 = (inp[3]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node16685 = (inp[8]) ? node16689 : node16686;
														assign node16686 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16689 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16692 = (inp[8]) ? node16708 : node16693;
												assign node16693 = (inp[15]) ? node16701 : node16694;
													assign node16694 = (inp[1]) ? node16698 : node16695;
														assign node16695 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16698 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16701 = (inp[3]) ? node16705 : node16702;
														assign node16702 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node16705 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16708 = (inp[0]) ? node16716 : node16709;
													assign node16709 = (inp[2]) ? node16713 : node16710;
														assign node16710 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16713 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16716 = (inp[1]) ? node16718 : 16'b0000000011111111;
														assign node16718 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node16721 = (inp[15]) ? node16751 : node16722;
											assign node16722 = (inp[1]) ? node16738 : node16723;
												assign node16723 = (inp[2]) ? node16731 : node16724;
													assign node16724 = (inp[0]) ? node16728 : node16725;
														assign node16725 = (inp[3]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node16728 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16731 = (inp[0]) ? node16735 : node16732;
														assign node16732 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16735 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node16738 = (inp[9]) ? node16744 : node16739;
													assign node16739 = (inp[0]) ? node16741 : 16'b0000000111111111;
														assign node16741 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16744 = (inp[3]) ? node16748 : node16745;
														assign node16745 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16748 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node16751 = (inp[0]) ? node16765 : node16752;
												assign node16752 = (inp[3]) ? node16758 : node16753;
													assign node16753 = (inp[1]) ? 16'b0000001111111111 : node16754;
														assign node16754 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node16758 = (inp[1]) ? node16762 : node16759;
														assign node16759 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16762 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node16765 = (inp[2]) ? node16773 : node16766;
													assign node16766 = (inp[8]) ? node16770 : node16767;
														assign node16767 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16770 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16773 = (inp[9]) ? node16777 : node16774;
														assign node16774 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16777 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node16780 = (inp[15]) ? node16904 : node16781;
									assign node16781 = (inp[9]) ? node16845 : node16782;
										assign node16782 = (inp[8]) ? node16814 : node16783;
											assign node16783 = (inp[14]) ? node16799 : node16784;
												assign node16784 = (inp[3]) ? node16792 : node16785;
													assign node16785 = (inp[2]) ? node16789 : node16786;
														assign node16786 = (inp[0]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node16789 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node16792 = (inp[2]) ? node16796 : node16793;
														assign node16793 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16796 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node16799 = (inp[0]) ? node16807 : node16800;
													assign node16800 = (inp[1]) ? node16804 : node16801;
														assign node16801 = (inp[7]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node16804 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16807 = (inp[3]) ? node16811 : node16808;
														assign node16808 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node16811 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16814 = (inp[1]) ? node16830 : node16815;
												assign node16815 = (inp[3]) ? node16823 : node16816;
													assign node16816 = (inp[14]) ? node16820 : node16817;
														assign node16817 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16820 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16823 = (inp[2]) ? node16827 : node16824;
														assign node16824 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16827 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16830 = (inp[0]) ? node16838 : node16831;
													assign node16831 = (inp[14]) ? node16835 : node16832;
														assign node16832 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16835 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16838 = (inp[3]) ? node16842 : node16839;
														assign node16839 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16842 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node16845 = (inp[7]) ? node16877 : node16846;
											assign node16846 = (inp[2]) ? node16862 : node16847;
												assign node16847 = (inp[0]) ? node16855 : node16848;
													assign node16848 = (inp[3]) ? node16852 : node16849;
														assign node16849 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node16852 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16855 = (inp[1]) ? node16859 : node16856;
														assign node16856 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16859 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16862 = (inp[8]) ? node16870 : node16863;
													assign node16863 = (inp[0]) ? node16867 : node16864;
														assign node16864 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node16867 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16870 = (inp[1]) ? node16874 : node16871;
														assign node16871 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16874 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node16877 = (inp[2]) ? node16891 : node16878;
												assign node16878 = (inp[8]) ? node16886 : node16879;
													assign node16879 = (inp[0]) ? node16883 : node16880;
														assign node16880 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node16883 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16886 = (inp[3]) ? 16'b0000000001111111 : node16887;
														assign node16887 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node16891 = (inp[1]) ? node16899 : node16892;
													assign node16892 = (inp[14]) ? node16896 : node16893;
														assign node16893 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node16896 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16899 = (inp[14]) ? node16901 : 16'b0000000001111111;
														assign node16901 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node16904 = (inp[9]) ? node16964 : node16905;
										assign node16905 = (inp[14]) ? node16935 : node16906;
											assign node16906 = (inp[2]) ? node16922 : node16907;
												assign node16907 = (inp[3]) ? node16915 : node16908;
													assign node16908 = (inp[7]) ? node16912 : node16909;
														assign node16909 = (inp[0]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node16912 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node16915 = (inp[8]) ? node16919 : node16916;
														assign node16916 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16919 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node16922 = (inp[8]) ? node16930 : node16923;
													assign node16923 = (inp[3]) ? node16927 : node16924;
														assign node16924 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16927 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16930 = (inp[7]) ? 16'b0000000011111111 : node16931;
														assign node16931 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node16935 = (inp[0]) ? node16949 : node16936;
												assign node16936 = (inp[2]) ? node16942 : node16937;
													assign node16937 = (inp[1]) ? node16939 : 16'b0000000111111111;
														assign node16939 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16942 = (inp[3]) ? node16946 : node16943;
														assign node16943 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node16946 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16949 = (inp[3]) ? node16957 : node16950;
													assign node16950 = (inp[8]) ? node16954 : node16951;
														assign node16951 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16954 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16957 = (inp[2]) ? node16961 : node16958;
														assign node16958 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node16961 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node16964 = (inp[1]) ? node16996 : node16965;
											assign node16965 = (inp[8]) ? node16981 : node16966;
												assign node16966 = (inp[7]) ? node16974 : node16967;
													assign node16967 = (inp[14]) ? node16971 : node16968;
														assign node16968 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node16971 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node16974 = (inp[14]) ? node16978 : node16975;
														assign node16975 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node16978 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node16981 = (inp[2]) ? node16989 : node16982;
													assign node16982 = (inp[7]) ? node16986 : node16983;
														assign node16983 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node16986 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node16989 = (inp[3]) ? node16993 : node16990;
														assign node16990 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node16993 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node16996 = (inp[3]) ? node17012 : node16997;
												assign node16997 = (inp[0]) ? node17005 : node16998;
													assign node16998 = (inp[14]) ? node17002 : node16999;
														assign node16999 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17002 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17005 = (inp[2]) ? node17009 : node17006;
														assign node17006 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17009 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node17012 = (inp[7]) ? node17020 : node17013;
													assign node17013 = (inp[0]) ? node17017 : node17014;
														assign node17014 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17017 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17020 = (inp[8]) ? node17022 : 16'b0000000001111111;
														assign node17022 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node17025 = (inp[3]) ? node17271 : node17026;
								assign node17026 = (inp[14]) ? node17148 : node17027;
									assign node17027 = (inp[7]) ? node17091 : node17028;
										assign node17028 = (inp[15]) ? node17060 : node17029;
											assign node17029 = (inp[1]) ? node17045 : node17030;
												assign node17030 = (inp[2]) ? node17038 : node17031;
													assign node17031 = (inp[8]) ? node17035 : node17032;
														assign node17032 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17035 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17038 = (inp[5]) ? node17042 : node17039;
														assign node17039 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17042 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17045 = (inp[2]) ? node17053 : node17046;
													assign node17046 = (inp[5]) ? node17050 : node17047;
														assign node17047 = (inp[8]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node17050 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17053 = (inp[9]) ? node17057 : node17054;
														assign node17054 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17057 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17060 = (inp[9]) ? node17076 : node17061;
												assign node17061 = (inp[0]) ? node17069 : node17062;
													assign node17062 = (inp[8]) ? node17066 : node17063;
														assign node17063 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17066 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node17069 = (inp[8]) ? node17073 : node17070;
														assign node17070 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17073 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node17076 = (inp[0]) ? node17084 : node17077;
													assign node17077 = (inp[8]) ? node17081 : node17078;
														assign node17078 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node17081 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node17084 = (inp[5]) ? node17088 : node17085;
														assign node17085 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17088 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
										assign node17091 = (inp[1]) ? node17121 : node17092;
											assign node17092 = (inp[5]) ? node17108 : node17093;
												assign node17093 = (inp[15]) ? node17101 : node17094;
													assign node17094 = (inp[0]) ? node17098 : node17095;
														assign node17095 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17098 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17101 = (inp[2]) ? node17105 : node17102;
														assign node17102 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17105 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node17108 = (inp[8]) ? node17116 : node17109;
													assign node17109 = (inp[15]) ? node17113 : node17110;
														assign node17110 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node17113 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17116 = (inp[15]) ? 16'b0000000011111111 : node17117;
														assign node17117 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17121 = (inp[9]) ? node17137 : node17122;
												assign node17122 = (inp[8]) ? node17130 : node17123;
													assign node17123 = (inp[0]) ? node17127 : node17124;
														assign node17124 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node17127 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17130 = (inp[2]) ? node17134 : node17131;
														assign node17131 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node17134 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17137 = (inp[15]) ? node17143 : node17138;
													assign node17138 = (inp[2]) ? node17140 : 16'b0000000111111111;
														assign node17140 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node17143 = (inp[5]) ? 16'b0000000000111111 : node17144;
														assign node17144 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
									assign node17148 = (inp[9]) ? node17208 : node17149;
										assign node17149 = (inp[7]) ? node17177 : node17150;
											assign node17150 = (inp[0]) ? node17164 : node17151;
												assign node17151 = (inp[1]) ? node17159 : node17152;
													assign node17152 = (inp[8]) ? node17156 : node17153;
														assign node17153 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17156 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17159 = (inp[15]) ? 16'b0000000111111111 : node17160;
														assign node17160 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
												assign node17164 = (inp[5]) ? node17170 : node17165;
													assign node17165 = (inp[2]) ? 16'b0000000111111111 : node17166;
														assign node17166 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17170 = (inp[15]) ? node17174 : node17171;
														assign node17171 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node17174 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node17177 = (inp[0]) ? node17193 : node17178;
												assign node17178 = (inp[2]) ? node17186 : node17179;
													assign node17179 = (inp[5]) ? node17183 : node17180;
														assign node17180 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17183 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17186 = (inp[5]) ? node17190 : node17187;
														assign node17187 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node17190 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17193 = (inp[15]) ? node17201 : node17194;
													assign node17194 = (inp[2]) ? node17198 : node17195;
														assign node17195 = (inp[8]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node17198 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17201 = (inp[8]) ? node17205 : node17202;
														assign node17202 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17205 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
										assign node17208 = (inp[8]) ? node17240 : node17209;
											assign node17209 = (inp[1]) ? node17225 : node17210;
												assign node17210 = (inp[2]) ? node17218 : node17211;
													assign node17211 = (inp[5]) ? node17215 : node17212;
														assign node17212 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17215 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17218 = (inp[7]) ? node17222 : node17219;
														assign node17219 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17222 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17225 = (inp[0]) ? node17233 : node17226;
													assign node17226 = (inp[5]) ? node17230 : node17227;
														assign node17227 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17230 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17233 = (inp[2]) ? node17237 : node17234;
														assign node17234 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node17237 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17240 = (inp[5]) ? node17256 : node17241;
												assign node17241 = (inp[0]) ? node17249 : node17242;
													assign node17242 = (inp[1]) ? node17246 : node17243;
														assign node17243 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17246 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17249 = (inp[2]) ? node17253 : node17250;
														assign node17250 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node17253 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17256 = (inp[1]) ? node17264 : node17257;
													assign node17257 = (inp[2]) ? node17261 : node17258;
														assign node17258 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node17261 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17264 = (inp[7]) ? node17268 : node17265;
														assign node17265 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17268 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node17271 = (inp[2]) ? node17391 : node17272;
									assign node17272 = (inp[8]) ? node17330 : node17273;
										assign node17273 = (inp[0]) ? node17299 : node17274;
											assign node17274 = (inp[14]) ? node17286 : node17275;
												assign node17275 = (inp[5]) ? node17283 : node17276;
													assign node17276 = (inp[1]) ? node17280 : node17277;
														assign node17277 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17280 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17283 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node17286 = (inp[15]) ? node17294 : node17287;
													assign node17287 = (inp[9]) ? node17291 : node17288;
														assign node17288 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17291 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17294 = (inp[1]) ? node17296 : 16'b0000000111111111;
														assign node17296 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node17299 = (inp[1]) ? node17315 : node17300;
												assign node17300 = (inp[5]) ? node17308 : node17301;
													assign node17301 = (inp[9]) ? node17305 : node17302;
														assign node17302 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node17305 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17308 = (inp[15]) ? node17312 : node17309;
														assign node17309 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node17312 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17315 = (inp[7]) ? node17323 : node17316;
													assign node17316 = (inp[15]) ? node17320 : node17317;
														assign node17317 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17320 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17323 = (inp[15]) ? node17327 : node17324;
														assign node17324 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17327 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node17330 = (inp[9]) ? node17360 : node17331;
											assign node17331 = (inp[14]) ? node17347 : node17332;
												assign node17332 = (inp[0]) ? node17340 : node17333;
													assign node17333 = (inp[1]) ? node17337 : node17334;
														assign node17334 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17337 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17340 = (inp[5]) ? node17344 : node17341;
														assign node17341 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17344 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17347 = (inp[15]) ? node17355 : node17348;
													assign node17348 = (inp[7]) ? node17352 : node17349;
														assign node17349 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17352 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17355 = (inp[1]) ? node17357 : 16'b0000000001111111;
														assign node17357 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17360 = (inp[5]) ? node17376 : node17361;
												assign node17361 = (inp[1]) ? node17369 : node17362;
													assign node17362 = (inp[0]) ? node17366 : node17363;
														assign node17363 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17366 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17369 = (inp[0]) ? node17373 : node17370;
														assign node17370 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17373 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17376 = (inp[15]) ? node17384 : node17377;
													assign node17377 = (inp[1]) ? node17381 : node17378;
														assign node17378 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17381 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17384 = (inp[7]) ? node17388 : node17385;
														assign node17385 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17388 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node17391 = (inp[9]) ? node17449 : node17392;
										assign node17392 = (inp[14]) ? node17418 : node17393;
											assign node17393 = (inp[7]) ? node17407 : node17394;
												assign node17394 = (inp[0]) ? node17400 : node17395;
													assign node17395 = (inp[15]) ? node17397 : 16'b0000000111111111;
														assign node17397 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17400 = (inp[5]) ? node17404 : node17401;
														assign node17401 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node17404 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17407 = (inp[15]) ? node17415 : node17408;
													assign node17408 = (inp[0]) ? node17412 : node17409;
														assign node17409 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17412 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17415 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17418 = (inp[0]) ? node17434 : node17419;
												assign node17419 = (inp[5]) ? node17427 : node17420;
													assign node17420 = (inp[7]) ? node17424 : node17421;
														assign node17421 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node17424 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17427 = (inp[15]) ? node17431 : node17428;
														assign node17428 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17431 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17434 = (inp[5]) ? node17442 : node17435;
													assign node17435 = (inp[7]) ? node17439 : node17436;
														assign node17436 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17439 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17442 = (inp[8]) ? node17446 : node17443;
														assign node17443 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17446 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node17449 = (inp[5]) ? node17481 : node17450;
											assign node17450 = (inp[1]) ? node17466 : node17451;
												assign node17451 = (inp[8]) ? node17459 : node17452;
													assign node17452 = (inp[14]) ? node17456 : node17453;
														assign node17453 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17456 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17459 = (inp[15]) ? node17463 : node17460;
														assign node17460 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node17463 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17466 = (inp[15]) ? node17474 : node17467;
													assign node17467 = (inp[8]) ? node17471 : node17468;
														assign node17468 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17471 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17474 = (inp[8]) ? node17478 : node17475;
														assign node17475 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17478 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node17481 = (inp[0]) ? node17491 : node17482;
												assign node17482 = (inp[14]) ? 16'b0000000000111111 : node17483;
													assign node17483 = (inp[15]) ? node17487 : node17484;
														assign node17484 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17487 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node17491 = (inp[1]) ? node17499 : node17492;
													assign node17492 = (inp[7]) ? node17496 : node17493;
														assign node17493 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17496 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node17499 = (inp[7]) ? node17503 : node17500;
														assign node17500 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node17503 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
					assign node17506 = (inp[2]) ? node18494 : node17507;
						assign node17507 = (inp[9]) ? node18001 : node17508;
							assign node17508 = (inp[8]) ? node17752 : node17509;
								assign node17509 = (inp[15]) ? node17635 : node17510;
									assign node17510 = (inp[4]) ? node17574 : node17511;
										assign node17511 = (inp[1]) ? node17543 : node17512;
											assign node17512 = (inp[0]) ? node17528 : node17513;
												assign node17513 = (inp[5]) ? node17521 : node17514;
													assign node17514 = (inp[3]) ? node17518 : node17515;
														assign node17515 = (inp[11]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node17518 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node17521 = (inp[11]) ? node17525 : node17522;
														assign node17522 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17525 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node17528 = (inp[14]) ? node17536 : node17529;
													assign node17529 = (inp[11]) ? node17533 : node17530;
														assign node17530 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17533 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17536 = (inp[11]) ? node17540 : node17537;
														assign node17537 = (inp[5]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node17540 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node17543 = (inp[7]) ? node17559 : node17544;
												assign node17544 = (inp[5]) ? node17552 : node17545;
													assign node17545 = (inp[0]) ? node17549 : node17546;
														assign node17546 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17549 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17552 = (inp[14]) ? node17556 : node17553;
														assign node17553 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17556 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17559 = (inp[3]) ? node17567 : node17560;
													assign node17560 = (inp[5]) ? node17564 : node17561;
														assign node17561 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17564 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17567 = (inp[5]) ? node17571 : node17568;
														assign node17568 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node17571 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node17574 = (inp[0]) ? node17606 : node17575;
											assign node17575 = (inp[11]) ? node17591 : node17576;
												assign node17576 = (inp[1]) ? node17584 : node17577;
													assign node17577 = (inp[14]) ? node17581 : node17578;
														assign node17578 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17581 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node17584 = (inp[7]) ? node17588 : node17585;
														assign node17585 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17588 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17591 = (inp[3]) ? node17599 : node17592;
													assign node17592 = (inp[5]) ? node17596 : node17593;
														assign node17593 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17596 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17599 = (inp[14]) ? node17603 : node17600;
														assign node17600 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17603 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17606 = (inp[1]) ? node17620 : node17607;
												assign node17607 = (inp[14]) ? node17615 : node17608;
													assign node17608 = (inp[7]) ? node17612 : node17609;
														assign node17609 = (inp[5]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node17612 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17615 = (inp[11]) ? 16'b0000000111111111 : node17616;
														assign node17616 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17620 = (inp[14]) ? node17628 : node17621;
													assign node17621 = (inp[11]) ? node17625 : node17622;
														assign node17622 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node17625 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17628 = (inp[5]) ? node17632 : node17629;
														assign node17629 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17632 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
									assign node17635 = (inp[11]) ? node17697 : node17636;
										assign node17636 = (inp[3]) ? node17666 : node17637;
											assign node17637 = (inp[0]) ? node17651 : node17638;
												assign node17638 = (inp[7]) ? node17644 : node17639;
													assign node17639 = (inp[1]) ? node17641 : 16'b0000111111111111;
														assign node17641 = (inp[4]) ? 16'b0000011111111111 : 16'b0000011111111111;
													assign node17644 = (inp[14]) ? node17648 : node17645;
														assign node17645 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17648 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17651 = (inp[7]) ? node17659 : node17652;
													assign node17652 = (inp[4]) ? node17656 : node17653;
														assign node17653 = (inp[1]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node17656 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17659 = (inp[5]) ? node17663 : node17660;
														assign node17660 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17663 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17666 = (inp[1]) ? node17682 : node17667;
												assign node17667 = (inp[14]) ? node17675 : node17668;
													assign node17668 = (inp[5]) ? node17672 : node17669;
														assign node17669 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17672 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17675 = (inp[4]) ? node17679 : node17676;
														assign node17676 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17679 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17682 = (inp[7]) ? node17690 : node17683;
													assign node17683 = (inp[5]) ? node17687 : node17684;
														assign node17684 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17687 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17690 = (inp[5]) ? node17694 : node17691;
														assign node17691 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17694 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node17697 = (inp[5]) ? node17725 : node17698;
											assign node17698 = (inp[3]) ? node17712 : node17699;
												assign node17699 = (inp[0]) ? node17705 : node17700;
													assign node17700 = (inp[7]) ? node17702 : 16'b0000011111111111;
														assign node17702 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17705 = (inp[1]) ? node17709 : node17706;
														assign node17706 = (inp[4]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node17709 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17712 = (inp[1]) ? node17720 : node17713;
													assign node17713 = (inp[7]) ? node17717 : node17714;
														assign node17714 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17717 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node17720 = (inp[4]) ? node17722 : 16'b0000000011111111;
														assign node17722 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17725 = (inp[4]) ? node17739 : node17726;
												assign node17726 = (inp[0]) ? node17734 : node17727;
													assign node17727 = (inp[7]) ? node17731 : node17728;
														assign node17728 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17731 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17734 = (inp[7]) ? 16'b0000000001111111 : node17735;
														assign node17735 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17739 = (inp[14]) ? node17747 : node17740;
													assign node17740 = (inp[7]) ? node17744 : node17741;
														assign node17741 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17744 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node17747 = (inp[7]) ? 16'b0000000001111111 : node17748;
														assign node17748 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node17752 = (inp[11]) ? node17878 : node17753;
									assign node17753 = (inp[14]) ? node17817 : node17754;
										assign node17754 = (inp[15]) ? node17786 : node17755;
											assign node17755 = (inp[7]) ? node17771 : node17756;
												assign node17756 = (inp[5]) ? node17764 : node17757;
													assign node17757 = (inp[4]) ? node17761 : node17758;
														assign node17758 = (inp[1]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node17761 = (inp[1]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node17764 = (inp[3]) ? node17768 : node17765;
														assign node17765 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17768 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node17771 = (inp[4]) ? node17779 : node17772;
													assign node17772 = (inp[0]) ? node17776 : node17773;
														assign node17773 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17776 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17779 = (inp[1]) ? node17783 : node17780;
														assign node17780 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17783 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node17786 = (inp[0]) ? node17802 : node17787;
												assign node17787 = (inp[1]) ? node17795 : node17788;
													assign node17788 = (inp[4]) ? node17792 : node17789;
														assign node17789 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17792 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17795 = (inp[3]) ? node17799 : node17796;
														assign node17796 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node17799 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node17802 = (inp[7]) ? node17810 : node17803;
													assign node17803 = (inp[5]) ? node17807 : node17804;
														assign node17804 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node17807 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17810 = (inp[4]) ? node17814 : node17811;
														assign node17811 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17814 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node17817 = (inp[4]) ? node17849 : node17818;
											assign node17818 = (inp[3]) ? node17834 : node17819;
												assign node17819 = (inp[7]) ? node17827 : node17820;
													assign node17820 = (inp[15]) ? node17824 : node17821;
														assign node17821 = (inp[5]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node17824 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17827 = (inp[5]) ? node17831 : node17828;
														assign node17828 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node17831 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17834 = (inp[5]) ? node17842 : node17835;
													assign node17835 = (inp[15]) ? node17839 : node17836;
														assign node17836 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17839 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node17842 = (inp[1]) ? node17846 : node17843;
														assign node17843 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17846 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node17849 = (inp[0]) ? node17865 : node17850;
												assign node17850 = (inp[1]) ? node17858 : node17851;
													assign node17851 = (inp[15]) ? node17855 : node17852;
														assign node17852 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17855 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17858 = (inp[3]) ? node17862 : node17859;
														assign node17859 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17862 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17865 = (inp[3]) ? node17873 : node17866;
													assign node17866 = (inp[5]) ? node17870 : node17867;
														assign node17867 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17870 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17873 = (inp[15]) ? 16'b0000000001111111 : node17874;
														assign node17874 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node17878 = (inp[7]) ? node17938 : node17879;
										assign node17879 = (inp[0]) ? node17911 : node17880;
											assign node17880 = (inp[3]) ? node17896 : node17881;
												assign node17881 = (inp[4]) ? node17889 : node17882;
													assign node17882 = (inp[15]) ? node17886 : node17883;
														assign node17883 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node17886 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node17889 = (inp[5]) ? node17893 : node17890;
														assign node17890 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17893 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node17896 = (inp[1]) ? node17904 : node17897;
													assign node17897 = (inp[5]) ? node17901 : node17898;
														assign node17898 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17901 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17904 = (inp[4]) ? node17908 : node17905;
														assign node17905 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17908 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node17911 = (inp[5]) ? node17925 : node17912;
												assign node17912 = (inp[14]) ? node17918 : node17913;
													assign node17913 = (inp[3]) ? node17915 : 16'b0000000111111111;
														assign node17915 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17918 = (inp[4]) ? node17922 : node17919;
														assign node17919 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17922 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node17925 = (inp[4]) ? node17933 : node17926;
													assign node17926 = (inp[15]) ? node17930 : node17927;
														assign node17927 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node17930 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17933 = (inp[3]) ? node17935 : 16'b0000000011111111;
														assign node17935 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node17938 = (inp[15]) ? node17970 : node17939;
											assign node17939 = (inp[3]) ? node17955 : node17940;
												assign node17940 = (inp[1]) ? node17948 : node17941;
													assign node17941 = (inp[4]) ? node17945 : node17942;
														assign node17942 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node17945 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node17948 = (inp[14]) ? node17952 : node17949;
														assign node17949 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17952 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node17955 = (inp[4]) ? node17963 : node17956;
													assign node17956 = (inp[5]) ? node17960 : node17957;
														assign node17957 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17960 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17963 = (inp[1]) ? node17967 : node17964;
														assign node17964 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17967 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node17970 = (inp[4]) ? node17986 : node17971;
												assign node17971 = (inp[1]) ? node17979 : node17972;
													assign node17972 = (inp[14]) ? node17976 : node17973;
														assign node17973 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node17976 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node17979 = (inp[0]) ? node17983 : node17980;
														assign node17980 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17983 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node17986 = (inp[0]) ? node17994 : node17987;
													assign node17987 = (inp[3]) ? node17991 : node17988;
														assign node17988 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node17991 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node17994 = (inp[14]) ? node17998 : node17995;
														assign node17995 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node17998 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
							assign node18001 = (inp[3]) ? node18245 : node18002;
								assign node18002 = (inp[4]) ? node18126 : node18003;
									assign node18003 = (inp[5]) ? node18067 : node18004;
										assign node18004 = (inp[1]) ? node18036 : node18005;
											assign node18005 = (inp[14]) ? node18021 : node18006;
												assign node18006 = (inp[8]) ? node18014 : node18007;
													assign node18007 = (inp[11]) ? node18011 : node18008;
														assign node18008 = (inp[15]) ? 16'b0000111111111111 : 16'b0000111111111111;
														assign node18011 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18014 = (inp[15]) ? node18018 : node18015;
														assign node18015 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18018 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18021 = (inp[7]) ? node18029 : node18022;
													assign node18022 = (inp[8]) ? node18026 : node18023;
														assign node18023 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18026 = (inp[15]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node18029 = (inp[15]) ? node18033 : node18030;
														assign node18030 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18033 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18036 = (inp[11]) ? node18052 : node18037;
												assign node18037 = (inp[14]) ? node18045 : node18038;
													assign node18038 = (inp[15]) ? node18042 : node18039;
														assign node18039 = (inp[7]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node18042 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18045 = (inp[8]) ? node18049 : node18046;
														assign node18046 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18049 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18052 = (inp[0]) ? node18060 : node18053;
													assign node18053 = (inp[15]) ? node18057 : node18054;
														assign node18054 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18057 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18060 = (inp[14]) ? node18064 : node18061;
														assign node18061 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18064 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node18067 = (inp[15]) ? node18097 : node18068;
											assign node18068 = (inp[8]) ? node18084 : node18069;
												assign node18069 = (inp[1]) ? node18077 : node18070;
													assign node18070 = (inp[14]) ? node18074 : node18071;
														assign node18071 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18074 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18077 = (inp[14]) ? node18081 : node18078;
														assign node18078 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node18081 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18084 = (inp[0]) ? node18092 : node18085;
													assign node18085 = (inp[14]) ? node18089 : node18086;
														assign node18086 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18089 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18092 = (inp[7]) ? node18094 : 16'b0000000011111111;
														assign node18094 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18097 = (inp[1]) ? node18113 : node18098;
												assign node18098 = (inp[11]) ? node18106 : node18099;
													assign node18099 = (inp[7]) ? node18103 : node18100;
														assign node18100 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node18103 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18106 = (inp[0]) ? node18110 : node18107;
														assign node18107 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node18110 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18113 = (inp[14]) ? node18119 : node18114;
													assign node18114 = (inp[11]) ? 16'b0000000011111111 : node18115;
														assign node18115 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18119 = (inp[11]) ? node18123 : node18120;
														assign node18120 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node18123 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node18126 = (inp[14]) ? node18186 : node18127;
										assign node18127 = (inp[15]) ? node18159 : node18128;
											assign node18128 = (inp[1]) ? node18144 : node18129;
												assign node18129 = (inp[11]) ? node18137 : node18130;
													assign node18130 = (inp[0]) ? node18134 : node18131;
														assign node18131 = (inp[8]) ? 16'b0000011111111111 : 16'b0000011111111111;
														assign node18134 = (inp[7]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node18137 = (inp[8]) ? node18141 : node18138;
														assign node18138 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18141 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18144 = (inp[7]) ? node18152 : node18145;
													assign node18145 = (inp[8]) ? node18149 : node18146;
														assign node18146 = (inp[0]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node18149 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18152 = (inp[11]) ? node18156 : node18153;
														assign node18153 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node18156 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18159 = (inp[5]) ? node18175 : node18160;
												assign node18160 = (inp[0]) ? node18168 : node18161;
													assign node18161 = (inp[8]) ? node18165 : node18162;
														assign node18162 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18165 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18168 = (inp[11]) ? node18172 : node18169;
														assign node18169 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18172 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18175 = (inp[0]) ? node18181 : node18176;
													assign node18176 = (inp[1]) ? node18178 : 16'b0000000011111111;
														assign node18178 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18181 = (inp[11]) ? node18183 : 16'b0000000001111111;
														assign node18183 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node18186 = (inp[11]) ? node18214 : node18187;
											assign node18187 = (inp[1]) ? node18199 : node18188;
												assign node18188 = (inp[5]) ? node18194 : node18189;
													assign node18189 = (inp[7]) ? node18191 : 16'b0000001111111111;
														assign node18191 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18194 = (inp[15]) ? 16'b0000000011111111 : node18195;
														assign node18195 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18199 = (inp[15]) ? node18207 : node18200;
													assign node18200 = (inp[7]) ? node18204 : node18201;
														assign node18201 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18204 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18207 = (inp[0]) ? node18211 : node18208;
														assign node18208 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18211 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node18214 = (inp[5]) ? node18230 : node18215;
												assign node18215 = (inp[8]) ? node18223 : node18216;
													assign node18216 = (inp[7]) ? node18220 : node18217;
														assign node18217 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18220 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18223 = (inp[15]) ? node18227 : node18224;
														assign node18224 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18227 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18230 = (inp[15]) ? node18238 : node18231;
													assign node18231 = (inp[7]) ? node18235 : node18232;
														assign node18232 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18235 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18238 = (inp[1]) ? node18242 : node18239;
														assign node18239 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18242 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node18245 = (inp[11]) ? node18369 : node18246;
									assign node18246 = (inp[7]) ? node18308 : node18247;
										assign node18247 = (inp[1]) ? node18277 : node18248;
											assign node18248 = (inp[4]) ? node18262 : node18249;
												assign node18249 = (inp[14]) ? node18255 : node18250;
													assign node18250 = (inp[15]) ? 16'b0000001111111111 : node18251;
														assign node18251 = (inp[0]) ? 16'b0000011111111111 : 16'b0000011111111111;
													assign node18255 = (inp[5]) ? node18259 : node18256;
														assign node18256 = (inp[8]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node18259 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18262 = (inp[0]) ? node18270 : node18263;
													assign node18263 = (inp[15]) ? node18267 : node18264;
														assign node18264 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18267 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18270 = (inp[14]) ? node18274 : node18271;
														assign node18271 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18274 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18277 = (inp[4]) ? node18293 : node18278;
												assign node18278 = (inp[14]) ? node18286 : node18279;
													assign node18279 = (inp[15]) ? node18283 : node18280;
														assign node18280 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18283 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18286 = (inp[8]) ? node18290 : node18287;
														assign node18287 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18290 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18293 = (inp[15]) ? node18301 : node18294;
													assign node18294 = (inp[5]) ? node18298 : node18295;
														assign node18295 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18298 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18301 = (inp[14]) ? node18305 : node18302;
														assign node18302 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18305 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node18308 = (inp[14]) ? node18340 : node18309;
											assign node18309 = (inp[1]) ? node18325 : node18310;
												assign node18310 = (inp[4]) ? node18318 : node18311;
													assign node18311 = (inp[5]) ? node18315 : node18312;
														assign node18312 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18315 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18318 = (inp[15]) ? node18322 : node18319;
														assign node18319 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18322 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18325 = (inp[8]) ? node18333 : node18326;
													assign node18326 = (inp[0]) ? node18330 : node18327;
														assign node18327 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18330 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node18333 = (inp[0]) ? node18337 : node18334;
														assign node18334 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node18337 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node18340 = (inp[4]) ? node18354 : node18341;
												assign node18341 = (inp[15]) ? node18347 : node18342;
													assign node18342 = (inp[1]) ? 16'b0000000001111111 : node18343;
														assign node18343 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node18347 = (inp[0]) ? node18351 : node18348;
														assign node18348 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18351 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18354 = (inp[1]) ? node18362 : node18355;
													assign node18355 = (inp[5]) ? node18359 : node18356;
														assign node18356 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18359 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node18362 = (inp[15]) ? node18366 : node18363;
														assign node18363 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node18366 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node18369 = (inp[5]) ? node18433 : node18370;
										assign node18370 = (inp[15]) ? node18402 : node18371;
											assign node18371 = (inp[14]) ? node18387 : node18372;
												assign node18372 = (inp[7]) ? node18380 : node18373;
													assign node18373 = (inp[1]) ? node18377 : node18374;
														assign node18374 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18377 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18380 = (inp[4]) ? node18384 : node18381;
														assign node18381 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18384 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18387 = (inp[0]) ? node18395 : node18388;
													assign node18388 = (inp[1]) ? node18392 : node18389;
														assign node18389 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18392 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18395 = (inp[7]) ? node18399 : node18396;
														assign node18396 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18399 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node18402 = (inp[4]) ? node18418 : node18403;
												assign node18403 = (inp[8]) ? node18411 : node18404;
													assign node18404 = (inp[1]) ? node18408 : node18405;
														assign node18405 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18408 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node18411 = (inp[7]) ? node18415 : node18412;
														assign node18412 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18415 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18418 = (inp[0]) ? node18426 : node18419;
													assign node18419 = (inp[14]) ? node18423 : node18420;
														assign node18420 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node18423 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18426 = (inp[1]) ? node18430 : node18427;
														assign node18427 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18430 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node18433 = (inp[7]) ? node18465 : node18434;
											assign node18434 = (inp[4]) ? node18450 : node18435;
												assign node18435 = (inp[8]) ? node18443 : node18436;
													assign node18436 = (inp[14]) ? node18440 : node18437;
														assign node18437 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node18440 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18443 = (inp[1]) ? node18447 : node18444;
														assign node18444 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18447 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node18450 = (inp[14]) ? node18458 : node18451;
													assign node18451 = (inp[15]) ? node18455 : node18452;
														assign node18452 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node18455 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18458 = (inp[0]) ? node18462 : node18459;
														assign node18459 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18462 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node18465 = (inp[1]) ? node18479 : node18466;
												assign node18466 = (inp[8]) ? node18472 : node18467;
													assign node18467 = (inp[0]) ? node18469 : 16'b0000000001111111;
														assign node18469 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18472 = (inp[0]) ? node18476 : node18473;
														assign node18473 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18476 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node18479 = (inp[14]) ? node18487 : node18480;
													assign node18480 = (inp[8]) ? node18484 : node18481;
														assign node18481 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18484 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node18487 = (inp[4]) ? node18491 : node18488;
														assign node18488 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node18491 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node18494 = (inp[8]) ? node18988 : node18495;
							assign node18495 = (inp[0]) ? node18741 : node18496;
								assign node18496 = (inp[15]) ? node18622 : node18497;
									assign node18497 = (inp[3]) ? node18559 : node18498;
										assign node18498 = (inp[9]) ? node18530 : node18499;
											assign node18499 = (inp[1]) ? node18515 : node18500;
												assign node18500 = (inp[4]) ? node18508 : node18501;
													assign node18501 = (inp[11]) ? node18505 : node18502;
														assign node18502 = (inp[5]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node18505 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node18508 = (inp[7]) ? node18512 : node18509;
														assign node18509 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18512 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node18515 = (inp[14]) ? node18523 : node18516;
													assign node18516 = (inp[11]) ? node18520 : node18517;
														assign node18517 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18520 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18523 = (inp[7]) ? node18527 : node18524;
														assign node18524 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18527 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node18530 = (inp[1]) ? node18546 : node18531;
												assign node18531 = (inp[14]) ? node18539 : node18532;
													assign node18532 = (inp[7]) ? node18536 : node18533;
														assign node18533 = (inp[5]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node18536 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18539 = (inp[4]) ? node18543 : node18540;
														assign node18540 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18543 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18546 = (inp[4]) ? node18554 : node18547;
													assign node18547 = (inp[14]) ? node18551 : node18548;
														assign node18548 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18551 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18554 = (inp[5]) ? 16'b0000000011111111 : node18555;
														assign node18555 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node18559 = (inp[7]) ? node18591 : node18560;
											assign node18560 = (inp[9]) ? node18576 : node18561;
												assign node18561 = (inp[11]) ? node18569 : node18562;
													assign node18562 = (inp[5]) ? node18566 : node18563;
														assign node18563 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18566 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18569 = (inp[4]) ? node18573 : node18570;
														assign node18570 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18573 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18576 = (inp[14]) ? node18584 : node18577;
													assign node18577 = (inp[1]) ? node18581 : node18578;
														assign node18578 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node18581 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18584 = (inp[11]) ? node18588 : node18585;
														assign node18585 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18588 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18591 = (inp[5]) ? node18607 : node18592;
												assign node18592 = (inp[4]) ? node18600 : node18593;
													assign node18593 = (inp[9]) ? node18597 : node18594;
														assign node18594 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18597 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18600 = (inp[14]) ? node18604 : node18601;
														assign node18601 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18604 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18607 = (inp[14]) ? node18615 : node18608;
													assign node18608 = (inp[4]) ? node18612 : node18609;
														assign node18609 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18612 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18615 = (inp[11]) ? node18619 : node18616;
														assign node18616 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18619 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node18622 = (inp[9]) ? node18682 : node18623;
										assign node18623 = (inp[3]) ? node18653 : node18624;
											assign node18624 = (inp[5]) ? node18638 : node18625;
												assign node18625 = (inp[4]) ? node18631 : node18626;
													assign node18626 = (inp[7]) ? node18628 : 16'b0000001111111111;
														assign node18628 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18631 = (inp[14]) ? node18635 : node18632;
														assign node18632 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18635 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node18638 = (inp[7]) ? node18646 : node18639;
													assign node18639 = (inp[11]) ? node18643 : node18640;
														assign node18640 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18643 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18646 = (inp[1]) ? node18650 : node18647;
														assign node18647 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18650 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18653 = (inp[1]) ? node18669 : node18654;
												assign node18654 = (inp[5]) ? node18662 : node18655;
													assign node18655 = (inp[7]) ? node18659 : node18656;
														assign node18656 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18659 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node18662 = (inp[7]) ? node18666 : node18663;
														assign node18663 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18666 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18669 = (inp[4]) ? node18677 : node18670;
													assign node18670 = (inp[5]) ? node18674 : node18671;
														assign node18671 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18674 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18677 = (inp[5]) ? 16'b0000000001111111 : node18678;
														assign node18678 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node18682 = (inp[1]) ? node18710 : node18683;
											assign node18683 = (inp[7]) ? node18699 : node18684;
												assign node18684 = (inp[14]) ? node18692 : node18685;
													assign node18685 = (inp[5]) ? node18689 : node18686;
														assign node18686 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18689 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18692 = (inp[4]) ? node18696 : node18693;
														assign node18693 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18696 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18699 = (inp[11]) ? node18705 : node18700;
													assign node18700 = (inp[3]) ? node18702 : 16'b0000000011111111;
														assign node18702 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18705 = (inp[5]) ? node18707 : 16'b0000000011111111;
														assign node18707 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node18710 = (inp[14]) ? node18726 : node18711;
												assign node18711 = (inp[4]) ? node18719 : node18712;
													assign node18712 = (inp[11]) ? node18716 : node18713;
														assign node18713 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18716 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18719 = (inp[5]) ? node18723 : node18720;
														assign node18720 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18723 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node18726 = (inp[5]) ? node18734 : node18727;
													assign node18727 = (inp[7]) ? node18731 : node18728;
														assign node18728 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node18731 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18734 = (inp[11]) ? node18738 : node18735;
														assign node18735 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18738 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node18741 = (inp[7]) ? node18867 : node18742;
									assign node18742 = (inp[14]) ? node18806 : node18743;
										assign node18743 = (inp[1]) ? node18775 : node18744;
											assign node18744 = (inp[3]) ? node18760 : node18745;
												assign node18745 = (inp[11]) ? node18753 : node18746;
													assign node18746 = (inp[9]) ? node18750 : node18747;
														assign node18747 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18750 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node18753 = (inp[4]) ? node18757 : node18754;
														assign node18754 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18757 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node18760 = (inp[15]) ? node18768 : node18761;
													assign node18761 = (inp[9]) ? node18765 : node18762;
														assign node18762 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18765 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18768 = (inp[4]) ? node18772 : node18769;
														assign node18769 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18772 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18775 = (inp[9]) ? node18791 : node18776;
												assign node18776 = (inp[4]) ? node18784 : node18777;
													assign node18777 = (inp[3]) ? node18781 : node18778;
														assign node18778 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18781 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18784 = (inp[5]) ? node18788 : node18785;
														assign node18785 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18788 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18791 = (inp[5]) ? node18799 : node18792;
													assign node18792 = (inp[3]) ? node18796 : node18793;
														assign node18793 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18796 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18799 = (inp[11]) ? node18803 : node18800;
														assign node18800 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18803 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node18806 = (inp[11]) ? node18836 : node18807;
											assign node18807 = (inp[9]) ? node18823 : node18808;
												assign node18808 = (inp[1]) ? node18816 : node18809;
													assign node18809 = (inp[5]) ? node18813 : node18810;
														assign node18810 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18813 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18816 = (inp[4]) ? node18820 : node18817;
														assign node18817 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18820 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node18823 = (inp[5]) ? node18829 : node18824;
													assign node18824 = (inp[4]) ? node18826 : 16'b0000000011111111;
														assign node18826 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18829 = (inp[1]) ? node18833 : node18830;
														assign node18830 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18833 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node18836 = (inp[15]) ? node18852 : node18837;
												assign node18837 = (inp[4]) ? node18845 : node18838;
													assign node18838 = (inp[3]) ? node18842 : node18839;
														assign node18839 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18842 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18845 = (inp[3]) ? node18849 : node18846;
														assign node18846 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18849 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18852 = (inp[1]) ? node18860 : node18853;
													assign node18853 = (inp[3]) ? node18857 : node18854;
														assign node18854 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18857 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node18860 = (inp[3]) ? node18864 : node18861;
														assign node18861 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node18864 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node18867 = (inp[3]) ? node18927 : node18868;
										assign node18868 = (inp[15]) ? node18898 : node18869;
											assign node18869 = (inp[1]) ? node18885 : node18870;
												assign node18870 = (inp[4]) ? node18878 : node18871;
													assign node18871 = (inp[9]) ? node18875 : node18872;
														assign node18872 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node18875 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node18878 = (inp[14]) ? node18882 : node18879;
														assign node18879 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18882 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node18885 = (inp[5]) ? node18893 : node18886;
													assign node18886 = (inp[11]) ? node18890 : node18887;
														assign node18887 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node18890 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18893 = (inp[11]) ? 16'b0000000001111111 : node18894;
														assign node18894 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node18898 = (inp[4]) ? node18914 : node18899;
												assign node18899 = (inp[14]) ? node18907 : node18900;
													assign node18900 = (inp[11]) ? node18904 : node18901;
														assign node18901 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18904 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18907 = (inp[9]) ? node18911 : node18908;
														assign node18908 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18911 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18914 = (inp[9]) ? node18922 : node18915;
													assign node18915 = (inp[5]) ? node18919 : node18916;
														assign node18916 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node18919 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node18922 = (inp[11]) ? node18924 : 16'b0000000000111111;
														assign node18924 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node18927 = (inp[1]) ? node18957 : node18928;
											assign node18928 = (inp[15]) ? node18944 : node18929;
												assign node18929 = (inp[14]) ? node18937 : node18930;
													assign node18930 = (inp[5]) ? node18934 : node18931;
														assign node18931 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node18934 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node18937 = (inp[5]) ? node18941 : node18938;
														assign node18938 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18941 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node18944 = (inp[4]) ? node18952 : node18945;
													assign node18945 = (inp[11]) ? node18949 : node18946;
														assign node18946 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18949 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node18952 = (inp[14]) ? node18954 : 16'b0000000000111111;
														assign node18954 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000111111;
											assign node18957 = (inp[14]) ? node18973 : node18958;
												assign node18958 = (inp[9]) ? node18966 : node18959;
													assign node18959 = (inp[4]) ? node18963 : node18960;
														assign node18960 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node18963 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node18966 = (inp[15]) ? node18970 : node18967;
														assign node18967 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node18970 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node18973 = (inp[11]) ? node18981 : node18974;
													assign node18974 = (inp[15]) ? node18978 : node18975;
														assign node18975 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node18978 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node18981 = (inp[5]) ? node18985 : node18982;
														assign node18982 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node18985 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node18988 = (inp[4]) ? node19236 : node18989;
								assign node18989 = (inp[14]) ? node19113 : node18990;
									assign node18990 = (inp[3]) ? node19054 : node18991;
										assign node18991 = (inp[1]) ? node19023 : node18992;
											assign node18992 = (inp[0]) ? node19008 : node18993;
												assign node18993 = (inp[5]) ? node19001 : node18994;
													assign node18994 = (inp[7]) ? node18998 : node18995;
														assign node18995 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node18998 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19001 = (inp[11]) ? node19005 : node19002;
														assign node19002 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19005 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19008 = (inp[9]) ? node19016 : node19009;
													assign node19009 = (inp[11]) ? node19013 : node19010;
														assign node19010 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19013 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19016 = (inp[15]) ? node19020 : node19017;
														assign node19017 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19020 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19023 = (inp[11]) ? node19039 : node19024;
												assign node19024 = (inp[15]) ? node19032 : node19025;
													assign node19025 = (inp[5]) ? node19029 : node19026;
														assign node19026 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19029 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19032 = (inp[7]) ? node19036 : node19033;
														assign node19033 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19036 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19039 = (inp[0]) ? node19047 : node19040;
													assign node19040 = (inp[15]) ? node19044 : node19041;
														assign node19041 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19044 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19047 = (inp[9]) ? node19051 : node19048;
														assign node19048 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19051 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node19054 = (inp[15]) ? node19084 : node19055;
											assign node19055 = (inp[9]) ? node19069 : node19056;
												assign node19056 = (inp[7]) ? node19064 : node19057;
													assign node19057 = (inp[5]) ? node19061 : node19058;
														assign node19058 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19061 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19064 = (inp[5]) ? 16'b0000000011111111 : node19065;
														assign node19065 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19069 = (inp[0]) ? node19077 : node19070;
													assign node19070 = (inp[7]) ? node19074 : node19071;
														assign node19071 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19074 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19077 = (inp[1]) ? node19081 : node19078;
														assign node19078 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node19081 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19084 = (inp[11]) ? node19098 : node19085;
												assign node19085 = (inp[5]) ? node19091 : node19086;
													assign node19086 = (inp[7]) ? node19088 : 16'b0000000111111111;
														assign node19088 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19091 = (inp[1]) ? node19095 : node19092;
														assign node19092 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19095 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19098 = (inp[5]) ? node19106 : node19099;
													assign node19099 = (inp[7]) ? node19103 : node19100;
														assign node19100 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19103 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19106 = (inp[1]) ? node19110 : node19107;
														assign node19107 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19110 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node19113 = (inp[0]) ? node19177 : node19114;
										assign node19114 = (inp[1]) ? node19146 : node19115;
											assign node19115 = (inp[11]) ? node19131 : node19116;
												assign node19116 = (inp[9]) ? node19124 : node19117;
													assign node19117 = (inp[7]) ? node19121 : node19118;
														assign node19118 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19121 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node19124 = (inp[5]) ? node19128 : node19125;
														assign node19125 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19128 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19131 = (inp[15]) ? node19139 : node19132;
													assign node19132 = (inp[9]) ? node19136 : node19133;
														assign node19133 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node19136 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19139 = (inp[9]) ? node19143 : node19140;
														assign node19140 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19143 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19146 = (inp[9]) ? node19162 : node19147;
												assign node19147 = (inp[3]) ? node19155 : node19148;
													assign node19148 = (inp[11]) ? node19152 : node19149;
														assign node19149 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19152 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19155 = (inp[7]) ? node19159 : node19156;
														assign node19156 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19159 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19162 = (inp[15]) ? node19170 : node19163;
													assign node19163 = (inp[3]) ? node19167 : node19164;
														assign node19164 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19167 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19170 = (inp[5]) ? node19174 : node19171;
														assign node19171 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19174 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node19177 = (inp[3]) ? node19207 : node19178;
											assign node19178 = (inp[7]) ? node19194 : node19179;
												assign node19179 = (inp[5]) ? node19187 : node19180;
													assign node19180 = (inp[9]) ? node19184 : node19181;
														assign node19181 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19184 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19187 = (inp[9]) ? node19191 : node19188;
														assign node19188 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19191 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node19194 = (inp[15]) ? node19200 : node19195;
													assign node19195 = (inp[11]) ? node19197 : 16'b0000000001111111;
														assign node19197 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19200 = (inp[5]) ? node19204 : node19201;
														assign node19201 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node19204 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node19207 = (inp[9]) ? node19223 : node19208;
												assign node19208 = (inp[15]) ? node19216 : node19209;
													assign node19209 = (inp[11]) ? node19213 : node19210;
														assign node19210 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19213 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19216 = (inp[1]) ? node19220 : node19217;
														assign node19217 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19220 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node19223 = (inp[15]) ? node19231 : node19224;
													assign node19224 = (inp[5]) ? node19228 : node19225;
														assign node19225 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19228 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node19231 = (inp[11]) ? node19233 : 16'b0000000000111111;
														assign node19233 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000001111;
								assign node19236 = (inp[11]) ? node19358 : node19237;
									assign node19237 = (inp[3]) ? node19299 : node19238;
										assign node19238 = (inp[1]) ? node19270 : node19239;
											assign node19239 = (inp[9]) ? node19255 : node19240;
												assign node19240 = (inp[7]) ? node19248 : node19241;
													assign node19241 = (inp[14]) ? node19245 : node19242;
														assign node19242 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node19245 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node19248 = (inp[5]) ? node19252 : node19249;
														assign node19249 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19252 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node19255 = (inp[0]) ? node19263 : node19256;
													assign node19256 = (inp[5]) ? node19260 : node19257;
														assign node19257 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19260 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node19263 = (inp[5]) ? node19267 : node19264;
														assign node19264 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19267 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19270 = (inp[5]) ? node19286 : node19271;
												assign node19271 = (inp[7]) ? node19279 : node19272;
													assign node19272 = (inp[15]) ? node19276 : node19273;
														assign node19273 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19276 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19279 = (inp[0]) ? node19283 : node19280;
														assign node19280 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19283 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19286 = (inp[14]) ? node19292 : node19287;
													assign node19287 = (inp[15]) ? 16'b0000000001111111 : node19288;
														assign node19288 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node19292 = (inp[0]) ? node19296 : node19293;
														assign node19293 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19296 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node19299 = (inp[1]) ? node19331 : node19300;
											assign node19300 = (inp[15]) ? node19316 : node19301;
												assign node19301 = (inp[0]) ? node19309 : node19302;
													assign node19302 = (inp[5]) ? node19306 : node19303;
														assign node19303 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19306 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19309 = (inp[5]) ? node19313 : node19310;
														assign node19310 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19313 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19316 = (inp[5]) ? node19324 : node19317;
													assign node19317 = (inp[9]) ? node19321 : node19318;
														assign node19318 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19321 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19324 = (inp[14]) ? node19328 : node19325;
														assign node19325 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19328 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node19331 = (inp[9]) ? node19345 : node19332;
												assign node19332 = (inp[0]) ? node19338 : node19333;
													assign node19333 = (inp[14]) ? 16'b0000000001111111 : node19334;
														assign node19334 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19338 = (inp[5]) ? node19342 : node19339;
														assign node19339 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19342 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node19345 = (inp[14]) ? node19351 : node19346;
													assign node19346 = (inp[0]) ? node19348 : 16'b0000000001111111;
														assign node19348 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
													assign node19351 = (inp[15]) ? node19355 : node19352;
														assign node19352 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node19355 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node19358 = (inp[7]) ? node19418 : node19359;
										assign node19359 = (inp[15]) ? node19387 : node19360;
											assign node19360 = (inp[14]) ? node19374 : node19361;
												assign node19361 = (inp[5]) ? node19367 : node19362;
													assign node19362 = (inp[3]) ? 16'b0000000011111111 : node19363;
														assign node19363 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node19367 = (inp[9]) ? node19371 : node19368;
														assign node19368 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19371 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19374 = (inp[1]) ? node19382 : node19375;
													assign node19375 = (inp[3]) ? node19379 : node19376;
														assign node19376 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node19379 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node19382 = (inp[0]) ? 16'b0000000000111111 : node19383;
														assign node19383 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19387 = (inp[14]) ? node19403 : node19388;
												assign node19388 = (inp[1]) ? node19396 : node19389;
													assign node19389 = (inp[5]) ? node19393 : node19390;
														assign node19390 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19393 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node19396 = (inp[0]) ? node19400 : node19397;
														assign node19397 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19400 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node19403 = (inp[5]) ? node19411 : node19404;
													assign node19404 = (inp[9]) ? node19408 : node19405;
														assign node19405 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node19408 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000011111;
													assign node19411 = (inp[0]) ? node19415 : node19412;
														assign node19412 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node19415 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node19418 = (inp[0]) ? node19448 : node19419;
											assign node19419 = (inp[1]) ? node19435 : node19420;
												assign node19420 = (inp[5]) ? node19428 : node19421;
													assign node19421 = (inp[15]) ? node19425 : node19422;
														assign node19422 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node19425 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19428 = (inp[3]) ? node19432 : node19429;
														assign node19429 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19432 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node19435 = (inp[5]) ? node19441 : node19436;
													assign node19436 = (inp[3]) ? node19438 : 16'b0000000000111111;
														assign node19438 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node19441 = (inp[14]) ? node19445 : node19442;
														assign node19442 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node19445 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node19448 = (inp[3]) ? node19464 : node19449;
												assign node19449 = (inp[1]) ? node19457 : node19450;
													assign node19450 = (inp[14]) ? node19454 : node19451;
														assign node19451 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19454 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node19457 = (inp[5]) ? node19461 : node19458;
														assign node19458 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node19461 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node19464 = (inp[5]) ? node19472 : node19465;
													assign node19465 = (inp[15]) ? node19469 : node19466;
														assign node19466 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node19469 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node19472 = (inp[14]) ? node19476 : node19473;
														assign node19473 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node19476 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
				assign node19479 = (inp[5]) ? node21419 : node19480;
					assign node19480 = (inp[8]) ? node20462 : node19481;
						assign node19481 = (inp[3]) ? node19973 : node19482;
							assign node19482 = (inp[1]) ? node19730 : node19483;
								assign node19483 = (inp[14]) ? node19605 : node19484;
									assign node19484 = (inp[4]) ? node19544 : node19485;
										assign node19485 = (inp[15]) ? node19515 : node19486;
											assign node19486 = (inp[9]) ? node19502 : node19487;
												assign node19487 = (inp[11]) ? node19495 : node19488;
													assign node19488 = (inp[13]) ? node19492 : node19489;
														assign node19489 = (inp[2]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node19492 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node19495 = (inp[2]) ? node19499 : node19496;
														assign node19496 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node19499 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node19502 = (inp[13]) ? node19510 : node19503;
													assign node19503 = (inp[0]) ? node19507 : node19504;
														assign node19504 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node19507 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19510 = (inp[11]) ? 16'b0000001111111111 : node19511;
														assign node19511 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
											assign node19515 = (inp[2]) ? node19529 : node19516;
												assign node19516 = (inp[11]) ? node19522 : node19517;
													assign node19517 = (inp[0]) ? 16'b0000011111111111 : node19518;
														assign node19518 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node19522 = (inp[13]) ? node19526 : node19523;
														assign node19523 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19526 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node19529 = (inp[11]) ? node19537 : node19530;
													assign node19530 = (inp[9]) ? node19534 : node19531;
														assign node19531 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19534 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19537 = (inp[7]) ? node19541 : node19538;
														assign node19538 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19541 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node19544 = (inp[7]) ? node19574 : node19545;
											assign node19545 = (inp[0]) ? node19559 : node19546;
												assign node19546 = (inp[13]) ? node19554 : node19547;
													assign node19547 = (inp[9]) ? node19551 : node19548;
														assign node19548 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node19551 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19554 = (inp[15]) ? node19556 : 16'b0000011111111111;
														assign node19556 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19559 = (inp[2]) ? node19567 : node19560;
													assign node19560 = (inp[13]) ? node19564 : node19561;
														assign node19561 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19564 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19567 = (inp[9]) ? node19571 : node19568;
														assign node19568 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19571 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node19574 = (inp[11]) ? node19590 : node19575;
												assign node19575 = (inp[0]) ? node19583 : node19576;
													assign node19576 = (inp[9]) ? node19580 : node19577;
														assign node19577 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19580 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19583 = (inp[2]) ? node19587 : node19584;
														assign node19584 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19587 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19590 = (inp[0]) ? node19598 : node19591;
													assign node19591 = (inp[9]) ? node19595 : node19592;
														assign node19592 = (inp[2]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node19595 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19598 = (inp[9]) ? node19602 : node19599;
														assign node19599 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19602 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node19605 = (inp[9]) ? node19667 : node19606;
										assign node19606 = (inp[7]) ? node19636 : node19607;
											assign node19607 = (inp[4]) ? node19623 : node19608;
												assign node19608 = (inp[15]) ? node19616 : node19609;
													assign node19609 = (inp[2]) ? node19613 : node19610;
														assign node19610 = (inp[11]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node19613 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19616 = (inp[11]) ? node19620 : node19617;
														assign node19617 = (inp[2]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node19620 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node19623 = (inp[13]) ? node19631 : node19624;
													assign node19624 = (inp[11]) ? node19628 : node19625;
														assign node19625 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node19628 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19631 = (inp[15]) ? 16'b0000000111111111 : node19632;
														assign node19632 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node19636 = (inp[2]) ? node19652 : node19637;
												assign node19637 = (inp[0]) ? node19645 : node19638;
													assign node19638 = (inp[15]) ? node19642 : node19639;
														assign node19639 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19642 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19645 = (inp[13]) ? node19649 : node19646;
														assign node19646 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19649 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19652 = (inp[4]) ? node19660 : node19653;
													assign node19653 = (inp[13]) ? node19657 : node19654;
														assign node19654 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19657 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19660 = (inp[11]) ? node19664 : node19661;
														assign node19661 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19664 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19667 = (inp[15]) ? node19699 : node19668;
											assign node19668 = (inp[2]) ? node19684 : node19669;
												assign node19669 = (inp[4]) ? node19677 : node19670;
													assign node19670 = (inp[0]) ? node19674 : node19671;
														assign node19671 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19674 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19677 = (inp[13]) ? node19681 : node19678;
														assign node19678 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19681 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19684 = (inp[13]) ? node19692 : node19685;
													assign node19685 = (inp[0]) ? node19689 : node19686;
														assign node19686 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19689 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19692 = (inp[11]) ? node19696 : node19693;
														assign node19693 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19696 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node19699 = (inp[7]) ? node19715 : node19700;
												assign node19700 = (inp[11]) ? node19708 : node19701;
													assign node19701 = (inp[0]) ? node19705 : node19702;
														assign node19702 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19705 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node19708 = (inp[0]) ? node19712 : node19709;
														assign node19709 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node19712 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node19715 = (inp[11]) ? node19723 : node19716;
													assign node19716 = (inp[2]) ? node19720 : node19717;
														assign node19717 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node19720 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19723 = (inp[0]) ? node19727 : node19724;
														assign node19724 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19727 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
								assign node19730 = (inp[0]) ? node19854 : node19731;
									assign node19731 = (inp[15]) ? node19793 : node19732;
										assign node19732 = (inp[11]) ? node19762 : node19733;
											assign node19733 = (inp[7]) ? node19747 : node19734;
												assign node19734 = (inp[9]) ? node19742 : node19735;
													assign node19735 = (inp[13]) ? node19739 : node19736;
														assign node19736 = (inp[2]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node19739 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19742 = (inp[14]) ? 16'b0000001111111111 : node19743;
														assign node19743 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node19747 = (inp[13]) ? node19755 : node19748;
													assign node19748 = (inp[14]) ? node19752 : node19749;
														assign node19749 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19752 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19755 = (inp[9]) ? node19759 : node19756;
														assign node19756 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node19759 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node19762 = (inp[7]) ? node19778 : node19763;
												assign node19763 = (inp[9]) ? node19771 : node19764;
													assign node19764 = (inp[14]) ? node19768 : node19765;
														assign node19765 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19768 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19771 = (inp[2]) ? node19775 : node19772;
														assign node19772 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19775 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node19778 = (inp[4]) ? node19786 : node19779;
													assign node19779 = (inp[13]) ? node19783 : node19780;
														assign node19780 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19783 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19786 = (inp[2]) ? node19790 : node19787;
														assign node19787 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node19790 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node19793 = (inp[4]) ? node19823 : node19794;
											assign node19794 = (inp[7]) ? node19810 : node19795;
												assign node19795 = (inp[14]) ? node19803 : node19796;
													assign node19796 = (inp[13]) ? node19800 : node19797;
														assign node19797 = (inp[9]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node19800 = (inp[11]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node19803 = (inp[9]) ? node19807 : node19804;
														assign node19804 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19807 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19810 = (inp[9]) ? node19818 : node19811;
													assign node19811 = (inp[11]) ? node19815 : node19812;
														assign node19812 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19815 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19818 = (inp[11]) ? 16'b0000000011111111 : node19819;
														assign node19819 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node19823 = (inp[13]) ? node19839 : node19824;
												assign node19824 = (inp[7]) ? node19832 : node19825;
													assign node19825 = (inp[9]) ? node19829 : node19826;
														assign node19826 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19829 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19832 = (inp[11]) ? node19836 : node19833;
														assign node19833 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19836 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node19839 = (inp[14]) ? node19847 : node19840;
													assign node19840 = (inp[7]) ? node19844 : node19841;
														assign node19841 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node19844 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19847 = (inp[9]) ? node19851 : node19848;
														assign node19848 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19851 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
									assign node19854 = (inp[7]) ? node19910 : node19855;
										assign node19855 = (inp[15]) ? node19883 : node19856;
											assign node19856 = (inp[13]) ? node19872 : node19857;
												assign node19857 = (inp[9]) ? node19865 : node19858;
													assign node19858 = (inp[11]) ? node19862 : node19859;
														assign node19859 = (inp[4]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node19862 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node19865 = (inp[11]) ? node19869 : node19866;
														assign node19866 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19869 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19872 = (inp[4]) ? node19876 : node19873;
													assign node19873 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node19876 = (inp[9]) ? node19880 : node19877;
														assign node19877 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19880 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node19883 = (inp[11]) ? node19897 : node19884;
												assign node19884 = (inp[4]) ? node19892 : node19885;
													assign node19885 = (inp[9]) ? node19889 : node19886;
														assign node19886 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19889 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19892 = (inp[2]) ? 16'b0000000011111111 : node19893;
														assign node19893 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node19897 = (inp[14]) ? node19903 : node19898;
													assign node19898 = (inp[2]) ? 16'b0000000011111111 : node19899;
														assign node19899 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node19903 = (inp[2]) ? node19907 : node19904;
														assign node19904 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19907 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node19910 = (inp[4]) ? node19942 : node19911;
											assign node19911 = (inp[13]) ? node19927 : node19912;
												assign node19912 = (inp[14]) ? node19920 : node19913;
													assign node19913 = (inp[9]) ? node19917 : node19914;
														assign node19914 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node19917 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node19920 = (inp[15]) ? node19924 : node19921;
														assign node19921 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19924 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node19927 = (inp[11]) ? node19935 : node19928;
													assign node19928 = (inp[14]) ? node19932 : node19929;
														assign node19929 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19932 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19935 = (inp[14]) ? node19939 : node19936;
														assign node19936 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node19939 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node19942 = (inp[15]) ? node19958 : node19943;
												assign node19943 = (inp[2]) ? node19951 : node19944;
													assign node19944 = (inp[11]) ? node19948 : node19945;
														assign node19945 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node19948 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node19951 = (inp[9]) ? node19955 : node19952;
														assign node19952 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node19955 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node19958 = (inp[9]) ? node19966 : node19959;
													assign node19959 = (inp[11]) ? node19963 : node19960;
														assign node19960 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node19963 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node19966 = (inp[11]) ? node19970 : node19967;
														assign node19967 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node19970 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
							assign node19973 = (inp[15]) ? node20217 : node19974;
								assign node19974 = (inp[11]) ? node20098 : node19975;
									assign node19975 = (inp[14]) ? node20037 : node19976;
										assign node19976 = (inp[2]) ? node20008 : node19977;
											assign node19977 = (inp[7]) ? node19993 : node19978;
												assign node19978 = (inp[9]) ? node19986 : node19979;
													assign node19979 = (inp[13]) ? node19983 : node19980;
														assign node19980 = (inp[0]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node19983 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node19986 = (inp[13]) ? node19990 : node19987;
														assign node19987 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19990 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
												assign node19993 = (inp[1]) ? node20001 : node19994;
													assign node19994 = (inp[13]) ? node19998 : node19995;
														assign node19995 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node19998 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20001 = (inp[9]) ? node20005 : node20002;
														assign node20002 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20005 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node20008 = (inp[4]) ? node20024 : node20009;
												assign node20009 = (inp[0]) ? node20017 : node20010;
													assign node20010 = (inp[9]) ? node20014 : node20011;
														assign node20011 = (inp[1]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node20014 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node20017 = (inp[7]) ? node20021 : node20018;
														assign node20018 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20021 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20024 = (inp[0]) ? node20030 : node20025;
													assign node20025 = (inp[13]) ? 16'b0000000111111111 : node20026;
														assign node20026 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20030 = (inp[7]) ? node20034 : node20031;
														assign node20031 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20034 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node20037 = (inp[1]) ? node20067 : node20038;
											assign node20038 = (inp[9]) ? node20054 : node20039;
												assign node20039 = (inp[2]) ? node20047 : node20040;
													assign node20040 = (inp[4]) ? node20044 : node20041;
														assign node20041 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20044 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20047 = (inp[13]) ? node20051 : node20048;
														assign node20048 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20051 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20054 = (inp[2]) ? node20062 : node20055;
													assign node20055 = (inp[0]) ? node20059 : node20056;
														assign node20056 = (inp[4]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node20059 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20062 = (inp[7]) ? node20064 : 16'b0000000011111111;
														assign node20064 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node20067 = (inp[4]) ? node20083 : node20068;
												assign node20068 = (inp[0]) ? node20076 : node20069;
													assign node20069 = (inp[13]) ? node20073 : node20070;
														assign node20070 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20073 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20076 = (inp[9]) ? node20080 : node20077;
														assign node20077 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20080 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20083 = (inp[9]) ? node20091 : node20084;
													assign node20084 = (inp[2]) ? node20088 : node20085;
														assign node20085 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node20088 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node20091 = (inp[2]) ? node20095 : node20092;
														assign node20092 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node20095 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node20098 = (inp[7]) ? node20156 : node20099;
										assign node20099 = (inp[1]) ? node20129 : node20100;
											assign node20100 = (inp[4]) ? node20116 : node20101;
												assign node20101 = (inp[2]) ? node20109 : node20102;
													assign node20102 = (inp[0]) ? node20106 : node20103;
														assign node20103 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20106 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20109 = (inp[0]) ? node20113 : node20110;
														assign node20110 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node20113 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node20116 = (inp[13]) ? node20124 : node20117;
													assign node20117 = (inp[14]) ? node20121 : node20118;
														assign node20118 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20121 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20124 = (inp[0]) ? 16'b0000000001111111 : node20125;
														assign node20125 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node20129 = (inp[2]) ? node20141 : node20130;
												assign node20130 = (inp[14]) ? node20136 : node20131;
													assign node20131 = (inp[4]) ? 16'b0000000111111111 : node20132;
														assign node20132 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20136 = (inp[4]) ? 16'b0000000011111111 : node20137;
														assign node20137 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20141 = (inp[13]) ? node20149 : node20142;
													assign node20142 = (inp[4]) ? node20146 : node20143;
														assign node20143 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20146 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20149 = (inp[4]) ? node20153 : node20150;
														assign node20150 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node20153 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node20156 = (inp[2]) ? node20186 : node20157;
											assign node20157 = (inp[14]) ? node20173 : node20158;
												assign node20158 = (inp[1]) ? node20166 : node20159;
													assign node20159 = (inp[0]) ? node20163 : node20160;
														assign node20160 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20163 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20166 = (inp[4]) ? node20170 : node20167;
														assign node20167 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20170 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20173 = (inp[0]) ? node20181 : node20174;
													assign node20174 = (inp[13]) ? node20178 : node20175;
														assign node20175 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node20178 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20181 = (inp[4]) ? node20183 : 16'b0000000001111111;
														assign node20183 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20186 = (inp[13]) ? node20202 : node20187;
												assign node20187 = (inp[4]) ? node20195 : node20188;
													assign node20188 = (inp[0]) ? node20192 : node20189;
														assign node20189 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20192 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20195 = (inp[9]) ? node20199 : node20196;
														assign node20196 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20199 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20202 = (inp[4]) ? node20210 : node20203;
													assign node20203 = (inp[9]) ? node20207 : node20204;
														assign node20204 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20207 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20210 = (inp[9]) ? node20214 : node20211;
														assign node20211 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node20214 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node20217 = (inp[4]) ? node20343 : node20218;
									assign node20218 = (inp[7]) ? node20280 : node20219;
										assign node20219 = (inp[2]) ? node20249 : node20220;
											assign node20220 = (inp[0]) ? node20234 : node20221;
												assign node20221 = (inp[13]) ? node20227 : node20222;
													assign node20222 = (inp[1]) ? 16'b0000001111111111 : node20223;
														assign node20223 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node20227 = (inp[14]) ? node20231 : node20228;
														assign node20228 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20231 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20234 = (inp[9]) ? node20242 : node20235;
													assign node20235 = (inp[1]) ? node20239 : node20236;
														assign node20236 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20239 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20242 = (inp[11]) ? node20246 : node20243;
														assign node20243 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20246 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20249 = (inp[9]) ? node20265 : node20250;
												assign node20250 = (inp[0]) ? node20258 : node20251;
													assign node20251 = (inp[11]) ? node20255 : node20252;
														assign node20252 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node20255 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20258 = (inp[13]) ? node20262 : node20259;
														assign node20259 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20262 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20265 = (inp[13]) ? node20273 : node20266;
													assign node20266 = (inp[14]) ? node20270 : node20267;
														assign node20267 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20270 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20273 = (inp[14]) ? node20277 : node20274;
														assign node20274 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20277 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node20280 = (inp[9]) ? node20312 : node20281;
											assign node20281 = (inp[0]) ? node20297 : node20282;
												assign node20282 = (inp[2]) ? node20290 : node20283;
													assign node20283 = (inp[14]) ? node20287 : node20284;
														assign node20284 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20287 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20290 = (inp[14]) ? node20294 : node20291;
														assign node20291 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20294 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20297 = (inp[1]) ? node20305 : node20298;
													assign node20298 = (inp[13]) ? node20302 : node20299;
														assign node20299 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20302 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node20305 = (inp[14]) ? node20309 : node20306;
														assign node20306 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20309 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node20312 = (inp[11]) ? node20328 : node20313;
												assign node20313 = (inp[0]) ? node20321 : node20314;
													assign node20314 = (inp[2]) ? node20318 : node20315;
														assign node20315 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20318 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20321 = (inp[14]) ? node20325 : node20322;
														assign node20322 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20325 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node20328 = (inp[13]) ? node20336 : node20329;
													assign node20329 = (inp[1]) ? node20333 : node20330;
														assign node20330 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node20333 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20336 = (inp[0]) ? node20340 : node20337;
														assign node20337 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20340 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node20343 = (inp[7]) ? node20407 : node20344;
										assign node20344 = (inp[14]) ? node20376 : node20345;
											assign node20345 = (inp[1]) ? node20361 : node20346;
												assign node20346 = (inp[11]) ? node20354 : node20347;
													assign node20347 = (inp[0]) ? node20351 : node20348;
														assign node20348 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20351 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20354 = (inp[0]) ? node20358 : node20355;
														assign node20355 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20358 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20361 = (inp[9]) ? node20369 : node20362;
													assign node20362 = (inp[11]) ? node20366 : node20363;
														assign node20363 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20366 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20369 = (inp[0]) ? node20373 : node20370;
														assign node20370 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20373 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20376 = (inp[0]) ? node20392 : node20377;
												assign node20377 = (inp[2]) ? node20385 : node20378;
													assign node20378 = (inp[9]) ? node20382 : node20379;
														assign node20379 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20382 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20385 = (inp[9]) ? node20389 : node20386;
														assign node20386 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20389 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20392 = (inp[11]) ? node20400 : node20393;
													assign node20393 = (inp[1]) ? node20397 : node20394;
														assign node20394 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20397 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20400 = (inp[2]) ? node20404 : node20401;
														assign node20401 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20404 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node20407 = (inp[1]) ? node20433 : node20408;
											assign node20408 = (inp[13]) ? node20418 : node20409;
												assign node20409 = (inp[2]) ? 16'b0000000001111111 : node20410;
													assign node20410 = (inp[14]) ? node20414 : node20411;
														assign node20411 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20414 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20418 = (inp[9]) ? node20426 : node20419;
													assign node20419 = (inp[11]) ? node20423 : node20420;
														assign node20420 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20423 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20426 = (inp[0]) ? node20430 : node20427;
														assign node20427 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20430 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node20433 = (inp[2]) ? node20449 : node20434;
												assign node20434 = (inp[14]) ? node20442 : node20435;
													assign node20435 = (inp[11]) ? node20439 : node20436;
														assign node20436 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20439 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20442 = (inp[11]) ? node20446 : node20443;
														assign node20443 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20446 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node20449 = (inp[9]) ? node20457 : node20450;
													assign node20450 = (inp[11]) ? node20454 : node20451;
														assign node20451 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20454 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20457 = (inp[13]) ? node20459 : 16'b0000000000011111;
														assign node20459 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
						assign node20462 = (inp[7]) ? node20942 : node20463;
							assign node20463 = (inp[15]) ? node20705 : node20464;
								assign node20464 = (inp[9]) ? node20588 : node20465;
									assign node20465 = (inp[0]) ? node20527 : node20466;
										assign node20466 = (inp[1]) ? node20498 : node20467;
											assign node20467 = (inp[11]) ? node20483 : node20468;
												assign node20468 = (inp[2]) ? node20476 : node20469;
													assign node20469 = (inp[3]) ? node20473 : node20470;
														assign node20470 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node20473 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node20476 = (inp[14]) ? node20480 : node20477;
														assign node20477 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20480 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node20483 = (inp[3]) ? node20491 : node20484;
													assign node20484 = (inp[4]) ? node20488 : node20485;
														assign node20485 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20488 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20491 = (inp[4]) ? node20495 : node20492;
														assign node20492 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20495 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
											assign node20498 = (inp[11]) ? node20514 : node20499;
												assign node20499 = (inp[3]) ? node20507 : node20500;
													assign node20500 = (inp[4]) ? node20504 : node20501;
														assign node20501 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20504 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20507 = (inp[13]) ? node20511 : node20508;
														assign node20508 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20511 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20514 = (inp[14]) ? node20522 : node20515;
													assign node20515 = (inp[4]) ? node20519 : node20516;
														assign node20516 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20519 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20522 = (inp[13]) ? 16'b0000000011111111 : node20523;
														assign node20523 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node20527 = (inp[3]) ? node20559 : node20528;
											assign node20528 = (inp[13]) ? node20544 : node20529;
												assign node20529 = (inp[14]) ? node20537 : node20530;
													assign node20530 = (inp[2]) ? node20534 : node20531;
														assign node20531 = (inp[4]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20534 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20537 = (inp[11]) ? node20541 : node20538;
														assign node20538 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20541 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20544 = (inp[1]) ? node20552 : node20545;
													assign node20545 = (inp[14]) ? node20549 : node20546;
														assign node20546 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20549 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20552 = (inp[14]) ? node20556 : node20553;
														assign node20553 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20556 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20559 = (inp[4]) ? node20573 : node20560;
												assign node20560 = (inp[1]) ? node20566 : node20561;
													assign node20561 = (inp[13]) ? 16'b0000000011111111 : node20562;
														assign node20562 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node20566 = (inp[2]) ? node20570 : node20567;
														assign node20567 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20570 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20573 = (inp[14]) ? node20581 : node20574;
													assign node20574 = (inp[1]) ? node20578 : node20575;
														assign node20575 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node20578 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20581 = (inp[13]) ? node20585 : node20582;
														assign node20582 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20585 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node20588 = (inp[1]) ? node20646 : node20589;
										assign node20589 = (inp[13]) ? node20615 : node20590;
											assign node20590 = (inp[4]) ? node20600 : node20591;
												assign node20591 = (inp[14]) ? 16'b0000000111111111 : node20592;
													assign node20592 = (inp[3]) ? node20596 : node20593;
														assign node20593 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20596 = (inp[2]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node20600 = (inp[2]) ? node20608 : node20601;
													assign node20601 = (inp[14]) ? node20605 : node20602;
														assign node20602 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20605 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20608 = (inp[11]) ? node20612 : node20609;
														assign node20609 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20612 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20615 = (inp[11]) ? node20631 : node20616;
												assign node20616 = (inp[3]) ? node20624 : node20617;
													assign node20617 = (inp[0]) ? node20621 : node20618;
														assign node20618 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20621 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20624 = (inp[14]) ? node20628 : node20625;
														assign node20625 = (inp[4]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node20628 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20631 = (inp[2]) ? node20639 : node20632;
													assign node20632 = (inp[14]) ? node20636 : node20633;
														assign node20633 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20636 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20639 = (inp[0]) ? node20643 : node20640;
														assign node20640 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node20643 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node20646 = (inp[11]) ? node20674 : node20647;
											assign node20647 = (inp[14]) ? node20659 : node20648;
												assign node20648 = (inp[3]) ? node20654 : node20649;
													assign node20649 = (inp[13]) ? 16'b0000000111111111 : node20650;
														assign node20650 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20654 = (inp[2]) ? 16'b0000000001111111 : node20655;
														assign node20655 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node20659 = (inp[2]) ? node20667 : node20660;
													assign node20660 = (inp[0]) ? node20664 : node20661;
														assign node20661 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20664 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20667 = (inp[13]) ? node20671 : node20668;
														assign node20668 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20671 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20674 = (inp[4]) ? node20690 : node20675;
												assign node20675 = (inp[13]) ? node20683 : node20676;
													assign node20676 = (inp[14]) ? node20680 : node20677;
														assign node20677 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20680 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20683 = (inp[0]) ? node20687 : node20684;
														assign node20684 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node20687 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20690 = (inp[3]) ? node20698 : node20691;
													assign node20691 = (inp[0]) ? node20695 : node20692;
														assign node20692 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20695 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20698 = (inp[2]) ? node20702 : node20699;
														assign node20699 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20702 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000111111;
								assign node20705 = (inp[0]) ? node20827 : node20706;
									assign node20706 = (inp[9]) ? node20766 : node20707;
										assign node20707 = (inp[1]) ? node20737 : node20708;
											assign node20708 = (inp[14]) ? node20722 : node20709;
												assign node20709 = (inp[13]) ? node20715 : node20710;
													assign node20710 = (inp[2]) ? node20712 : 16'b0000001111111111;
														assign node20712 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20715 = (inp[3]) ? node20719 : node20716;
														assign node20716 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20719 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20722 = (inp[4]) ? node20730 : node20723;
													assign node20723 = (inp[2]) ? node20727 : node20724;
														assign node20724 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20727 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20730 = (inp[13]) ? node20734 : node20731;
														assign node20731 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20734 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20737 = (inp[11]) ? node20751 : node20738;
												assign node20738 = (inp[13]) ? node20744 : node20739;
													assign node20739 = (inp[14]) ? node20741 : 16'b0000000111111111;
														assign node20741 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20744 = (inp[2]) ? node20748 : node20745;
														assign node20745 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20748 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node20751 = (inp[13]) ? node20759 : node20752;
													assign node20752 = (inp[2]) ? node20756 : node20753;
														assign node20753 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20756 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20759 = (inp[4]) ? node20763 : node20760;
														assign node20760 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20763 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node20766 = (inp[13]) ? node20798 : node20767;
											assign node20767 = (inp[2]) ? node20783 : node20768;
												assign node20768 = (inp[1]) ? node20776 : node20769;
													assign node20769 = (inp[3]) ? node20773 : node20770;
														assign node20770 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20773 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20776 = (inp[4]) ? node20780 : node20777;
														assign node20777 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20780 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node20783 = (inp[3]) ? node20791 : node20784;
													assign node20784 = (inp[11]) ? node20788 : node20785;
														assign node20785 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20788 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20791 = (inp[14]) ? node20795 : node20792;
														assign node20792 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20795 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20798 = (inp[4]) ? node20814 : node20799;
												assign node20799 = (inp[3]) ? node20807 : node20800;
													assign node20800 = (inp[1]) ? node20804 : node20801;
														assign node20801 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20804 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20807 = (inp[14]) ? node20811 : node20808;
														assign node20808 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20811 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20814 = (inp[2]) ? node20822 : node20815;
													assign node20815 = (inp[11]) ? node20819 : node20816;
														assign node20816 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node20819 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node20822 = (inp[14]) ? node20824 : 16'b0000000000111111;
														assign node20824 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node20827 = (inp[11]) ? node20887 : node20828;
										assign node20828 = (inp[4]) ? node20858 : node20829;
											assign node20829 = (inp[1]) ? node20843 : node20830;
												assign node20830 = (inp[13]) ? node20838 : node20831;
													assign node20831 = (inp[9]) ? node20835 : node20832;
														assign node20832 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20835 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20838 = (inp[2]) ? node20840 : 16'b0000000111111111;
														assign node20840 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20843 = (inp[14]) ? node20851 : node20844;
													assign node20844 = (inp[2]) ? node20848 : node20845;
														assign node20845 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20848 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20851 = (inp[13]) ? node20855 : node20852;
														assign node20852 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20855 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node20858 = (inp[13]) ? node20874 : node20859;
												assign node20859 = (inp[9]) ? node20867 : node20860;
													assign node20860 = (inp[14]) ? node20864 : node20861;
														assign node20861 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20864 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node20867 = (inp[3]) ? node20871 : node20868;
														assign node20868 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node20871 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node20874 = (inp[3]) ? node20882 : node20875;
													assign node20875 = (inp[2]) ? node20879 : node20876;
														assign node20876 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node20879 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node20882 = (inp[14]) ? node20884 : 16'b0000000000111111;
														assign node20884 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node20887 = (inp[14]) ? node20913 : node20888;
											assign node20888 = (inp[2]) ? node20900 : node20889;
												assign node20889 = (inp[3]) ? node20895 : node20890;
													assign node20890 = (inp[4]) ? 16'b0000000011111111 : node20891;
														assign node20891 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20895 = (inp[9]) ? 16'b0000000000111111 : node20896;
														assign node20896 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20900 = (inp[3]) ? node20906 : node20901;
													assign node20901 = (inp[9]) ? node20903 : 16'b0000000001111111;
														assign node20903 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node20906 = (inp[13]) ? node20910 : node20907;
														assign node20907 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20910 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node20913 = (inp[13]) ? node20927 : node20914;
												assign node20914 = (inp[2]) ? node20920 : node20915;
													assign node20915 = (inp[4]) ? node20917 : 16'b0000000001111111;
														assign node20917 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node20920 = (inp[3]) ? node20924 : node20921;
														assign node20921 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20924 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node20927 = (inp[9]) ? node20935 : node20928;
													assign node20928 = (inp[4]) ? node20932 : node20929;
														assign node20929 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node20932 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node20935 = (inp[2]) ? node20939 : node20936;
														assign node20936 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node20939 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000011111;
							assign node20942 = (inp[9]) ? node21182 : node20943;
								assign node20943 = (inp[2]) ? node21065 : node20944;
									assign node20944 = (inp[3]) ? node21004 : node20945;
										assign node20945 = (inp[13]) ? node20977 : node20946;
											assign node20946 = (inp[1]) ? node20962 : node20947;
												assign node20947 = (inp[15]) ? node20955 : node20948;
													assign node20948 = (inp[11]) ? node20952 : node20949;
														assign node20949 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node20952 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node20955 = (inp[11]) ? node20959 : node20956;
														assign node20956 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node20959 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node20962 = (inp[4]) ? node20970 : node20963;
													assign node20963 = (inp[11]) ? node20967 : node20964;
														assign node20964 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20967 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20970 = (inp[11]) ? node20974 : node20971;
														assign node20971 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node20974 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node20977 = (inp[1]) ? node20991 : node20978;
												assign node20978 = (inp[0]) ? node20986 : node20979;
													assign node20979 = (inp[15]) ? node20983 : node20980;
														assign node20980 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node20983 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node20986 = (inp[15]) ? node20988 : 16'b0000000011111111;
														assign node20988 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node20991 = (inp[14]) ? node20997 : node20992;
													assign node20992 = (inp[0]) ? node20994 : 16'b0000000011111111;
														assign node20994 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node20997 = (inp[15]) ? node21001 : node20998;
														assign node20998 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21001 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node21004 = (inp[4]) ? node21034 : node21005;
											assign node21005 = (inp[11]) ? node21021 : node21006;
												assign node21006 = (inp[14]) ? node21014 : node21007;
													assign node21007 = (inp[13]) ? node21011 : node21008;
														assign node21008 = (inp[15]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node21011 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21014 = (inp[0]) ? node21018 : node21015;
														assign node21015 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21018 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21021 = (inp[14]) ? node21027 : node21022;
													assign node21022 = (inp[13]) ? 16'b0000000001111111 : node21023;
														assign node21023 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21027 = (inp[1]) ? node21031 : node21028;
														assign node21028 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21031 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21034 = (inp[1]) ? node21050 : node21035;
												assign node21035 = (inp[14]) ? node21043 : node21036;
													assign node21036 = (inp[13]) ? node21040 : node21037;
														assign node21037 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21040 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21043 = (inp[15]) ? node21047 : node21044;
														assign node21044 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21047 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21050 = (inp[11]) ? node21058 : node21051;
													assign node21051 = (inp[15]) ? node21055 : node21052;
														assign node21052 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21055 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21058 = (inp[14]) ? node21062 : node21059;
														assign node21059 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21062 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node21065 = (inp[0]) ? node21127 : node21066;
										assign node21066 = (inp[15]) ? node21096 : node21067;
											assign node21067 = (inp[4]) ? node21083 : node21068;
												assign node21068 = (inp[14]) ? node21076 : node21069;
													assign node21069 = (inp[1]) ? node21073 : node21070;
														assign node21070 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21073 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21076 = (inp[1]) ? node21080 : node21077;
														assign node21077 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21080 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21083 = (inp[13]) ? node21089 : node21084;
													assign node21084 = (inp[11]) ? 16'b0000000011111111 : node21085;
														assign node21085 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21089 = (inp[11]) ? node21093 : node21090;
														assign node21090 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21093 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21096 = (inp[3]) ? node21112 : node21097;
												assign node21097 = (inp[14]) ? node21105 : node21098;
													assign node21098 = (inp[4]) ? node21102 : node21099;
														assign node21099 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node21102 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21105 = (inp[11]) ? node21109 : node21106;
														assign node21106 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21109 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21112 = (inp[13]) ? node21120 : node21113;
													assign node21113 = (inp[11]) ? node21117 : node21114;
														assign node21114 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21117 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node21120 = (inp[4]) ? node21124 : node21121;
														assign node21121 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node21124 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node21127 = (inp[13]) ? node21157 : node21128;
											assign node21128 = (inp[3]) ? node21142 : node21129;
												assign node21129 = (inp[14]) ? node21137 : node21130;
													assign node21130 = (inp[11]) ? node21134 : node21131;
														assign node21131 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21134 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21137 = (inp[11]) ? node21139 : 16'b0000000001111111;
														assign node21139 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node21142 = (inp[1]) ? node21150 : node21143;
													assign node21143 = (inp[15]) ? node21147 : node21144;
														assign node21144 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21147 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21150 = (inp[11]) ? node21154 : node21151;
														assign node21151 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node21154 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21157 = (inp[1]) ? node21171 : node21158;
												assign node21158 = (inp[4]) ? node21166 : node21159;
													assign node21159 = (inp[11]) ? node21163 : node21160;
														assign node21160 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21163 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node21166 = (inp[3]) ? node21168 : 16'b0000000000111111;
														assign node21168 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21171 = (inp[3]) ? node21177 : node21172;
													assign node21172 = (inp[15]) ? node21174 : 16'b0000000000111111;
														assign node21174 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21177 = (inp[4]) ? 16'b0000000000001111 : node21178;
														assign node21178 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node21182 = (inp[1]) ? node21300 : node21183;
									assign node21183 = (inp[4]) ? node21237 : node21184;
										assign node21184 = (inp[13]) ? node21210 : node21185;
											assign node21185 = (inp[0]) ? node21199 : node21186;
												assign node21186 = (inp[3]) ? node21194 : node21187;
													assign node21187 = (inp[15]) ? node21191 : node21188;
														assign node21188 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node21191 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node21194 = (inp[11]) ? 16'b0000000011111111 : node21195;
														assign node21195 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
												assign node21199 = (inp[3]) ? node21205 : node21200;
													assign node21200 = (inp[11]) ? node21202 : 16'b0000000011111111;
														assign node21202 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node21205 = (inp[2]) ? 16'b0000000001111111 : node21206;
														assign node21206 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21210 = (inp[11]) ? node21224 : node21211;
												assign node21211 = (inp[3]) ? node21219 : node21212;
													assign node21212 = (inp[14]) ? node21216 : node21213;
														assign node21213 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21216 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21219 = (inp[0]) ? 16'b0000000000111111 : node21220;
														assign node21220 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21224 = (inp[3]) ? node21232 : node21225;
													assign node21225 = (inp[2]) ? node21229 : node21226;
														assign node21226 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21229 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21232 = (inp[2]) ? 16'b0000000000011111 : node21233;
														assign node21233 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node21237 = (inp[3]) ? node21269 : node21238;
											assign node21238 = (inp[2]) ? node21254 : node21239;
												assign node21239 = (inp[15]) ? node21247 : node21240;
													assign node21240 = (inp[13]) ? node21244 : node21241;
														assign node21241 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21244 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node21247 = (inp[14]) ? node21251 : node21248;
														assign node21248 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21251 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21254 = (inp[15]) ? node21262 : node21255;
													assign node21255 = (inp[14]) ? node21259 : node21256;
														assign node21256 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21259 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21262 = (inp[11]) ? node21266 : node21263;
														assign node21263 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21266 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node21269 = (inp[0]) ? node21285 : node21270;
												assign node21270 = (inp[14]) ? node21278 : node21271;
													assign node21271 = (inp[15]) ? node21275 : node21272;
														assign node21272 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21275 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21278 = (inp[2]) ? node21282 : node21279;
														assign node21279 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node21282 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21285 = (inp[11]) ? node21293 : node21286;
													assign node21286 = (inp[14]) ? node21290 : node21287;
														assign node21287 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node21290 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node21293 = (inp[13]) ? node21297 : node21294;
														assign node21294 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21297 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node21300 = (inp[11]) ? node21360 : node21301;
										assign node21301 = (inp[13]) ? node21333 : node21302;
											assign node21302 = (inp[14]) ? node21318 : node21303;
												assign node21303 = (inp[3]) ? node21311 : node21304;
													assign node21304 = (inp[0]) ? node21308 : node21305;
														assign node21305 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21308 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21311 = (inp[15]) ? node21315 : node21312;
														assign node21312 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21315 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node21318 = (inp[0]) ? node21326 : node21319;
													assign node21319 = (inp[15]) ? node21323 : node21320;
														assign node21320 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21323 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21326 = (inp[4]) ? node21330 : node21327;
														assign node21327 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21330 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21333 = (inp[15]) ? node21349 : node21334;
												assign node21334 = (inp[2]) ? node21342 : node21335;
													assign node21335 = (inp[14]) ? node21339 : node21336;
														assign node21336 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node21339 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21342 = (inp[3]) ? node21346 : node21343;
														assign node21343 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21346 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21349 = (inp[0]) ? node21355 : node21350;
													assign node21350 = (inp[4]) ? node21352 : 16'b0000000000111111;
														assign node21352 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21355 = (inp[4]) ? node21357 : 16'b0000000000011111;
														assign node21357 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000111111;
										assign node21360 = (inp[4]) ? node21390 : node21361;
											assign node21361 = (inp[14]) ? node21375 : node21362;
												assign node21362 = (inp[3]) ? node21370 : node21363;
													assign node21363 = (inp[0]) ? node21367 : node21364;
														assign node21364 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21367 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21370 = (inp[2]) ? node21372 : 16'b0000000000111111;
														assign node21372 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node21375 = (inp[15]) ? node21383 : node21376;
													assign node21376 = (inp[2]) ? node21380 : node21377;
														assign node21377 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node21380 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21383 = (inp[2]) ? node21387 : node21384;
														assign node21384 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21387 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node21390 = (inp[3]) ? node21404 : node21391;
												assign node21391 = (inp[13]) ? node21397 : node21392;
													assign node21392 = (inp[14]) ? node21394 : 16'b0000000000111111;
														assign node21394 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21397 = (inp[15]) ? node21401 : node21398;
														assign node21398 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21401 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node21404 = (inp[15]) ? node21412 : node21405;
													assign node21405 = (inp[0]) ? node21409 : node21406;
														assign node21406 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21409 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000011111;
													assign node21412 = (inp[2]) ? node21416 : node21413;
														assign node21413 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node21416 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000001111;
					assign node21419 = (inp[11]) ? node22403 : node21420;
						assign node21420 = (inp[8]) ? node21906 : node21421;
							assign node21421 = (inp[0]) ? node21663 : node21422;
								assign node21422 = (inp[9]) ? node21544 : node21423;
									assign node21423 = (inp[7]) ? node21481 : node21424;
										assign node21424 = (inp[15]) ? node21452 : node21425;
											assign node21425 = (inp[3]) ? node21439 : node21426;
												assign node21426 = (inp[4]) ? node21434 : node21427;
													assign node21427 = (inp[2]) ? node21431 : node21428;
														assign node21428 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node21431 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node21434 = (inp[1]) ? 16'b0000001111111111 : node21435;
														assign node21435 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node21439 = (inp[1]) ? node21447 : node21440;
													assign node21440 = (inp[4]) ? node21444 : node21441;
														assign node21441 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21444 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21447 = (inp[14]) ? node21449 : 16'b0000001111111111;
														assign node21449 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node21452 = (inp[1]) ? node21468 : node21453;
												assign node21453 = (inp[2]) ? node21461 : node21454;
													assign node21454 = (inp[14]) ? node21458 : node21455;
														assign node21455 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21458 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21461 = (inp[4]) ? node21465 : node21462;
														assign node21462 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node21465 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21468 = (inp[3]) ? node21476 : node21469;
													assign node21469 = (inp[2]) ? node21473 : node21470;
														assign node21470 = (inp[14]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node21473 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node21476 = (inp[2]) ? node21478 : 16'b0000000011111111;
														assign node21478 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
										assign node21481 = (inp[3]) ? node21513 : node21482;
											assign node21482 = (inp[2]) ? node21498 : node21483;
												assign node21483 = (inp[4]) ? node21491 : node21484;
													assign node21484 = (inp[1]) ? node21488 : node21485;
														assign node21485 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21488 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21491 = (inp[13]) ? node21495 : node21492;
														assign node21492 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21495 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21498 = (inp[15]) ? node21506 : node21499;
													assign node21499 = (inp[4]) ? node21503 : node21500;
														assign node21500 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21503 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21506 = (inp[14]) ? node21510 : node21507;
														assign node21507 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21510 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21513 = (inp[15]) ? node21529 : node21514;
												assign node21514 = (inp[4]) ? node21522 : node21515;
													assign node21515 = (inp[1]) ? node21519 : node21516;
														assign node21516 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21519 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node21522 = (inp[13]) ? node21526 : node21523;
														assign node21523 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21526 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21529 = (inp[2]) ? node21537 : node21530;
													assign node21530 = (inp[1]) ? node21534 : node21531;
														assign node21531 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node21534 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21537 = (inp[13]) ? node21541 : node21538;
														assign node21538 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21541 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node21544 = (inp[15]) ? node21606 : node21545;
										assign node21545 = (inp[7]) ? node21577 : node21546;
											assign node21546 = (inp[3]) ? node21562 : node21547;
												assign node21547 = (inp[2]) ? node21555 : node21548;
													assign node21548 = (inp[1]) ? node21552 : node21549;
														assign node21549 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21552 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21555 = (inp[14]) ? node21559 : node21556;
														assign node21556 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21559 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21562 = (inp[2]) ? node21570 : node21563;
													assign node21563 = (inp[1]) ? node21567 : node21564;
														assign node21564 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21567 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21570 = (inp[4]) ? node21574 : node21571;
														assign node21571 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21574 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21577 = (inp[13]) ? node21591 : node21578;
												assign node21578 = (inp[1]) ? node21584 : node21579;
													assign node21579 = (inp[14]) ? node21581 : 16'b0000000111111111;
														assign node21581 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21584 = (inp[3]) ? node21588 : node21585;
														assign node21585 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21588 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21591 = (inp[4]) ? node21599 : node21592;
													assign node21592 = (inp[1]) ? node21596 : node21593;
														assign node21593 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21596 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21599 = (inp[14]) ? node21603 : node21600;
														assign node21600 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21603 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node21606 = (inp[14]) ? node21636 : node21607;
											assign node21607 = (inp[13]) ? node21621 : node21608;
												assign node21608 = (inp[4]) ? node21614 : node21609;
													assign node21609 = (inp[7]) ? 16'b0000000111111111 : node21610;
														assign node21610 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21614 = (inp[7]) ? node21618 : node21615;
														assign node21615 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21618 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21621 = (inp[3]) ? node21629 : node21622;
													assign node21622 = (inp[2]) ? node21626 : node21623;
														assign node21623 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21626 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21629 = (inp[1]) ? node21633 : node21630;
														assign node21630 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21633 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21636 = (inp[4]) ? node21652 : node21637;
												assign node21637 = (inp[2]) ? node21645 : node21638;
													assign node21638 = (inp[13]) ? node21642 : node21639;
														assign node21639 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node21642 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21645 = (inp[3]) ? node21649 : node21646;
														assign node21646 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21649 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21652 = (inp[2]) ? node21660 : node21653;
													assign node21653 = (inp[7]) ? node21657 : node21654;
														assign node21654 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21657 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21660 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node21663 = (inp[13]) ? node21787 : node21664;
									assign node21664 = (inp[15]) ? node21726 : node21665;
										assign node21665 = (inp[2]) ? node21697 : node21666;
											assign node21666 = (inp[1]) ? node21682 : node21667;
												assign node21667 = (inp[7]) ? node21675 : node21668;
													assign node21668 = (inp[4]) ? node21672 : node21669;
														assign node21669 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21672 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21675 = (inp[14]) ? node21679 : node21676;
														assign node21676 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21679 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21682 = (inp[4]) ? node21690 : node21683;
													assign node21683 = (inp[7]) ? node21687 : node21684;
														assign node21684 = (inp[3]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node21687 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21690 = (inp[7]) ? node21694 : node21691;
														assign node21691 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21694 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21697 = (inp[3]) ? node21713 : node21698;
												assign node21698 = (inp[1]) ? node21706 : node21699;
													assign node21699 = (inp[9]) ? node21703 : node21700;
														assign node21700 = (inp[4]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21703 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21706 = (inp[4]) ? node21710 : node21707;
														assign node21707 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21710 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21713 = (inp[1]) ? node21721 : node21714;
													assign node21714 = (inp[14]) ? node21718 : node21715;
														assign node21715 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21718 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21721 = (inp[7]) ? 16'b0000000001111111 : node21722;
														assign node21722 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node21726 = (inp[14]) ? node21756 : node21727;
											assign node21727 = (inp[1]) ? node21741 : node21728;
												assign node21728 = (inp[2]) ? node21736 : node21729;
													assign node21729 = (inp[7]) ? node21733 : node21730;
														assign node21730 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21733 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21736 = (inp[7]) ? 16'b0000000001111111 : node21737;
														assign node21737 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node21741 = (inp[7]) ? node21749 : node21742;
													assign node21742 = (inp[9]) ? node21746 : node21743;
														assign node21743 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21746 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21749 = (inp[4]) ? node21753 : node21750;
														assign node21750 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21753 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21756 = (inp[9]) ? node21772 : node21757;
												assign node21757 = (inp[3]) ? node21765 : node21758;
													assign node21758 = (inp[7]) ? node21762 : node21759;
														assign node21759 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21762 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21765 = (inp[1]) ? node21769 : node21766;
														assign node21766 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21769 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21772 = (inp[2]) ? node21780 : node21773;
													assign node21773 = (inp[7]) ? node21777 : node21774;
														assign node21774 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21777 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21780 = (inp[1]) ? node21784 : node21781;
														assign node21781 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21784 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
									assign node21787 = (inp[9]) ? node21845 : node21788;
										assign node21788 = (inp[7]) ? node21816 : node21789;
											assign node21789 = (inp[14]) ? node21803 : node21790;
												assign node21790 = (inp[15]) ? node21796 : node21791;
													assign node21791 = (inp[3]) ? 16'b0000000111111111 : node21792;
														assign node21792 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21796 = (inp[1]) ? node21800 : node21797;
														assign node21797 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21800 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21803 = (inp[1]) ? node21809 : node21804;
													assign node21804 = (inp[3]) ? node21806 : 16'b0000000111111111;
														assign node21806 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21809 = (inp[4]) ? node21813 : node21810;
														assign node21810 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node21813 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node21816 = (inp[1]) ? node21832 : node21817;
												assign node21817 = (inp[2]) ? node21825 : node21818;
													assign node21818 = (inp[14]) ? node21822 : node21819;
														assign node21819 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21822 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21825 = (inp[3]) ? node21829 : node21826;
														assign node21826 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21829 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node21832 = (inp[4]) ? node21840 : node21833;
													assign node21833 = (inp[2]) ? node21837 : node21834;
														assign node21834 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21837 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21840 = (inp[3]) ? node21842 : 16'b0000000000111111;
														assign node21842 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node21845 = (inp[15]) ? node21877 : node21846;
											assign node21846 = (inp[2]) ? node21862 : node21847;
												assign node21847 = (inp[4]) ? node21855 : node21848;
													assign node21848 = (inp[14]) ? node21852 : node21849;
														assign node21849 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node21852 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21855 = (inp[1]) ? node21859 : node21856;
														assign node21856 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node21859 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node21862 = (inp[14]) ? node21870 : node21863;
													assign node21863 = (inp[1]) ? node21867 : node21864;
														assign node21864 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21867 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21870 = (inp[1]) ? node21874 : node21871;
														assign node21871 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node21874 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node21877 = (inp[3]) ? node21893 : node21878;
												assign node21878 = (inp[1]) ? node21886 : node21879;
													assign node21879 = (inp[4]) ? node21883 : node21880;
														assign node21880 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21883 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node21886 = (inp[14]) ? node21890 : node21887;
														assign node21887 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node21890 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node21893 = (inp[14]) ? node21899 : node21894;
													assign node21894 = (inp[7]) ? node21896 : 16'b0000000000111111;
														assign node21896 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node21899 = (inp[4]) ? node21903 : node21900;
														assign node21900 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node21903 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node21906 = (inp[2]) ? node22156 : node21907;
								assign node21907 = (inp[4]) ? node22031 : node21908;
									assign node21908 = (inp[15]) ? node21968 : node21909;
										assign node21909 = (inp[14]) ? node21939 : node21910;
											assign node21910 = (inp[13]) ? node21924 : node21911;
												assign node21911 = (inp[7]) ? node21919 : node21912;
													assign node21912 = (inp[1]) ? node21916 : node21913;
														assign node21913 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node21916 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node21919 = (inp[0]) ? 16'b0000000111111111 : node21920;
														assign node21920 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node21924 = (inp[1]) ? node21932 : node21925;
													assign node21925 = (inp[7]) ? node21929 : node21926;
														assign node21926 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node21929 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node21932 = (inp[3]) ? node21936 : node21933;
														assign node21933 = (inp[0]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node21936 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node21939 = (inp[3]) ? node21955 : node21940;
												assign node21940 = (inp[7]) ? node21948 : node21941;
													assign node21941 = (inp[13]) ? node21945 : node21942;
														assign node21942 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node21945 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21948 = (inp[9]) ? node21952 : node21949;
														assign node21949 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21952 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node21955 = (inp[0]) ? node21963 : node21956;
													assign node21956 = (inp[13]) ? node21960 : node21957;
														assign node21957 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21960 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21963 = (inp[13]) ? 16'b0000000001111111 : node21964;
														assign node21964 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node21968 = (inp[14]) ? node22000 : node21969;
											assign node21969 = (inp[1]) ? node21985 : node21970;
												assign node21970 = (inp[0]) ? node21978 : node21971;
													assign node21971 = (inp[13]) ? node21975 : node21972;
														assign node21972 = (inp[9]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node21975 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node21978 = (inp[3]) ? node21982 : node21979;
														assign node21979 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node21982 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node21985 = (inp[13]) ? node21993 : node21986;
													assign node21986 = (inp[3]) ? node21990 : node21987;
														assign node21987 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node21990 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node21993 = (inp[9]) ? node21997 : node21994;
														assign node21994 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node21997 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22000 = (inp[3]) ? node22016 : node22001;
												assign node22001 = (inp[1]) ? node22009 : node22002;
													assign node22002 = (inp[13]) ? node22006 : node22003;
														assign node22003 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22006 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22009 = (inp[13]) ? node22013 : node22010;
														assign node22010 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22013 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22016 = (inp[7]) ? node22024 : node22017;
													assign node22017 = (inp[1]) ? node22021 : node22018;
														assign node22018 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node22021 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22024 = (inp[9]) ? node22028 : node22025;
														assign node22025 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22028 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node22031 = (inp[13]) ? node22095 : node22032;
										assign node22032 = (inp[1]) ? node22064 : node22033;
											assign node22033 = (inp[14]) ? node22049 : node22034;
												assign node22034 = (inp[0]) ? node22042 : node22035;
													assign node22035 = (inp[7]) ? node22039 : node22036;
														assign node22036 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node22039 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22042 = (inp[9]) ? node22046 : node22043;
														assign node22043 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22046 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22049 = (inp[9]) ? node22057 : node22050;
													assign node22050 = (inp[3]) ? node22054 : node22051;
														assign node22051 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22054 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22057 = (inp[7]) ? node22061 : node22058;
														assign node22058 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node22061 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node22064 = (inp[15]) ? node22080 : node22065;
												assign node22065 = (inp[7]) ? node22073 : node22066;
													assign node22066 = (inp[3]) ? node22070 : node22067;
														assign node22067 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22070 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node22073 = (inp[3]) ? node22077 : node22074;
														assign node22074 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22077 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22080 = (inp[9]) ? node22088 : node22081;
													assign node22081 = (inp[3]) ? node22085 : node22082;
														assign node22082 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node22085 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22088 = (inp[3]) ? node22092 : node22089;
														assign node22089 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22092 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node22095 = (inp[0]) ? node22125 : node22096;
											assign node22096 = (inp[15]) ? node22110 : node22097;
												assign node22097 = (inp[1]) ? node22105 : node22098;
													assign node22098 = (inp[9]) ? node22102 : node22099;
														assign node22099 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22102 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22105 = (inp[9]) ? 16'b0000000000111111 : node22106;
														assign node22106 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22110 = (inp[3]) ? node22118 : node22111;
													assign node22111 = (inp[1]) ? node22115 : node22112;
														assign node22112 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22115 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22118 = (inp[7]) ? node22122 : node22119;
														assign node22119 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22122 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22125 = (inp[9]) ? node22141 : node22126;
												assign node22126 = (inp[14]) ? node22134 : node22127;
													assign node22127 = (inp[7]) ? node22131 : node22128;
														assign node22128 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node22131 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22134 = (inp[1]) ? node22138 : node22135;
														assign node22135 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node22138 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node22141 = (inp[14]) ? node22149 : node22142;
													assign node22142 = (inp[15]) ? node22146 : node22143;
														assign node22143 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22146 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22149 = (inp[3]) ? node22153 : node22150;
														assign node22150 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22153 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node22156 = (inp[7]) ? node22278 : node22157;
									assign node22157 = (inp[9]) ? node22217 : node22158;
										assign node22158 = (inp[1]) ? node22186 : node22159;
											assign node22159 = (inp[13]) ? node22173 : node22160;
												assign node22160 = (inp[14]) ? node22168 : node22161;
													assign node22161 = (inp[0]) ? node22165 : node22162;
														assign node22162 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22165 = (inp[4]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22168 = (inp[3]) ? node22170 : 16'b0000000111111111;
														assign node22170 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22173 = (inp[15]) ? node22181 : node22174;
													assign node22174 = (inp[0]) ? node22178 : node22175;
														assign node22175 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22178 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22181 = (inp[4]) ? node22183 : 16'b0000000001111111;
														assign node22183 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22186 = (inp[0]) ? node22202 : node22187;
												assign node22187 = (inp[14]) ? node22195 : node22188;
													assign node22188 = (inp[4]) ? node22192 : node22189;
														assign node22189 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22192 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22195 = (inp[13]) ? node22199 : node22196;
														assign node22196 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22199 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22202 = (inp[15]) ? node22210 : node22203;
													assign node22203 = (inp[3]) ? node22207 : node22204;
														assign node22204 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node22207 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22210 = (inp[4]) ? node22214 : node22211;
														assign node22211 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22214 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node22217 = (inp[14]) ? node22247 : node22218;
											assign node22218 = (inp[13]) ? node22234 : node22219;
												assign node22219 = (inp[15]) ? node22227 : node22220;
													assign node22220 = (inp[4]) ? node22224 : node22221;
														assign node22221 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22224 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22227 = (inp[0]) ? node22231 : node22228;
														assign node22228 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22231 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22234 = (inp[4]) ? node22242 : node22235;
													assign node22235 = (inp[15]) ? node22239 : node22236;
														assign node22236 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node22239 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node22242 = (inp[0]) ? 16'b0000000000111111 : node22243;
														assign node22243 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22247 = (inp[4]) ? node22263 : node22248;
												assign node22248 = (inp[15]) ? node22256 : node22249;
													assign node22249 = (inp[1]) ? node22253 : node22250;
														assign node22250 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22253 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22256 = (inp[13]) ? node22260 : node22257;
														assign node22257 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22260 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22263 = (inp[1]) ? node22271 : node22264;
													assign node22264 = (inp[0]) ? node22268 : node22265;
														assign node22265 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node22268 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22271 = (inp[15]) ? node22275 : node22272;
														assign node22272 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22275 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node22278 = (inp[0]) ? node22342 : node22279;
										assign node22279 = (inp[13]) ? node22311 : node22280;
											assign node22280 = (inp[14]) ? node22296 : node22281;
												assign node22281 = (inp[15]) ? node22289 : node22282;
													assign node22282 = (inp[4]) ? node22286 : node22283;
														assign node22283 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22286 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22289 = (inp[1]) ? node22293 : node22290;
														assign node22290 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22293 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22296 = (inp[4]) ? node22304 : node22297;
													assign node22297 = (inp[1]) ? node22301 : node22298;
														assign node22298 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22301 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22304 = (inp[1]) ? node22308 : node22305;
														assign node22305 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22308 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22311 = (inp[3]) ? node22327 : node22312;
												assign node22312 = (inp[4]) ? node22320 : node22313;
													assign node22313 = (inp[15]) ? node22317 : node22314;
														assign node22314 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22317 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node22320 = (inp[9]) ? node22324 : node22321;
														assign node22321 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22324 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22327 = (inp[9]) ? node22335 : node22328;
													assign node22328 = (inp[14]) ? node22332 : node22329;
														assign node22329 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node22332 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22335 = (inp[14]) ? node22339 : node22336;
														assign node22336 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node22339 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node22342 = (inp[9]) ? node22372 : node22343;
											assign node22343 = (inp[3]) ? node22357 : node22344;
												assign node22344 = (inp[13]) ? node22350 : node22345;
													assign node22345 = (inp[14]) ? node22347 : 16'b0000000001111111;
														assign node22347 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22350 = (inp[4]) ? node22354 : node22351;
														assign node22351 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22354 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node22357 = (inp[4]) ? node22365 : node22358;
													assign node22358 = (inp[15]) ? node22362 : node22359;
														assign node22359 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22362 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22365 = (inp[15]) ? node22369 : node22366;
														assign node22366 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22369 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node22372 = (inp[14]) ? node22388 : node22373;
												assign node22373 = (inp[15]) ? node22381 : node22374;
													assign node22374 = (inp[4]) ? node22378 : node22375;
														assign node22375 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22378 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22381 = (inp[4]) ? node22385 : node22382;
														assign node22382 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22385 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000011111;
												assign node22388 = (inp[4]) ? node22396 : node22389;
													assign node22389 = (inp[15]) ? node22393 : node22390;
														assign node22390 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node22393 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node22396 = (inp[3]) ? node22400 : node22397;
														assign node22397 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node22400 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
						assign node22403 = (inp[3]) ? node22897 : node22404;
							assign node22404 = (inp[15]) ? node22650 : node22405;
								assign node22405 = (inp[4]) ? node22531 : node22406;
									assign node22406 = (inp[9]) ? node22468 : node22407;
										assign node22407 = (inp[0]) ? node22437 : node22408;
											assign node22408 = (inp[13]) ? node22424 : node22409;
												assign node22409 = (inp[2]) ? node22417 : node22410;
													assign node22410 = (inp[8]) ? node22414 : node22411;
														assign node22411 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node22414 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22417 = (inp[1]) ? node22421 : node22418;
														assign node22418 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22421 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node22424 = (inp[1]) ? node22432 : node22425;
													assign node22425 = (inp[8]) ? node22429 : node22426;
														assign node22426 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22429 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22432 = (inp[14]) ? 16'b0000000011111111 : node22433;
														assign node22433 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
											assign node22437 = (inp[7]) ? node22453 : node22438;
												assign node22438 = (inp[2]) ? node22446 : node22439;
													assign node22439 = (inp[8]) ? node22443 : node22440;
														assign node22440 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22443 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22446 = (inp[8]) ? node22450 : node22447;
														assign node22447 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22450 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node22453 = (inp[13]) ? node22461 : node22454;
													assign node22454 = (inp[8]) ? node22458 : node22455;
														assign node22455 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22458 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node22461 = (inp[14]) ? node22465 : node22462;
														assign node22462 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22465 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node22468 = (inp[8]) ? node22500 : node22469;
											assign node22469 = (inp[7]) ? node22485 : node22470;
												assign node22470 = (inp[0]) ? node22478 : node22471;
													assign node22471 = (inp[1]) ? node22475 : node22472;
														assign node22472 = (inp[14]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node22475 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22478 = (inp[13]) ? node22482 : node22479;
														assign node22479 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node22482 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22485 = (inp[14]) ? node22493 : node22486;
													assign node22486 = (inp[1]) ? node22490 : node22487;
														assign node22487 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node22490 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22493 = (inp[0]) ? node22497 : node22494;
														assign node22494 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22497 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22500 = (inp[2]) ? node22516 : node22501;
												assign node22501 = (inp[14]) ? node22509 : node22502;
													assign node22502 = (inp[7]) ? node22506 : node22503;
														assign node22503 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22506 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node22509 = (inp[7]) ? node22513 : node22510;
														assign node22510 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22513 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22516 = (inp[0]) ? node22524 : node22517;
													assign node22517 = (inp[1]) ? node22521 : node22518;
														assign node22518 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node22521 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22524 = (inp[1]) ? node22528 : node22525;
														assign node22525 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22528 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node22531 = (inp[13]) ? node22591 : node22532;
										assign node22532 = (inp[7]) ? node22562 : node22533;
											assign node22533 = (inp[14]) ? node22547 : node22534;
												assign node22534 = (inp[1]) ? node22540 : node22535;
													assign node22535 = (inp[9]) ? 16'b0000000111111111 : node22536;
														assign node22536 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node22540 = (inp[0]) ? node22544 : node22541;
														assign node22541 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22544 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node22547 = (inp[2]) ? node22555 : node22548;
													assign node22548 = (inp[8]) ? node22552 : node22549;
														assign node22549 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node22552 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22555 = (inp[8]) ? node22559 : node22556;
														assign node22556 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node22559 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22562 = (inp[1]) ? node22576 : node22563;
												assign node22563 = (inp[2]) ? node22569 : node22564;
													assign node22564 = (inp[9]) ? 16'b0000000011111111 : node22565;
														assign node22565 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22569 = (inp[14]) ? node22573 : node22570;
														assign node22570 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22573 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node22576 = (inp[14]) ? node22584 : node22577;
													assign node22577 = (inp[2]) ? node22581 : node22578;
														assign node22578 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22581 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22584 = (inp[9]) ? node22588 : node22585;
														assign node22585 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22588 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node22591 = (inp[9]) ? node22621 : node22592;
											assign node22592 = (inp[2]) ? node22608 : node22593;
												assign node22593 = (inp[1]) ? node22601 : node22594;
													assign node22594 = (inp[14]) ? node22598 : node22595;
														assign node22595 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22598 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22601 = (inp[14]) ? node22605 : node22602;
														assign node22602 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22605 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22608 = (inp[1]) ? node22614 : node22609;
													assign node22609 = (inp[0]) ? node22611 : 16'b0000000001111111;
														assign node22611 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22614 = (inp[0]) ? node22618 : node22615;
														assign node22615 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22618 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22621 = (inp[8]) ? node22637 : node22622;
												assign node22622 = (inp[1]) ? node22630 : node22623;
													assign node22623 = (inp[0]) ? node22627 : node22624;
														assign node22624 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22627 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22630 = (inp[14]) ? node22634 : node22631;
														assign node22631 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22634 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22637 = (inp[1]) ? node22643 : node22638;
													assign node22638 = (inp[2]) ? node22640 : 16'b0000000001111111;
														assign node22640 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
													assign node22643 = (inp[2]) ? node22647 : node22644;
														assign node22644 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22647 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node22650 = (inp[7]) ? node22772 : node22651;
									assign node22651 = (inp[2]) ? node22709 : node22652;
										assign node22652 = (inp[13]) ? node22682 : node22653;
											assign node22653 = (inp[4]) ? node22667 : node22654;
												assign node22654 = (inp[0]) ? node22660 : node22655;
													assign node22655 = (inp[9]) ? node22657 : 16'b0000001111111111;
														assign node22657 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22660 = (inp[9]) ? node22664 : node22661;
														assign node22661 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22664 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22667 = (inp[0]) ? node22675 : node22668;
													assign node22668 = (inp[14]) ? node22672 : node22669;
														assign node22669 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22672 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node22675 = (inp[1]) ? node22679 : node22676;
														assign node22676 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22679 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node22682 = (inp[1]) ? node22698 : node22683;
												assign node22683 = (inp[4]) ? node22691 : node22684;
													assign node22684 = (inp[0]) ? node22688 : node22685;
														assign node22685 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22688 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22691 = (inp[8]) ? node22695 : node22692;
														assign node22692 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22695 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22698 = (inp[0]) ? node22704 : node22699;
													assign node22699 = (inp[4]) ? node22701 : 16'b0000000001111111;
														assign node22701 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22704 = (inp[4]) ? 16'b0000000000011111 : node22705;
														assign node22705 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node22709 = (inp[9]) ? node22741 : node22710;
											assign node22710 = (inp[4]) ? node22726 : node22711;
												assign node22711 = (inp[1]) ? node22719 : node22712;
													assign node22712 = (inp[13]) ? node22716 : node22713;
														assign node22713 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22716 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22719 = (inp[0]) ? node22723 : node22720;
														assign node22720 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22723 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22726 = (inp[0]) ? node22734 : node22727;
													assign node22727 = (inp[13]) ? node22731 : node22728;
														assign node22728 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22731 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22734 = (inp[14]) ? node22738 : node22735;
														assign node22735 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22738 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22741 = (inp[1]) ? node22757 : node22742;
												assign node22742 = (inp[14]) ? node22750 : node22743;
													assign node22743 = (inp[0]) ? node22747 : node22744;
														assign node22744 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node22747 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22750 = (inp[4]) ? node22754 : node22751;
														assign node22751 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22754 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22757 = (inp[8]) ? node22765 : node22758;
													assign node22758 = (inp[13]) ? node22762 : node22759;
														assign node22759 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node22762 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22765 = (inp[14]) ? node22769 : node22766;
														assign node22766 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node22769 = (inp[13]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node22772 = (inp[0]) ? node22836 : node22773;
										assign node22773 = (inp[14]) ? node22805 : node22774;
											assign node22774 = (inp[8]) ? node22790 : node22775;
												assign node22775 = (inp[4]) ? node22783 : node22776;
													assign node22776 = (inp[1]) ? node22780 : node22777;
														assign node22777 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22780 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22783 = (inp[1]) ? node22787 : node22784;
														assign node22784 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22787 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22790 = (inp[13]) ? node22798 : node22791;
													assign node22791 = (inp[2]) ? node22795 : node22792;
														assign node22792 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node22795 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22798 = (inp[9]) ? node22802 : node22799;
														assign node22799 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22802 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22805 = (inp[2]) ? node22821 : node22806;
												assign node22806 = (inp[4]) ? node22814 : node22807;
													assign node22807 = (inp[8]) ? node22811 : node22808;
														assign node22808 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22811 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22814 = (inp[13]) ? node22818 : node22815;
														assign node22815 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22818 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node22821 = (inp[1]) ? node22829 : node22822;
													assign node22822 = (inp[9]) ? node22826 : node22823;
														assign node22823 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node22826 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node22829 = (inp[9]) ? node22833 : node22830;
														assign node22830 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22833 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node22836 = (inp[2]) ? node22868 : node22837;
											assign node22837 = (inp[4]) ? node22853 : node22838;
												assign node22838 = (inp[9]) ? node22846 : node22839;
													assign node22839 = (inp[14]) ? node22843 : node22840;
														assign node22840 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22843 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22846 = (inp[1]) ? node22850 : node22847;
														assign node22847 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node22850 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node22853 = (inp[13]) ? node22861 : node22854;
													assign node22854 = (inp[8]) ? node22858 : node22855;
														assign node22855 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node22858 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node22861 = (inp[14]) ? node22865 : node22862;
														assign node22862 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22865 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node22868 = (inp[1]) ? node22882 : node22869;
												assign node22869 = (inp[13]) ? node22875 : node22870;
													assign node22870 = (inp[4]) ? node22872 : 16'b0000000000111111;
														assign node22872 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000011111;
													assign node22875 = (inp[9]) ? node22879 : node22876;
														assign node22876 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node22879 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node22882 = (inp[14]) ? node22890 : node22883;
													assign node22883 = (inp[8]) ? node22887 : node22884;
														assign node22884 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node22887 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node22890 = (inp[9]) ? node22894 : node22891;
														assign node22891 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node22894 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node22897 = (inp[15]) ? node23143 : node22898;
								assign node22898 = (inp[14]) ? node23018 : node22899;
									assign node22899 = (inp[7]) ? node22957 : node22900;
										assign node22900 = (inp[1]) ? node22930 : node22901;
											assign node22901 = (inp[4]) ? node22917 : node22902;
												assign node22902 = (inp[8]) ? node22910 : node22903;
													assign node22903 = (inp[0]) ? node22907 : node22904;
														assign node22904 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node22907 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22910 = (inp[2]) ? node22914 : node22911;
														assign node22911 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22914 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node22917 = (inp[0]) ? node22923 : node22918;
													assign node22918 = (inp[2]) ? 16'b0000000011111111 : node22919;
														assign node22919 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node22923 = (inp[13]) ? node22927 : node22924;
														assign node22924 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22927 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node22930 = (inp[9]) ? node22946 : node22931;
												assign node22931 = (inp[0]) ? node22939 : node22932;
													assign node22932 = (inp[13]) ? node22936 : node22933;
														assign node22933 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node22936 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22939 = (inp[13]) ? node22943 : node22940;
														assign node22940 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node22943 = (inp[4]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node22946 = (inp[13]) ? node22952 : node22947;
													assign node22947 = (inp[2]) ? 16'b0000000000111111 : node22948;
														assign node22948 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node22952 = (inp[4]) ? node22954 : 16'b0000000000111111;
														assign node22954 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node22957 = (inp[1]) ? node22989 : node22958;
											assign node22958 = (inp[2]) ? node22974 : node22959;
												assign node22959 = (inp[4]) ? node22967 : node22960;
													assign node22960 = (inp[13]) ? node22964 : node22961;
														assign node22961 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node22964 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node22967 = (inp[13]) ? node22971 : node22968;
														assign node22968 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node22971 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node22974 = (inp[0]) ? node22982 : node22975;
													assign node22975 = (inp[9]) ? node22979 : node22976;
														assign node22976 = (inp[4]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22979 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node22982 = (inp[13]) ? node22986 : node22983;
														assign node22983 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node22986 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node22989 = (inp[9]) ? node23005 : node22990;
												assign node22990 = (inp[2]) ? node22998 : node22991;
													assign node22991 = (inp[0]) ? node22995 : node22992;
														assign node22992 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node22995 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node22998 = (inp[4]) ? node23002 : node22999;
														assign node22999 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23002 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node23005 = (inp[8]) ? node23011 : node23006;
													assign node23006 = (inp[2]) ? 16'b0000000000011111 : node23007;
														assign node23007 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node23011 = (inp[4]) ? node23015 : node23012;
														assign node23012 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node23015 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node23018 = (inp[8]) ? node23082 : node23019;
										assign node23019 = (inp[4]) ? node23051 : node23020;
											assign node23020 = (inp[2]) ? node23036 : node23021;
												assign node23021 = (inp[9]) ? node23029 : node23022;
													assign node23022 = (inp[7]) ? node23026 : node23023;
														assign node23023 = (inp[1]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node23026 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23029 = (inp[1]) ? node23033 : node23030;
														assign node23030 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23033 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23036 = (inp[7]) ? node23044 : node23037;
													assign node23037 = (inp[0]) ? node23041 : node23038;
														assign node23038 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23041 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23044 = (inp[9]) ? node23048 : node23045;
														assign node23045 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23048 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node23051 = (inp[13]) ? node23067 : node23052;
												assign node23052 = (inp[9]) ? node23060 : node23053;
													assign node23053 = (inp[0]) ? node23057 : node23054;
														assign node23054 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node23057 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23060 = (inp[1]) ? node23064 : node23061;
														assign node23061 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23064 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23067 = (inp[1]) ? node23075 : node23068;
													assign node23068 = (inp[2]) ? node23072 : node23069;
														assign node23069 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23072 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23075 = (inp[2]) ? node23079 : node23076;
														assign node23076 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node23079 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node23082 = (inp[0]) ? node23112 : node23083;
											assign node23083 = (inp[9]) ? node23097 : node23084;
												assign node23084 = (inp[1]) ? node23090 : node23085;
													assign node23085 = (inp[7]) ? node23087 : 16'b0000000001111111;
														assign node23087 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node23090 = (inp[4]) ? node23094 : node23091;
														assign node23091 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node23094 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23097 = (inp[7]) ? node23105 : node23098;
													assign node23098 = (inp[4]) ? node23102 : node23099;
														assign node23099 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node23102 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23105 = (inp[2]) ? node23109 : node23106;
														assign node23106 = (inp[4]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23109 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000001111;
											assign node23112 = (inp[13]) ? node23128 : node23113;
												assign node23113 = (inp[1]) ? node23121 : node23114;
													assign node23114 = (inp[9]) ? node23118 : node23115;
														assign node23115 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node23118 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23121 = (inp[2]) ? node23125 : node23122;
														assign node23122 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23125 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node23128 = (inp[1]) ? node23136 : node23129;
													assign node23129 = (inp[9]) ? node23133 : node23130;
														assign node23130 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23133 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23136 = (inp[4]) ? node23140 : node23137;
														assign node23137 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node23140 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000000111;
								assign node23143 = (inp[2]) ? node23265 : node23144;
									assign node23144 = (inp[0]) ? node23208 : node23145;
										assign node23145 = (inp[9]) ? node23177 : node23146;
											assign node23146 = (inp[7]) ? node23162 : node23147;
												assign node23147 = (inp[4]) ? node23155 : node23148;
													assign node23148 = (inp[14]) ? node23152 : node23149;
														assign node23149 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23152 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23155 = (inp[1]) ? node23159 : node23156;
														assign node23156 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node23159 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23162 = (inp[4]) ? node23170 : node23163;
													assign node23163 = (inp[14]) ? node23167 : node23164;
														assign node23164 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node23167 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23170 = (inp[14]) ? node23174 : node23171;
														assign node23171 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23174 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node23177 = (inp[7]) ? node23193 : node23178;
												assign node23178 = (inp[1]) ? node23186 : node23179;
													assign node23179 = (inp[4]) ? node23183 : node23180;
														assign node23180 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23183 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23186 = (inp[8]) ? node23190 : node23187;
														assign node23187 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23190 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23193 = (inp[4]) ? node23201 : node23194;
													assign node23194 = (inp[13]) ? node23198 : node23195;
														assign node23195 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node23198 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23201 = (inp[8]) ? node23205 : node23202;
														assign node23202 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23205 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node23208 = (inp[13]) ? node23238 : node23209;
											assign node23209 = (inp[8]) ? node23223 : node23210;
												assign node23210 = (inp[4]) ? node23216 : node23211;
													assign node23211 = (inp[9]) ? node23213 : 16'b0000000011111111;
														assign node23213 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23216 = (inp[7]) ? node23220 : node23217;
														assign node23217 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23220 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23223 = (inp[4]) ? node23231 : node23224;
													assign node23224 = (inp[1]) ? node23228 : node23225;
														assign node23225 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23228 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23231 = (inp[7]) ? node23235 : node23232;
														assign node23232 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23235 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node23238 = (inp[1]) ? node23250 : node23239;
												assign node23239 = (inp[7]) ? node23245 : node23240;
													assign node23240 = (inp[4]) ? node23242 : 16'b0000000000111111;
														assign node23242 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node23245 = (inp[14]) ? node23247 : 16'b0000000000111111;
														assign node23247 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node23250 = (inp[9]) ? node23258 : node23251;
													assign node23251 = (inp[8]) ? node23255 : node23252;
														assign node23252 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23255 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000011111;
													assign node23258 = (inp[7]) ? node23262 : node23259;
														assign node23259 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node23262 = (inp[4]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node23265 = (inp[14]) ? node23325 : node23266;
										assign node23266 = (inp[13]) ? node23296 : node23267;
											assign node23267 = (inp[9]) ? node23281 : node23268;
												assign node23268 = (inp[4]) ? node23274 : node23269;
													assign node23269 = (inp[8]) ? node23271 : 16'b0000000011111111;
														assign node23271 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node23274 = (inp[0]) ? node23278 : node23275;
														assign node23275 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23278 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node23281 = (inp[4]) ? node23289 : node23282;
													assign node23282 = (inp[1]) ? node23286 : node23283;
														assign node23283 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23286 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23289 = (inp[8]) ? node23293 : node23290;
														assign node23290 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23293 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node23296 = (inp[1]) ? node23312 : node23297;
												assign node23297 = (inp[4]) ? node23305 : node23298;
													assign node23298 = (inp[7]) ? node23302 : node23299;
														assign node23299 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node23302 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23305 = (inp[9]) ? node23309 : node23306;
														assign node23306 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23309 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node23312 = (inp[9]) ? node23318 : node23313;
													assign node23313 = (inp[7]) ? node23315 : 16'b0000000000011111;
														assign node23315 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23318 = (inp[7]) ? node23322 : node23319;
														assign node23319 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node23322 = (inp[8]) ? 16'b0000000000000011 : 16'b0000000000000111;
										assign node23325 = (inp[1]) ? node23357 : node23326;
											assign node23326 = (inp[8]) ? node23342 : node23327;
												assign node23327 = (inp[0]) ? node23335 : node23328;
													assign node23328 = (inp[4]) ? node23332 : node23329;
														assign node23329 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node23332 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node23335 = (inp[13]) ? node23339 : node23336;
														assign node23336 = (inp[4]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node23339 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node23342 = (inp[13]) ? node23350 : node23343;
													assign node23343 = (inp[4]) ? node23347 : node23344;
														assign node23344 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node23347 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node23350 = (inp[0]) ? node23354 : node23351;
														assign node23351 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node23354 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node23357 = (inp[9]) ? node23373 : node23358;
												assign node23358 = (inp[4]) ? node23366 : node23359;
													assign node23359 = (inp[8]) ? node23363 : node23360;
														assign node23360 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node23363 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000011111;
													assign node23366 = (inp[7]) ? node23370 : node23367;
														assign node23367 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node23370 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node23373 = (inp[4]) ? node23381 : node23374;
													assign node23374 = (inp[7]) ? node23378 : node23375;
														assign node23375 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node23378 = (inp[8]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node23381 = (inp[0]) ? node23385 : node23382;
														assign node23382 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000000111;
														assign node23385 = (inp[13]) ? 16'b0000000000000011 : 16'b0000000000000111;
			assign node23388 = (inp[4]) ? node27208 : node23389;
				assign node23389 = (inp[2]) ? node25293 : node23390;
					assign node23390 = (inp[8]) ? node24336 : node23391;
						assign node23391 = (inp[0]) ? node23873 : node23392;
							assign node23392 = (inp[9]) ? node23634 : node23393;
								assign node23393 = (inp[14]) ? node23513 : node23394;
									assign node23394 = (inp[1]) ? node23456 : node23395;
										assign node23395 = (inp[11]) ? node23427 : node23396;
											assign node23396 = (inp[15]) ? node23412 : node23397;
												assign node23397 = (inp[7]) ? node23405 : node23398;
													assign node23398 = (inp[5]) ? node23402 : node23399;
														assign node23399 = (inp[3]) ? 16'b0000111111111111 : 16'b0001111111111111;
														assign node23402 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
													assign node23405 = (inp[12]) ? node23409 : node23406;
														assign node23406 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node23409 = (inp[3]) ? 16'b0000000111111111 : 16'b0000011111111111;
												assign node23412 = (inp[13]) ? node23420 : node23413;
													assign node23413 = (inp[3]) ? node23417 : node23414;
														assign node23414 = (inp[7]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node23417 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node23420 = (inp[5]) ? node23424 : node23421;
														assign node23421 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23424 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node23427 = (inp[12]) ? node23443 : node23428;
												assign node23428 = (inp[5]) ? node23436 : node23429;
													assign node23429 = (inp[7]) ? node23433 : node23430;
														assign node23430 = (inp[3]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node23433 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node23436 = (inp[15]) ? node23440 : node23437;
														assign node23437 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23440 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node23443 = (inp[15]) ? node23451 : node23444;
													assign node23444 = (inp[7]) ? node23448 : node23445;
														assign node23445 = (inp[13]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node23448 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23451 = (inp[5]) ? node23453 : 16'b0000000111111111;
														assign node23453 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
										assign node23456 = (inp[7]) ? node23484 : node23457;
											assign node23457 = (inp[3]) ? node23469 : node23458;
												assign node23458 = (inp[12]) ? node23462 : node23459;
													assign node23459 = (inp[15]) ? 16'b0000111111111111 : 16'b0000011111111111;
													assign node23462 = (inp[5]) ? node23466 : node23463;
														assign node23463 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23466 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node23469 = (inp[5]) ? node23477 : node23470;
													assign node23470 = (inp[12]) ? node23474 : node23471;
														assign node23471 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23474 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23477 = (inp[12]) ? node23481 : node23478;
														assign node23478 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23481 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
											assign node23484 = (inp[5]) ? node23500 : node23485;
												assign node23485 = (inp[13]) ? node23493 : node23486;
													assign node23486 = (inp[15]) ? node23490 : node23487;
														assign node23487 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23490 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23493 = (inp[15]) ? node23497 : node23494;
														assign node23494 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node23497 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23500 = (inp[13]) ? node23508 : node23501;
													assign node23501 = (inp[11]) ? node23505 : node23502;
														assign node23502 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23505 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node23508 = (inp[15]) ? node23510 : 16'b0000000011111111;
														assign node23510 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node23513 = (inp[11]) ? node23575 : node23514;
										assign node23514 = (inp[13]) ? node23544 : node23515;
											assign node23515 = (inp[7]) ? node23531 : node23516;
												assign node23516 = (inp[3]) ? node23524 : node23517;
													assign node23517 = (inp[5]) ? node23521 : node23518;
														assign node23518 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node23521 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node23524 = (inp[15]) ? node23528 : node23525;
														assign node23525 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23528 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node23531 = (inp[15]) ? node23537 : node23532;
													assign node23532 = (inp[5]) ? 16'b0000000111111111 : node23533;
														assign node23533 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node23537 = (inp[1]) ? node23541 : node23538;
														assign node23538 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23541 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node23544 = (inp[7]) ? node23560 : node23545;
												assign node23545 = (inp[12]) ? node23553 : node23546;
													assign node23546 = (inp[15]) ? node23550 : node23547;
														assign node23547 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23550 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23553 = (inp[5]) ? node23557 : node23554;
														assign node23554 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23557 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23560 = (inp[15]) ? node23568 : node23561;
													assign node23561 = (inp[1]) ? node23565 : node23562;
														assign node23562 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node23565 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23568 = (inp[5]) ? node23572 : node23569;
														assign node23569 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23572 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node23575 = (inp[5]) ? node23607 : node23576;
											assign node23576 = (inp[3]) ? node23592 : node23577;
												assign node23577 = (inp[13]) ? node23585 : node23578;
													assign node23578 = (inp[1]) ? node23582 : node23579;
														assign node23579 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23582 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23585 = (inp[12]) ? node23589 : node23586;
														assign node23586 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23589 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node23592 = (inp[12]) ? node23600 : node23593;
													assign node23593 = (inp[1]) ? node23597 : node23594;
														assign node23594 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node23597 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23600 = (inp[7]) ? node23604 : node23601;
														assign node23601 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23604 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node23607 = (inp[1]) ? node23623 : node23608;
												assign node23608 = (inp[3]) ? node23616 : node23609;
													assign node23609 = (inp[7]) ? node23613 : node23610;
														assign node23610 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23613 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23616 = (inp[13]) ? node23620 : node23617;
														assign node23617 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node23620 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23623 = (inp[13]) ? node23629 : node23624;
													assign node23624 = (inp[7]) ? 16'b0000000011111111 : node23625;
														assign node23625 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23629 = (inp[12]) ? 16'b0000000001111111 : node23630;
														assign node23630 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
								assign node23634 = (inp[7]) ? node23748 : node23635;
									assign node23635 = (inp[1]) ? node23687 : node23636;
										assign node23636 = (inp[12]) ? node23662 : node23637;
											assign node23637 = (inp[5]) ? node23647 : node23638;
												assign node23638 = (inp[14]) ? 16'b0000001111111111 : node23639;
													assign node23639 = (inp[11]) ? node23643 : node23640;
														assign node23640 = (inp[13]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node23643 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
												assign node23647 = (inp[11]) ? node23655 : node23648;
													assign node23648 = (inp[13]) ? node23652 : node23649;
														assign node23649 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23652 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23655 = (inp[3]) ? node23659 : node23656;
														assign node23656 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node23659 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node23662 = (inp[11]) ? node23678 : node23663;
												assign node23663 = (inp[14]) ? node23671 : node23664;
													assign node23664 = (inp[13]) ? node23668 : node23665;
														assign node23665 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23668 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23671 = (inp[5]) ? node23675 : node23672;
														assign node23672 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23675 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23678 = (inp[15]) ? node23680 : 16'b0000000111111111;
													assign node23680 = (inp[13]) ? node23684 : node23681;
														assign node23681 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node23684 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node23687 = (inp[13]) ? node23719 : node23688;
											assign node23688 = (inp[12]) ? node23704 : node23689;
												assign node23689 = (inp[3]) ? node23697 : node23690;
													assign node23690 = (inp[14]) ? node23694 : node23691;
														assign node23691 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23694 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23697 = (inp[15]) ? node23701 : node23698;
														assign node23698 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node23701 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23704 = (inp[5]) ? node23712 : node23705;
													assign node23705 = (inp[11]) ? node23709 : node23706;
														assign node23706 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23709 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23712 = (inp[14]) ? node23716 : node23713;
														assign node23713 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23716 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node23719 = (inp[11]) ? node23735 : node23720;
												assign node23720 = (inp[3]) ? node23728 : node23721;
													assign node23721 = (inp[12]) ? node23725 : node23722;
														assign node23722 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23725 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23728 = (inp[12]) ? node23732 : node23729;
														assign node23729 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23732 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23735 = (inp[12]) ? node23743 : node23736;
													assign node23736 = (inp[3]) ? node23740 : node23737;
														assign node23737 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23740 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23743 = (inp[5]) ? node23745 : 16'b0000000011111111;
														assign node23745 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node23748 = (inp[5]) ? node23810 : node23749;
										assign node23749 = (inp[13]) ? node23781 : node23750;
											assign node23750 = (inp[15]) ? node23766 : node23751;
												assign node23751 = (inp[14]) ? node23759 : node23752;
													assign node23752 = (inp[3]) ? node23756 : node23753;
														assign node23753 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23756 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23759 = (inp[1]) ? node23763 : node23760;
														assign node23760 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23763 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23766 = (inp[3]) ? node23774 : node23767;
													assign node23767 = (inp[14]) ? node23771 : node23768;
														assign node23768 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node23771 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23774 = (inp[12]) ? node23778 : node23775;
														assign node23775 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23778 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node23781 = (inp[14]) ? node23795 : node23782;
												assign node23782 = (inp[12]) ? node23790 : node23783;
													assign node23783 = (inp[1]) ? node23787 : node23784;
														assign node23784 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23787 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23790 = (inp[15]) ? 16'b0000000011111111 : node23791;
														assign node23791 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node23795 = (inp[12]) ? node23803 : node23796;
													assign node23796 = (inp[3]) ? node23800 : node23797;
														assign node23797 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node23800 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23803 = (inp[3]) ? node23807 : node23804;
														assign node23804 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23807 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node23810 = (inp[11]) ? node23842 : node23811;
											assign node23811 = (inp[13]) ? node23827 : node23812;
												assign node23812 = (inp[14]) ? node23820 : node23813;
													assign node23813 = (inp[3]) ? node23817 : node23814;
														assign node23814 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23817 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23820 = (inp[1]) ? node23824 : node23821;
														assign node23821 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23824 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23827 = (inp[1]) ? node23835 : node23828;
													assign node23828 = (inp[14]) ? node23832 : node23829;
														assign node23829 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node23832 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23835 = (inp[3]) ? node23839 : node23836;
														assign node23836 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23839 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node23842 = (inp[1]) ? node23858 : node23843;
												assign node23843 = (inp[12]) ? node23851 : node23844;
													assign node23844 = (inp[3]) ? node23848 : node23845;
														assign node23845 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node23848 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23851 = (inp[15]) ? node23855 : node23852;
														assign node23852 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23855 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node23858 = (inp[3]) ? node23866 : node23859;
													assign node23859 = (inp[13]) ? node23863 : node23860;
														assign node23860 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23863 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node23866 = (inp[15]) ? node23870 : node23867;
														assign node23867 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node23870 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
							assign node23873 = (inp[15]) ? node24107 : node23874;
								assign node23874 = (inp[12]) ? node23992 : node23875;
									assign node23875 = (inp[1]) ? node23937 : node23876;
										assign node23876 = (inp[11]) ? node23906 : node23877;
											assign node23877 = (inp[7]) ? node23893 : node23878;
												assign node23878 = (inp[13]) ? node23886 : node23879;
													assign node23879 = (inp[9]) ? node23883 : node23880;
														assign node23880 = (inp[14]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node23883 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node23886 = (inp[5]) ? node23890 : node23887;
														assign node23887 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23890 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node23893 = (inp[14]) ? node23901 : node23894;
													assign node23894 = (inp[13]) ? node23898 : node23895;
														assign node23895 = (inp[9]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node23898 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23901 = (inp[9]) ? 16'b0000000111111111 : node23902;
														assign node23902 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node23906 = (inp[7]) ? node23922 : node23907;
												assign node23907 = (inp[3]) ? node23915 : node23908;
													assign node23908 = (inp[14]) ? node23912 : node23909;
														assign node23909 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23912 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23915 = (inp[13]) ? node23919 : node23916;
														assign node23916 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23919 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node23922 = (inp[3]) ? node23930 : node23923;
													assign node23923 = (inp[5]) ? node23927 : node23924;
														assign node23924 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node23927 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23930 = (inp[13]) ? node23934 : node23931;
														assign node23931 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23934 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node23937 = (inp[13]) ? node23967 : node23938;
											assign node23938 = (inp[5]) ? node23954 : node23939;
												assign node23939 = (inp[3]) ? node23947 : node23940;
													assign node23940 = (inp[7]) ? node23944 : node23941;
														assign node23941 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node23944 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node23947 = (inp[14]) ? node23951 : node23948;
														assign node23948 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23951 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
												assign node23954 = (inp[9]) ? node23962 : node23955;
													assign node23955 = (inp[3]) ? node23959 : node23956;
														assign node23956 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node23959 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node23962 = (inp[11]) ? node23964 : 16'b0000000111111111;
														assign node23964 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node23967 = (inp[9]) ? node23977 : node23968;
												assign node23968 = (inp[7]) ? node23970 : 16'b0000000111111111;
													assign node23970 = (inp[3]) ? node23974 : node23971;
														assign node23971 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node23974 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node23977 = (inp[5]) ? node23985 : node23978;
													assign node23978 = (inp[3]) ? node23982 : node23979;
														assign node23979 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node23982 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node23985 = (inp[11]) ? node23989 : node23986;
														assign node23986 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node23989 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node23992 = (inp[14]) ? node24050 : node23993;
										assign node23993 = (inp[3]) ? node24021 : node23994;
											assign node23994 = (inp[13]) ? node24008 : node23995;
												assign node23995 = (inp[5]) ? node24003 : node23996;
													assign node23996 = (inp[9]) ? node24000 : node23997;
														assign node23997 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node24000 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24003 = (inp[9]) ? 16'b0000000011111111 : node24004;
														assign node24004 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node24008 = (inp[1]) ? node24016 : node24009;
													assign node24009 = (inp[11]) ? node24013 : node24010;
														assign node24010 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node24013 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24016 = (inp[5]) ? 16'b0000000011111111 : node24017;
														assign node24017 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node24021 = (inp[1]) ? node24037 : node24022;
												assign node24022 = (inp[5]) ? node24030 : node24023;
													assign node24023 = (inp[9]) ? node24027 : node24024;
														assign node24024 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24027 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24030 = (inp[11]) ? node24034 : node24031;
														assign node24031 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24034 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24037 = (inp[11]) ? node24045 : node24038;
													assign node24038 = (inp[13]) ? node24042 : node24039;
														assign node24039 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24042 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24045 = (inp[7]) ? 16'b0000000001111111 : node24046;
														assign node24046 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node24050 = (inp[7]) ? node24078 : node24051;
											assign node24051 = (inp[3]) ? node24065 : node24052;
												assign node24052 = (inp[1]) ? node24060 : node24053;
													assign node24053 = (inp[13]) ? node24057 : node24054;
														assign node24054 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24057 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node24060 = (inp[11]) ? node24062 : 16'b0000000111111111;
														assign node24062 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24065 = (inp[11]) ? node24073 : node24066;
													assign node24066 = (inp[1]) ? node24070 : node24067;
														assign node24067 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24070 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node24073 = (inp[9]) ? node24075 : 16'b0000000001111111;
														assign node24075 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node24078 = (inp[11]) ? node24094 : node24079;
												assign node24079 = (inp[3]) ? node24087 : node24080;
													assign node24080 = (inp[13]) ? node24084 : node24081;
														assign node24081 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node24084 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24087 = (inp[5]) ? node24091 : node24088;
														assign node24088 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24091 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24094 = (inp[13]) ? node24100 : node24095;
													assign node24095 = (inp[3]) ? 16'b0000000000111111 : node24096;
														assign node24096 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24100 = (inp[9]) ? node24104 : node24101;
														assign node24101 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node24104 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node24107 = (inp[7]) ? node24223 : node24108;
									assign node24108 = (inp[12]) ? node24168 : node24109;
										assign node24109 = (inp[3]) ? node24141 : node24110;
											assign node24110 = (inp[14]) ? node24126 : node24111;
												assign node24111 = (inp[9]) ? node24119 : node24112;
													assign node24112 = (inp[11]) ? node24116 : node24113;
														assign node24113 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node24116 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24119 = (inp[1]) ? node24123 : node24120;
														assign node24120 = (inp[5]) ? 16'b0000001111111111 : 16'b0000000111111111;
														assign node24123 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node24126 = (inp[13]) ? node24134 : node24127;
													assign node24127 = (inp[1]) ? node24131 : node24128;
														assign node24128 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24131 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24134 = (inp[1]) ? node24138 : node24135;
														assign node24135 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24138 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node24141 = (inp[5]) ? node24155 : node24142;
												assign node24142 = (inp[9]) ? node24148 : node24143;
													assign node24143 = (inp[14]) ? 16'b0000000011111111 : node24144;
														assign node24144 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24148 = (inp[11]) ? node24152 : node24149;
														assign node24149 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24152 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24155 = (inp[13]) ? node24161 : node24156;
													assign node24156 = (inp[11]) ? 16'b0000000011111111 : node24157;
														assign node24157 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24161 = (inp[1]) ? node24165 : node24162;
														assign node24162 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node24165 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node24168 = (inp[1]) ? node24198 : node24169;
											assign node24169 = (inp[13]) ? node24185 : node24170;
												assign node24170 = (inp[5]) ? node24178 : node24171;
													assign node24171 = (inp[11]) ? node24175 : node24172;
														assign node24172 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24175 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24178 = (inp[9]) ? node24182 : node24179;
														assign node24179 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24182 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24185 = (inp[9]) ? node24193 : node24186;
													assign node24186 = (inp[3]) ? node24190 : node24187;
														assign node24187 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24190 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24193 = (inp[11]) ? node24195 : 16'b0000000001111111;
														assign node24195 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node24198 = (inp[11]) ? node24212 : node24199;
												assign node24199 = (inp[9]) ? node24205 : node24200;
													assign node24200 = (inp[14]) ? node24202 : 16'b0000000011111111;
														assign node24202 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24205 = (inp[3]) ? node24209 : node24206;
														assign node24206 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24209 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24212 = (inp[9]) ? node24218 : node24213;
													assign node24213 = (inp[14]) ? node24215 : 16'b0000000001111111;
														assign node24215 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24218 = (inp[5]) ? 16'b0000000000111111 : node24219;
														assign node24219 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node24223 = (inp[14]) ? node24279 : node24224;
										assign node24224 = (inp[13]) ? node24250 : node24225;
											assign node24225 = (inp[3]) ? node24237 : node24226;
												assign node24226 = (inp[9]) ? node24232 : node24227;
													assign node24227 = (inp[12]) ? node24229 : 16'b0000000111111111;
														assign node24229 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24232 = (inp[5]) ? 16'b0000000011111111 : node24233;
														assign node24233 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node24237 = (inp[11]) ? node24245 : node24238;
													assign node24238 = (inp[12]) ? node24242 : node24239;
														assign node24239 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24242 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24245 = (inp[1]) ? 16'b0000000000111111 : node24246;
														assign node24246 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node24250 = (inp[11]) ? node24266 : node24251;
												assign node24251 = (inp[3]) ? node24259 : node24252;
													assign node24252 = (inp[5]) ? node24256 : node24253;
														assign node24253 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24256 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24259 = (inp[9]) ? node24263 : node24260;
														assign node24260 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24263 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24266 = (inp[1]) ? node24274 : node24267;
													assign node24267 = (inp[3]) ? node24271 : node24268;
														assign node24268 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node24271 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24274 = (inp[5]) ? node24276 : 16'b0000000000111111;
														assign node24276 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node24279 = (inp[1]) ? node24309 : node24280;
											assign node24280 = (inp[5]) ? node24294 : node24281;
												assign node24281 = (inp[3]) ? node24287 : node24282;
													assign node24282 = (inp[12]) ? 16'b0000000011111111 : node24283;
														assign node24283 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24287 = (inp[12]) ? node24291 : node24288;
														assign node24288 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24291 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24294 = (inp[3]) ? node24302 : node24295;
													assign node24295 = (inp[9]) ? node24299 : node24296;
														assign node24296 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24299 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node24302 = (inp[11]) ? node24306 : node24303;
														assign node24303 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node24306 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node24309 = (inp[12]) ? node24323 : node24310;
												assign node24310 = (inp[13]) ? node24316 : node24311;
													assign node24311 = (inp[9]) ? node24313 : 16'b0000000001111111;
														assign node24313 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24316 = (inp[3]) ? node24320 : node24317;
														assign node24317 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node24320 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node24323 = (inp[9]) ? node24329 : node24324;
													assign node24324 = (inp[13]) ? 16'b0000000000111111 : node24325;
														assign node24325 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node24329 = (inp[3]) ? node24333 : node24330;
														assign node24330 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node24333 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000011111;
						assign node24336 = (inp[1]) ? node24824 : node24337;
							assign node24337 = (inp[7]) ? node24579 : node24338;
								assign node24338 = (inp[3]) ? node24460 : node24339;
									assign node24339 = (inp[14]) ? node24401 : node24340;
										assign node24340 = (inp[5]) ? node24370 : node24341;
											assign node24341 = (inp[13]) ? node24357 : node24342;
												assign node24342 = (inp[9]) ? node24350 : node24343;
													assign node24343 = (inp[0]) ? node24347 : node24344;
														assign node24344 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node24347 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node24350 = (inp[11]) ? node24354 : node24351;
														assign node24351 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node24354 = (inp[12]) ? 16'b0000000011111111 : 16'b0000001111111111;
												assign node24357 = (inp[0]) ? node24365 : node24358;
													assign node24358 = (inp[9]) ? node24362 : node24359;
														assign node24359 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node24362 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24365 = (inp[9]) ? 16'b0000000111111111 : node24366;
														assign node24366 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node24370 = (inp[0]) ? node24386 : node24371;
												assign node24371 = (inp[11]) ? node24379 : node24372;
													assign node24372 = (inp[13]) ? node24376 : node24373;
														assign node24373 = (inp[15]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node24376 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24379 = (inp[13]) ? node24383 : node24380;
														assign node24380 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24383 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node24386 = (inp[13]) ? node24394 : node24387;
													assign node24387 = (inp[9]) ? node24391 : node24388;
														assign node24388 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24391 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24394 = (inp[11]) ? node24398 : node24395;
														assign node24395 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node24398 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node24401 = (inp[15]) ? node24431 : node24402;
											assign node24402 = (inp[0]) ? node24416 : node24403;
												assign node24403 = (inp[5]) ? node24411 : node24404;
													assign node24404 = (inp[12]) ? node24408 : node24405;
														assign node24405 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node24408 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24411 = (inp[12]) ? 16'b0000000011111111 : node24412;
														assign node24412 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node24416 = (inp[13]) ? node24424 : node24417;
													assign node24417 = (inp[11]) ? node24421 : node24418;
														assign node24418 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24421 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24424 = (inp[5]) ? node24428 : node24425;
														assign node24425 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24428 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node24431 = (inp[11]) ? node24447 : node24432;
												assign node24432 = (inp[5]) ? node24440 : node24433;
													assign node24433 = (inp[9]) ? node24437 : node24434;
														assign node24434 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24437 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24440 = (inp[12]) ? node24444 : node24441;
														assign node24441 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24444 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node24447 = (inp[13]) ? node24455 : node24448;
													assign node24448 = (inp[0]) ? node24452 : node24449;
														assign node24449 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24452 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24455 = (inp[12]) ? node24457 : 16'b0000000001111111;
														assign node24457 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
									assign node24460 = (inp[15]) ? node24516 : node24461;
										assign node24461 = (inp[13]) ? node24491 : node24462;
											assign node24462 = (inp[9]) ? node24478 : node24463;
												assign node24463 = (inp[12]) ? node24471 : node24464;
													assign node24464 = (inp[11]) ? node24468 : node24465;
														assign node24465 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node24468 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node24471 = (inp[14]) ? node24475 : node24472;
														assign node24472 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24475 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node24478 = (inp[14]) ? node24484 : node24479;
													assign node24479 = (inp[5]) ? node24481 : 16'b0000001111111111;
														assign node24481 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24484 = (inp[5]) ? node24488 : node24485;
														assign node24485 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24488 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node24491 = (inp[12]) ? node24501 : node24492;
												assign node24492 = (inp[11]) ? node24494 : 16'b0000000111111111;
													assign node24494 = (inp[9]) ? node24498 : node24495;
														assign node24495 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24498 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24501 = (inp[14]) ? node24509 : node24502;
													assign node24502 = (inp[0]) ? node24506 : node24503;
														assign node24503 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24506 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24509 = (inp[11]) ? node24513 : node24510;
														assign node24510 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24513 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node24516 = (inp[5]) ? node24548 : node24517;
											assign node24517 = (inp[0]) ? node24533 : node24518;
												assign node24518 = (inp[9]) ? node24526 : node24519;
													assign node24519 = (inp[12]) ? node24523 : node24520;
														assign node24520 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24523 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24526 = (inp[11]) ? node24530 : node24527;
														assign node24527 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24530 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node24533 = (inp[13]) ? node24541 : node24534;
													assign node24534 = (inp[11]) ? node24538 : node24535;
														assign node24535 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node24538 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24541 = (inp[11]) ? node24545 : node24542;
														assign node24542 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node24545 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node24548 = (inp[11]) ? node24564 : node24549;
												assign node24549 = (inp[13]) ? node24557 : node24550;
													assign node24550 = (inp[14]) ? node24554 : node24551;
														assign node24551 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24554 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24557 = (inp[14]) ? node24561 : node24558;
														assign node24558 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24561 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24564 = (inp[14]) ? node24572 : node24565;
													assign node24565 = (inp[9]) ? node24569 : node24566;
														assign node24566 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node24569 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24572 = (inp[9]) ? node24576 : node24573;
														assign node24573 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node24576 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node24579 = (inp[14]) ? node24705 : node24580;
									assign node24580 = (inp[5]) ? node24642 : node24581;
										assign node24581 = (inp[13]) ? node24613 : node24582;
											assign node24582 = (inp[11]) ? node24598 : node24583;
												assign node24583 = (inp[12]) ? node24591 : node24584;
													assign node24584 = (inp[15]) ? node24588 : node24585;
														assign node24585 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node24588 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node24591 = (inp[15]) ? node24595 : node24592;
														assign node24592 = (inp[9]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node24595 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node24598 = (inp[15]) ? node24606 : node24599;
													assign node24599 = (inp[9]) ? node24603 : node24600;
														assign node24600 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24603 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24606 = (inp[12]) ? node24610 : node24607;
														assign node24607 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node24610 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node24613 = (inp[15]) ? node24629 : node24614;
												assign node24614 = (inp[0]) ? node24622 : node24615;
													assign node24615 = (inp[3]) ? node24619 : node24616;
														assign node24616 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24619 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24622 = (inp[12]) ? node24626 : node24623;
														assign node24623 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24626 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24629 = (inp[3]) ? node24637 : node24630;
													assign node24630 = (inp[9]) ? node24634 : node24631;
														assign node24631 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24634 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24637 = (inp[11]) ? node24639 : 16'b0000000001111111;
														assign node24639 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
										assign node24642 = (inp[0]) ? node24674 : node24643;
											assign node24643 = (inp[13]) ? node24659 : node24644;
												assign node24644 = (inp[15]) ? node24652 : node24645;
													assign node24645 = (inp[3]) ? node24649 : node24646;
														assign node24646 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24649 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24652 = (inp[11]) ? node24656 : node24653;
														assign node24653 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24656 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24659 = (inp[15]) ? node24667 : node24660;
													assign node24660 = (inp[12]) ? node24664 : node24661;
														assign node24661 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24664 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24667 = (inp[9]) ? node24671 : node24668;
														assign node24668 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24671 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node24674 = (inp[13]) ? node24690 : node24675;
												assign node24675 = (inp[12]) ? node24683 : node24676;
													assign node24676 = (inp[9]) ? node24680 : node24677;
														assign node24677 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24680 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24683 = (inp[3]) ? node24687 : node24684;
														assign node24684 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24687 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24690 = (inp[15]) ? node24698 : node24691;
													assign node24691 = (inp[12]) ? node24695 : node24692;
														assign node24692 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node24695 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node24698 = (inp[11]) ? node24702 : node24699;
														assign node24699 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node24702 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node24705 = (inp[3]) ? node24767 : node24706;
										assign node24706 = (inp[9]) ? node24736 : node24707;
											assign node24707 = (inp[15]) ? node24723 : node24708;
												assign node24708 = (inp[5]) ? node24716 : node24709;
													assign node24709 = (inp[0]) ? node24713 : node24710;
														assign node24710 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24713 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node24716 = (inp[12]) ? node24720 : node24717;
														assign node24717 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24720 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node24723 = (inp[12]) ? node24729 : node24724;
													assign node24724 = (inp[11]) ? node24726 : 16'b0000000011111111;
														assign node24726 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24729 = (inp[13]) ? node24733 : node24730;
														assign node24730 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000001111111;
														assign node24733 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node24736 = (inp[12]) ? node24752 : node24737;
												assign node24737 = (inp[0]) ? node24745 : node24738;
													assign node24738 = (inp[13]) ? node24742 : node24739;
														assign node24739 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node24742 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24745 = (inp[5]) ? node24749 : node24746;
														assign node24746 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24749 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24752 = (inp[13]) ? node24760 : node24753;
													assign node24753 = (inp[15]) ? node24757 : node24754;
														assign node24754 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24757 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24760 = (inp[0]) ? node24764 : node24761;
														assign node24761 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24764 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node24767 = (inp[13]) ? node24797 : node24768;
											assign node24768 = (inp[12]) ? node24782 : node24769;
												assign node24769 = (inp[15]) ? node24777 : node24770;
													assign node24770 = (inp[5]) ? node24774 : node24771;
														assign node24771 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24774 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24777 = (inp[9]) ? 16'b0000000000111111 : node24778;
														assign node24778 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24782 = (inp[15]) ? node24790 : node24783;
													assign node24783 = (inp[5]) ? node24787 : node24784;
														assign node24784 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24787 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24790 = (inp[9]) ? node24794 : node24791;
														assign node24791 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24794 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node24797 = (inp[9]) ? node24813 : node24798;
												assign node24798 = (inp[15]) ? node24806 : node24799;
													assign node24799 = (inp[5]) ? node24803 : node24800;
														assign node24800 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node24803 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node24806 = (inp[5]) ? node24810 : node24807;
														assign node24807 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node24810 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node24813 = (inp[12]) ? node24819 : node24814;
													assign node24814 = (inp[11]) ? node24816 : 16'b0000000000111111;
														assign node24816 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node24819 = (inp[5]) ? node24821 : 16'b0000000000011111;
														assign node24821 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node24824 = (inp[5]) ? node25054 : node24825;
								assign node24825 = (inp[12]) ? node24937 : node24826;
									assign node24826 = (inp[11]) ? node24882 : node24827;
										assign node24827 = (inp[0]) ? node24853 : node24828;
											assign node24828 = (inp[3]) ? node24840 : node24829;
												assign node24829 = (inp[15]) ? node24835 : node24830;
													assign node24830 = (inp[14]) ? 16'b0000000111111111 : node24831;
														assign node24831 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node24835 = (inp[13]) ? 16'b0000000111111111 : node24836;
														assign node24836 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000111111111;
												assign node24840 = (inp[7]) ? node24848 : node24841;
													assign node24841 = (inp[9]) ? node24845 : node24842;
														assign node24842 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24845 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24848 = (inp[13]) ? 16'b0000000011111111 : node24849;
														assign node24849 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node24853 = (inp[13]) ? node24869 : node24854;
												assign node24854 = (inp[7]) ? node24862 : node24855;
													assign node24855 = (inp[14]) ? node24859 : node24856;
														assign node24856 = (inp[9]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node24859 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24862 = (inp[14]) ? node24866 : node24863;
														assign node24863 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24866 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24869 = (inp[9]) ? node24877 : node24870;
													assign node24870 = (inp[7]) ? node24874 : node24871;
														assign node24871 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24874 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24877 = (inp[3]) ? 16'b0000000001111111 : node24878;
														assign node24878 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node24882 = (inp[9]) ? node24910 : node24883;
											assign node24883 = (inp[15]) ? node24897 : node24884;
												assign node24884 = (inp[3]) ? node24890 : node24885;
													assign node24885 = (inp[14]) ? node24887 : 16'b0000001111111111;
														assign node24887 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24890 = (inp[0]) ? node24894 : node24891;
														assign node24891 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24894 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node24897 = (inp[0]) ? node24905 : node24898;
													assign node24898 = (inp[13]) ? node24902 : node24899;
														assign node24899 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24902 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node24905 = (inp[13]) ? node24907 : 16'b0000000001111111;
														assign node24907 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node24910 = (inp[15]) ? node24926 : node24911;
												assign node24911 = (inp[3]) ? node24919 : node24912;
													assign node24912 = (inp[7]) ? node24916 : node24913;
														assign node24913 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node24916 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24919 = (inp[0]) ? node24923 : node24920;
														assign node24920 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node24923 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24926 = (inp[13]) ? node24932 : node24927;
													assign node24927 = (inp[3]) ? 16'b0000000000111111 : node24928;
														assign node24928 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node24932 = (inp[14]) ? 16'b0000000000111111 : node24933;
														assign node24933 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node24937 = (inp[0]) ? node25001 : node24938;
										assign node24938 = (inp[3]) ? node24970 : node24939;
											assign node24939 = (inp[11]) ? node24955 : node24940;
												assign node24940 = (inp[7]) ? node24948 : node24941;
													assign node24941 = (inp[13]) ? node24945 : node24942;
														assign node24942 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node24945 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node24948 = (inp[15]) ? node24952 : node24949;
														assign node24949 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24952 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node24955 = (inp[9]) ? node24963 : node24956;
													assign node24956 = (inp[13]) ? node24960 : node24957;
														assign node24957 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24960 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24963 = (inp[7]) ? node24967 : node24964;
														assign node24964 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node24967 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node24970 = (inp[13]) ? node24986 : node24971;
												assign node24971 = (inp[11]) ? node24979 : node24972;
													assign node24972 = (inp[7]) ? node24976 : node24973;
														assign node24973 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node24976 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node24979 = (inp[15]) ? node24983 : node24980;
														assign node24980 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24983 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node24986 = (inp[15]) ? node24994 : node24987;
													assign node24987 = (inp[9]) ? node24991 : node24988;
														assign node24988 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node24991 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node24994 = (inp[9]) ? node24998 : node24995;
														assign node24995 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node24998 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node25001 = (inp[11]) ? node25027 : node25002;
											assign node25002 = (inp[14]) ? node25014 : node25003;
												assign node25003 = (inp[9]) ? node25007 : node25004;
													assign node25004 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25007 = (inp[3]) ? node25011 : node25008;
														assign node25008 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node25011 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node25014 = (inp[13]) ? node25020 : node25015;
													assign node25015 = (inp[7]) ? node25017 : 16'b0000000001111111;
														assign node25017 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25020 = (inp[7]) ? node25024 : node25021;
														assign node25021 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25024 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node25027 = (inp[15]) ? node25041 : node25028;
												assign node25028 = (inp[9]) ? node25034 : node25029;
													assign node25029 = (inp[14]) ? node25031 : 16'b0000000011111111;
														assign node25031 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25034 = (inp[14]) ? node25038 : node25035;
														assign node25035 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25038 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node25041 = (inp[9]) ? node25049 : node25042;
													assign node25042 = (inp[7]) ? node25046 : node25043;
														assign node25043 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25046 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node25049 = (inp[13]) ? 16'b0000000000001111 : node25050;
														assign node25050 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node25054 = (inp[3]) ? node25174 : node25055;
									assign node25055 = (inp[13]) ? node25115 : node25056;
										assign node25056 = (inp[15]) ? node25084 : node25057;
											assign node25057 = (inp[0]) ? node25071 : node25058;
												assign node25058 = (inp[9]) ? node25064 : node25059;
													assign node25059 = (inp[14]) ? 16'b0000000111111111 : node25060;
														assign node25060 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25064 = (inp[11]) ? node25068 : node25065;
														assign node25065 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25068 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node25071 = (inp[11]) ? node25079 : node25072;
													assign node25072 = (inp[14]) ? node25076 : node25073;
														assign node25073 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25076 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25079 = (inp[14]) ? 16'b0000000000111111 : node25080;
														assign node25080 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000011111111;
											assign node25084 = (inp[14]) ? node25100 : node25085;
												assign node25085 = (inp[0]) ? node25093 : node25086;
													assign node25086 = (inp[11]) ? node25090 : node25087;
														assign node25087 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25090 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25093 = (inp[11]) ? node25097 : node25094;
														assign node25094 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node25097 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node25100 = (inp[12]) ? node25108 : node25101;
													assign node25101 = (inp[0]) ? node25105 : node25102;
														assign node25102 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25105 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25108 = (inp[11]) ? node25112 : node25109;
														assign node25109 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25112 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node25115 = (inp[0]) ? node25145 : node25116;
											assign node25116 = (inp[7]) ? node25132 : node25117;
												assign node25117 = (inp[12]) ? node25125 : node25118;
													assign node25118 = (inp[11]) ? node25122 : node25119;
														assign node25119 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25122 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25125 = (inp[11]) ? node25129 : node25126;
														assign node25126 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25129 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node25132 = (inp[9]) ? node25138 : node25133;
													assign node25133 = (inp[14]) ? 16'b0000000001111111 : node25134;
														assign node25134 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node25138 = (inp[12]) ? node25142 : node25139;
														assign node25139 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25142 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node25145 = (inp[9]) ? node25161 : node25146;
												assign node25146 = (inp[15]) ? node25154 : node25147;
													assign node25147 = (inp[14]) ? node25151 : node25148;
														assign node25148 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25151 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25154 = (inp[11]) ? node25158 : node25155;
														assign node25155 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25158 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node25161 = (inp[14]) ? node25169 : node25162;
													assign node25162 = (inp[12]) ? node25166 : node25163;
														assign node25163 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25166 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node25169 = (inp[7]) ? node25171 : 16'b0000000000011111;
														assign node25171 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node25174 = (inp[13]) ? node25236 : node25175;
										assign node25175 = (inp[7]) ? node25207 : node25176;
											assign node25176 = (inp[9]) ? node25192 : node25177;
												assign node25177 = (inp[0]) ? node25185 : node25178;
													assign node25178 = (inp[14]) ? node25182 : node25179;
														assign node25179 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node25182 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25185 = (inp[14]) ? node25189 : node25186;
														assign node25186 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25189 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node25192 = (inp[15]) ? node25200 : node25193;
													assign node25193 = (inp[11]) ? node25197 : node25194;
														assign node25194 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25197 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node25200 = (inp[12]) ? node25204 : node25201;
														assign node25201 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node25204 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node25207 = (inp[0]) ? node25221 : node25208;
												assign node25208 = (inp[11]) ? node25214 : node25209;
													assign node25209 = (inp[9]) ? node25211 : 16'b0000000001111111;
														assign node25211 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25214 = (inp[12]) ? node25218 : node25215;
														assign node25215 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25218 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node25221 = (inp[12]) ? node25229 : node25222;
													assign node25222 = (inp[14]) ? node25226 : node25223;
														assign node25223 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25226 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node25229 = (inp[14]) ? node25233 : node25230;
														assign node25230 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node25233 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node25236 = (inp[0]) ? node25262 : node25237;
											assign node25237 = (inp[7]) ? node25251 : node25238;
												assign node25238 = (inp[14]) ? node25246 : node25239;
													assign node25239 = (inp[11]) ? node25243 : node25240;
														assign node25240 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node25243 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25246 = (inp[9]) ? 16'b0000000000111111 : node25247;
														assign node25247 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node25251 = (inp[11]) ? node25257 : node25252;
													assign node25252 = (inp[12]) ? node25254 : 16'b0000000000111111;
														assign node25254 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node25257 = (inp[15]) ? 16'b0000000000011111 : node25258;
														assign node25258 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node25262 = (inp[7]) ? node25278 : node25263;
												assign node25263 = (inp[11]) ? node25271 : node25264;
													assign node25264 = (inp[12]) ? node25268 : node25265;
														assign node25265 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25268 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node25271 = (inp[15]) ? node25275 : node25272;
														assign node25272 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node25275 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node25278 = (inp[14]) ? node25286 : node25279;
													assign node25279 = (inp[12]) ? node25283 : node25280;
														assign node25280 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node25283 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node25286 = (inp[11]) ? node25290 : node25287;
														assign node25287 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000011111;
														assign node25290 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
					assign node25293 = (inp[3]) ? node26253 : node25294;
						assign node25294 = (inp[1]) ? node25776 : node25295;
							assign node25295 = (inp[15]) ? node25535 : node25296;
								assign node25296 = (inp[0]) ? node25414 : node25297;
									assign node25297 = (inp[7]) ? node25355 : node25298;
										assign node25298 = (inp[9]) ? node25326 : node25299;
											assign node25299 = (inp[11]) ? node25315 : node25300;
												assign node25300 = (inp[8]) ? node25308 : node25301;
													assign node25301 = (inp[14]) ? node25305 : node25302;
														assign node25302 = (inp[12]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node25305 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node25308 = (inp[5]) ? node25312 : node25309;
														assign node25309 = (inp[12]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25312 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node25315 = (inp[14]) ? node25321 : node25316;
													assign node25316 = (inp[5]) ? 16'b0000001111111111 : node25317;
														assign node25317 = (inp[13]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node25321 = (inp[12]) ? 16'b0000000111111111 : node25322;
														assign node25322 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
											assign node25326 = (inp[13]) ? node25340 : node25327;
												assign node25327 = (inp[11]) ? node25333 : node25328;
													assign node25328 = (inp[14]) ? node25330 : 16'b0000001111111111;
														assign node25330 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25333 = (inp[5]) ? node25337 : node25334;
														assign node25334 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node25337 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25340 = (inp[12]) ? node25348 : node25341;
													assign node25341 = (inp[8]) ? node25345 : node25342;
														assign node25342 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25345 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25348 = (inp[5]) ? node25352 : node25349;
														assign node25349 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25352 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node25355 = (inp[13]) ? node25385 : node25356;
											assign node25356 = (inp[11]) ? node25372 : node25357;
												assign node25357 = (inp[14]) ? node25365 : node25358;
													assign node25358 = (inp[12]) ? node25362 : node25359;
														assign node25359 = (inp[8]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25362 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25365 = (inp[8]) ? node25369 : node25366;
														assign node25366 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25369 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25372 = (inp[5]) ? node25380 : node25373;
													assign node25373 = (inp[9]) ? node25377 : node25374;
														assign node25374 = (inp[8]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25377 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node25380 = (inp[12]) ? node25382 : 16'b0000000111111111;
														assign node25382 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25385 = (inp[11]) ? node25401 : node25386;
												assign node25386 = (inp[9]) ? node25394 : node25387;
													assign node25387 = (inp[8]) ? node25391 : node25388;
														assign node25388 = (inp[5]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node25391 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25394 = (inp[8]) ? node25398 : node25395;
														assign node25395 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25398 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25401 = (inp[8]) ? node25409 : node25402;
													assign node25402 = (inp[14]) ? node25406 : node25403;
														assign node25403 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25406 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25409 = (inp[9]) ? 16'b0000000000111111 : node25410;
														assign node25410 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
									assign node25414 = (inp[8]) ? node25476 : node25415;
										assign node25415 = (inp[5]) ? node25445 : node25416;
											assign node25416 = (inp[9]) ? node25430 : node25417;
												assign node25417 = (inp[7]) ? node25425 : node25418;
													assign node25418 = (inp[11]) ? node25422 : node25419;
														assign node25419 = (inp[14]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25422 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25425 = (inp[11]) ? 16'b0000000011111111 : node25426;
														assign node25426 = (inp[14]) ? 16'b0000000111111111 : 16'b0000000111111111;
												assign node25430 = (inp[14]) ? node25438 : node25431;
													assign node25431 = (inp[11]) ? node25435 : node25432;
														assign node25432 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25435 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25438 = (inp[7]) ? node25442 : node25439;
														assign node25439 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25442 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25445 = (inp[13]) ? node25461 : node25446;
												assign node25446 = (inp[12]) ? node25454 : node25447;
													assign node25447 = (inp[11]) ? node25451 : node25448;
														assign node25448 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25451 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25454 = (inp[9]) ? node25458 : node25455;
														assign node25455 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25458 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25461 = (inp[11]) ? node25469 : node25462;
													assign node25462 = (inp[14]) ? node25466 : node25463;
														assign node25463 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node25466 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25469 = (inp[14]) ? node25473 : node25470;
														assign node25470 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node25473 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node25476 = (inp[7]) ? node25508 : node25477;
											assign node25477 = (inp[9]) ? node25493 : node25478;
												assign node25478 = (inp[14]) ? node25486 : node25479;
													assign node25479 = (inp[12]) ? node25483 : node25480;
														assign node25480 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25483 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25486 = (inp[11]) ? node25490 : node25487;
														assign node25487 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25490 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25493 = (inp[13]) ? node25501 : node25494;
													assign node25494 = (inp[12]) ? node25498 : node25495;
														assign node25495 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node25498 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node25501 = (inp[5]) ? node25505 : node25502;
														assign node25502 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25505 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node25508 = (inp[5]) ? node25520 : node25509;
												assign node25509 = (inp[12]) ? node25515 : node25510;
													assign node25510 = (inp[14]) ? node25512 : 16'b0000000111111111;
														assign node25512 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25515 = (inp[11]) ? 16'b0000000001111111 : node25516;
														assign node25516 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25520 = (inp[13]) ? node25528 : node25521;
													assign node25521 = (inp[14]) ? node25525 : node25522;
														assign node25522 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25525 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node25528 = (inp[11]) ? node25532 : node25529;
														assign node25529 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25532 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
								assign node25535 = (inp[13]) ? node25651 : node25536;
									assign node25536 = (inp[8]) ? node25596 : node25537;
										assign node25537 = (inp[7]) ? node25565 : node25538;
											assign node25538 = (inp[5]) ? node25552 : node25539;
												assign node25539 = (inp[0]) ? node25547 : node25540;
													assign node25540 = (inp[14]) ? node25544 : node25541;
														assign node25541 = (inp[9]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25544 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25547 = (inp[14]) ? 16'b0000000011111111 : node25548;
														assign node25548 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node25552 = (inp[11]) ? node25558 : node25553;
													assign node25553 = (inp[0]) ? 16'b0000000011111111 : node25554;
														assign node25554 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node25558 = (inp[14]) ? node25562 : node25559;
														assign node25559 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25562 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25565 = (inp[11]) ? node25581 : node25566;
												assign node25566 = (inp[14]) ? node25574 : node25567;
													assign node25567 = (inp[5]) ? node25571 : node25568;
														assign node25568 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25571 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25574 = (inp[9]) ? node25578 : node25575;
														assign node25575 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25578 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25581 = (inp[12]) ? node25589 : node25582;
													assign node25582 = (inp[5]) ? node25586 : node25583;
														assign node25583 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25586 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25589 = (inp[9]) ? node25593 : node25590;
														assign node25590 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25593 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node25596 = (inp[12]) ? node25626 : node25597;
											assign node25597 = (inp[0]) ? node25613 : node25598;
												assign node25598 = (inp[11]) ? node25606 : node25599;
													assign node25599 = (inp[9]) ? node25603 : node25600;
														assign node25600 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25603 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25606 = (inp[5]) ? node25610 : node25607;
														assign node25607 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25610 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25613 = (inp[9]) ? node25619 : node25614;
													assign node25614 = (inp[14]) ? 16'b0000000001111111 : node25615;
														assign node25615 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25619 = (inp[7]) ? node25623 : node25620;
														assign node25620 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25623 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node25626 = (inp[7]) ? node25636 : node25627;
												assign node25627 = (inp[9]) ? node25629 : 16'b0000000011111111;
													assign node25629 = (inp[11]) ? node25633 : node25630;
														assign node25630 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25633 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node25636 = (inp[5]) ? node25644 : node25637;
													assign node25637 = (inp[0]) ? node25641 : node25638;
														assign node25638 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node25641 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25644 = (inp[11]) ? node25648 : node25645;
														assign node25645 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25648 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node25651 = (inp[12]) ? node25713 : node25652;
										assign node25652 = (inp[9]) ? node25682 : node25653;
											assign node25653 = (inp[0]) ? node25667 : node25654;
												assign node25654 = (inp[7]) ? node25662 : node25655;
													assign node25655 = (inp[14]) ? node25659 : node25656;
														assign node25656 = (inp[8]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node25659 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25662 = (inp[8]) ? node25664 : 16'b0000000011111111;
														assign node25664 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25667 = (inp[14]) ? node25675 : node25668;
													assign node25668 = (inp[5]) ? node25672 : node25669;
														assign node25669 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25672 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25675 = (inp[7]) ? node25679 : node25676;
														assign node25676 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node25679 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node25682 = (inp[11]) ? node25698 : node25683;
												assign node25683 = (inp[5]) ? node25691 : node25684;
													assign node25684 = (inp[7]) ? node25688 : node25685;
														assign node25685 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25688 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25691 = (inp[8]) ? node25695 : node25692;
														assign node25692 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node25695 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node25698 = (inp[14]) ? node25706 : node25699;
													assign node25699 = (inp[0]) ? node25703 : node25700;
														assign node25700 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25703 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25706 = (inp[7]) ? node25710 : node25707;
														assign node25707 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25710 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node25713 = (inp[7]) ? node25745 : node25714;
											assign node25714 = (inp[8]) ? node25730 : node25715;
												assign node25715 = (inp[0]) ? node25723 : node25716;
													assign node25716 = (inp[9]) ? node25720 : node25717;
														assign node25717 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25720 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25723 = (inp[14]) ? node25727 : node25724;
														assign node25724 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25727 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node25730 = (inp[5]) ? node25738 : node25731;
													assign node25731 = (inp[11]) ? node25735 : node25732;
														assign node25732 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25735 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25738 = (inp[9]) ? node25742 : node25739;
														assign node25739 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25742 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node25745 = (inp[14]) ? node25761 : node25746;
												assign node25746 = (inp[0]) ? node25754 : node25747;
													assign node25747 = (inp[9]) ? node25751 : node25748;
														assign node25748 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25751 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25754 = (inp[8]) ? node25758 : node25755;
														assign node25755 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25758 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node25761 = (inp[5]) ? node25769 : node25762;
													assign node25762 = (inp[8]) ? node25766 : node25763;
														assign node25763 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25766 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node25769 = (inp[0]) ? node25773 : node25770;
														assign node25770 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node25773 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
							assign node25776 = (inp[5]) ? node26014 : node25777;
								assign node25777 = (inp[8]) ? node25893 : node25778;
									assign node25778 = (inp[11]) ? node25832 : node25779;
										assign node25779 = (inp[9]) ? node25809 : node25780;
											assign node25780 = (inp[15]) ? node25796 : node25781;
												assign node25781 = (inp[0]) ? node25789 : node25782;
													assign node25782 = (inp[14]) ? node25786 : node25783;
														assign node25783 = (inp[7]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node25786 = (inp[12]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node25789 = (inp[12]) ? node25793 : node25790;
														assign node25790 = (inp[7]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node25793 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node25796 = (inp[13]) ? node25804 : node25797;
													assign node25797 = (inp[7]) ? node25801 : node25798;
														assign node25798 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25801 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25804 = (inp[14]) ? node25806 : 16'b0000000011111111;
														assign node25806 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node25809 = (inp[12]) ? node25825 : node25810;
												assign node25810 = (inp[7]) ? node25818 : node25811;
													assign node25811 = (inp[14]) ? node25815 : node25812;
														assign node25812 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25815 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25818 = (inp[13]) ? node25822 : node25819;
														assign node25819 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node25822 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25825 = (inp[14]) ? node25827 : 16'b0000000011111111;
													assign node25827 = (inp[13]) ? 16'b0000000001111111 : node25828;
														assign node25828 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node25832 = (inp[13]) ? node25864 : node25833;
											assign node25833 = (inp[7]) ? node25849 : node25834;
												assign node25834 = (inp[0]) ? node25842 : node25835;
													assign node25835 = (inp[15]) ? node25839 : node25836;
														assign node25836 = (inp[9]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node25839 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25842 = (inp[12]) ? node25846 : node25843;
														assign node25843 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25846 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25849 = (inp[15]) ? node25857 : node25850;
													assign node25850 = (inp[9]) ? node25854 : node25851;
														assign node25851 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25854 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25857 = (inp[14]) ? node25861 : node25858;
														assign node25858 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25861 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node25864 = (inp[12]) ? node25880 : node25865;
												assign node25865 = (inp[0]) ? node25873 : node25866;
													assign node25866 = (inp[9]) ? node25870 : node25867;
														assign node25867 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25870 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25873 = (inp[15]) ? node25877 : node25874;
														assign node25874 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25877 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node25880 = (inp[14]) ? node25888 : node25881;
													assign node25881 = (inp[0]) ? node25885 : node25882;
														assign node25882 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node25885 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node25888 = (inp[7]) ? node25890 : 16'b0000000000111111;
														assign node25890 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000011111;
									assign node25893 = (inp[7]) ? node25953 : node25894;
										assign node25894 = (inp[15]) ? node25922 : node25895;
											assign node25895 = (inp[12]) ? node25909 : node25896;
												assign node25896 = (inp[13]) ? node25902 : node25897;
													assign node25897 = (inp[0]) ? node25899 : 16'b0000001111111111;
														assign node25899 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node25902 = (inp[0]) ? node25906 : node25903;
														assign node25903 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25906 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node25909 = (inp[9]) ? node25915 : node25910;
													assign node25910 = (inp[13]) ? node25912 : 16'b0000000111111111;
														assign node25912 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25915 = (inp[13]) ? node25919 : node25916;
														assign node25916 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25919 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node25922 = (inp[9]) ? node25938 : node25923;
												assign node25923 = (inp[12]) ? node25931 : node25924;
													assign node25924 = (inp[14]) ? node25928 : node25925;
														assign node25925 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25928 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25931 = (inp[0]) ? node25935 : node25932;
														assign node25932 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25935 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node25938 = (inp[0]) ? node25946 : node25939;
													assign node25939 = (inp[14]) ? node25943 : node25940;
														assign node25940 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node25943 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25946 = (inp[13]) ? node25950 : node25947;
														assign node25947 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25950 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node25953 = (inp[13]) ? node25985 : node25954;
											assign node25954 = (inp[0]) ? node25970 : node25955;
												assign node25955 = (inp[15]) ? node25963 : node25956;
													assign node25956 = (inp[14]) ? node25960 : node25957;
														assign node25957 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node25960 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node25963 = (inp[14]) ? node25967 : node25964;
														assign node25964 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25967 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node25970 = (inp[14]) ? node25978 : node25971;
													assign node25971 = (inp[12]) ? node25975 : node25972;
														assign node25972 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25975 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node25978 = (inp[15]) ? node25982 : node25979;
														assign node25979 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25982 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node25985 = (inp[9]) ? node26001 : node25986;
												assign node25986 = (inp[15]) ? node25994 : node25987;
													assign node25987 = (inp[11]) ? node25991 : node25988;
														assign node25988 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node25991 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node25994 = (inp[11]) ? node25998 : node25995;
														assign node25995 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node25998 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26001 = (inp[15]) ? node26009 : node26002;
													assign node26002 = (inp[11]) ? node26006 : node26003;
														assign node26003 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26006 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26009 = (inp[0]) ? node26011 : 16'b0000000000011111;
														assign node26011 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000011111;
								assign node26014 = (inp[12]) ? node26134 : node26015;
									assign node26015 = (inp[7]) ? node26075 : node26016;
										assign node26016 = (inp[14]) ? node26044 : node26017;
											assign node26017 = (inp[11]) ? node26031 : node26018;
												assign node26018 = (inp[13]) ? node26026 : node26019;
													assign node26019 = (inp[8]) ? node26023 : node26020;
														assign node26020 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26023 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26026 = (inp[8]) ? 16'b0000000011111111 : node26027;
														assign node26027 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node26031 = (inp[15]) ? node26039 : node26032;
													assign node26032 = (inp[13]) ? node26036 : node26033;
														assign node26033 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26036 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node26039 = (inp[9]) ? node26041 : 16'b0000000001111111;
														assign node26041 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node26044 = (inp[9]) ? node26060 : node26045;
												assign node26045 = (inp[8]) ? node26053 : node26046;
													assign node26046 = (inp[11]) ? node26050 : node26047;
														assign node26047 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26050 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26053 = (inp[0]) ? node26057 : node26054;
														assign node26054 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26057 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26060 = (inp[13]) ? node26068 : node26061;
													assign node26061 = (inp[0]) ? node26065 : node26062;
														assign node26062 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node26065 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node26068 = (inp[8]) ? node26072 : node26069;
														assign node26069 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26072 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node26075 = (inp[8]) ? node26107 : node26076;
											assign node26076 = (inp[14]) ? node26092 : node26077;
												assign node26077 = (inp[13]) ? node26085 : node26078;
													assign node26078 = (inp[9]) ? node26082 : node26079;
														assign node26079 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26082 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26085 = (inp[9]) ? node26089 : node26086;
														assign node26086 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node26089 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26092 = (inp[9]) ? node26100 : node26093;
													assign node26093 = (inp[15]) ? node26097 : node26094;
														assign node26094 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26097 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26100 = (inp[0]) ? node26104 : node26101;
														assign node26101 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26104 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node26107 = (inp[15]) ? node26123 : node26108;
												assign node26108 = (inp[11]) ? node26116 : node26109;
													assign node26109 = (inp[9]) ? node26113 : node26110;
														assign node26110 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node26113 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26116 = (inp[9]) ? node26120 : node26117;
														assign node26117 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26120 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26123 = (inp[14]) ? node26129 : node26124;
													assign node26124 = (inp[0]) ? node26126 : 16'b0000000001111111;
														assign node26126 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26129 = (inp[0]) ? 16'b0000000000001111 : node26130;
														assign node26130 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000011111;
									assign node26134 = (inp[0]) ? node26194 : node26135;
										assign node26135 = (inp[8]) ? node26165 : node26136;
											assign node26136 = (inp[9]) ? node26150 : node26137;
												assign node26137 = (inp[15]) ? node26145 : node26138;
													assign node26138 = (inp[14]) ? node26142 : node26139;
														assign node26139 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26142 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node26145 = (inp[7]) ? node26147 : 16'b0000000001111111;
														assign node26147 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node26150 = (inp[13]) ? node26158 : node26151;
													assign node26151 = (inp[14]) ? node26155 : node26152;
														assign node26152 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26155 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26158 = (inp[7]) ? node26162 : node26159;
														assign node26159 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26162 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node26165 = (inp[9]) ? node26179 : node26166;
												assign node26166 = (inp[11]) ? node26172 : node26167;
													assign node26167 = (inp[15]) ? 16'b0000000001111111 : node26168;
														assign node26168 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26172 = (inp[14]) ? node26176 : node26173;
														assign node26173 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26176 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26179 = (inp[13]) ? node26187 : node26180;
													assign node26180 = (inp[14]) ? node26184 : node26181;
														assign node26181 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26184 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26187 = (inp[7]) ? node26191 : node26188;
														assign node26188 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node26191 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node26194 = (inp[8]) ? node26226 : node26195;
											assign node26195 = (inp[13]) ? node26211 : node26196;
												assign node26196 = (inp[14]) ? node26204 : node26197;
													assign node26197 = (inp[15]) ? node26201 : node26198;
														assign node26198 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26201 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node26204 = (inp[11]) ? node26208 : node26205;
														assign node26205 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26208 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node26211 = (inp[7]) ? node26219 : node26212;
													assign node26212 = (inp[9]) ? node26216 : node26213;
														assign node26213 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26216 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26219 = (inp[9]) ? node26223 : node26220;
														assign node26220 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node26223 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node26226 = (inp[13]) ? node26240 : node26227;
												assign node26227 = (inp[11]) ? node26235 : node26228;
													assign node26228 = (inp[7]) ? node26232 : node26229;
														assign node26229 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node26232 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000011111;
													assign node26235 = (inp[15]) ? node26237 : 16'b0000000000011111;
														assign node26237 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node26240 = (inp[14]) ? node26246 : node26241;
													assign node26241 = (inp[11]) ? node26243 : 16'b0000000000111111;
														assign node26243 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node26246 = (inp[11]) ? node26250 : node26247;
														assign node26247 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node26250 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000000111;
						assign node26253 = (inp[9]) ? node26727 : node26254;
							assign node26254 = (inp[1]) ? node26486 : node26255;
								assign node26255 = (inp[0]) ? node26369 : node26256;
									assign node26256 = (inp[5]) ? node26316 : node26257;
										assign node26257 = (inp[14]) ? node26287 : node26258;
											assign node26258 = (inp[11]) ? node26272 : node26259;
												assign node26259 = (inp[8]) ? node26267 : node26260;
													assign node26260 = (inp[12]) ? node26264 : node26261;
														assign node26261 = (inp[15]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node26264 = (inp[7]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node26267 = (inp[15]) ? 16'b0000000111111111 : node26268;
														assign node26268 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node26272 = (inp[13]) ? node26280 : node26273;
													assign node26273 = (inp[8]) ? node26277 : node26274;
														assign node26274 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26277 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node26280 = (inp[12]) ? node26284 : node26281;
														assign node26281 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26284 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node26287 = (inp[8]) ? node26301 : node26288;
												assign node26288 = (inp[13]) ? node26296 : node26289;
													assign node26289 = (inp[12]) ? node26293 : node26290;
														assign node26290 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26293 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26296 = (inp[15]) ? 16'b0000000011111111 : node26297;
														assign node26297 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node26301 = (inp[7]) ? node26309 : node26302;
													assign node26302 = (inp[15]) ? node26306 : node26303;
														assign node26303 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26306 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26309 = (inp[12]) ? node26313 : node26310;
														assign node26310 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node26313 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node26316 = (inp[13]) ? node26342 : node26317;
											assign node26317 = (inp[11]) ? node26333 : node26318;
												assign node26318 = (inp[12]) ? node26326 : node26319;
													assign node26319 = (inp[14]) ? node26323 : node26320;
														assign node26320 = (inp[7]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26323 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node26326 = (inp[15]) ? node26330 : node26327;
														assign node26327 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26330 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26333 = (inp[12]) ? 16'b0000000001111111 : node26334;
													assign node26334 = (inp[7]) ? node26338 : node26335;
														assign node26335 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26338 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node26342 = (inp[8]) ? node26356 : node26343;
												assign node26343 = (inp[14]) ? node26349 : node26344;
													assign node26344 = (inp[15]) ? node26346 : 16'b0000000111111111;
														assign node26346 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26349 = (inp[7]) ? node26353 : node26350;
														assign node26350 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26353 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26356 = (inp[15]) ? node26362 : node26357;
													assign node26357 = (inp[11]) ? 16'b0000000001111111 : node26358;
														assign node26358 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node26362 = (inp[12]) ? node26366 : node26363;
														assign node26363 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26366 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node26369 = (inp[7]) ? node26431 : node26370;
										assign node26370 = (inp[5]) ? node26400 : node26371;
											assign node26371 = (inp[11]) ? node26387 : node26372;
												assign node26372 = (inp[14]) ? node26380 : node26373;
													assign node26373 = (inp[8]) ? node26377 : node26374;
														assign node26374 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26377 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26380 = (inp[8]) ? node26384 : node26381;
														assign node26381 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node26384 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26387 = (inp[13]) ? node26395 : node26388;
													assign node26388 = (inp[15]) ? node26392 : node26389;
														assign node26389 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26392 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node26395 = (inp[15]) ? 16'b0000000001111111 : node26396;
														assign node26396 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node26400 = (inp[14]) ? node26416 : node26401;
												assign node26401 = (inp[13]) ? node26409 : node26402;
													assign node26402 = (inp[15]) ? node26406 : node26403;
														assign node26403 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26406 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26409 = (inp[15]) ? node26413 : node26410;
														assign node26410 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26413 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node26416 = (inp[12]) ? node26424 : node26417;
													assign node26417 = (inp[11]) ? node26421 : node26418;
														assign node26418 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node26421 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26424 = (inp[8]) ? node26428 : node26425;
														assign node26425 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26428 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node26431 = (inp[8]) ? node26457 : node26432;
											assign node26432 = (inp[12]) ? node26446 : node26433;
												assign node26433 = (inp[11]) ? node26441 : node26434;
													assign node26434 = (inp[13]) ? node26438 : node26435;
														assign node26435 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26438 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node26441 = (inp[14]) ? 16'b0000000001111111 : node26442;
														assign node26442 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26446 = (inp[15]) ? node26452 : node26447;
													assign node26447 = (inp[11]) ? node26449 : 16'b0000000011111111;
														assign node26449 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26452 = (inp[13]) ? 16'b0000000000111111 : node26453;
														assign node26453 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node26457 = (inp[14]) ? node26471 : node26458;
												assign node26458 = (inp[13]) ? node26464 : node26459;
													assign node26459 = (inp[12]) ? 16'b0000000000011111 : node26460;
														assign node26460 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26464 = (inp[15]) ? node26468 : node26465;
														assign node26465 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26468 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26471 = (inp[15]) ? node26479 : node26472;
													assign node26472 = (inp[13]) ? node26476 : node26473;
														assign node26473 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26476 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26479 = (inp[11]) ? node26483 : node26480;
														assign node26480 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node26483 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node26486 = (inp[5]) ? node26606 : node26487;
									assign node26487 = (inp[14]) ? node26549 : node26488;
										assign node26488 = (inp[0]) ? node26520 : node26489;
											assign node26489 = (inp[11]) ? node26505 : node26490;
												assign node26490 = (inp[13]) ? node26498 : node26491;
													assign node26491 = (inp[15]) ? node26495 : node26492;
														assign node26492 = (inp[12]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26495 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26498 = (inp[8]) ? node26502 : node26499;
														assign node26499 = (inp[7]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26502 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node26505 = (inp[15]) ? node26513 : node26506;
													assign node26506 = (inp[7]) ? node26510 : node26507;
														assign node26507 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26510 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26513 = (inp[8]) ? node26517 : node26514;
														assign node26514 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26517 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node26520 = (inp[13]) ? node26534 : node26521;
												assign node26521 = (inp[12]) ? node26529 : node26522;
													assign node26522 = (inp[7]) ? node26526 : node26523;
														assign node26523 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26526 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26529 = (inp[7]) ? 16'b0000000001111111 : node26530;
														assign node26530 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26534 = (inp[15]) ? node26542 : node26535;
													assign node26535 = (inp[11]) ? node26539 : node26536;
														assign node26536 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node26539 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26542 = (inp[11]) ? node26546 : node26543;
														assign node26543 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26546 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000111111;
										assign node26549 = (inp[13]) ? node26579 : node26550;
											assign node26550 = (inp[8]) ? node26564 : node26551;
												assign node26551 = (inp[7]) ? node26557 : node26552;
													assign node26552 = (inp[11]) ? 16'b0000000011111111 : node26553;
														assign node26553 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node26557 = (inp[11]) ? node26561 : node26558;
														assign node26558 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26561 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26564 = (inp[7]) ? node26572 : node26565;
													assign node26565 = (inp[15]) ? node26569 : node26566;
														assign node26566 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26569 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26572 = (inp[0]) ? node26576 : node26573;
														assign node26573 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26576 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node26579 = (inp[8]) ? node26593 : node26580;
												assign node26580 = (inp[12]) ? node26588 : node26581;
													assign node26581 = (inp[11]) ? node26585 : node26582;
														assign node26582 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26585 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26588 = (inp[7]) ? 16'b0000000000111111 : node26589;
														assign node26589 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node26593 = (inp[15]) ? node26601 : node26594;
													assign node26594 = (inp[0]) ? node26598 : node26595;
														assign node26595 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26598 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26601 = (inp[7]) ? node26603 : 16'b0000000000011111;
														assign node26603 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node26606 = (inp[11]) ? node26666 : node26607;
										assign node26607 = (inp[8]) ? node26637 : node26608;
											assign node26608 = (inp[14]) ? node26624 : node26609;
												assign node26609 = (inp[7]) ? node26617 : node26610;
													assign node26610 = (inp[15]) ? node26614 : node26611;
														assign node26611 = (inp[12]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26614 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node26617 = (inp[13]) ? node26621 : node26618;
														assign node26618 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26621 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26624 = (inp[0]) ? node26632 : node26625;
													assign node26625 = (inp[13]) ? node26629 : node26626;
														assign node26626 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26629 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node26632 = (inp[12]) ? 16'b0000000000111111 : node26633;
														assign node26633 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node26637 = (inp[12]) ? node26651 : node26638;
												assign node26638 = (inp[15]) ? node26644 : node26639;
													assign node26639 = (inp[14]) ? 16'b0000000000111111 : node26640;
														assign node26640 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26644 = (inp[13]) ? node26648 : node26645;
														assign node26645 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26648 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26651 = (inp[14]) ? node26659 : node26652;
													assign node26652 = (inp[7]) ? node26656 : node26653;
														assign node26653 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node26656 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26659 = (inp[15]) ? node26663 : node26660;
														assign node26660 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node26663 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node26666 = (inp[14]) ? node26696 : node26667;
											assign node26667 = (inp[0]) ? node26681 : node26668;
												assign node26668 = (inp[13]) ? node26674 : node26669;
													assign node26669 = (inp[15]) ? 16'b0000000000111111 : node26670;
														assign node26670 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26674 = (inp[12]) ? node26678 : node26675;
														assign node26675 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26678 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26681 = (inp[13]) ? node26689 : node26682;
													assign node26682 = (inp[15]) ? node26686 : node26683;
														assign node26683 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26686 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26689 = (inp[15]) ? node26693 : node26690;
														assign node26690 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node26693 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node26696 = (inp[8]) ? node26712 : node26697;
												assign node26697 = (inp[13]) ? node26705 : node26698;
													assign node26698 = (inp[12]) ? node26702 : node26699;
														assign node26699 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26702 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26705 = (inp[12]) ? node26709 : node26706;
														assign node26706 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node26709 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node26712 = (inp[12]) ? node26720 : node26713;
													assign node26713 = (inp[0]) ? node26717 : node26714;
														assign node26714 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node26717 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node26720 = (inp[15]) ? node26724 : node26721;
														assign node26721 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node26724 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node26727 = (inp[7]) ? node26973 : node26728;
								assign node26728 = (inp[15]) ? node26852 : node26729;
									assign node26729 = (inp[1]) ? node26791 : node26730;
										assign node26730 = (inp[12]) ? node26762 : node26731;
											assign node26731 = (inp[5]) ? node26747 : node26732;
												assign node26732 = (inp[0]) ? node26740 : node26733;
													assign node26733 = (inp[13]) ? node26737 : node26734;
														assign node26734 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node26737 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node26740 = (inp[14]) ? node26744 : node26741;
														assign node26741 = (inp[8]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node26744 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26747 = (inp[13]) ? node26755 : node26748;
													assign node26748 = (inp[14]) ? node26752 : node26749;
														assign node26749 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26752 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26755 = (inp[0]) ? node26759 : node26756;
														assign node26756 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26759 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node26762 = (inp[14]) ? node26776 : node26763;
												assign node26763 = (inp[0]) ? node26771 : node26764;
													assign node26764 = (inp[8]) ? node26768 : node26765;
														assign node26765 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node26768 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26771 = (inp[11]) ? 16'b0000000001111111 : node26772;
														assign node26772 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node26776 = (inp[11]) ? node26784 : node26777;
													assign node26777 = (inp[13]) ? node26781 : node26778;
														assign node26778 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26781 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26784 = (inp[13]) ? node26788 : node26785;
														assign node26785 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node26788 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node26791 = (inp[11]) ? node26821 : node26792;
											assign node26792 = (inp[13]) ? node26808 : node26793;
												assign node26793 = (inp[12]) ? node26801 : node26794;
													assign node26794 = (inp[5]) ? node26798 : node26795;
														assign node26795 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node26798 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26801 = (inp[0]) ? node26805 : node26802;
														assign node26802 = (inp[8]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26805 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node26808 = (inp[0]) ? node26814 : node26809;
													assign node26809 = (inp[8]) ? node26811 : 16'b0000000001111111;
														assign node26811 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26814 = (inp[5]) ? node26818 : node26815;
														assign node26815 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node26818 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node26821 = (inp[14]) ? node26837 : node26822;
												assign node26822 = (inp[5]) ? node26830 : node26823;
													assign node26823 = (inp[0]) ? node26827 : node26824;
														assign node26824 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26827 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26830 = (inp[0]) ? node26834 : node26831;
														assign node26831 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26834 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26837 = (inp[5]) ? node26845 : node26838;
													assign node26838 = (inp[12]) ? node26842 : node26839;
														assign node26839 = (inp[8]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26842 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node26845 = (inp[13]) ? node26849 : node26846;
														assign node26846 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node26849 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000001111;
									assign node26852 = (inp[11]) ? node26916 : node26853;
										assign node26853 = (inp[8]) ? node26885 : node26854;
											assign node26854 = (inp[13]) ? node26870 : node26855;
												assign node26855 = (inp[0]) ? node26863 : node26856;
													assign node26856 = (inp[1]) ? node26860 : node26857;
														assign node26857 = (inp[5]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node26860 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node26863 = (inp[12]) ? node26867 : node26864;
														assign node26864 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26867 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26870 = (inp[0]) ? node26878 : node26871;
													assign node26871 = (inp[12]) ? node26875 : node26872;
														assign node26872 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node26875 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26878 = (inp[1]) ? node26882 : node26879;
														assign node26879 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node26882 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node26885 = (inp[14]) ? node26901 : node26886;
												assign node26886 = (inp[12]) ? node26894 : node26887;
													assign node26887 = (inp[0]) ? node26891 : node26888;
														assign node26888 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node26891 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node26894 = (inp[1]) ? node26898 : node26895;
														assign node26895 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26898 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26901 = (inp[13]) ? node26909 : node26902;
													assign node26902 = (inp[12]) ? node26906 : node26903;
														assign node26903 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node26906 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26909 = (inp[12]) ? node26913 : node26910;
														assign node26910 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node26913 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node26916 = (inp[14]) ? node26944 : node26917;
											assign node26917 = (inp[5]) ? node26931 : node26918;
												assign node26918 = (inp[8]) ? node26926 : node26919;
													assign node26919 = (inp[12]) ? node26923 : node26920;
														assign node26920 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26923 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node26926 = (inp[12]) ? node26928 : 16'b0000000000111111;
														assign node26928 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node26931 = (inp[8]) ? node26937 : node26932;
													assign node26932 = (inp[1]) ? node26934 : 16'b0000000000111111;
														assign node26934 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26937 = (inp[1]) ? node26941 : node26938;
														assign node26938 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node26941 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node26944 = (inp[13]) ? node26960 : node26945;
												assign node26945 = (inp[1]) ? node26953 : node26946;
													assign node26946 = (inp[0]) ? node26950 : node26947;
														assign node26947 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node26950 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node26953 = (inp[8]) ? node26957 : node26954;
														assign node26954 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node26957 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000011111;
												assign node26960 = (inp[5]) ? node26966 : node26961;
													assign node26961 = (inp[8]) ? node26963 : 16'b0000000000011111;
														assign node26963 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node26966 = (inp[8]) ? node26970 : node26967;
														assign node26967 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node26970 = (inp[12]) ? 16'b0000000000000011 : 16'b0000000000001111;
								assign node26973 = (inp[13]) ? node27087 : node26974;
									assign node26974 = (inp[0]) ? node27034 : node26975;
										assign node26975 = (inp[1]) ? node27005 : node26976;
											assign node26976 = (inp[14]) ? node26992 : node26977;
												assign node26977 = (inp[8]) ? node26985 : node26978;
													assign node26978 = (inp[15]) ? node26982 : node26979;
														assign node26979 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node26982 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node26985 = (inp[11]) ? node26989 : node26986;
														assign node26986 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node26989 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node26992 = (inp[5]) ? node27000 : node26993;
													assign node26993 = (inp[12]) ? node26997 : node26994;
														assign node26994 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node26997 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27000 = (inp[8]) ? 16'b0000000000011111 : node27001;
														assign node27001 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27005 = (inp[12]) ? node27019 : node27006;
												assign node27006 = (inp[8]) ? node27014 : node27007;
													assign node27007 = (inp[14]) ? node27011 : node27008;
														assign node27008 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27011 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27014 = (inp[5]) ? 16'b0000000000011111 : node27015;
														assign node27015 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27019 = (inp[15]) ? node27027 : node27020;
													assign node27020 = (inp[14]) ? node27024 : node27021;
														assign node27021 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27024 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27027 = (inp[11]) ? node27031 : node27028;
														assign node27028 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node27031 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node27034 = (inp[8]) ? node27058 : node27035;
											assign node27035 = (inp[12]) ? node27047 : node27036;
												assign node27036 = (inp[5]) ? node27042 : node27037;
													assign node27037 = (inp[1]) ? 16'b0000000001111111 : node27038;
														assign node27038 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27042 = (inp[11]) ? 16'b0000000000011111 : node27043;
														assign node27043 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27047 = (inp[1]) ? node27053 : node27048;
													assign node27048 = (inp[11]) ? node27050 : 16'b0000000001111111;
														assign node27050 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27053 = (inp[15]) ? 16'b0000000000011111 : node27054;
														assign node27054 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node27058 = (inp[15]) ? node27074 : node27059;
												assign node27059 = (inp[12]) ? node27067 : node27060;
													assign node27060 = (inp[11]) ? node27064 : node27061;
														assign node27061 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27064 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27067 = (inp[1]) ? node27071 : node27068;
														assign node27068 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node27071 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node27074 = (inp[14]) ? node27080 : node27075;
													assign node27075 = (inp[1]) ? 16'b0000000000001111 : node27076;
														assign node27076 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27080 = (inp[11]) ? node27084 : node27081;
														assign node27081 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node27084 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node27087 = (inp[14]) ? node27149 : node27088;
										assign node27088 = (inp[0]) ? node27118 : node27089;
											assign node27089 = (inp[15]) ? node27103 : node27090;
												assign node27090 = (inp[5]) ? node27096 : node27091;
													assign node27091 = (inp[8]) ? 16'b0000000000111111 : node27092;
														assign node27092 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27096 = (inp[12]) ? node27100 : node27097;
														assign node27097 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27100 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node27103 = (inp[12]) ? node27111 : node27104;
													assign node27104 = (inp[1]) ? node27108 : node27105;
														assign node27105 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27108 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27111 = (inp[11]) ? node27115 : node27112;
														assign node27112 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node27115 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node27118 = (inp[12]) ? node27134 : node27119;
												assign node27119 = (inp[8]) ? node27127 : node27120;
													assign node27120 = (inp[15]) ? node27124 : node27121;
														assign node27121 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27124 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27127 = (inp[11]) ? node27131 : node27128;
														assign node27128 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node27131 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node27134 = (inp[11]) ? node27142 : node27135;
													assign node27135 = (inp[15]) ? node27139 : node27136;
														assign node27136 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node27139 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node27142 = (inp[1]) ? node27146 : node27143;
														assign node27143 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node27146 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node27149 = (inp[5]) ? node27181 : node27150;
											assign node27150 = (inp[11]) ? node27166 : node27151;
												assign node27151 = (inp[1]) ? node27159 : node27152;
													assign node27152 = (inp[8]) ? node27156 : node27153;
														assign node27153 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node27156 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node27159 = (inp[0]) ? node27163 : node27160;
														assign node27160 = (inp[8]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node27163 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node27166 = (inp[1]) ? node27174 : node27167;
													assign node27167 = (inp[0]) ? node27171 : node27168;
														assign node27168 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node27171 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node27174 = (inp[0]) ? node27178 : node27175;
														assign node27175 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node27178 = (inp[8]) ? 16'b0000000000000011 : 16'b0000000000001111;
											assign node27181 = (inp[0]) ? node27195 : node27182;
												assign node27182 = (inp[12]) ? node27188 : node27183;
													assign node27183 = (inp[15]) ? node27185 : 16'b0000000000011111;
														assign node27185 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node27188 = (inp[15]) ? node27192 : node27189;
														assign node27189 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node27192 = (inp[11]) ? 16'b0000000000000011 : 16'b0000000000000111;
												assign node27195 = (inp[11]) ? node27203 : node27196;
													assign node27196 = (inp[1]) ? node27200 : node27197;
														assign node27197 = (inp[8]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node27200 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000000111;
													assign node27203 = (inp[8]) ? node27205 : 16'b0000000000000111;
														assign node27205 = (inp[15]) ? 16'b0000000000000001 : 16'b0000000000000111;
				assign node27208 = (inp[8]) ? node29136 : node27209;
					assign node27209 = (inp[12]) ? node28171 : node27210;
						assign node27210 = (inp[9]) ? node27686 : node27211;
							assign node27211 = (inp[7]) ? node27451 : node27212;
								assign node27212 = (inp[11]) ? node27330 : node27213;
									assign node27213 = (inp[1]) ? node27275 : node27214;
										assign node27214 = (inp[13]) ? node27246 : node27215;
											assign node27215 = (inp[14]) ? node27231 : node27216;
												assign node27216 = (inp[3]) ? node27224 : node27217;
													assign node27217 = (inp[2]) ? node27221 : node27218;
														assign node27218 = (inp[15]) ? 16'b0000011111111111 : 16'b0000111111111111;
														assign node27221 = (inp[5]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node27224 = (inp[2]) ? node27228 : node27225;
														assign node27225 = (inp[0]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node27228 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node27231 = (inp[2]) ? node27239 : node27232;
													assign node27232 = (inp[0]) ? node27236 : node27233;
														assign node27233 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node27236 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27239 = (inp[5]) ? node27243 : node27240;
														assign node27240 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27243 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node27246 = (inp[15]) ? node27260 : node27247;
												assign node27247 = (inp[2]) ? node27255 : node27248;
													assign node27248 = (inp[14]) ? node27252 : node27249;
														assign node27249 = (inp[3]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node27252 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27255 = (inp[14]) ? node27257 : 16'b0000001111111111;
														assign node27257 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27260 = (inp[0]) ? node27268 : node27261;
													assign node27261 = (inp[5]) ? node27265 : node27262;
														assign node27262 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node27265 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27268 = (inp[14]) ? node27272 : node27269;
														assign node27269 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27272 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node27275 = (inp[2]) ? node27301 : node27276;
											assign node27276 = (inp[5]) ? node27290 : node27277;
												assign node27277 = (inp[0]) ? node27285 : node27278;
													assign node27278 = (inp[15]) ? node27282 : node27279;
														assign node27279 = (inp[3]) ? 16'b0000001111111111 : 16'b0000001111111111;
														assign node27282 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
													assign node27285 = (inp[3]) ? 16'b0000000111111111 : node27286;
														assign node27286 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node27290 = (inp[13]) ? node27296 : node27291;
													assign node27291 = (inp[0]) ? node27293 : 16'b0000001111111111;
														assign node27293 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27296 = (inp[3]) ? 16'b0000000001111111 : node27297;
														assign node27297 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
											assign node27301 = (inp[15]) ? node27317 : node27302;
												assign node27302 = (inp[0]) ? node27310 : node27303;
													assign node27303 = (inp[3]) ? node27307 : node27304;
														assign node27304 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27307 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27310 = (inp[14]) ? node27314 : node27311;
														assign node27311 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27314 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27317 = (inp[13]) ? node27325 : node27318;
													assign node27318 = (inp[3]) ? node27322 : node27319;
														assign node27319 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27322 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27325 = (inp[0]) ? 16'b0000000000111111 : node27326;
														assign node27326 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node27330 = (inp[0]) ? node27390 : node27331;
										assign node27331 = (inp[14]) ? node27361 : node27332;
											assign node27332 = (inp[5]) ? node27348 : node27333;
												assign node27333 = (inp[3]) ? node27341 : node27334;
													assign node27334 = (inp[1]) ? node27338 : node27335;
														assign node27335 = (inp[2]) ? 16'b0000001111111111 : 16'b0000111111111111;
														assign node27338 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27341 = (inp[1]) ? node27345 : node27342;
														assign node27342 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27345 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node27348 = (inp[1]) ? node27354 : node27349;
													assign node27349 = (inp[15]) ? 16'b0000000111111111 : node27350;
														assign node27350 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27354 = (inp[15]) ? node27358 : node27355;
														assign node27355 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27358 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000001111111;
											assign node27361 = (inp[2]) ? node27375 : node27362;
												assign node27362 = (inp[13]) ? node27368 : node27363;
													assign node27363 = (inp[3]) ? node27365 : 16'b0000001111111111;
														assign node27365 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27368 = (inp[1]) ? node27372 : node27369;
														assign node27369 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27372 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27375 = (inp[5]) ? node27383 : node27376;
													assign node27376 = (inp[3]) ? node27380 : node27377;
														assign node27377 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27380 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27383 = (inp[15]) ? node27387 : node27384;
														assign node27384 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27387 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node27390 = (inp[3]) ? node27420 : node27391;
											assign node27391 = (inp[14]) ? node27405 : node27392;
												assign node27392 = (inp[5]) ? node27400 : node27393;
													assign node27393 = (inp[15]) ? node27397 : node27394;
														assign node27394 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27397 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27400 = (inp[2]) ? node27402 : 16'b0000000011111111;
														assign node27402 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27405 = (inp[15]) ? node27413 : node27406;
													assign node27406 = (inp[13]) ? node27410 : node27407;
														assign node27407 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27410 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27413 = (inp[2]) ? node27417 : node27414;
														assign node27414 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27417 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node27420 = (inp[1]) ? node27436 : node27421;
												assign node27421 = (inp[5]) ? node27429 : node27422;
													assign node27422 = (inp[15]) ? node27426 : node27423;
														assign node27423 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27426 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
													assign node27429 = (inp[14]) ? node27433 : node27430;
														assign node27430 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node27433 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000111111;
												assign node27436 = (inp[14]) ? node27444 : node27437;
													assign node27437 = (inp[13]) ? node27441 : node27438;
														assign node27438 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node27441 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27444 = (inp[2]) ? node27448 : node27445;
														assign node27445 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node27448 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000011111;
								assign node27451 = (inp[5]) ? node27573 : node27452;
									assign node27452 = (inp[13]) ? node27514 : node27453;
										assign node27453 = (inp[3]) ? node27483 : node27454;
											assign node27454 = (inp[15]) ? node27468 : node27455;
												assign node27455 = (inp[14]) ? node27463 : node27456;
													assign node27456 = (inp[11]) ? node27460 : node27457;
														assign node27457 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node27460 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27463 = (inp[1]) ? 16'b0000000111111111 : node27464;
														assign node27464 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
												assign node27468 = (inp[2]) ? node27476 : node27469;
													assign node27469 = (inp[11]) ? node27473 : node27470;
														assign node27470 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27473 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27476 = (inp[1]) ? node27480 : node27477;
														assign node27477 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27480 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node27483 = (inp[0]) ? node27499 : node27484;
												assign node27484 = (inp[11]) ? node27492 : node27485;
													assign node27485 = (inp[14]) ? node27489 : node27486;
														assign node27486 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27489 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27492 = (inp[1]) ? node27496 : node27493;
														assign node27493 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27496 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27499 = (inp[15]) ? node27507 : node27500;
													assign node27500 = (inp[1]) ? node27504 : node27501;
														assign node27501 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27504 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27507 = (inp[14]) ? node27511 : node27508;
														assign node27508 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27511 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node27514 = (inp[14]) ? node27546 : node27515;
											assign node27515 = (inp[2]) ? node27531 : node27516;
												assign node27516 = (inp[11]) ? node27524 : node27517;
													assign node27517 = (inp[15]) ? node27521 : node27518;
														assign node27518 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node27521 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27524 = (inp[0]) ? node27528 : node27525;
														assign node27525 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27528 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27531 = (inp[15]) ? node27539 : node27532;
													assign node27532 = (inp[1]) ? node27536 : node27533;
														assign node27533 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node27536 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27539 = (inp[0]) ? node27543 : node27540;
														assign node27540 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node27543 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27546 = (inp[11]) ? node27562 : node27547;
												assign node27547 = (inp[1]) ? node27555 : node27548;
													assign node27548 = (inp[15]) ? node27552 : node27549;
														assign node27549 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27552 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27555 = (inp[2]) ? node27559 : node27556;
														assign node27556 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27559 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node27562 = (inp[3]) ? node27568 : node27563;
													assign node27563 = (inp[1]) ? node27565 : 16'b0000000001111111;
														assign node27565 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27568 = (inp[2]) ? 16'b0000000000011111 : node27569;
														assign node27569 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
									assign node27573 = (inp[15]) ? node27637 : node27574;
										assign node27574 = (inp[1]) ? node27606 : node27575;
											assign node27575 = (inp[11]) ? node27591 : node27576;
												assign node27576 = (inp[14]) ? node27584 : node27577;
													assign node27577 = (inp[13]) ? node27581 : node27578;
														assign node27578 = (inp[3]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27581 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27584 = (inp[0]) ? node27588 : node27585;
														assign node27585 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27588 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node27591 = (inp[2]) ? node27599 : node27592;
													assign node27592 = (inp[3]) ? node27596 : node27593;
														assign node27593 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node27596 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27599 = (inp[3]) ? node27603 : node27600;
														assign node27600 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27603 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27606 = (inp[11]) ? node27622 : node27607;
												assign node27607 = (inp[3]) ? node27615 : node27608;
													assign node27608 = (inp[2]) ? node27612 : node27609;
														assign node27609 = (inp[14]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node27612 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27615 = (inp[2]) ? node27619 : node27616;
														assign node27616 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27619 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27622 = (inp[0]) ? node27630 : node27623;
													assign node27623 = (inp[3]) ? node27627 : node27624;
														assign node27624 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27627 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node27630 = (inp[2]) ? node27634 : node27631;
														assign node27631 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27634 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node27637 = (inp[14]) ? node27665 : node27638;
											assign node27638 = (inp[2]) ? node27652 : node27639;
												assign node27639 = (inp[13]) ? node27647 : node27640;
													assign node27640 = (inp[1]) ? node27644 : node27641;
														assign node27641 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27644 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27647 = (inp[3]) ? node27649 : 16'b0000000011111111;
														assign node27649 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node27652 = (inp[11]) ? node27660 : node27653;
													assign node27653 = (inp[0]) ? node27657 : node27654;
														assign node27654 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node27657 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27660 = (inp[13]) ? 16'b0000000000011111 : node27661;
														assign node27661 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27665 = (inp[1]) ? node27677 : node27666;
												assign node27666 = (inp[0]) ? node27672 : node27667;
													assign node27667 = (inp[3]) ? node27669 : 16'b0000000011111111;
														assign node27669 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node27672 = (inp[3]) ? node27674 : 16'b0000000000111111;
														assign node27674 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node27677 = (inp[3]) ? 16'b0000000000011111 : node27678;
													assign node27678 = (inp[2]) ? node27682 : node27679;
														assign node27679 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node27682 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000111111;
							assign node27686 = (inp[14]) ? node27926 : node27687;
								assign node27687 = (inp[15]) ? node27803 : node27688;
									assign node27688 = (inp[5]) ? node27744 : node27689;
										assign node27689 = (inp[0]) ? node27717 : node27690;
											assign node27690 = (inp[7]) ? node27704 : node27691;
												assign node27691 = (inp[11]) ? node27699 : node27692;
													assign node27692 = (inp[1]) ? node27696 : node27693;
														assign node27693 = (inp[2]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node27696 = (inp[13]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node27699 = (inp[2]) ? node27701 : 16'b0000001111111111;
														assign node27701 = (inp[3]) ? 16'b0000000111111111 : 16'b0000000111111111;
												assign node27704 = (inp[2]) ? node27710 : node27705;
													assign node27705 = (inp[13]) ? node27707 : 16'b0000000111111111;
														assign node27707 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27710 = (inp[11]) ? node27714 : node27711;
														assign node27711 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27714 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node27717 = (inp[2]) ? node27731 : node27718;
												assign node27718 = (inp[3]) ? node27724 : node27719;
													assign node27719 = (inp[13]) ? 16'b0000000111111111 : node27720;
														assign node27720 = (inp[1]) ? 16'b0000000111111111 : 16'b0000011111111111;
													assign node27724 = (inp[1]) ? node27728 : node27725;
														assign node27725 = (inp[13]) ? 16'b0000000011111111 : 16'b0000001111111111;
														assign node27728 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27731 = (inp[11]) ? node27739 : node27732;
													assign node27732 = (inp[3]) ? node27736 : node27733;
														assign node27733 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27736 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27739 = (inp[3]) ? node27741 : 16'b0000000001111111;
														assign node27741 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node27744 = (inp[2]) ? node27776 : node27745;
											assign node27745 = (inp[11]) ? node27761 : node27746;
												assign node27746 = (inp[0]) ? node27754 : node27747;
													assign node27747 = (inp[3]) ? node27751 : node27748;
														assign node27748 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27751 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27754 = (inp[7]) ? node27758 : node27755;
														assign node27755 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27758 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27761 = (inp[3]) ? node27769 : node27762;
													assign node27762 = (inp[7]) ? node27766 : node27763;
														assign node27763 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27766 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27769 = (inp[13]) ? node27773 : node27770;
														assign node27770 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27773 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27776 = (inp[11]) ? node27790 : node27777;
												assign node27777 = (inp[0]) ? node27785 : node27778;
													assign node27778 = (inp[13]) ? node27782 : node27779;
														assign node27779 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27782 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27785 = (inp[7]) ? 16'b0000000000111111 : node27786;
														assign node27786 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27790 = (inp[1]) ? node27798 : node27791;
													assign node27791 = (inp[7]) ? node27795 : node27792;
														assign node27792 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node27795 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node27798 = (inp[3]) ? 16'b0000000000011111 : node27799;
														assign node27799 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node27803 = (inp[1]) ? node27867 : node27804;
										assign node27804 = (inp[2]) ? node27836 : node27805;
											assign node27805 = (inp[3]) ? node27821 : node27806;
												assign node27806 = (inp[13]) ? node27814 : node27807;
													assign node27807 = (inp[11]) ? node27811 : node27808;
														assign node27808 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27811 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27814 = (inp[0]) ? node27818 : node27815;
														assign node27815 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node27818 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node27821 = (inp[13]) ? node27829 : node27822;
													assign node27822 = (inp[5]) ? node27826 : node27823;
														assign node27823 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27826 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27829 = (inp[11]) ? node27833 : node27830;
														assign node27830 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node27833 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27836 = (inp[5]) ? node27852 : node27837;
												assign node27837 = (inp[7]) ? node27845 : node27838;
													assign node27838 = (inp[0]) ? node27842 : node27839;
														assign node27839 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27842 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27845 = (inp[0]) ? node27849 : node27846;
														assign node27846 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27849 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27852 = (inp[3]) ? node27860 : node27853;
													assign node27853 = (inp[7]) ? node27857 : node27854;
														assign node27854 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27857 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27860 = (inp[7]) ? node27864 : node27861;
														assign node27861 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27864 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node27867 = (inp[7]) ? node27895 : node27868;
											assign node27868 = (inp[3]) ? node27882 : node27869;
												assign node27869 = (inp[2]) ? node27875 : node27870;
													assign node27870 = (inp[0]) ? 16'b0000000011111111 : node27871;
														assign node27871 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27875 = (inp[11]) ? node27879 : node27876;
														assign node27876 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27879 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27882 = (inp[0]) ? node27890 : node27883;
													assign node27883 = (inp[11]) ? node27887 : node27884;
														assign node27884 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27887 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27890 = (inp[2]) ? 16'b0000000000111111 : node27891;
														assign node27891 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node27895 = (inp[3]) ? node27911 : node27896;
												assign node27896 = (inp[11]) ? node27904 : node27897;
													assign node27897 = (inp[0]) ? node27901 : node27898;
														assign node27898 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node27901 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27904 = (inp[0]) ? node27908 : node27905;
														assign node27905 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node27908 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node27911 = (inp[0]) ? node27919 : node27912;
													assign node27912 = (inp[11]) ? node27916 : node27913;
														assign node27913 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27916 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node27919 = (inp[13]) ? node27923 : node27920;
														assign node27920 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node27923 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000001111;
								assign node27926 = (inp[1]) ? node28048 : node27927;
									assign node27927 = (inp[11]) ? node27989 : node27928;
										assign node27928 = (inp[7]) ? node27958 : node27929;
											assign node27929 = (inp[2]) ? node27945 : node27930;
												assign node27930 = (inp[3]) ? node27938 : node27931;
													assign node27931 = (inp[13]) ? node27935 : node27932;
														assign node27932 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node27935 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node27938 = (inp[5]) ? node27942 : node27939;
														assign node27939 = (inp[13]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27942 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node27945 = (inp[0]) ? node27951 : node27946;
													assign node27946 = (inp[3]) ? node27948 : 16'b0000000111111111;
														assign node27948 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27951 = (inp[15]) ? node27955 : node27952;
														assign node27952 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node27955 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node27958 = (inp[13]) ? node27974 : node27959;
												assign node27959 = (inp[3]) ? node27967 : node27960;
													assign node27960 = (inp[15]) ? node27964 : node27961;
														assign node27961 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node27964 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27967 = (inp[15]) ? node27971 : node27968;
														assign node27968 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27971 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node27974 = (inp[2]) ? node27982 : node27975;
													assign node27975 = (inp[5]) ? node27979 : node27976;
														assign node27976 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node27979 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node27982 = (inp[15]) ? node27986 : node27983;
														assign node27983 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node27986 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node27989 = (inp[3]) ? node28019 : node27990;
											assign node27990 = (inp[15]) ? node28004 : node27991;
												assign node27991 = (inp[13]) ? node27997 : node27992;
													assign node27992 = (inp[0]) ? node27994 : 16'b0000000111111111;
														assign node27994 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node27997 = (inp[2]) ? node28001 : node27998;
														assign node27998 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node28001 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28004 = (inp[0]) ? node28012 : node28005;
													assign node28005 = (inp[13]) ? node28009 : node28006;
														assign node28006 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28009 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28012 = (inp[2]) ? node28016 : node28013;
														assign node28013 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28016 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node28019 = (inp[5]) ? node28035 : node28020;
												assign node28020 = (inp[0]) ? node28028 : node28021;
													assign node28021 = (inp[7]) ? node28025 : node28022;
														assign node28022 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28025 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28028 = (inp[15]) ? node28032 : node28029;
														assign node28029 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28032 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28035 = (inp[7]) ? node28043 : node28036;
													assign node28036 = (inp[2]) ? node28040 : node28037;
														assign node28037 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28040 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28043 = (inp[13]) ? node28045 : 16'b0000000000011111;
														assign node28045 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000011111;
									assign node28048 = (inp[3]) ? node28112 : node28049;
										assign node28049 = (inp[0]) ? node28081 : node28050;
											assign node28050 = (inp[13]) ? node28066 : node28051;
												assign node28051 = (inp[11]) ? node28059 : node28052;
													assign node28052 = (inp[7]) ? node28056 : node28053;
														assign node28053 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node28056 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28059 = (inp[2]) ? node28063 : node28060;
														assign node28060 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28063 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28066 = (inp[11]) ? node28074 : node28067;
													assign node28067 = (inp[7]) ? node28071 : node28068;
														assign node28068 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node28071 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28074 = (inp[15]) ? node28078 : node28075;
														assign node28075 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28078 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node28081 = (inp[5]) ? node28097 : node28082;
												assign node28082 = (inp[15]) ? node28090 : node28083;
													assign node28083 = (inp[2]) ? node28087 : node28084;
														assign node28084 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node28087 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28090 = (inp[11]) ? node28094 : node28091;
														assign node28091 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28094 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28097 = (inp[15]) ? node28105 : node28098;
													assign node28098 = (inp[11]) ? node28102 : node28099;
														assign node28099 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28102 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28105 = (inp[7]) ? node28109 : node28106;
														assign node28106 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node28109 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node28112 = (inp[7]) ? node28140 : node28113;
											assign node28113 = (inp[5]) ? node28129 : node28114;
												assign node28114 = (inp[11]) ? node28122 : node28115;
													assign node28115 = (inp[13]) ? node28119 : node28116;
														assign node28116 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28119 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28122 = (inp[0]) ? node28126 : node28123;
														assign node28123 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28126 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28129 = (inp[0]) ? node28135 : node28130;
													assign node28130 = (inp[11]) ? 16'b0000000000011111 : node28131;
														assign node28131 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28135 = (inp[13]) ? node28137 : 16'b0000000000111111;
														assign node28137 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node28140 = (inp[2]) ? node28156 : node28141;
												assign node28141 = (inp[5]) ? node28149 : node28142;
													assign node28142 = (inp[13]) ? node28146 : node28143;
														assign node28143 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28146 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28149 = (inp[15]) ? node28153 : node28150;
														assign node28150 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28153 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node28156 = (inp[0]) ? node28164 : node28157;
													assign node28157 = (inp[11]) ? node28161 : node28158;
														assign node28158 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28161 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node28164 = (inp[11]) ? node28168 : node28165;
														assign node28165 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node28168 = (inp[15]) ? 16'b0000000000000011 : 16'b0000000000001111;
						assign node28171 = (inp[13]) ? node28651 : node28172;
							assign node28172 = (inp[11]) ? node28406 : node28173;
								assign node28173 = (inp[7]) ? node28289 : node28174;
									assign node28174 = (inp[15]) ? node28234 : node28175;
										assign node28175 = (inp[3]) ? node28203 : node28176;
											assign node28176 = (inp[0]) ? node28190 : node28177;
												assign node28177 = (inp[2]) ? node28183 : node28178;
													assign node28178 = (inp[9]) ? 16'b0000001111111111 : node28179;
														assign node28179 = (inp[1]) ? 16'b0000001111111111 : 16'b0000011111111111;
													assign node28183 = (inp[1]) ? node28187 : node28184;
														assign node28184 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node28187 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node28190 = (inp[2]) ? node28198 : node28191;
													assign node28191 = (inp[9]) ? node28195 : node28192;
														assign node28192 = (inp[5]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node28195 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28198 = (inp[5]) ? node28200 : 16'b0000000111111111;
														assign node28200 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node28203 = (inp[1]) ? node28219 : node28204;
												assign node28204 = (inp[2]) ? node28212 : node28205;
													assign node28205 = (inp[9]) ? node28209 : node28206;
														assign node28206 = (inp[0]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node28209 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28212 = (inp[0]) ? node28216 : node28213;
														assign node28213 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28216 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28219 = (inp[9]) ? node28227 : node28220;
													assign node28220 = (inp[0]) ? node28224 : node28221;
														assign node28221 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28224 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28227 = (inp[2]) ? node28231 : node28228;
														assign node28228 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28231 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
										assign node28234 = (inp[9]) ? node28262 : node28235;
											assign node28235 = (inp[5]) ? node28249 : node28236;
												assign node28236 = (inp[3]) ? node28242 : node28237;
													assign node28237 = (inp[1]) ? 16'b0000000111111111 : node28238;
														assign node28238 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node28242 = (inp[0]) ? node28246 : node28243;
														assign node28243 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node28246 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000001111111;
												assign node28249 = (inp[14]) ? node28257 : node28250;
													assign node28250 = (inp[3]) ? node28254 : node28251;
														assign node28251 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28254 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000111111111;
													assign node28257 = (inp[2]) ? 16'b0000000001111111 : node28258;
														assign node28258 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node28262 = (inp[0]) ? node28276 : node28263;
												assign node28263 = (inp[1]) ? node28271 : node28264;
													assign node28264 = (inp[5]) ? node28268 : node28265;
														assign node28265 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28268 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28271 = (inp[14]) ? 16'b0000000001111111 : node28272;
														assign node28272 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28276 = (inp[3]) ? node28284 : node28277;
													assign node28277 = (inp[1]) ? node28281 : node28278;
														assign node28278 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node28281 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28284 = (inp[5]) ? 16'b0000000000111111 : node28285;
														assign node28285 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
									assign node28289 = (inp[1]) ? node28349 : node28290;
										assign node28290 = (inp[3]) ? node28320 : node28291;
											assign node28291 = (inp[14]) ? node28305 : node28292;
												assign node28292 = (inp[0]) ? node28300 : node28293;
													assign node28293 = (inp[9]) ? node28297 : node28294;
														assign node28294 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node28297 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28300 = (inp[2]) ? node28302 : 16'b0000000111111111;
														assign node28302 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node28305 = (inp[2]) ? node28313 : node28306;
													assign node28306 = (inp[15]) ? node28310 : node28307;
														assign node28307 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28310 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28313 = (inp[0]) ? node28317 : node28314;
														assign node28314 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28317 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node28320 = (inp[2]) ? node28334 : node28321;
												assign node28321 = (inp[9]) ? node28329 : node28322;
													assign node28322 = (inp[15]) ? node28326 : node28323;
														assign node28323 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28326 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28329 = (inp[14]) ? node28331 : 16'b0000000001111111;
														assign node28331 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node28334 = (inp[14]) ? node28342 : node28335;
													assign node28335 = (inp[0]) ? node28339 : node28336;
														assign node28336 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node28339 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28342 = (inp[0]) ? node28346 : node28343;
														assign node28343 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28346 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000111111;
										assign node28349 = (inp[9]) ? node28377 : node28350;
											assign node28350 = (inp[5]) ? node28364 : node28351;
												assign node28351 = (inp[0]) ? node28359 : node28352;
													assign node28352 = (inp[14]) ? node28356 : node28353;
														assign node28353 = (inp[3]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28356 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28359 = (inp[3]) ? 16'b0000000001111111 : node28360;
														assign node28360 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node28364 = (inp[15]) ? node28370 : node28365;
													assign node28365 = (inp[0]) ? 16'b0000000001111111 : node28366;
														assign node28366 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28370 = (inp[2]) ? node28374 : node28371;
														assign node28371 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28374 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node28377 = (inp[15]) ? node28391 : node28378;
												assign node28378 = (inp[14]) ? node28386 : node28379;
													assign node28379 = (inp[3]) ? node28383 : node28380;
														assign node28380 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28383 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node28386 = (inp[2]) ? node28388 : 16'b0000000000111111;
														assign node28388 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node28391 = (inp[5]) ? node28399 : node28392;
													assign node28392 = (inp[2]) ? node28396 : node28393;
														assign node28393 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28396 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28399 = (inp[2]) ? node28403 : node28400;
														assign node28400 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node28403 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node28406 = (inp[3]) ? node28528 : node28407;
									assign node28407 = (inp[7]) ? node28471 : node28408;
										assign node28408 = (inp[5]) ? node28440 : node28409;
											assign node28409 = (inp[9]) ? node28425 : node28410;
												assign node28410 = (inp[15]) ? node28418 : node28411;
													assign node28411 = (inp[14]) ? node28415 : node28412;
														assign node28412 = (inp[1]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node28415 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28418 = (inp[2]) ? node28422 : node28419;
														assign node28419 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28422 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28425 = (inp[1]) ? node28433 : node28426;
													assign node28426 = (inp[15]) ? node28430 : node28427;
														assign node28427 = (inp[0]) ? 16'b0000000111111111 : 16'b0000000011111111;
														assign node28430 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28433 = (inp[14]) ? node28437 : node28434;
														assign node28434 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28437 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node28440 = (inp[15]) ? node28456 : node28441;
												assign node28441 = (inp[1]) ? node28449 : node28442;
													assign node28442 = (inp[2]) ? node28446 : node28443;
														assign node28443 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node28446 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28449 = (inp[2]) ? node28453 : node28450;
														assign node28450 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28453 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28456 = (inp[1]) ? node28464 : node28457;
													assign node28457 = (inp[2]) ? node28461 : node28458;
														assign node28458 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28461 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28464 = (inp[0]) ? node28468 : node28465;
														assign node28465 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28468 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node28471 = (inp[0]) ? node28503 : node28472;
											assign node28472 = (inp[2]) ? node28488 : node28473;
												assign node28473 = (inp[1]) ? node28481 : node28474;
													assign node28474 = (inp[15]) ? node28478 : node28475;
														assign node28475 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node28478 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28481 = (inp[15]) ? node28485 : node28482;
														assign node28482 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node28485 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28488 = (inp[14]) ? node28496 : node28489;
													assign node28489 = (inp[1]) ? node28493 : node28490;
														assign node28490 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28493 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28496 = (inp[9]) ? node28500 : node28497;
														assign node28497 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28500 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node28503 = (inp[9]) ? node28515 : node28504;
												assign node28504 = (inp[15]) ? node28510 : node28505;
													assign node28505 = (inp[1]) ? 16'b0000000000111111 : node28506;
														assign node28506 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28510 = (inp[2]) ? 16'b0000000000111111 : node28511;
														assign node28511 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28515 = (inp[14]) ? node28521 : node28516;
													assign node28516 = (inp[5]) ? 16'b0000000000111111 : node28517;
														assign node28517 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28521 = (inp[2]) ? node28525 : node28522;
														assign node28522 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node28525 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node28528 = (inp[0]) ? node28588 : node28529;
										assign node28529 = (inp[14]) ? node28557 : node28530;
											assign node28530 = (inp[1]) ? node28544 : node28531;
												assign node28531 = (inp[7]) ? node28539 : node28532;
													assign node28532 = (inp[9]) ? node28536 : node28533;
														assign node28533 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28536 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28539 = (inp[2]) ? node28541 : 16'b0000000011111111;
														assign node28541 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28544 = (inp[15]) ? node28550 : node28545;
													assign node28545 = (inp[9]) ? 16'b0000000001111111 : node28546;
														assign node28546 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28550 = (inp[5]) ? node28554 : node28551;
														assign node28551 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28554 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node28557 = (inp[9]) ? node28573 : node28558;
												assign node28558 = (inp[5]) ? node28566 : node28559;
													assign node28559 = (inp[7]) ? node28563 : node28560;
														assign node28560 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28563 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28566 = (inp[7]) ? node28570 : node28567;
														assign node28567 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28570 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28573 = (inp[5]) ? node28581 : node28574;
													assign node28574 = (inp[7]) ? node28578 : node28575;
														assign node28575 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28578 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28581 = (inp[7]) ? node28585 : node28582;
														assign node28582 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28585 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node28588 = (inp[14]) ? node28620 : node28589;
											assign node28589 = (inp[1]) ? node28605 : node28590;
												assign node28590 = (inp[5]) ? node28598 : node28591;
													assign node28591 = (inp[7]) ? node28595 : node28592;
														assign node28592 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28595 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28598 = (inp[9]) ? node28602 : node28599;
														assign node28599 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28602 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28605 = (inp[7]) ? node28613 : node28606;
													assign node28606 = (inp[9]) ? node28610 : node28607;
														assign node28607 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28610 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28613 = (inp[15]) ? node28617 : node28614;
														assign node28614 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28617 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node28620 = (inp[5]) ? node28636 : node28621;
												assign node28621 = (inp[15]) ? node28629 : node28622;
													assign node28622 = (inp[1]) ? node28626 : node28623;
														assign node28623 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28626 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node28629 = (inp[2]) ? node28633 : node28630;
														assign node28630 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28633 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node28636 = (inp[9]) ? node28644 : node28637;
													assign node28637 = (inp[15]) ? node28641 : node28638;
														assign node28638 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node28641 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node28644 = (inp[7]) ? node28648 : node28645;
														assign node28645 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node28648 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node28651 = (inp[1]) ? node28891 : node28652;
								assign node28652 = (inp[14]) ? node28770 : node28653;
									assign node28653 = (inp[7]) ? node28711 : node28654;
										assign node28654 = (inp[9]) ? node28682 : node28655;
											assign node28655 = (inp[15]) ? node28669 : node28656;
												assign node28656 = (inp[2]) ? node28662 : node28657;
													assign node28657 = (inp[5]) ? node28659 : 16'b0000000111111111;
														assign node28659 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node28662 = (inp[3]) ? node28666 : node28663;
														assign node28663 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28666 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28669 = (inp[0]) ? node28675 : node28670;
													assign node28670 = (inp[3]) ? node28672 : 16'b0000000111111111;
														assign node28672 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28675 = (inp[2]) ? node28679 : node28676;
														assign node28676 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28679 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node28682 = (inp[3]) ? node28696 : node28683;
												assign node28683 = (inp[0]) ? node28691 : node28684;
													assign node28684 = (inp[2]) ? node28688 : node28685;
														assign node28685 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28688 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28691 = (inp[11]) ? 16'b0000000000111111 : node28692;
														assign node28692 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node28696 = (inp[2]) ? node28704 : node28697;
													assign node28697 = (inp[5]) ? node28701 : node28698;
														assign node28698 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28701 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28704 = (inp[15]) ? node28708 : node28705;
														assign node28705 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node28708 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node28711 = (inp[15]) ? node28741 : node28712;
											assign node28712 = (inp[11]) ? node28726 : node28713;
												assign node28713 = (inp[5]) ? node28721 : node28714;
													assign node28714 = (inp[0]) ? node28718 : node28715;
														assign node28715 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28718 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28721 = (inp[9]) ? 16'b0000000000111111 : node28722;
														assign node28722 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node28726 = (inp[5]) ? node28734 : node28727;
													assign node28727 = (inp[0]) ? node28731 : node28728;
														assign node28728 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node28731 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28734 = (inp[2]) ? node28738 : node28735;
														assign node28735 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28738 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node28741 = (inp[5]) ? node28757 : node28742;
												assign node28742 = (inp[2]) ? node28750 : node28743;
													assign node28743 = (inp[9]) ? node28747 : node28744;
														assign node28744 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node28747 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node28750 = (inp[3]) ? node28754 : node28751;
														assign node28751 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28754 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28757 = (inp[0]) ? node28763 : node28758;
													assign node28758 = (inp[9]) ? node28760 : 16'b0000000001111111;
														assign node28760 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28763 = (inp[9]) ? node28767 : node28764;
														assign node28764 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28767 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000011111;
									assign node28770 = (inp[5]) ? node28830 : node28771;
										assign node28771 = (inp[0]) ? node28801 : node28772;
											assign node28772 = (inp[11]) ? node28786 : node28773;
												assign node28773 = (inp[15]) ? node28779 : node28774;
													assign node28774 = (inp[7]) ? node28776 : 16'b0000000011111111;
														assign node28776 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28779 = (inp[3]) ? node28783 : node28780;
														assign node28780 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28783 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28786 = (inp[15]) ? node28794 : node28787;
													assign node28787 = (inp[2]) ? node28791 : node28788;
														assign node28788 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28791 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28794 = (inp[3]) ? node28798 : node28795;
														assign node28795 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28798 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node28801 = (inp[7]) ? node28815 : node28802;
												assign node28802 = (inp[11]) ? node28808 : node28803;
													assign node28803 = (inp[15]) ? node28805 : 16'b0000000011111111;
														assign node28805 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28808 = (inp[9]) ? node28812 : node28809;
														assign node28809 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28812 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28815 = (inp[3]) ? node28823 : node28816;
													assign node28816 = (inp[11]) ? node28820 : node28817;
														assign node28817 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28820 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28823 = (inp[15]) ? node28827 : node28824;
														assign node28824 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28827 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node28830 = (inp[9]) ? node28860 : node28831;
											assign node28831 = (inp[3]) ? node28845 : node28832;
												assign node28832 = (inp[15]) ? node28838 : node28833;
													assign node28833 = (inp[0]) ? node28835 : 16'b0000000011111111;
														assign node28835 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28838 = (inp[7]) ? node28842 : node28839;
														assign node28839 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28842 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28845 = (inp[11]) ? node28853 : node28846;
													assign node28846 = (inp[2]) ? node28850 : node28847;
														assign node28847 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node28850 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28853 = (inp[2]) ? node28857 : node28854;
														assign node28854 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28857 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000001111;
											assign node28860 = (inp[11]) ? node28876 : node28861;
												assign node28861 = (inp[3]) ? node28869 : node28862;
													assign node28862 = (inp[0]) ? node28866 : node28863;
														assign node28863 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28866 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28869 = (inp[0]) ? node28873 : node28870;
														assign node28870 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28873 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node28876 = (inp[15]) ? node28884 : node28877;
													assign node28877 = (inp[7]) ? node28881 : node28878;
														assign node28878 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node28881 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node28884 = (inp[2]) ? node28888 : node28885;
														assign node28885 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node28888 = (inp[3]) ? 16'b0000000000000011 : 16'b0000000000001111;
								assign node28891 = (inp[0]) ? node29013 : node28892;
									assign node28892 = (inp[15]) ? node28952 : node28893;
										assign node28893 = (inp[5]) ? node28923 : node28894;
											assign node28894 = (inp[3]) ? node28910 : node28895;
												assign node28895 = (inp[7]) ? node28903 : node28896;
													assign node28896 = (inp[14]) ? node28900 : node28897;
														assign node28897 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node28900 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node28903 = (inp[9]) ? node28907 : node28904;
														assign node28904 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28907 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28910 = (inp[2]) ? node28918 : node28911;
													assign node28911 = (inp[11]) ? node28915 : node28912;
														assign node28912 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node28915 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28918 = (inp[9]) ? 16'b0000000000111111 : node28919;
														assign node28919 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node28923 = (inp[14]) ? node28937 : node28924;
												assign node28924 = (inp[9]) ? node28932 : node28925;
													assign node28925 = (inp[2]) ? node28929 : node28926;
														assign node28926 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node28929 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28932 = (inp[3]) ? 16'b0000000000011111 : node28933;
														assign node28933 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node28937 = (inp[2]) ? node28945 : node28938;
													assign node28938 = (inp[3]) ? node28942 : node28939;
														assign node28939 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node28942 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28945 = (inp[7]) ? node28949 : node28946;
														assign node28946 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28949 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000001111;
										assign node28952 = (inp[7]) ? node28984 : node28953;
											assign node28953 = (inp[14]) ? node28969 : node28954;
												assign node28954 = (inp[11]) ? node28962 : node28955;
													assign node28955 = (inp[3]) ? node28959 : node28956;
														assign node28956 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node28959 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node28962 = (inp[5]) ? node28966 : node28963;
														assign node28963 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000000111111;
														assign node28966 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28969 = (inp[2]) ? node28977 : node28970;
													assign node28970 = (inp[5]) ? node28974 : node28971;
														assign node28971 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28974 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28977 = (inp[3]) ? node28981 : node28978;
														assign node28978 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node28981 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node28984 = (inp[11]) ? node28998 : node28985;
												assign node28985 = (inp[5]) ? node28993 : node28986;
													assign node28986 = (inp[2]) ? node28990 : node28987;
														assign node28987 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node28990 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node28993 = (inp[9]) ? 16'b0000000000001111 : node28994;
														assign node28994 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node28998 = (inp[2]) ? node29006 : node28999;
													assign node28999 = (inp[9]) ? node29003 : node29000;
														assign node29000 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node29003 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node29006 = (inp[5]) ? node29010 : node29007;
														assign node29007 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node29010 = (inp[3]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node29013 = (inp[9]) ? node29075 : node29014;
										assign node29014 = (inp[11]) ? node29044 : node29015;
											assign node29015 = (inp[2]) ? node29031 : node29016;
												assign node29016 = (inp[14]) ? node29024 : node29017;
													assign node29017 = (inp[5]) ? node29021 : node29018;
														assign node29018 = (inp[3]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29021 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node29024 = (inp[7]) ? node29028 : node29025;
														assign node29025 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29028 = (inp[3]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29031 = (inp[5]) ? node29039 : node29032;
													assign node29032 = (inp[15]) ? node29036 : node29033;
														assign node29033 = (inp[3]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29036 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node29039 = (inp[14]) ? node29041 : 16'b0000000000011111;
														assign node29041 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node29044 = (inp[2]) ? node29060 : node29045;
												assign node29045 = (inp[14]) ? node29053 : node29046;
													assign node29046 = (inp[3]) ? node29050 : node29047;
														assign node29047 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29050 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29053 = (inp[3]) ? node29057 : node29054;
														assign node29054 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29057 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node29060 = (inp[7]) ? node29068 : node29061;
													assign node29061 = (inp[5]) ? node29065 : node29062;
														assign node29062 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29065 = (inp[3]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node29068 = (inp[15]) ? node29072 : node29069;
														assign node29069 = (inp[14]) ? 16'b0000000000000111 : 16'b0000000000011111;
														assign node29072 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node29075 = (inp[3]) ? node29105 : node29076;
											assign node29076 = (inp[14]) ? node29090 : node29077;
												assign node29077 = (inp[5]) ? node29085 : node29078;
													assign node29078 = (inp[15]) ? node29082 : node29079;
														assign node29079 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29082 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29085 = (inp[7]) ? 16'b0000000000001111 : node29086;
														assign node29086 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29090 = (inp[15]) ? node29098 : node29091;
													assign node29091 = (inp[7]) ? node29095 : node29092;
														assign node29092 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29095 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node29098 = (inp[11]) ? node29102 : node29099;
														assign node29099 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node29102 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node29105 = (inp[11]) ? node29121 : node29106;
												assign node29106 = (inp[14]) ? node29114 : node29107;
													assign node29107 = (inp[7]) ? node29111 : node29108;
														assign node29108 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29111 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000011111;
													assign node29114 = (inp[2]) ? node29118 : node29115;
														assign node29115 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node29118 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node29121 = (inp[14]) ? node29129 : node29122;
													assign node29122 = (inp[7]) ? node29126 : node29123;
														assign node29123 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node29126 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node29129 = (inp[5]) ? node29133 : node29130;
														assign node29130 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node29133 = (inp[7]) ? 16'b0000000000000011 : 16'b0000000000000111;
					assign node29136 = (inp[3]) ? node30110 : node29137;
						assign node29137 = (inp[9]) ? node29625 : node29138;
							assign node29138 = (inp[7]) ? node29382 : node29139;
								assign node29139 = (inp[12]) ? node29257 : node29140;
									assign node29140 = (inp[1]) ? node29200 : node29141;
										assign node29141 = (inp[13]) ? node29173 : node29142;
											assign node29142 = (inp[2]) ? node29158 : node29143;
												assign node29143 = (inp[14]) ? node29151 : node29144;
													assign node29144 = (inp[0]) ? node29148 : node29145;
														assign node29145 = (inp[11]) ? 16'b0000001111111111 : 16'b0000011111111111;
														assign node29148 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node29151 = (inp[5]) ? node29155 : node29152;
														assign node29152 = (inp[0]) ? 16'b0000000111111111 : 16'b0000011111111111;
														assign node29155 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node29158 = (inp[5]) ? node29166 : node29159;
													assign node29159 = (inp[14]) ? node29163 : node29160;
														assign node29160 = (inp[11]) ? 16'b0000000111111111 : 16'b0000000111111111;
														assign node29163 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29166 = (inp[15]) ? node29170 : node29167;
														assign node29167 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29170 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
											assign node29173 = (inp[5]) ? node29189 : node29174;
												assign node29174 = (inp[0]) ? node29182 : node29175;
													assign node29175 = (inp[2]) ? node29179 : node29176;
														assign node29176 = (inp[15]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29179 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29182 = (inp[15]) ? node29186 : node29183;
														assign node29183 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29186 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29189 = (inp[11]) ? node29195 : node29190;
													assign node29190 = (inp[0]) ? node29192 : 16'b0000000011111111;
														assign node29192 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
													assign node29195 = (inp[14]) ? 16'b0000000001111111 : node29196;
														assign node29196 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
										assign node29200 = (inp[11]) ? node29228 : node29201;
											assign node29201 = (inp[14]) ? node29215 : node29202;
												assign node29202 = (inp[13]) ? node29208 : node29203;
													assign node29203 = (inp[0]) ? 16'b0000000111111111 : node29204;
														assign node29204 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
													assign node29208 = (inp[5]) ? node29212 : node29209;
														assign node29209 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29212 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29215 = (inp[0]) ? node29221 : node29216;
													assign node29216 = (inp[13]) ? node29218 : 16'b0000000011111111;
														assign node29218 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29221 = (inp[5]) ? node29225 : node29222;
														assign node29222 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29225 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node29228 = (inp[5]) ? node29242 : node29229;
												assign node29229 = (inp[14]) ? node29235 : node29230;
													assign node29230 = (inp[0]) ? node29232 : 16'b0000000011111111;
														assign node29232 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29235 = (inp[0]) ? node29239 : node29236;
														assign node29236 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29239 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29242 = (inp[14]) ? node29250 : node29243;
													assign node29243 = (inp[0]) ? node29247 : node29244;
														assign node29244 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29247 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29250 = (inp[15]) ? node29254 : node29251;
														assign node29251 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29254 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
									assign node29257 = (inp[15]) ? node29319 : node29258;
										assign node29258 = (inp[13]) ? node29290 : node29259;
											assign node29259 = (inp[0]) ? node29275 : node29260;
												assign node29260 = (inp[11]) ? node29268 : node29261;
													assign node29261 = (inp[5]) ? node29265 : node29262;
														assign node29262 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29265 = (inp[1]) ? 16'b0000000111111111 : 16'b0000000111111111;
													assign node29268 = (inp[2]) ? node29272 : node29269;
														assign node29269 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29272 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node29275 = (inp[11]) ? node29283 : node29276;
													assign node29276 = (inp[2]) ? node29280 : node29277;
														assign node29277 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29280 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000011111111;
													assign node29283 = (inp[1]) ? node29287 : node29284;
														assign node29284 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29287 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000001111111;
											assign node29290 = (inp[0]) ? node29304 : node29291;
												assign node29291 = (inp[5]) ? node29297 : node29292;
													assign node29292 = (inp[11]) ? node29294 : 16'b0000000011111111;
														assign node29294 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29297 = (inp[2]) ? node29301 : node29298;
														assign node29298 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29301 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29304 = (inp[14]) ? node29312 : node29305;
													assign node29305 = (inp[5]) ? node29309 : node29306;
														assign node29306 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29309 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29312 = (inp[2]) ? node29316 : node29313;
														assign node29313 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29316 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node29319 = (inp[0]) ? node29351 : node29320;
											assign node29320 = (inp[2]) ? node29336 : node29321;
												assign node29321 = (inp[11]) ? node29329 : node29322;
													assign node29322 = (inp[5]) ? node29326 : node29323;
														assign node29323 = (inp[14]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29326 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29329 = (inp[13]) ? node29333 : node29330;
														assign node29330 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29333 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29336 = (inp[14]) ? node29344 : node29337;
													assign node29337 = (inp[1]) ? node29341 : node29338;
														assign node29338 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29341 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29344 = (inp[13]) ? node29348 : node29345;
														assign node29345 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29348 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node29351 = (inp[1]) ? node29367 : node29352;
												assign node29352 = (inp[11]) ? node29360 : node29353;
													assign node29353 = (inp[13]) ? node29357 : node29354;
														assign node29354 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29357 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node29360 = (inp[5]) ? node29364 : node29361;
														assign node29361 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node29364 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29367 = (inp[2]) ? node29375 : node29368;
													assign node29368 = (inp[14]) ? node29372 : node29369;
														assign node29369 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node29372 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29375 = (inp[13]) ? node29379 : node29376;
														assign node29376 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node29379 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
								assign node29382 = (inp[13]) ? node29502 : node29383;
									assign node29383 = (inp[0]) ? node29441 : node29384;
										assign node29384 = (inp[5]) ? node29414 : node29385;
											assign node29385 = (inp[14]) ? node29399 : node29386;
												assign node29386 = (inp[12]) ? node29394 : node29387;
													assign node29387 = (inp[2]) ? node29391 : node29388;
														assign node29388 = (inp[11]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29391 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29394 = (inp[2]) ? 16'b0000000011111111 : node29395;
														assign node29395 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node29399 = (inp[12]) ? node29407 : node29400;
													assign node29400 = (inp[15]) ? node29404 : node29401;
														assign node29401 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29404 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29407 = (inp[11]) ? node29411 : node29408;
														assign node29408 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29411 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node29414 = (inp[12]) ? node29430 : node29415;
												assign node29415 = (inp[2]) ? node29423 : node29416;
													assign node29416 = (inp[11]) ? node29420 : node29417;
														assign node29417 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29420 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29423 = (inp[1]) ? node29427 : node29424;
														assign node29424 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29427 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29430 = (inp[11]) ? node29436 : node29431;
													assign node29431 = (inp[14]) ? node29433 : 16'b0000000001111111;
														assign node29433 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29436 = (inp[14]) ? 16'b0000000000111111 : node29437;
														assign node29437 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
										assign node29441 = (inp[14]) ? node29471 : node29442;
											assign node29442 = (inp[2]) ? node29456 : node29443;
												assign node29443 = (inp[11]) ? node29449 : node29444;
													assign node29444 = (inp[1]) ? node29446 : 16'b0000000111111111;
														assign node29446 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29449 = (inp[12]) ? node29453 : node29450;
														assign node29450 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29453 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node29456 = (inp[11]) ? node29464 : node29457;
													assign node29457 = (inp[12]) ? node29461 : node29458;
														assign node29458 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29461 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29464 = (inp[1]) ? node29468 : node29465;
														assign node29465 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29468 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node29471 = (inp[5]) ? node29487 : node29472;
												assign node29472 = (inp[11]) ? node29480 : node29473;
													assign node29473 = (inp[15]) ? node29477 : node29474;
														assign node29474 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29477 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29480 = (inp[15]) ? node29484 : node29481;
														assign node29481 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29484 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node29487 = (inp[2]) ? node29495 : node29488;
													assign node29488 = (inp[11]) ? node29492 : node29489;
														assign node29489 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29492 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29495 = (inp[1]) ? node29499 : node29496;
														assign node29496 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29499 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000001111;
									assign node29502 = (inp[1]) ? node29564 : node29503;
										assign node29503 = (inp[11]) ? node29535 : node29504;
											assign node29504 = (inp[12]) ? node29520 : node29505;
												assign node29505 = (inp[0]) ? node29513 : node29506;
													assign node29506 = (inp[15]) ? node29510 : node29507;
														assign node29507 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29510 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29513 = (inp[5]) ? node29517 : node29514;
														assign node29514 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29517 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29520 = (inp[2]) ? node29528 : node29521;
													assign node29521 = (inp[5]) ? node29525 : node29522;
														assign node29522 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29525 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29528 = (inp[14]) ? node29532 : node29529;
														assign node29529 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29532 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
											assign node29535 = (inp[5]) ? node29551 : node29536;
												assign node29536 = (inp[12]) ? node29544 : node29537;
													assign node29537 = (inp[14]) ? node29541 : node29538;
														assign node29538 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node29541 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29544 = (inp[14]) ? node29548 : node29545;
														assign node29545 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29548 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29551 = (inp[0]) ? node29559 : node29552;
													assign node29552 = (inp[12]) ? node29556 : node29553;
														assign node29553 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node29556 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29559 = (inp[2]) ? 16'b0000000000011111 : node29560;
														assign node29560 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node29564 = (inp[5]) ? node29596 : node29565;
											assign node29565 = (inp[15]) ? node29581 : node29566;
												assign node29566 = (inp[2]) ? node29574 : node29567;
													assign node29567 = (inp[14]) ? node29571 : node29568;
														assign node29568 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node29571 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29574 = (inp[11]) ? node29578 : node29575;
														assign node29575 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29578 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29581 = (inp[11]) ? node29589 : node29582;
													assign node29582 = (inp[12]) ? node29586 : node29583;
														assign node29583 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29586 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
													assign node29589 = (inp[14]) ? node29593 : node29590;
														assign node29590 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29593 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node29596 = (inp[11]) ? node29612 : node29597;
												assign node29597 = (inp[2]) ? node29605 : node29598;
													assign node29598 = (inp[0]) ? node29602 : node29599;
														assign node29599 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29602 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29605 = (inp[12]) ? node29609 : node29606;
														assign node29606 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29609 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node29612 = (inp[0]) ? node29618 : node29613;
													assign node29613 = (inp[15]) ? 16'b0000000000001111 : node29614;
														assign node29614 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node29618 = (inp[15]) ? node29622 : node29619;
														assign node29619 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node29622 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
							assign node29625 = (inp[1]) ? node29867 : node29626;
								assign node29626 = (inp[7]) ? node29748 : node29627;
									assign node29627 = (inp[11]) ? node29687 : node29628;
										assign node29628 = (inp[13]) ? node29656 : node29629;
											assign node29629 = (inp[14]) ? node29645 : node29630;
												assign node29630 = (inp[15]) ? node29638 : node29631;
													assign node29631 = (inp[5]) ? node29635 : node29632;
														assign node29632 = (inp[2]) ? 16'b0000000111111111 : 16'b0000001111111111;
														assign node29635 = (inp[2]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node29638 = (inp[2]) ? node29642 : node29639;
														assign node29639 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29642 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
												assign node29645 = (inp[15]) ? node29653 : node29646;
													assign node29646 = (inp[12]) ? node29650 : node29647;
														assign node29647 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node29650 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29653 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000000111111;
											assign node29656 = (inp[0]) ? node29672 : node29657;
												assign node29657 = (inp[15]) ? node29665 : node29658;
													assign node29658 = (inp[2]) ? node29662 : node29659;
														assign node29659 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29662 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29665 = (inp[5]) ? node29669 : node29666;
														assign node29666 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29669 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29672 = (inp[14]) ? node29680 : node29673;
													assign node29673 = (inp[15]) ? node29677 : node29674;
														assign node29674 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29677 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29680 = (inp[5]) ? node29684 : node29681;
														assign node29681 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29684 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
										assign node29687 = (inp[13]) ? node29717 : node29688;
											assign node29688 = (inp[5]) ? node29702 : node29689;
												assign node29689 = (inp[0]) ? node29697 : node29690;
													assign node29690 = (inp[2]) ? node29694 : node29691;
														assign node29691 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29694 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29697 = (inp[15]) ? node29699 : 16'b0000000011111111;
														assign node29699 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29702 = (inp[12]) ? node29710 : node29703;
													assign node29703 = (inp[14]) ? node29707 : node29704;
														assign node29704 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node29707 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29710 = (inp[15]) ? node29714 : node29711;
														assign node29711 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29714 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node29717 = (inp[2]) ? node29733 : node29718;
												assign node29718 = (inp[15]) ? node29726 : node29719;
													assign node29719 = (inp[5]) ? node29723 : node29720;
														assign node29720 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node29723 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29726 = (inp[5]) ? node29730 : node29727;
														assign node29727 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29730 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29733 = (inp[14]) ? node29741 : node29734;
													assign node29734 = (inp[0]) ? node29738 : node29735;
														assign node29735 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node29738 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29741 = (inp[0]) ? node29745 : node29742;
														assign node29742 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29745 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node29748 = (inp[13]) ? node29812 : node29749;
										assign node29749 = (inp[14]) ? node29781 : node29750;
											assign node29750 = (inp[5]) ? node29766 : node29751;
												assign node29751 = (inp[0]) ? node29759 : node29752;
													assign node29752 = (inp[2]) ? node29756 : node29753;
														assign node29753 = (inp[15]) ? 16'b0000000011111111 : 16'b0000000011111111;
														assign node29756 = (inp[15]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29759 = (inp[12]) ? node29763 : node29760;
														assign node29760 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29763 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node29766 = (inp[0]) ? node29774 : node29767;
													assign node29767 = (inp[15]) ? node29771 : node29768;
														assign node29768 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29771 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node29774 = (inp[2]) ? node29778 : node29775;
														assign node29775 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29778 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node29781 = (inp[15]) ? node29797 : node29782;
												assign node29782 = (inp[0]) ? node29790 : node29783;
													assign node29783 = (inp[12]) ? node29787 : node29784;
														assign node29784 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node29787 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29790 = (inp[11]) ? node29794 : node29791;
														assign node29791 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29794 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29797 = (inp[12]) ? node29805 : node29798;
													assign node29798 = (inp[5]) ? node29802 : node29799;
														assign node29799 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29802 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29805 = (inp[11]) ? node29809 : node29806;
														assign node29806 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29809 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node29812 = (inp[2]) ? node29844 : node29813;
											assign node29813 = (inp[11]) ? node29829 : node29814;
												assign node29814 = (inp[5]) ? node29822 : node29815;
													assign node29815 = (inp[15]) ? node29819 : node29816;
														assign node29816 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29819 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29822 = (inp[14]) ? node29826 : node29823;
														assign node29823 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node29826 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29829 = (inp[14]) ? node29837 : node29830;
													assign node29830 = (inp[0]) ? node29834 : node29831;
														assign node29831 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29834 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29837 = (inp[0]) ? node29841 : node29838;
														assign node29838 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29841 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000001111;
											assign node29844 = (inp[14]) ? node29856 : node29845;
												assign node29845 = (inp[0]) ? node29849 : node29846;
													assign node29846 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29849 = (inp[12]) ? node29853 : node29850;
														assign node29850 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29853 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node29856 = (inp[12]) ? node29862 : node29857;
													assign node29857 = (inp[5]) ? 16'b0000000000001111 : node29858;
														assign node29858 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29862 = (inp[5]) ? node29864 : 16'b0000000000001111;
														assign node29864 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
								assign node29867 = (inp[13]) ? node29989 : node29868;
									assign node29868 = (inp[12]) ? node29930 : node29869;
										assign node29869 = (inp[5]) ? node29901 : node29870;
											assign node29870 = (inp[2]) ? node29886 : node29871;
												assign node29871 = (inp[7]) ? node29879 : node29872;
													assign node29872 = (inp[14]) ? node29876 : node29873;
														assign node29873 = (inp[0]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node29876 = (inp[11]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node29879 = (inp[15]) ? node29883 : node29880;
														assign node29880 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29883 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000001111111;
												assign node29886 = (inp[11]) ? node29894 : node29887;
													assign node29887 = (inp[0]) ? node29891 : node29888;
														assign node29888 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29891 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29894 = (inp[15]) ? node29898 : node29895;
														assign node29895 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29898 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node29901 = (inp[15]) ? node29915 : node29902;
												assign node29902 = (inp[14]) ? node29908 : node29903;
													assign node29903 = (inp[0]) ? node29905 : 16'b0000000011111111;
														assign node29905 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node29908 = (inp[7]) ? node29912 : node29909;
														assign node29909 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node29912 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000111111;
												assign node29915 = (inp[11]) ? node29923 : node29916;
													assign node29916 = (inp[7]) ? node29920 : node29917;
														assign node29917 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29920 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29923 = (inp[14]) ? node29927 : node29924;
														assign node29924 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29927 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node29930 = (inp[11]) ? node29960 : node29931;
											assign node29931 = (inp[15]) ? node29947 : node29932;
												assign node29932 = (inp[2]) ? node29940 : node29933;
													assign node29933 = (inp[7]) ? node29937 : node29934;
														assign node29934 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29937 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
													assign node29940 = (inp[0]) ? node29944 : node29941;
														assign node29941 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29944 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node29947 = (inp[7]) ? node29955 : node29948;
													assign node29948 = (inp[0]) ? node29952 : node29949;
														assign node29949 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node29952 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29955 = (inp[0]) ? node29957 : 16'b0000000000011111;
														assign node29957 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node29960 = (inp[14]) ? node29976 : node29961;
												assign node29961 = (inp[2]) ? node29969 : node29962;
													assign node29962 = (inp[5]) ? node29966 : node29963;
														assign node29963 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node29966 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node29969 = (inp[7]) ? node29973 : node29970;
														assign node29970 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node29973 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node29976 = (inp[7]) ? node29982 : node29977;
													assign node29977 = (inp[2]) ? node29979 : 16'b0000000000011111;
														assign node29979 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node29982 = (inp[15]) ? node29986 : node29983;
														assign node29983 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node29986 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node29989 = (inp[5]) ? node30053 : node29990;
										assign node29990 = (inp[2]) ? node30022 : node29991;
											assign node29991 = (inp[11]) ? node30007 : node29992;
												assign node29992 = (inp[0]) ? node30000 : node29993;
													assign node29993 = (inp[12]) ? node29997 : node29994;
														assign node29994 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node29997 = (inp[15]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30000 = (inp[14]) ? node30004 : node30001;
														assign node30001 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30004 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30007 = (inp[0]) ? node30015 : node30008;
													assign node30008 = (inp[7]) ? node30012 : node30009;
														assign node30009 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30012 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30015 = (inp[15]) ? node30019 : node30016;
														assign node30016 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30019 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node30022 = (inp[0]) ? node30038 : node30023;
												assign node30023 = (inp[7]) ? node30031 : node30024;
													assign node30024 = (inp[14]) ? node30028 : node30025;
														assign node30025 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node30028 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30031 = (inp[12]) ? node30035 : node30032;
														assign node30032 = (inp[15]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30035 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30038 = (inp[11]) ? node30046 : node30039;
													assign node30039 = (inp[7]) ? node30043 : node30040;
														assign node30040 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30043 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30046 = (inp[14]) ? node30050 : node30047;
														assign node30047 = (inp[15]) ? 16'b0000000000001111 : 16'b0000000000111111;
														assign node30050 = (inp[15]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node30053 = (inp[14]) ? node30079 : node30054;
											assign node30054 = (inp[15]) ? node30064 : node30055;
												assign node30055 = (inp[12]) ? node30059 : node30056;
													assign node30056 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30059 = (inp[7]) ? 16'b0000000000011111 : node30060;
														assign node30060 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30064 = (inp[7]) ? node30072 : node30065;
													assign node30065 = (inp[0]) ? node30069 : node30066;
														assign node30066 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30069 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30072 = (inp[12]) ? node30076 : node30073;
														assign node30073 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30076 = (inp[11]) ? 16'b0000000000000011 : 16'b0000000000001111;
											assign node30079 = (inp[15]) ? node30095 : node30080;
												assign node30080 = (inp[12]) ? node30088 : node30081;
													assign node30081 = (inp[7]) ? node30085 : node30082;
														assign node30082 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node30085 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30088 = (inp[0]) ? node30092 : node30089;
														assign node30089 = (inp[11]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30092 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node30095 = (inp[0]) ? node30103 : node30096;
													assign node30096 = (inp[11]) ? node30100 : node30097;
														assign node30097 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30100 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000000111;
													assign node30103 = (inp[12]) ? node30107 : node30104;
														assign node30104 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node30107 = (inp[7]) ? 16'b0000000000000011 : 16'b0000000000000111;
						assign node30110 = (inp[15]) ? node30586 : node30111;
							assign node30111 = (inp[0]) ? node30351 : node30112;
								assign node30112 = (inp[12]) ? node30228 : node30113;
									assign node30113 = (inp[5]) ? node30173 : node30114;
										assign node30114 = (inp[13]) ? node30142 : node30115;
											assign node30115 = (inp[11]) ? node30127 : node30116;
												assign node30116 = (inp[7]) ? node30122 : node30117;
													assign node30117 = (inp[2]) ? node30119 : 16'b0000001111111111;
														assign node30119 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node30122 = (inp[1]) ? 16'b0000000011111111 : node30123;
														assign node30123 = (inp[14]) ? 16'b0000000011111111 : 16'b0000000111111111;
												assign node30127 = (inp[9]) ? node30135 : node30128;
													assign node30128 = (inp[14]) ? node30132 : node30129;
														assign node30129 = (inp[1]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30132 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30135 = (inp[14]) ? node30139 : node30136;
														assign node30136 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30139 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000001111111;
											assign node30142 = (inp[1]) ? node30158 : node30143;
												assign node30143 = (inp[11]) ? node30151 : node30144;
													assign node30144 = (inp[2]) ? node30148 : node30145;
														assign node30145 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node30148 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30151 = (inp[14]) ? node30155 : node30152;
														assign node30152 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30155 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30158 = (inp[11]) ? node30166 : node30159;
													assign node30159 = (inp[14]) ? node30163 : node30160;
														assign node30160 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30163 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30166 = (inp[14]) ? node30170 : node30167;
														assign node30167 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30170 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000011111;
										assign node30173 = (inp[11]) ? node30203 : node30174;
											assign node30174 = (inp[7]) ? node30190 : node30175;
												assign node30175 = (inp[2]) ? node30183 : node30176;
													assign node30176 = (inp[13]) ? node30180 : node30177;
														assign node30177 = (inp[9]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30180 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30183 = (inp[9]) ? node30187 : node30184;
														assign node30184 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30187 = (inp[1]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node30190 = (inp[2]) ? node30198 : node30191;
													assign node30191 = (inp[14]) ? node30195 : node30192;
														assign node30192 = (inp[9]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node30195 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30198 = (inp[1]) ? node30200 : 16'b0000000000111111;
														assign node30200 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
											assign node30203 = (inp[13]) ? node30217 : node30204;
												assign node30204 = (inp[1]) ? node30210 : node30205;
													assign node30205 = (inp[2]) ? node30207 : 16'b0000000001111111;
														assign node30207 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30210 = (inp[9]) ? node30214 : node30211;
														assign node30211 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node30214 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30217 = (inp[9]) ? node30223 : node30218;
													assign node30218 = (inp[1]) ? node30220 : 16'b0000000000111111;
														assign node30220 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30223 = (inp[1]) ? node30225 : 16'b0000000000011111;
														assign node30225 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
									assign node30228 = (inp[11]) ? node30290 : node30229;
										assign node30229 = (inp[2]) ? node30261 : node30230;
											assign node30230 = (inp[7]) ? node30246 : node30231;
												assign node30231 = (inp[14]) ? node30239 : node30232;
													assign node30232 = (inp[1]) ? node30236 : node30233;
														assign node30233 = (inp[5]) ? 16'b0000000011111111 : 16'b0000000111111111;
														assign node30236 = (inp[13]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30239 = (inp[9]) ? node30243 : node30240;
														assign node30240 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30243 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000001111111;
												assign node30246 = (inp[13]) ? node30254 : node30247;
													assign node30247 = (inp[5]) ? node30251 : node30248;
														assign node30248 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30251 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node30254 = (inp[14]) ? node30258 : node30255;
														assign node30255 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30258 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30261 = (inp[1]) ? node30275 : node30262;
												assign node30262 = (inp[13]) ? node30268 : node30263;
													assign node30263 = (inp[14]) ? node30265 : 16'b0000000001111111;
														assign node30265 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30268 = (inp[9]) ? node30272 : node30269;
														assign node30269 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node30272 = (inp[14]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30275 = (inp[9]) ? node30283 : node30276;
													assign node30276 = (inp[7]) ? node30280 : node30277;
														assign node30277 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node30280 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30283 = (inp[13]) ? node30287 : node30284;
														assign node30284 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node30287 = (inp[14]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node30290 = (inp[1]) ? node30320 : node30291;
											assign node30291 = (inp[2]) ? node30305 : node30292;
												assign node30292 = (inp[7]) ? node30300 : node30293;
													assign node30293 = (inp[13]) ? node30297 : node30294;
														assign node30294 = (inp[14]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node30297 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30300 = (inp[5]) ? node30302 : 16'b0000000000111111;
														assign node30302 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
												assign node30305 = (inp[9]) ? node30313 : node30306;
													assign node30306 = (inp[7]) ? node30310 : node30307;
														assign node30307 = (inp[14]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30310 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30313 = (inp[14]) ? node30317 : node30314;
														assign node30314 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30317 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node30320 = (inp[9]) ? node30336 : node30321;
												assign node30321 = (inp[5]) ? node30329 : node30322;
													assign node30322 = (inp[2]) ? node30326 : node30323;
														assign node30323 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30326 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node30329 = (inp[14]) ? node30333 : node30330;
														assign node30330 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30333 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30336 = (inp[7]) ? node30344 : node30337;
													assign node30337 = (inp[14]) ? node30341 : node30338;
														assign node30338 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30341 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30344 = (inp[14]) ? node30348 : node30345;
														assign node30345 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node30348 = (inp[2]) ? 16'b0000000000000011 : 16'b0000000000001111;
								assign node30351 = (inp[14]) ? node30471 : node30352;
									assign node30352 = (inp[1]) ? node30410 : node30353;
										assign node30353 = (inp[13]) ? node30381 : node30354;
											assign node30354 = (inp[12]) ? node30366 : node30355;
												assign node30355 = (inp[5]) ? node30361 : node30356;
													assign node30356 = (inp[9]) ? 16'b0000000011111111 : node30357;
														assign node30357 = (inp[11]) ? 16'b0000000011111111 : 16'b0000000111111111;
													assign node30361 = (inp[9]) ? node30363 : 16'b0000000011111111;
														assign node30363 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000000111111;
												assign node30366 = (inp[7]) ? node30374 : node30367;
													assign node30367 = (inp[5]) ? node30371 : node30368;
														assign node30368 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30371 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30374 = (inp[9]) ? node30378 : node30375;
														assign node30375 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30378 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30381 = (inp[12]) ? node30397 : node30382;
												assign node30382 = (inp[9]) ? node30390 : node30383;
													assign node30383 = (inp[2]) ? node30387 : node30384;
														assign node30384 = (inp[7]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node30387 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30390 = (inp[2]) ? node30394 : node30391;
														assign node30391 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30394 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30397 = (inp[2]) ? node30405 : node30398;
													assign node30398 = (inp[5]) ? node30402 : node30399;
														assign node30399 = (inp[11]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30402 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30405 = (inp[7]) ? node30407 : 16'b0000000000011111;
														assign node30407 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node30410 = (inp[2]) ? node30442 : node30411;
											assign node30411 = (inp[11]) ? node30427 : node30412;
												assign node30412 = (inp[5]) ? node30420 : node30413;
													assign node30413 = (inp[9]) ? node30417 : node30414;
														assign node30414 = (inp[12]) ? 16'b0000000001111111 : 16'b0000000111111111;
														assign node30417 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30420 = (inp[12]) ? node30424 : node30421;
														assign node30421 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30424 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30427 = (inp[9]) ? node30435 : node30428;
													assign node30428 = (inp[13]) ? node30432 : node30429;
														assign node30429 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node30432 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30435 = (inp[12]) ? node30439 : node30436;
														assign node30436 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30439 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node30442 = (inp[9]) ? node30458 : node30443;
												assign node30443 = (inp[11]) ? node30451 : node30444;
													assign node30444 = (inp[13]) ? node30448 : node30445;
														assign node30445 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node30448 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30451 = (inp[12]) ? node30455 : node30452;
														assign node30452 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30455 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30458 = (inp[12]) ? node30464 : node30459;
													assign node30459 = (inp[13]) ? node30461 : 16'b0000000000111111;
														assign node30461 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30464 = (inp[7]) ? node30468 : node30465;
														assign node30465 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30468 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
									assign node30471 = (inp[11]) ? node30527 : node30472;
										assign node30472 = (inp[12]) ? node30496 : node30473;
											assign node30473 = (inp[5]) ? node30483 : node30474;
												assign node30474 = (inp[1]) ? node30476 : 16'b0000000001111111;
													assign node30476 = (inp[13]) ? node30480 : node30477;
														assign node30477 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30480 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30483 = (inp[9]) ? node30489 : node30484;
													assign node30484 = (inp[1]) ? node30486 : 16'b0000000001111111;
														assign node30486 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30489 = (inp[2]) ? node30493 : node30490;
														assign node30490 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30493 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node30496 = (inp[2]) ? node30512 : node30497;
												assign node30497 = (inp[7]) ? node30505 : node30498;
													assign node30498 = (inp[1]) ? node30502 : node30499;
														assign node30499 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node30502 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node30505 = (inp[13]) ? node30509 : node30506;
														assign node30506 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node30509 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30512 = (inp[5]) ? node30520 : node30513;
													assign node30513 = (inp[13]) ? node30517 : node30514;
														assign node30514 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30517 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000011111;
													assign node30520 = (inp[1]) ? node30524 : node30521;
														assign node30521 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30524 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node30527 = (inp[9]) ? node30557 : node30528;
											assign node30528 = (inp[12]) ? node30542 : node30529;
												assign node30529 = (inp[1]) ? node30535 : node30530;
													assign node30530 = (inp[5]) ? node30532 : 16'b0000000001111111;
														assign node30532 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000111111;
													assign node30535 = (inp[2]) ? node30539 : node30536;
														assign node30536 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30539 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30542 = (inp[7]) ? node30550 : node30543;
													assign node30543 = (inp[13]) ? node30547 : node30544;
														assign node30544 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30547 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30550 = (inp[2]) ? node30554 : node30551;
														assign node30551 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30554 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000011111;
											assign node30557 = (inp[12]) ? node30573 : node30558;
												assign node30558 = (inp[7]) ? node30566 : node30559;
													assign node30559 = (inp[5]) ? node30563 : node30560;
														assign node30560 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30563 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30566 = (inp[5]) ? node30570 : node30567;
														assign node30567 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30570 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node30573 = (inp[2]) ? node30579 : node30574;
													assign node30574 = (inp[13]) ? node30576 : 16'b0000000000011111;
														assign node30576 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node30579 = (inp[5]) ? node30583 : node30580;
														assign node30580 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node30583 = (inp[1]) ? 16'b0000000000000011 : 16'b0000000000000111;
							assign node30586 = (inp[14]) ? node30820 : node30587;
								assign node30587 = (inp[12]) ? node30709 : node30588;
									assign node30588 = (inp[9]) ? node30646 : node30589;
										assign node30589 = (inp[11]) ? node30615 : node30590;
											assign node30590 = (inp[5]) ? node30600 : node30591;
												assign node30591 = (inp[2]) ? node30593 : 16'b0000000011111111;
													assign node30593 = (inp[7]) ? node30597 : node30594;
														assign node30594 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30597 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000011111111;
												assign node30600 = (inp[7]) ? node30608 : node30601;
													assign node30601 = (inp[2]) ? node30605 : node30602;
														assign node30602 = (inp[0]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30605 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30608 = (inp[2]) ? node30612 : node30609;
														assign node30609 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30612 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30615 = (inp[13]) ? node30631 : node30616;
												assign node30616 = (inp[1]) ? node30624 : node30617;
													assign node30617 = (inp[5]) ? node30621 : node30618;
														assign node30618 = (inp[0]) ? 16'b0000000000111111 : 16'b0000000011111111;
														assign node30621 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30624 = (inp[2]) ? node30628 : node30625;
														assign node30625 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30628 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000011111;
												assign node30631 = (inp[0]) ? node30639 : node30632;
													assign node30632 = (inp[1]) ? node30636 : node30633;
														assign node30633 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30636 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000011111;
													assign node30639 = (inp[5]) ? node30643 : node30640;
														assign node30640 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30643 = (inp[7]) ? 16'b0000000000000111 : 16'b0000000000011111;
										assign node30646 = (inp[5]) ? node30678 : node30647;
											assign node30647 = (inp[7]) ? node30663 : node30648;
												assign node30648 = (inp[0]) ? node30656 : node30649;
													assign node30649 = (inp[11]) ? node30653 : node30650;
														assign node30650 = (inp[2]) ? 16'b0000000001111111 : 16'b0000000011111111;
														assign node30653 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
													assign node30656 = (inp[1]) ? node30660 : node30657;
														assign node30657 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30660 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30663 = (inp[2]) ? node30671 : node30664;
													assign node30664 = (inp[1]) ? node30668 : node30665;
														assign node30665 = (inp[13]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30668 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30671 = (inp[1]) ? node30675 : node30672;
														assign node30672 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node30675 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node30678 = (inp[1]) ? node30694 : node30679;
												assign node30679 = (inp[11]) ? node30687 : node30680;
													assign node30680 = (inp[13]) ? node30684 : node30681;
														assign node30681 = (inp[7]) ? 16'b0000000000111111 : 16'b0000000000111111;
														assign node30684 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30687 = (inp[13]) ? node30691 : node30688;
														assign node30688 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node30691 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000001111;
												assign node30694 = (inp[0]) ? node30702 : node30695;
													assign node30695 = (inp[11]) ? node30699 : node30696;
														assign node30696 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30699 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30702 = (inp[7]) ? node30706 : node30703;
														assign node30703 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000001111;
														assign node30706 = (inp[2]) ? 16'b0000000000000011 : 16'b0000000000001111;
									assign node30709 = (inp[11]) ? node30765 : node30710;
										assign node30710 = (inp[1]) ? node30742 : node30711;
											assign node30711 = (inp[9]) ? node30727 : node30712;
												assign node30712 = (inp[13]) ? node30720 : node30713;
													assign node30713 = (inp[7]) ? node30717 : node30714;
														assign node30714 = (inp[5]) ? 16'b0000000001111111 : 16'b0000000001111111;
														assign node30717 = (inp[2]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node30720 = (inp[0]) ? node30724 : node30721;
														assign node30721 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30724 = (inp[7]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30727 = (inp[7]) ? node30735 : node30728;
													assign node30728 = (inp[13]) ? node30732 : node30729;
														assign node30729 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30732 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30735 = (inp[13]) ? node30739 : node30736;
														assign node30736 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node30739 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
											assign node30742 = (inp[0]) ? node30756 : node30743;
												assign node30743 = (inp[2]) ? node30751 : node30744;
													assign node30744 = (inp[7]) ? node30748 : node30745;
														assign node30745 = (inp[9]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node30748 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30751 = (inp[13]) ? node30753 : 16'b0000000000011111;
														assign node30753 = (inp[7]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30756 = (inp[5]) ? node30758 : 16'b0000000000011111;
													assign node30758 = (inp[9]) ? node30762 : node30759;
														assign node30759 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30762 = (inp[2]) ? 16'b0000000000000111 : 16'b0000000000001111;
										assign node30765 = (inp[13]) ? node30793 : node30766;
											assign node30766 = (inp[9]) ? node30778 : node30767;
												assign node30767 = (inp[5]) ? node30773 : node30768;
													assign node30768 = (inp[0]) ? node30770 : 16'b0000000001111111;
														assign node30770 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30773 = (inp[2]) ? 16'b0000000000011111 : node30774;
														assign node30774 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30778 = (inp[2]) ? node30786 : node30779;
													assign node30779 = (inp[7]) ? node30783 : node30780;
														assign node30780 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node30783 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30786 = (inp[5]) ? node30790 : node30787;
														assign node30787 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30790 = (inp[1]) ? 16'b0000000000000011 : 16'b0000000000001111;
											assign node30793 = (inp[7]) ? node30809 : node30794;
												assign node30794 = (inp[9]) ? node30802 : node30795;
													assign node30795 = (inp[5]) ? node30799 : node30796;
														assign node30796 = (inp[2]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30799 = (inp[2]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30802 = (inp[2]) ? node30806 : node30803;
														assign node30803 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30806 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node30809 = (inp[1]) ? node30815 : node30810;
													assign node30810 = (inp[5]) ? node30812 : 16'b0000000000011111;
														assign node30812 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node30815 = (inp[0]) ? node30817 : 16'b0000000000000111;
														assign node30817 = (inp[9]) ? 16'b0000000000000011 : 16'b0000000000000111;
								assign node30820 = (inp[2]) ? node30938 : node30821;
									assign node30821 = (inp[7]) ? node30877 : node30822;
										assign node30822 = (inp[12]) ? node30848 : node30823;
											assign node30823 = (inp[0]) ? node30835 : node30824;
												assign node30824 = (inp[9]) ? node30828 : node30825;
													assign node30825 = (inp[1]) ? 16'b0000000001111111 : 16'b0000000011111111;
													assign node30828 = (inp[11]) ? node30832 : node30829;
														assign node30829 = (inp[5]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30832 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
												assign node30835 = (inp[1]) ? node30843 : node30836;
													assign node30836 = (inp[11]) ? node30840 : node30837;
														assign node30837 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30840 = (inp[9]) ? 16'b0000000000111111 : 16'b0000000000111111;
													assign node30843 = (inp[9]) ? 16'b0000000000011111 : node30844;
														assign node30844 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
											assign node30848 = (inp[11]) ? node30864 : node30849;
												assign node30849 = (inp[9]) ? node30857 : node30850;
													assign node30850 = (inp[5]) ? node30854 : node30851;
														assign node30851 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node30854 = (inp[13]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30857 = (inp[1]) ? node30861 : node30858;
														assign node30858 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000001111111;
														assign node30861 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30864 = (inp[5]) ? node30872 : node30865;
													assign node30865 = (inp[13]) ? node30869 : node30866;
														assign node30866 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node30869 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30872 = (inp[0]) ? 16'b0000000000001111 : node30873;
														assign node30873 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
										assign node30877 = (inp[9]) ? node30907 : node30878;
											assign node30878 = (inp[13]) ? node30894 : node30879;
												assign node30879 = (inp[11]) ? node30887 : node30880;
													assign node30880 = (inp[0]) ? node30884 : node30881;
														assign node30881 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30884 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30887 = (inp[1]) ? node30891 : node30888;
														assign node30888 = (inp[12]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30891 = (inp[5]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30894 = (inp[12]) ? node30900 : node30895;
													assign node30895 = (inp[1]) ? 16'b0000000000011111 : node30896;
														assign node30896 = (inp[0]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30900 = (inp[11]) ? node30904 : node30901;
														assign node30901 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30904 = (inp[0]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node30907 = (inp[0]) ? node30923 : node30908;
												assign node30908 = (inp[11]) ? node30916 : node30909;
													assign node30909 = (inp[12]) ? node30913 : node30910;
														assign node30910 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000011111;
														assign node30913 = (inp[13]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30916 = (inp[1]) ? node30920 : node30917;
														assign node30917 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30920 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node30923 = (inp[13]) ? node30931 : node30924;
													assign node30924 = (inp[5]) ? node30928 : node30925;
														assign node30925 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30928 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node30931 = (inp[1]) ? node30935 : node30932;
														assign node30932 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node30935 = (inp[11]) ? 16'b0000000000000011 : 16'b0000000000000111;
									assign node30938 = (inp[13]) ? node30998 : node30939;
										assign node30939 = (inp[11]) ? node30969 : node30940;
											assign node30940 = (inp[0]) ? node30954 : node30941;
												assign node30941 = (inp[5]) ? node30949 : node30942;
													assign node30942 = (inp[9]) ? node30946 : node30943;
														assign node30943 = (inp[12]) ? 16'b0000000000111111 : 16'b0000000001111111;
														assign node30946 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
													assign node30949 = (inp[7]) ? node30951 : 16'b0000000000111111;
														assign node30951 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
												assign node30954 = (inp[7]) ? node30962 : node30955;
													assign node30955 = (inp[12]) ? node30959 : node30956;
														assign node30956 = (inp[5]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30959 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000011111;
													assign node30962 = (inp[1]) ? node30966 : node30963;
														assign node30963 = (inp[12]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30966 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000001111;
											assign node30969 = (inp[9]) ? node30983 : node30970;
												assign node30970 = (inp[7]) ? node30978 : node30971;
													assign node30971 = (inp[12]) ? node30975 : node30972;
														assign node30972 = (inp[1]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node30975 = (inp[1]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node30978 = (inp[0]) ? node30980 : 16'b0000000000011111;
														assign node30980 = (inp[12]) ? 16'b0000000000000011 : 16'b0000000000001111;
												assign node30983 = (inp[5]) ? node30991 : node30984;
													assign node30984 = (inp[12]) ? node30988 : node30985;
														assign node30985 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node30988 = (inp[1]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node30991 = (inp[1]) ? node30995 : node30992;
														assign node30992 = (inp[12]) ? 16'b0000000000000111 : 16'b0000000000000111;
														assign node30995 = (inp[7]) ? 16'b0000000000000011 : 16'b0000000000000111;
										assign node30998 = (inp[7]) ? node31030 : node30999;
											assign node30999 = (inp[1]) ? node31015 : node31000;
												assign node31000 = (inp[5]) ? node31008 : node31001;
													assign node31001 = (inp[12]) ? node31005 : node31002;
														assign node31002 = (inp[11]) ? 16'b0000000000011111 : 16'b0000000000111111;
														assign node31005 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
													assign node31008 = (inp[9]) ? node31012 : node31009;
														assign node31009 = (inp[0]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node31012 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
												assign node31015 = (inp[0]) ? node31023 : node31016;
													assign node31016 = (inp[12]) ? node31020 : node31017;
														assign node31017 = (inp[9]) ? 16'b0000000000001111 : 16'b0000000000011111;
														assign node31020 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node31023 = (inp[9]) ? node31027 : node31024;
														assign node31024 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node31027 = (inp[11]) ? 16'b0000000000000011 : 16'b0000000000000111;
											assign node31030 = (inp[0]) ? node31044 : node31031;
												assign node31031 = (inp[12]) ? node31037 : node31032;
													assign node31032 = (inp[5]) ? node31034 : 16'b0000000000011111;
														assign node31034 = (inp[9]) ? 16'b0000000000000111 : 16'b0000000000001111;
													assign node31037 = (inp[1]) ? node31041 : node31038;
														assign node31038 = (inp[11]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node31041 = (inp[5]) ? 16'b0000000000000011 : 16'b0000000000000111;
												assign node31044 = (inp[9]) ? node31052 : node31045;
													assign node31045 = (inp[12]) ? node31049 : node31046;
														assign node31046 = (inp[5]) ? 16'b0000000000000111 : 16'b0000000000001111;
														assign node31049 = (inp[11]) ? 16'b0000000000000011 : 16'b0000000000000111;
													assign node31052 = (inp[11]) ? node31056 : node31053;
														assign node31053 = (inp[12]) ? 16'b0000000000000011 : 16'b0000000000000111;
														assign node31056 = (inp[12]) ? 16'b0000000000000001 : 16'b0000000000000001;

endmodule