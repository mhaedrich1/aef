module dtc_split875_bm97 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node3;
	wire [3-1:0] node4;
	wire [3-1:0] node5;
	wire [3-1:0] node7;
	wire [3-1:0] node8;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node13;
	wire [3-1:0] node17;
	wire [3-1:0] node18;
	wire [3-1:0] node19;
	wire [3-1:0] node21;
	wire [3-1:0] node23;
	wire [3-1:0] node26;
	wire [3-1:0] node27;
	wire [3-1:0] node29;
	wire [3-1:0] node33;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node46;
	wire [3-1:0] node47;
	wire [3-1:0] node49;
	wire [3-1:0] node51;
	wire [3-1:0] node53;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node59;
	wire [3-1:0] node61;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node77;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node82;
	wire [3-1:0] node84;
	wire [3-1:0] node87;
	wire [3-1:0] node88;
	wire [3-1:0] node90;
	wire [3-1:0] node93;
	wire [3-1:0] node94;
	wire [3-1:0] node97;
	wire [3-1:0] node99;
	wire [3-1:0] node102;
	wire [3-1:0] node103;
	wire [3-1:0] node104;
	wire [3-1:0] node107;
	wire [3-1:0] node109;
	wire [3-1:0] node111;
	wire [3-1:0] node112;
	wire [3-1:0] node114;
	wire [3-1:0] node116;
	wire [3-1:0] node118;
	wire [3-1:0] node120;
	wire [3-1:0] node123;
	wire [3-1:0] node124;
	wire [3-1:0] node125;
	wire [3-1:0] node127;
	wire [3-1:0] node131;
	wire [3-1:0] node133;
	wire [3-1:0] node135;
	wire [3-1:0] node138;
	wire [3-1:0] node139;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node144;
	wire [3-1:0] node146;
	wire [3-1:0] node148;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node154;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node160;
	wire [3-1:0] node162;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node169;
	wire [3-1:0] node170;
	wire [3-1:0] node175;
	wire [3-1:0] node177;
	wire [3-1:0] node179;
	wire [3-1:0] node180;
	wire [3-1:0] node182;
	wire [3-1:0] node184;
	wire [3-1:0] node187;
	wire [3-1:0] node189;
	wire [3-1:0] node191;
	wire [3-1:0] node194;
	wire [3-1:0] node195;
	wire [3-1:0] node197;
	wire [3-1:0] node199;
	wire [3-1:0] node200;
	wire [3-1:0] node202;
	wire [3-1:0] node204;
	wire [3-1:0] node207;
	wire [3-1:0] node209;
	wire [3-1:0] node211;
	wire [3-1:0] node213;

	assign outp = (inp[9]) ? node46 : node1;
		assign node1 = (inp[3]) ? node3 : 3'b000;
			assign node3 = (inp[7]) ? 3'b000 : node4;
				assign node4 = (inp[6]) ? 3'b000 : node5;
					assign node5 = (inp[4]) ? node7 : 3'b100;
						assign node7 = (inp[11]) ? node17 : node8;
							assign node8 = (inp[8]) ? 3'b100 : node9;
								assign node9 = (inp[10]) ? node11 : 3'b100;
									assign node11 = (inp[2]) ? node13 : 3'b000;
										assign node13 = (inp[1]) ? 3'b100 : 3'b000;
							assign node17 = (inp[5]) ? node33 : node18;
								assign node18 = (inp[10]) ? node26 : node19;
									assign node19 = (inp[1]) ? node21 : 3'b100;
										assign node21 = (inp[2]) ? node23 : 3'b100;
											assign node23 = (inp[0]) ? 3'b000 : 3'b100;
									assign node26 = (inp[8]) ? 3'b000 : node27;
										assign node27 = (inp[0]) ? node29 : 3'b100;
											assign node29 = (inp[1]) ? 3'b000 : 3'b100;
								assign node33 = (inp[0]) ? 3'b000 : node34;
									assign node34 = (inp[10]) ? node40 : node35;
										assign node35 = (inp[2]) ? node37 : 3'b000;
											assign node37 = (inp[8]) ? 3'b100 : 3'b000;
										assign node40 = (inp[8]) ? 3'b000 : 3'b100;
		assign node46 = (inp[3]) ? node102 : node47;
			assign node47 = (inp[6]) ? node49 : 3'b000;
				assign node49 = (inp[7]) ? node51 : 3'b001;
					assign node51 = (inp[10]) ? node53 : 3'b000;
						assign node53 = (inp[4]) ? node77 : node54;
							assign node54 = (inp[11]) ? node56 : 3'b000;
								assign node56 = (inp[8]) ? node64 : node57;
									assign node57 = (inp[5]) ? node59 : 3'b000;
										assign node59 = (inp[0]) ? node61 : 3'b001;
											assign node61 = (inp[1]) ? 3'b101 : 3'b001;
									assign node64 = (inp[5]) ? node72 : node65;
										assign node65 = (inp[2]) ? node67 : 3'b100;
											assign node67 = (inp[1]) ? node69 : 3'b100;
												assign node69 = (inp[0]) ? 3'b101 : 3'b100;
										assign node72 = (inp[2]) ? node74 : 3'b101;
											assign node74 = (inp[0]) ? 3'b101 : 3'b100;
							assign node77 = (inp[11]) ? node79 : 3'b100;
								assign node79 = (inp[5]) ? node87 : node80;
									assign node80 = (inp[8]) ? node82 : 3'b000;
										assign node82 = (inp[2]) ? node84 : 3'b100;
											assign node84 = (inp[1]) ? 3'b110 : 3'b100;
									assign node87 = (inp[8]) ? node93 : node88;
										assign node88 = (inp[0]) ? node90 : 3'b010;
											assign node90 = (inp[1]) ? 3'b110 : 3'b010;
										assign node93 = (inp[0]) ? node97 : node94;
											assign node94 = (inp[2]) ? 3'b100 : 3'b110;
											assign node97 = (inp[2]) ? node99 : 3'b110;
												assign node99 = (inp[1]) ? 3'b010 : 3'b110;
			assign node102 = (inp[4]) ? node138 : node103;
				assign node103 = (inp[7]) ? node107 : node104;
					assign node104 = (inp[6]) ? 3'b110 : 3'b000;
					assign node107 = (inp[6]) ? node109 : 3'b110;
						assign node109 = (inp[10]) ? node111 : 3'b000;
							assign node111 = (inp[5]) ? node123 : node112;
								assign node112 = (inp[2]) ? node114 : 3'b010;
									assign node114 = (inp[8]) ? node116 : 3'b010;
										assign node116 = (inp[0]) ? node118 : 3'b010;
											assign node118 = (inp[1]) ? node120 : 3'b010;
												assign node120 = (inp[11]) ? 3'b100 : 3'b000;
								assign node123 = (inp[11]) ? node131 : node124;
									assign node124 = (inp[0]) ? 3'b000 : node125;
										assign node125 = (inp[2]) ? node127 : 3'b000;
											assign node127 = (inp[8]) ? 3'b010 : 3'b000;
									assign node131 = (inp[8]) ? node133 : 3'b100;
										assign node133 = (inp[2]) ? node135 : 3'b100;
											assign node135 = (inp[0]) ? 3'b100 : 3'b010;
				assign node138 = (inp[6]) ? node194 : node139;
					assign node139 = (inp[7]) ? node175 : node140;
						assign node140 = (inp[10]) ? node158 : node141;
							assign node141 = (inp[11]) ? node143 : 3'b010;
								assign node143 = (inp[5]) ? node151 : node144;
									assign node144 = (inp[8]) ? node146 : 3'b010;
										assign node146 = (inp[2]) ? node148 : 3'b010;
											assign node148 = (inp[1]) ? 3'b110 : 3'b010;
									assign node151 = (inp[0]) ? 3'b110 : node152;
										assign node152 = (inp[8]) ? node154 : 3'b110;
											assign node154 = (inp[2]) ? 3'b010 : 3'b110;
							assign node158 = (inp[11]) ? node166 : node159;
								assign node159 = (inp[8]) ? 3'b001 : node160;
									assign node160 = (inp[1]) ? node162 : 3'b101;
										assign node162 = (inp[2]) ? 3'b001 : 3'b101;
								assign node166 = (inp[8]) ? 3'b101 : node167;
									assign node167 = (inp[0]) ? node169 : 3'b011;
										assign node169 = (inp[1]) ? 3'b101 : node170;
											assign node170 = (inp[5]) ? 3'b101 : 3'b011;
						assign node175 = (inp[11]) ? node177 : 3'b001;
							assign node177 = (inp[10]) ? node179 : 3'b001;
								assign node179 = (inp[8]) ? node187 : node180;
									assign node180 = (inp[1]) ? node182 : 3'b001;
										assign node182 = (inp[0]) ? node184 : 3'b001;
											assign node184 = (inp[5]) ? 3'b110 : 3'b001;
									assign node187 = (inp[0]) ? node189 : 3'b110;
										assign node189 = (inp[1]) ? node191 : 3'b110;
											assign node191 = (inp[2]) ? 3'b001 : 3'b110;
					assign node194 = (inp[7]) ? 3'b000 : node195;
						assign node195 = (inp[11]) ? node197 : 3'b000;
							assign node197 = (inp[10]) ? node199 : 3'b000;
								assign node199 = (inp[8]) ? node207 : node200;
									assign node200 = (inp[1]) ? node202 : 3'b010;
										assign node202 = (inp[5]) ? node204 : 3'b010;
											assign node204 = (inp[0]) ? 3'b100 : 3'b010;
									assign node207 = (inp[1]) ? node209 : 3'b100;
										assign node209 = (inp[2]) ? node211 : 3'b100;
											assign node211 = (inp[0]) ? node213 : 3'b100;
												assign node213 = (inp[5]) ? 3'b000 : 3'b100;

endmodule