module dtc_split33_bm85 (
	input  wire [12-1:0] inp,
	output wire [3-1:0] outp
);

	wire [3-1:0] node1;
	wire [3-1:0] node2;
	wire [3-1:0] node4;
	wire [3-1:0] node6;
	wire [3-1:0] node7;
	wire [3-1:0] node9;
	wire [3-1:0] node11;
	wire [3-1:0] node12;
	wire [3-1:0] node13;
	wire [3-1:0] node14;
	wire [3-1:0] node17;
	wire [3-1:0] node22;
	wire [3-1:0] node23;
	wire [3-1:0] node24;
	wire [3-1:0] node25;
	wire [3-1:0] node28;
	wire [3-1:0] node29;
	wire [3-1:0] node34;
	wire [3-1:0] node35;
	wire [3-1:0] node36;
	wire [3-1:0] node37;
	wire [3-1:0] node40;
	wire [3-1:0] node43;
	wire [3-1:0] node45;
	wire [3-1:0] node47;
	wire [3-1:0] node48;
	wire [3-1:0] node51;
	wire [3-1:0] node54;
	wire [3-1:0] node56;
	wire [3-1:0] node57;
	wire [3-1:0] node58;
	wire [3-1:0] node64;
	wire [3-1:0] node65;
	wire [3-1:0] node66;
	wire [3-1:0] node67;
	wire [3-1:0] node69;
	wire [3-1:0] node71;
	wire [3-1:0] node72;
	wire [3-1:0] node74;
	wire [3-1:0] node78;
	wire [3-1:0] node79;
	wire [3-1:0] node80;
	wire [3-1:0] node81;
	wire [3-1:0] node83;
	wire [3-1:0] node85;
	wire [3-1:0] node86;
	wire [3-1:0] node89;
	wire [3-1:0] node90;
	wire [3-1:0] node94;
	wire [3-1:0] node95;
	wire [3-1:0] node98;
	wire [3-1:0] node99;
	wire [3-1:0] node104;
	wire [3-1:0] node105;
	wire [3-1:0] node106;
	wire [3-1:0] node107;
	wire [3-1:0] node108;
	wire [3-1:0] node109;
	wire [3-1:0] node110;
	wire [3-1:0] node117;
	wire [3-1:0] node118;
	wire [3-1:0] node119;
	wire [3-1:0] node122;
	wire [3-1:0] node125;
	wire [3-1:0] node126;
	wire [3-1:0] node127;
	wire [3-1:0] node128;
	wire [3-1:0] node134;
	wire [3-1:0] node135;
	wire [3-1:0] node136;
	wire [3-1:0] node140;
	wire [3-1:0] node141;
	wire [3-1:0] node143;
	wire [3-1:0] node146;
	wire [3-1:0] node147;
	wire [3-1:0] node151;
	wire [3-1:0] node152;
	wire [3-1:0] node153;
	wire [3-1:0] node154;
	wire [3-1:0] node155;
	wire [3-1:0] node157;
	wire [3-1:0] node158;
	wire [3-1:0] node159;
	wire [3-1:0] node163;
	wire [3-1:0] node166;
	wire [3-1:0] node167;
	wire [3-1:0] node170;
	wire [3-1:0] node171;
	wire [3-1:0] node175;
	wire [3-1:0] node176;
	wire [3-1:0] node178;
	wire [3-1:0] node179;
	wire [3-1:0] node183;
	wire [3-1:0] node184;
	wire [3-1:0] node185;
	wire [3-1:0] node187;
	wire [3-1:0] node190;
	wire [3-1:0] node192;
	wire [3-1:0] node195;
	wire [3-1:0] node198;
	wire [3-1:0] node200;
	wire [3-1:0] node201;
	wire [3-1:0] node203;
	wire [3-1:0] node204;
	wire [3-1:0] node205;
	wire [3-1:0] node208;
	wire [3-1:0] node212;
	wire [3-1:0] node213;
	wire [3-1:0] node214;
	wire [3-1:0] node219;
	wire [3-1:0] node221;
	wire [3-1:0] node222;
	wire [3-1:0] node223;
	wire [3-1:0] node225;
	wire [3-1:0] node227;
	wire [3-1:0] node230;
	wire [3-1:0] node231;
	wire [3-1:0] node232;
	wire [3-1:0] node235;
	wire [3-1:0] node236;
	wire [3-1:0] node240;
	wire [3-1:0] node241;
	wire [3-1:0] node245;
	wire [3-1:0] node246;
	wire [3-1:0] node247;
	wire [3-1:0] node250;
	wire [3-1:0] node251;
	wire [3-1:0] node255;
	wire [3-1:0] node256;
	wire [3-1:0] node259;
	wire [3-1:0] node260;
	wire [3-1:0] node262;
	wire [3-1:0] node265;
	wire [3-1:0] node268;
	wire [3-1:0] node270;
	wire [3-1:0] node272;
	wire [3-1:0] node273;
	wire [3-1:0] node274;
	wire [3-1:0] node276;
	wire [3-1:0] node278;
	wire [3-1:0] node279;
	wire [3-1:0] node280;
	wire [3-1:0] node284;
	wire [3-1:0] node285;
	wire [3-1:0] node289;
	wire [3-1:0] node290;
	wire [3-1:0] node291;
	wire [3-1:0] node294;
	wire [3-1:0] node297;
	wire [3-1:0] node298;
	wire [3-1:0] node300;
	wire [3-1:0] node303;
	wire [3-1:0] node304;
	wire [3-1:0] node308;
	wire [3-1:0] node309;
	wire [3-1:0] node311;
	wire [3-1:0] node313;
	wire [3-1:0] node315;
	wire [3-1:0] node318;
	wire [3-1:0] node320;
	wire [3-1:0] node322;
	wire [3-1:0] node323;

	assign outp = (inp[0]) ? node64 : node1;
		assign node1 = (inp[6]) ? 3'b000 : node2;
			assign node2 = (inp[3]) ? node4 : 3'b000;
				assign node4 = (inp[9]) ? node6 : 3'b000;
					assign node6 = (inp[4]) ? node22 : node7;
						assign node7 = (inp[2]) ? node9 : 3'b000;
							assign node9 = (inp[1]) ? node11 : 3'b000;
								assign node11 = (inp[7]) ? 3'b000 : node12;
									assign node12 = (inp[5]) ? 3'b100 : node13;
										assign node13 = (inp[8]) ? node17 : node14;
											assign node14 = (inp[10]) ? 3'b100 : 3'b000;
											assign node17 = (inp[10]) ? 3'b000 : 3'b100;
						assign node22 = (inp[1]) ? node34 : node23;
							assign node23 = (inp[7]) ? 3'b000 : node24;
								assign node24 = (inp[10]) ? node28 : node25;
									assign node25 = (inp[8]) ? 3'b011 : 3'b010;
									assign node28 = (inp[2]) ? 3'b000 : node29;
										assign node29 = (inp[11]) ? 3'b010 : 3'b000;
							assign node34 = (inp[7]) ? node54 : node35;
								assign node35 = (inp[5]) ? node43 : node36;
									assign node36 = (inp[11]) ? node40 : node37;
										assign node37 = (inp[2]) ? 3'b101 : 3'b110;
										assign node40 = (inp[10]) ? 3'b110 : 3'b010;
									assign node43 = (inp[2]) ? node45 : 3'b001;
										assign node45 = (inp[11]) ? node47 : 3'b101;
											assign node47 = (inp[8]) ? node51 : node48;
												assign node48 = (inp[10]) ? 3'b011 : 3'b101;
												assign node51 = (inp[10]) ? 3'b101 : 3'b001;
								assign node54 = (inp[10]) ? node56 : 3'b100;
									assign node56 = (inp[8]) ? 3'b000 : node57;
										assign node57 = (inp[11]) ? 3'b010 : node58;
											assign node58 = (inp[5]) ? 3'b010 : 3'b110;
		assign node64 = (inp[6]) ? node268 : node65;
			assign node65 = (inp[3]) ? node151 : node66;
				assign node66 = (inp[4]) ? node78 : node67;
					assign node67 = (inp[11]) ? node69 : 3'b000;
						assign node69 = (inp[5]) ? node71 : 3'b000;
							assign node71 = (inp[8]) ? 3'b000 : node72;
								assign node72 = (inp[9]) ? node74 : 3'b000;
									assign node74 = (inp[10]) ? 3'b100 : 3'b000;
					assign node78 = (inp[9]) ? node104 : node79;
						assign node79 = (inp[7]) ? 3'b100 : node80;
							assign node80 = (inp[5]) ? node94 : node81;
								assign node81 = (inp[2]) ? node83 : 3'b100;
									assign node83 = (inp[11]) ? node85 : 3'b100;
										assign node85 = (inp[1]) ? node89 : node86;
											assign node86 = (inp[8]) ? 3'b000 : 3'b100;
											assign node89 = (inp[8]) ? 3'b100 : node90;
												assign node90 = (inp[10]) ? 3'b100 : 3'b000;
								assign node94 = (inp[1]) ? node98 : node95;
									assign node95 = (inp[2]) ? 3'b100 : 3'b000;
									assign node98 = (inp[8]) ? 3'b100 : node99;
										assign node99 = (inp[10]) ? 3'b000 : 3'b100;
						assign node104 = (inp[2]) ? node134 : node105;
							assign node105 = (inp[11]) ? node117 : node106;
								assign node106 = (inp[10]) ? 3'b000 : node107;
									assign node107 = (inp[8]) ? 3'b000 : node108;
										assign node108 = (inp[7]) ? 3'b100 : node109;
											assign node109 = (inp[1]) ? 3'b000 : node110;
												assign node110 = (inp[5]) ? 3'b000 : 3'b100;
								assign node117 = (inp[8]) ? node125 : node118;
									assign node118 = (inp[10]) ? node122 : node119;
										assign node119 = (inp[1]) ? 3'b100 : 3'b000;
										assign node122 = (inp[1]) ? 3'b000 : 3'b100;
									assign node125 = (inp[1]) ? 3'b100 : node126;
										assign node126 = (inp[5]) ? 3'b000 : node127;
											assign node127 = (inp[10]) ? 3'b100 : node128;
												assign node128 = (inp[7]) ? 3'b000 : 3'b100;
							assign node134 = (inp[1]) ? node140 : node135;
								assign node135 = (inp[5]) ? 3'b100 : node136;
									assign node136 = (inp[7]) ? 3'b000 : 3'b100;
								assign node140 = (inp[7]) ? node146 : node141;
									assign node141 = (inp[10]) ? node143 : 3'b110;
										assign node143 = (inp[5]) ? 3'b001 : 3'b010;
									assign node146 = (inp[10]) ? 3'b100 : node147;
										assign node147 = (inp[8]) ? 3'b000 : 3'b100;
				assign node151 = (inp[7]) ? node219 : node152;
					assign node152 = (inp[4]) ? node198 : node153;
						assign node153 = (inp[9]) ? node175 : node154;
							assign node154 = (inp[5]) ? node166 : node155;
								assign node155 = (inp[11]) ? node157 : 3'b001;
									assign node157 = (inp[2]) ? node163 : node158;
										assign node158 = (inp[10]) ? 3'b101 : node159;
											assign node159 = (inp[8]) ? 3'b001 : 3'b101;
										assign node163 = (inp[1]) ? 3'b101 : 3'b001;
								assign node166 = (inp[2]) ? node170 : node167;
									assign node167 = (inp[1]) ? 3'b101 : 3'b001;
									assign node170 = (inp[8]) ? 3'b101 : node171;
										assign node171 = (inp[10]) ? 3'b101 : 3'b001;
							assign node175 = (inp[1]) ? node183 : node176;
								assign node176 = (inp[5]) ? node178 : 3'b010;
									assign node178 = (inp[11]) ? 3'b001 : node179;
										assign node179 = (inp[2]) ? 3'b010 : 3'b110;
								assign node183 = (inp[10]) ? node195 : node184;
									assign node184 = (inp[5]) ? node190 : node185;
										assign node185 = (inp[2]) ? node187 : 3'b011;
											assign node187 = (inp[8]) ? 3'b001 : 3'b101;
										assign node190 = (inp[2]) ? node192 : 3'b101;
											assign node192 = (inp[8]) ? 3'b111 : 3'b011;
									assign node195 = (inp[2]) ? 3'b111 : 3'b101;
						assign node198 = (inp[9]) ? node200 : 3'b111;
							assign node200 = (inp[2]) ? node212 : node201;
								assign node201 = (inp[5]) ? node203 : 3'b001;
									assign node203 = (inp[1]) ? 3'b111 : node204;
										assign node204 = (inp[10]) ? node208 : node205;
											assign node205 = (inp[11]) ? 3'b011 : 3'b101;
											assign node208 = (inp[11]) ? 3'b111 : 3'b011;
								assign node212 = (inp[1]) ? 3'b111 : node213;
									assign node213 = (inp[5]) ? 3'b111 : node214;
										assign node214 = (inp[10]) ? 3'b111 : 3'b101;
					assign node219 = (inp[9]) ? node221 : 3'b001;
						assign node221 = (inp[8]) ? node245 : node222;
							assign node222 = (inp[4]) ? node230 : node223;
								assign node223 = (inp[10]) ? node225 : 3'b010;
									assign node225 = (inp[1]) ? node227 : 3'b110;
										assign node227 = (inp[2]) ? 3'b110 : 3'b101;
								assign node230 = (inp[1]) ? node240 : node231;
									assign node231 = (inp[5]) ? node235 : node232;
										assign node232 = (inp[2]) ? 3'b001 : 3'b100;
										assign node235 = (inp[10]) ? 3'b101 : node236;
											assign node236 = (inp[2]) ? 3'b101 : 3'b001;
									assign node240 = (inp[2]) ? 3'b111 : node241;
										assign node241 = (inp[5]) ? 3'b011 : 3'b001;
							assign node245 = (inp[10]) ? node255 : node246;
								assign node246 = (inp[4]) ? node250 : node247;
									assign node247 = (inp[2]) ? 3'b110 : 3'b101;
									assign node250 = (inp[2]) ? 3'b001 : node251;
										assign node251 = (inp[1]) ? 3'b001 : 3'b100;
								assign node255 = (inp[4]) ? node259 : node256;
									assign node256 = (inp[1]) ? 3'b010 : 3'b001;
									assign node259 = (inp[2]) ? node265 : node260;
										assign node260 = (inp[11]) ? node262 : 3'b101;
											assign node262 = (inp[5]) ? 3'b011 : 3'b001;
										assign node265 = (inp[11]) ? 3'b111 : 3'b011;
			assign node268 = (inp[9]) ? node270 : 3'b000;
				assign node270 = (inp[3]) ? node272 : 3'b000;
					assign node272 = (inp[7]) ? node308 : node273;
						assign node273 = (inp[4]) ? node289 : node274;
							assign node274 = (inp[1]) ? node276 : 3'b000;
								assign node276 = (inp[2]) ? node278 : 3'b000;
									assign node278 = (inp[11]) ? node284 : node279;
										assign node279 = (inp[10]) ? 3'b100 : node280;
											assign node280 = (inp[5]) ? 3'b000 : 3'b100;
										assign node284 = (inp[8]) ? 3'b100 : node285;
											assign node285 = (inp[10]) ? 3'b110 : 3'b010;
							assign node289 = (inp[1]) ? node297 : node290;
								assign node290 = (inp[8]) ? node294 : node291;
									assign node291 = (inp[10]) ? 3'b110 : 3'b100;
									assign node294 = (inp[10]) ? 3'b010 : 3'b000;
								assign node297 = (inp[10]) ? node303 : node298;
									assign node298 = (inp[8]) ? node300 : 3'b110;
										assign node300 = (inp[2]) ? 3'b110 : 3'b010;
									assign node303 = (inp[2]) ? 3'b111 : node304;
										assign node304 = (inp[8]) ? 3'b101 : 3'b001;
						assign node308 = (inp[10]) ? node318 : node309;
							assign node309 = (inp[1]) ? node311 : 3'b000;
								assign node311 = (inp[5]) ? node313 : 3'b000;
									assign node313 = (inp[8]) ? node315 : 3'b000;
										assign node315 = (inp[2]) ? 3'b100 : 3'b000;
							assign node318 = (inp[2]) ? node320 : 3'b000;
								assign node320 = (inp[4]) ? node322 : 3'b000;
									assign node322 = (inp[8]) ? 3'b010 : node323;
										assign node323 = (inp[5]) ? 3'b110 : 3'b010;

endmodule