module dtc_split33_bm23 (
	input  wire [12-1:0] inp,
	output wire [12-1:0] outp
);

	wire [12-1:0] node1;
	wire [12-1:0] node2;
	wire [12-1:0] node3;
	wire [12-1:0] node4;
	wire [12-1:0] node5;
	wire [12-1:0] node6;
	wire [12-1:0] node7;
	wire [12-1:0] node8;
	wire [12-1:0] node9;
	wire [12-1:0] node12;
	wire [12-1:0] node15;
	wire [12-1:0] node16;
	wire [12-1:0] node19;
	wire [12-1:0] node22;
	wire [12-1:0] node23;
	wire [12-1:0] node24;
	wire [12-1:0] node28;
	wire [12-1:0] node29;
	wire [12-1:0] node32;
	wire [12-1:0] node35;
	wire [12-1:0] node36;
	wire [12-1:0] node37;
	wire [12-1:0] node39;
	wire [12-1:0] node42;
	wire [12-1:0] node43;
	wire [12-1:0] node46;
	wire [12-1:0] node49;
	wire [12-1:0] node50;
	wire [12-1:0] node51;
	wire [12-1:0] node54;
	wire [12-1:0] node57;
	wire [12-1:0] node58;
	wire [12-1:0] node61;
	wire [12-1:0] node64;
	wire [12-1:0] node65;
	wire [12-1:0] node66;
	wire [12-1:0] node67;
	wire [12-1:0] node69;
	wire [12-1:0] node72;
	wire [12-1:0] node74;
	wire [12-1:0] node77;
	wire [12-1:0] node78;
	wire [12-1:0] node80;
	wire [12-1:0] node83;
	wire [12-1:0] node84;
	wire [12-1:0] node88;
	wire [12-1:0] node89;
	wire [12-1:0] node90;
	wire [12-1:0] node93;
	wire [12-1:0] node94;
	wire [12-1:0] node98;
	wire [12-1:0] node99;
	wire [12-1:0] node100;
	wire [12-1:0] node104;
	wire [12-1:0] node107;
	wire [12-1:0] node108;
	wire [12-1:0] node109;
	wire [12-1:0] node110;
	wire [12-1:0] node111;
	wire [12-1:0] node112;
	wire [12-1:0] node115;
	wire [12-1:0] node118;
	wire [12-1:0] node119;
	wire [12-1:0] node122;
	wire [12-1:0] node125;
	wire [12-1:0] node126;
	wire [12-1:0] node127;
	wire [12-1:0] node130;
	wire [12-1:0] node133;
	wire [12-1:0] node135;
	wire [12-1:0] node138;
	wire [12-1:0] node139;
	wire [12-1:0] node140;
	wire [12-1:0] node142;
	wire [12-1:0] node145;
	wire [12-1:0] node147;
	wire [12-1:0] node150;
	wire [12-1:0] node152;
	wire [12-1:0] node153;
	wire [12-1:0] node157;
	wire [12-1:0] node158;
	wire [12-1:0] node159;
	wire [12-1:0] node160;
	wire [12-1:0] node163;
	wire [12-1:0] node164;
	wire [12-1:0] node167;
	wire [12-1:0] node170;
	wire [12-1:0] node171;
	wire [12-1:0] node172;
	wire [12-1:0] node175;
	wire [12-1:0] node179;
	wire [12-1:0] node180;
	wire [12-1:0] node181;
	wire [12-1:0] node184;
	wire [12-1:0] node185;
	wire [12-1:0] node188;
	wire [12-1:0] node191;
	wire [12-1:0] node192;
	wire [12-1:0] node193;
	wire [12-1:0] node196;
	wire [12-1:0] node199;
	wire [12-1:0] node200;
	wire [12-1:0] node204;
	wire [12-1:0] node205;
	wire [12-1:0] node206;
	wire [12-1:0] node207;
	wire [12-1:0] node208;
	wire [12-1:0] node209;
	wire [12-1:0] node210;
	wire [12-1:0] node213;
	wire [12-1:0] node216;
	wire [12-1:0] node217;
	wire [12-1:0] node221;
	wire [12-1:0] node222;
	wire [12-1:0] node223;
	wire [12-1:0] node226;
	wire [12-1:0] node229;
	wire [12-1:0] node230;
	wire [12-1:0] node234;
	wire [12-1:0] node235;
	wire [12-1:0] node236;
	wire [12-1:0] node238;
	wire [12-1:0] node241;
	wire [12-1:0] node242;
	wire [12-1:0] node246;
	wire [12-1:0] node247;
	wire [12-1:0] node248;
	wire [12-1:0] node252;
	wire [12-1:0] node253;
	wire [12-1:0] node256;
	wire [12-1:0] node259;
	wire [12-1:0] node260;
	wire [12-1:0] node261;
	wire [12-1:0] node262;
	wire [12-1:0] node263;
	wire [12-1:0] node266;
	wire [12-1:0] node269;
	wire [12-1:0] node271;
	wire [12-1:0] node274;
	wire [12-1:0] node275;
	wire [12-1:0] node277;
	wire [12-1:0] node280;
	wire [12-1:0] node282;
	wire [12-1:0] node285;
	wire [12-1:0] node286;
	wire [12-1:0] node287;
	wire [12-1:0] node289;
	wire [12-1:0] node292;
	wire [12-1:0] node293;
	wire [12-1:0] node296;
	wire [12-1:0] node299;
	wire [12-1:0] node300;
	wire [12-1:0] node301;
	wire [12-1:0] node305;
	wire [12-1:0] node306;
	wire [12-1:0] node310;
	wire [12-1:0] node311;
	wire [12-1:0] node312;
	wire [12-1:0] node313;
	wire [12-1:0] node314;
	wire [12-1:0] node315;
	wire [12-1:0] node318;
	wire [12-1:0] node321;
	wire [12-1:0] node322;
	wire [12-1:0] node326;
	wire [12-1:0] node327;
	wire [12-1:0] node328;
	wire [12-1:0] node332;
	wire [12-1:0] node334;
	wire [12-1:0] node337;
	wire [12-1:0] node338;
	wire [12-1:0] node339;
	wire [12-1:0] node340;
	wire [12-1:0] node343;
	wire [12-1:0] node346;
	wire [12-1:0] node348;
	wire [12-1:0] node351;
	wire [12-1:0] node352;
	wire [12-1:0] node355;
	wire [12-1:0] node357;
	wire [12-1:0] node360;
	wire [12-1:0] node361;
	wire [12-1:0] node362;
	wire [12-1:0] node363;
	wire [12-1:0] node364;
	wire [12-1:0] node369;
	wire [12-1:0] node370;
	wire [12-1:0] node371;
	wire [12-1:0] node374;
	wire [12-1:0] node377;
	wire [12-1:0] node378;
	wire [12-1:0] node381;
	wire [12-1:0] node384;
	wire [12-1:0] node385;
	wire [12-1:0] node386;
	wire [12-1:0] node387;
	wire [12-1:0] node390;
	wire [12-1:0] node393;
	wire [12-1:0] node394;
	wire [12-1:0] node397;
	wire [12-1:0] node400;
	wire [12-1:0] node401;
	wire [12-1:0] node402;
	wire [12-1:0] node406;
	wire [12-1:0] node408;
	wire [12-1:0] node411;
	wire [12-1:0] node412;
	wire [12-1:0] node413;
	wire [12-1:0] node414;
	wire [12-1:0] node415;
	wire [12-1:0] node416;
	wire [12-1:0] node417;
	wire [12-1:0] node418;
	wire [12-1:0] node421;
	wire [12-1:0] node424;
	wire [12-1:0] node425;
	wire [12-1:0] node429;
	wire [12-1:0] node430;
	wire [12-1:0] node432;
	wire [12-1:0] node435;
	wire [12-1:0] node436;
	wire [12-1:0] node440;
	wire [12-1:0] node441;
	wire [12-1:0] node442;
	wire [12-1:0] node443;
	wire [12-1:0] node446;
	wire [12-1:0] node449;
	wire [12-1:0] node451;
	wire [12-1:0] node454;
	wire [12-1:0] node455;
	wire [12-1:0] node456;
	wire [12-1:0] node460;
	wire [12-1:0] node461;
	wire [12-1:0] node464;
	wire [12-1:0] node467;
	wire [12-1:0] node468;
	wire [12-1:0] node469;
	wire [12-1:0] node472;
	wire [12-1:0] node473;
	wire [12-1:0] node474;
	wire [12-1:0] node477;
	wire [12-1:0] node480;
	wire [12-1:0] node482;
	wire [12-1:0] node485;
	wire [12-1:0] node486;
	wire [12-1:0] node487;
	wire [12-1:0] node488;
	wire [12-1:0] node491;
	wire [12-1:0] node494;
	wire [12-1:0] node495;
	wire [12-1:0] node498;
	wire [12-1:0] node501;
	wire [12-1:0] node502;
	wire [12-1:0] node503;
	wire [12-1:0] node506;
	wire [12-1:0] node509;
	wire [12-1:0] node511;
	wire [12-1:0] node514;
	wire [12-1:0] node515;
	wire [12-1:0] node516;
	wire [12-1:0] node517;
	wire [12-1:0] node518;
	wire [12-1:0] node519;
	wire [12-1:0] node523;
	wire [12-1:0] node524;
	wire [12-1:0] node527;
	wire [12-1:0] node530;
	wire [12-1:0] node531;
	wire [12-1:0] node532;
	wire [12-1:0] node535;
	wire [12-1:0] node538;
	wire [12-1:0] node540;
	wire [12-1:0] node543;
	wire [12-1:0] node544;
	wire [12-1:0] node545;
	wire [12-1:0] node547;
	wire [12-1:0] node550;
	wire [12-1:0] node551;
	wire [12-1:0] node554;
	wire [12-1:0] node557;
	wire [12-1:0] node558;
	wire [12-1:0] node559;
	wire [12-1:0] node562;
	wire [12-1:0] node565;
	wire [12-1:0] node567;
	wire [12-1:0] node570;
	wire [12-1:0] node571;
	wire [12-1:0] node572;
	wire [12-1:0] node573;
	wire [12-1:0] node574;
	wire [12-1:0] node577;
	wire [12-1:0] node580;
	wire [12-1:0] node581;
	wire [12-1:0] node585;
	wire [12-1:0] node586;
	wire [12-1:0] node587;
	wire [12-1:0] node591;
	wire [12-1:0] node593;
	wire [12-1:0] node596;
	wire [12-1:0] node597;
	wire [12-1:0] node598;
	wire [12-1:0] node599;
	wire [12-1:0] node602;
	wire [12-1:0] node606;
	wire [12-1:0] node607;
	wire [12-1:0] node609;
	wire [12-1:0] node612;
	wire [12-1:0] node613;
	wire [12-1:0] node617;
	wire [12-1:0] node618;
	wire [12-1:0] node619;
	wire [12-1:0] node620;
	wire [12-1:0] node621;
	wire [12-1:0] node622;
	wire [12-1:0] node623;
	wire [12-1:0] node627;
	wire [12-1:0] node629;
	wire [12-1:0] node632;
	wire [12-1:0] node633;
	wire [12-1:0] node634;
	wire [12-1:0] node637;
	wire [12-1:0] node640;
	wire [12-1:0] node641;
	wire [12-1:0] node644;
	wire [12-1:0] node647;
	wire [12-1:0] node648;
	wire [12-1:0] node649;
	wire [12-1:0] node651;
	wire [12-1:0] node654;
	wire [12-1:0] node657;
	wire [12-1:0] node658;
	wire [12-1:0] node659;
	wire [12-1:0] node662;
	wire [12-1:0] node665;
	wire [12-1:0] node666;
	wire [12-1:0] node669;
	wire [12-1:0] node672;
	wire [12-1:0] node673;
	wire [12-1:0] node674;
	wire [12-1:0] node675;
	wire [12-1:0] node676;
	wire [12-1:0] node679;
	wire [12-1:0] node682;
	wire [12-1:0] node683;
	wire [12-1:0] node686;
	wire [12-1:0] node689;
	wire [12-1:0] node690;
	wire [12-1:0] node691;
	wire [12-1:0] node694;
	wire [12-1:0] node697;
	wire [12-1:0] node698;
	wire [12-1:0] node702;
	wire [12-1:0] node703;
	wire [12-1:0] node704;
	wire [12-1:0] node705;
	wire [12-1:0] node708;
	wire [12-1:0] node711;
	wire [12-1:0] node712;
	wire [12-1:0] node715;
	wire [12-1:0] node718;
	wire [12-1:0] node719;
	wire [12-1:0] node720;
	wire [12-1:0] node723;
	wire [12-1:0] node726;
	wire [12-1:0] node728;
	wire [12-1:0] node731;
	wire [12-1:0] node732;
	wire [12-1:0] node733;
	wire [12-1:0] node734;
	wire [12-1:0] node735;
	wire [12-1:0] node736;
	wire [12-1:0] node739;
	wire [12-1:0] node742;
	wire [12-1:0] node743;
	wire [12-1:0] node747;
	wire [12-1:0] node748;
	wire [12-1:0] node749;
	wire [12-1:0] node752;
	wire [12-1:0] node755;
	wire [12-1:0] node756;
	wire [12-1:0] node759;
	wire [12-1:0] node762;
	wire [12-1:0] node763;
	wire [12-1:0] node764;
	wire [12-1:0] node765;
	wire [12-1:0] node768;
	wire [12-1:0] node771;
	wire [12-1:0] node772;
	wire [12-1:0] node775;
	wire [12-1:0] node778;
	wire [12-1:0] node779;
	wire [12-1:0] node780;
	wire [12-1:0] node784;
	wire [12-1:0] node785;
	wire [12-1:0] node788;
	wire [12-1:0] node791;
	wire [12-1:0] node792;
	wire [12-1:0] node793;
	wire [12-1:0] node794;
	wire [12-1:0] node796;
	wire [12-1:0] node799;
	wire [12-1:0] node802;
	wire [12-1:0] node803;
	wire [12-1:0] node805;
	wire [12-1:0] node808;
	wire [12-1:0] node809;
	wire [12-1:0] node812;
	wire [12-1:0] node815;
	wire [12-1:0] node816;
	wire [12-1:0] node817;
	wire [12-1:0] node820;
	wire [12-1:0] node821;
	wire [12-1:0] node825;
	wire [12-1:0] node826;
	wire [12-1:0] node827;
	wire [12-1:0] node831;
	wire [12-1:0] node832;
	wire [12-1:0] node835;
	wire [12-1:0] node838;
	wire [12-1:0] node839;
	wire [12-1:0] node840;
	wire [12-1:0] node841;
	wire [12-1:0] node842;
	wire [12-1:0] node843;
	wire [12-1:0] node844;
	wire [12-1:0] node845;
	wire [12-1:0] node847;
	wire [12-1:0] node850;
	wire [12-1:0] node851;
	wire [12-1:0] node854;
	wire [12-1:0] node857;
	wire [12-1:0] node858;
	wire [12-1:0] node859;
	wire [12-1:0] node863;
	wire [12-1:0] node864;
	wire [12-1:0] node867;
	wire [12-1:0] node870;
	wire [12-1:0] node871;
	wire [12-1:0] node872;
	wire [12-1:0] node873;
	wire [12-1:0] node877;
	wire [12-1:0] node878;
	wire [12-1:0] node881;
	wire [12-1:0] node884;
	wire [12-1:0] node885;
	wire [12-1:0] node886;
	wire [12-1:0] node889;
	wire [12-1:0] node892;
	wire [12-1:0] node893;
	wire [12-1:0] node897;
	wire [12-1:0] node898;
	wire [12-1:0] node899;
	wire [12-1:0] node900;
	wire [12-1:0] node901;
	wire [12-1:0] node905;
	wire [12-1:0] node906;
	wire [12-1:0] node910;
	wire [12-1:0] node911;
	wire [12-1:0] node912;
	wire [12-1:0] node915;
	wire [12-1:0] node918;
	wire [12-1:0] node919;
	wire [12-1:0] node923;
	wire [12-1:0] node924;
	wire [12-1:0] node925;
	wire [12-1:0] node926;
	wire [12-1:0] node930;
	wire [12-1:0] node931;
	wire [12-1:0] node934;
	wire [12-1:0] node937;
	wire [12-1:0] node939;
	wire [12-1:0] node940;
	wire [12-1:0] node943;
	wire [12-1:0] node946;
	wire [12-1:0] node947;
	wire [12-1:0] node948;
	wire [12-1:0] node949;
	wire [12-1:0] node950;
	wire [12-1:0] node951;
	wire [12-1:0] node955;
	wire [12-1:0] node956;
	wire [12-1:0] node960;
	wire [12-1:0] node961;
	wire [12-1:0] node962;
	wire [12-1:0] node965;
	wire [12-1:0] node968;
	wire [12-1:0] node969;
	wire [12-1:0] node972;
	wire [12-1:0] node975;
	wire [12-1:0] node976;
	wire [12-1:0] node977;
	wire [12-1:0] node979;
	wire [12-1:0] node982;
	wire [12-1:0] node983;
	wire [12-1:0] node987;
	wire [12-1:0] node988;
	wire [12-1:0] node989;
	wire [12-1:0] node992;
	wire [12-1:0] node996;
	wire [12-1:0] node997;
	wire [12-1:0] node998;
	wire [12-1:0] node999;
	wire [12-1:0] node1001;
	wire [12-1:0] node1004;
	wire [12-1:0] node1005;
	wire [12-1:0] node1008;
	wire [12-1:0] node1011;
	wire [12-1:0] node1012;
	wire [12-1:0] node1014;
	wire [12-1:0] node1017;
	wire [12-1:0] node1018;
	wire [12-1:0] node1022;
	wire [12-1:0] node1023;
	wire [12-1:0] node1024;
	wire [12-1:0] node1027;
	wire [12-1:0] node1028;
	wire [12-1:0] node1031;
	wire [12-1:0] node1034;
	wire [12-1:0] node1035;
	wire [12-1:0] node1038;
	wire [12-1:0] node1039;
	wire [12-1:0] node1042;
	wire [12-1:0] node1045;
	wire [12-1:0] node1046;
	wire [12-1:0] node1047;
	wire [12-1:0] node1048;
	wire [12-1:0] node1049;
	wire [12-1:0] node1050;
	wire [12-1:0] node1051;
	wire [12-1:0] node1054;
	wire [12-1:0] node1057;
	wire [12-1:0] node1059;
	wire [12-1:0] node1062;
	wire [12-1:0] node1063;
	wire [12-1:0] node1064;
	wire [12-1:0] node1068;
	wire [12-1:0] node1069;
	wire [12-1:0] node1072;
	wire [12-1:0] node1075;
	wire [12-1:0] node1076;
	wire [12-1:0] node1077;
	wire [12-1:0] node1078;
	wire [12-1:0] node1082;
	wire [12-1:0] node1083;
	wire [12-1:0] node1087;
	wire [12-1:0] node1088;
	wire [12-1:0] node1090;
	wire [12-1:0] node1093;
	wire [12-1:0] node1096;
	wire [12-1:0] node1097;
	wire [12-1:0] node1098;
	wire [12-1:0] node1099;
	wire [12-1:0] node1102;
	wire [12-1:0] node1103;
	wire [12-1:0] node1106;
	wire [12-1:0] node1109;
	wire [12-1:0] node1110;
	wire [12-1:0] node1111;
	wire [12-1:0] node1114;
	wire [12-1:0] node1117;
	wire [12-1:0] node1119;
	wire [12-1:0] node1122;
	wire [12-1:0] node1123;
	wire [12-1:0] node1124;
	wire [12-1:0] node1126;
	wire [12-1:0] node1129;
	wire [12-1:0] node1131;
	wire [12-1:0] node1134;
	wire [12-1:0] node1135;
	wire [12-1:0] node1136;
	wire [12-1:0] node1139;
	wire [12-1:0] node1143;
	wire [12-1:0] node1144;
	wire [12-1:0] node1145;
	wire [12-1:0] node1146;
	wire [12-1:0] node1147;
	wire [12-1:0] node1148;
	wire [12-1:0] node1151;
	wire [12-1:0] node1154;
	wire [12-1:0] node1155;
	wire [12-1:0] node1158;
	wire [12-1:0] node1161;
	wire [12-1:0] node1162;
	wire [12-1:0] node1163;
	wire [12-1:0] node1166;
	wire [12-1:0] node1169;
	wire [12-1:0] node1171;
	wire [12-1:0] node1174;
	wire [12-1:0] node1175;
	wire [12-1:0] node1176;
	wire [12-1:0] node1177;
	wire [12-1:0] node1180;
	wire [12-1:0] node1183;
	wire [12-1:0] node1184;
	wire [12-1:0] node1188;
	wire [12-1:0] node1189;
	wire [12-1:0] node1190;
	wire [12-1:0] node1193;
	wire [12-1:0] node1196;
	wire [12-1:0] node1197;
	wire [12-1:0] node1200;
	wire [12-1:0] node1203;
	wire [12-1:0] node1204;
	wire [12-1:0] node1205;
	wire [12-1:0] node1206;
	wire [12-1:0] node1208;
	wire [12-1:0] node1211;
	wire [12-1:0] node1212;
	wire [12-1:0] node1215;
	wire [12-1:0] node1218;
	wire [12-1:0] node1219;
	wire [12-1:0] node1220;
	wire [12-1:0] node1223;
	wire [12-1:0] node1226;
	wire [12-1:0] node1227;
	wire [12-1:0] node1230;
	wire [12-1:0] node1233;
	wire [12-1:0] node1234;
	wire [12-1:0] node1235;
	wire [12-1:0] node1236;
	wire [12-1:0] node1239;
	wire [12-1:0] node1242;
	wire [12-1:0] node1245;
	wire [12-1:0] node1246;
	wire [12-1:0] node1248;
	wire [12-1:0] node1251;
	wire [12-1:0] node1252;
	wire [12-1:0] node1255;
	wire [12-1:0] node1258;
	wire [12-1:0] node1259;
	wire [12-1:0] node1260;
	wire [12-1:0] node1261;
	wire [12-1:0] node1262;
	wire [12-1:0] node1263;
	wire [12-1:0] node1264;
	wire [12-1:0] node1265;
	wire [12-1:0] node1269;
	wire [12-1:0] node1270;
	wire [12-1:0] node1273;
	wire [12-1:0] node1276;
	wire [12-1:0] node1278;
	wire [12-1:0] node1279;
	wire [12-1:0] node1282;
	wire [12-1:0] node1285;
	wire [12-1:0] node1286;
	wire [12-1:0] node1287;
	wire [12-1:0] node1288;
	wire [12-1:0] node1293;
	wire [12-1:0] node1294;
	wire [12-1:0] node1297;
	wire [12-1:0] node1298;
	wire [12-1:0] node1301;
	wire [12-1:0] node1304;
	wire [12-1:0] node1305;
	wire [12-1:0] node1306;
	wire [12-1:0] node1307;
	wire [12-1:0] node1308;
	wire [12-1:0] node1312;
	wire [12-1:0] node1313;
	wire [12-1:0] node1316;
	wire [12-1:0] node1319;
	wire [12-1:0] node1320;
	wire [12-1:0] node1321;
	wire [12-1:0] node1324;
	wire [12-1:0] node1327;
	wire [12-1:0] node1329;
	wire [12-1:0] node1332;
	wire [12-1:0] node1333;
	wire [12-1:0] node1334;
	wire [12-1:0] node1338;
	wire [12-1:0] node1339;
	wire [12-1:0] node1341;
	wire [12-1:0] node1344;
	wire [12-1:0] node1345;
	wire [12-1:0] node1348;
	wire [12-1:0] node1351;
	wire [12-1:0] node1352;
	wire [12-1:0] node1353;
	wire [12-1:0] node1354;
	wire [12-1:0] node1355;
	wire [12-1:0] node1356;
	wire [12-1:0] node1359;
	wire [12-1:0] node1362;
	wire [12-1:0] node1365;
	wire [12-1:0] node1367;
	wire [12-1:0] node1368;
	wire [12-1:0] node1372;
	wire [12-1:0] node1373;
	wire [12-1:0] node1374;
	wire [12-1:0] node1375;
	wire [12-1:0] node1378;
	wire [12-1:0] node1381;
	wire [12-1:0] node1383;
	wire [12-1:0] node1386;
	wire [12-1:0] node1387;
	wire [12-1:0] node1389;
	wire [12-1:0] node1392;
	wire [12-1:0] node1393;
	wire [12-1:0] node1396;
	wire [12-1:0] node1399;
	wire [12-1:0] node1400;
	wire [12-1:0] node1401;
	wire [12-1:0] node1402;
	wire [12-1:0] node1404;
	wire [12-1:0] node1407;
	wire [12-1:0] node1408;
	wire [12-1:0] node1411;
	wire [12-1:0] node1414;
	wire [12-1:0] node1416;
	wire [12-1:0] node1417;
	wire [12-1:0] node1421;
	wire [12-1:0] node1422;
	wire [12-1:0] node1423;
	wire [12-1:0] node1424;
	wire [12-1:0] node1427;
	wire [12-1:0] node1430;
	wire [12-1:0] node1431;
	wire [12-1:0] node1434;
	wire [12-1:0] node1437;
	wire [12-1:0] node1438;
	wire [12-1:0] node1439;
	wire [12-1:0] node1442;
	wire [12-1:0] node1445;
	wire [12-1:0] node1447;
	wire [12-1:0] node1450;
	wire [12-1:0] node1451;
	wire [12-1:0] node1452;
	wire [12-1:0] node1453;
	wire [12-1:0] node1454;
	wire [12-1:0] node1455;
	wire [12-1:0] node1456;
	wire [12-1:0] node1461;
	wire [12-1:0] node1462;
	wire [12-1:0] node1463;
	wire [12-1:0] node1466;
	wire [12-1:0] node1470;
	wire [12-1:0] node1471;
	wire [12-1:0] node1472;
	wire [12-1:0] node1473;
	wire [12-1:0] node1476;
	wire [12-1:0] node1479;
	wire [12-1:0] node1482;
	wire [12-1:0] node1483;
	wire [12-1:0] node1485;
	wire [12-1:0] node1488;
	wire [12-1:0] node1489;
	wire [12-1:0] node1492;
	wire [12-1:0] node1495;
	wire [12-1:0] node1496;
	wire [12-1:0] node1497;
	wire [12-1:0] node1498;
	wire [12-1:0] node1500;
	wire [12-1:0] node1503;
	wire [12-1:0] node1505;
	wire [12-1:0] node1508;
	wire [12-1:0] node1509;
	wire [12-1:0] node1510;
	wire [12-1:0] node1513;
	wire [12-1:0] node1516;
	wire [12-1:0] node1519;
	wire [12-1:0] node1520;
	wire [12-1:0] node1521;
	wire [12-1:0] node1522;
	wire [12-1:0] node1525;
	wire [12-1:0] node1528;
	wire [12-1:0] node1529;
	wire [12-1:0] node1532;
	wire [12-1:0] node1535;
	wire [12-1:0] node1536;
	wire [12-1:0] node1538;
	wire [12-1:0] node1541;
	wire [12-1:0] node1544;
	wire [12-1:0] node1545;
	wire [12-1:0] node1546;
	wire [12-1:0] node1547;
	wire [12-1:0] node1548;
	wire [12-1:0] node1549;
	wire [12-1:0] node1553;
	wire [12-1:0] node1555;
	wire [12-1:0] node1558;
	wire [12-1:0] node1559;
	wire [12-1:0] node1560;
	wire [12-1:0] node1564;
	wire [12-1:0] node1565;
	wire [12-1:0] node1569;
	wire [12-1:0] node1570;
	wire [12-1:0] node1571;
	wire [12-1:0] node1573;
	wire [12-1:0] node1576;
	wire [12-1:0] node1577;
	wire [12-1:0] node1581;
	wire [12-1:0] node1582;
	wire [12-1:0] node1583;
	wire [12-1:0] node1586;
	wire [12-1:0] node1589;
	wire [12-1:0] node1590;
	wire [12-1:0] node1593;
	wire [12-1:0] node1596;
	wire [12-1:0] node1597;
	wire [12-1:0] node1598;
	wire [12-1:0] node1599;
	wire [12-1:0] node1600;
	wire [12-1:0] node1603;
	wire [12-1:0] node1606;
	wire [12-1:0] node1607;
	wire [12-1:0] node1611;
	wire [12-1:0] node1612;
	wire [12-1:0] node1615;
	wire [12-1:0] node1617;
	wire [12-1:0] node1620;
	wire [12-1:0] node1621;
	wire [12-1:0] node1622;
	wire [12-1:0] node1624;
	wire [12-1:0] node1627;
	wire [12-1:0] node1628;
	wire [12-1:0] node1631;
	wire [12-1:0] node1634;
	wire [12-1:0] node1635;
	wire [12-1:0] node1637;
	wire [12-1:0] node1640;
	wire [12-1:0] node1641;
	wire [12-1:0] node1644;

	assign outp = (inp[7]) ? node838 : node1;
		assign node1 = (inp[0]) ? node411 : node2;
			assign node2 = (inp[1]) ? node204 : node3;
				assign node3 = (inp[3]) ? node107 : node4;
					assign node4 = (inp[9]) ? node64 : node5;
						assign node5 = (inp[2]) ? node35 : node6;
							assign node6 = (inp[10]) ? node22 : node7;
								assign node7 = (inp[11]) ? node15 : node8;
									assign node8 = (inp[4]) ? node12 : node9;
										assign node9 = (inp[5]) ? 12'b001111111111 : 12'b011111111111;
										assign node12 = (inp[6]) ? 12'b000111111111 : 12'b001111111111;
									assign node15 = (inp[4]) ? node19 : node16;
										assign node16 = (inp[6]) ? 12'b000111111111 : 12'b001111111111;
										assign node19 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
								assign node22 = (inp[11]) ? node28 : node23;
									assign node23 = (inp[4]) ? 12'b000111111111 : node24;
										assign node24 = (inp[6]) ? 12'b000111111111 : 12'b001111111111;
									assign node28 = (inp[6]) ? node32 : node29;
										assign node29 = (inp[8]) ? 12'b000011111111 : 12'b000111111111;
										assign node32 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
							assign node35 = (inp[6]) ? node49 : node36;
								assign node36 = (inp[4]) ? node42 : node37;
									assign node37 = (inp[10]) ? node39 : 12'b001111111111;
										assign node39 = (inp[8]) ? 12'b000011111111 : 12'b000111111111;
									assign node42 = (inp[5]) ? node46 : node43;
										assign node43 = (inp[8]) ? 12'b000011111111 : 12'b000011111111;
										assign node46 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
								assign node49 = (inp[11]) ? node57 : node50;
									assign node50 = (inp[10]) ? node54 : node51;
										assign node51 = (inp[8]) ? 12'b000111111111 : 12'b000011111111;
										assign node54 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node57 = (inp[5]) ? node61 : node58;
										assign node58 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
										assign node61 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
						assign node64 = (inp[8]) ? node88 : node65;
							assign node65 = (inp[10]) ? node77 : node66;
								assign node66 = (inp[6]) ? node72 : node67;
									assign node67 = (inp[2]) ? node69 : 12'b000111111111;
										assign node69 = (inp[11]) ? 12'b000011111111 : 12'b000111111111;
									assign node72 = (inp[2]) ? node74 : 12'b000111111111;
										assign node74 = (inp[4]) ? 12'b000001111111 : 12'b000001111111;
								assign node77 = (inp[4]) ? node83 : node78;
									assign node78 = (inp[11]) ? node80 : 12'b000111111111;
										assign node80 = (inp[5]) ? 12'b000000111111 : 12'b000011111111;
									assign node83 = (inp[6]) ? 12'b000001111111 : node84;
										assign node84 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
							assign node88 = (inp[11]) ? node98 : node89;
								assign node89 = (inp[6]) ? node93 : node90;
									assign node90 = (inp[10]) ? 12'b000111111111 : 12'b000011111111;
									assign node93 = (inp[5]) ? 12'b000001111111 : node94;
										assign node94 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
								assign node98 = (inp[10]) ? node104 : node99;
									assign node99 = (inp[4]) ? 12'b000001111111 : node100;
										assign node100 = (inp[6]) ? 12'b000001111111 : 12'b000011111111;
									assign node104 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
					assign node107 = (inp[9]) ? node157 : node108;
						assign node108 = (inp[8]) ? node138 : node109;
							assign node109 = (inp[4]) ? node125 : node110;
								assign node110 = (inp[11]) ? node118 : node111;
									assign node111 = (inp[2]) ? node115 : node112;
										assign node112 = (inp[5]) ? 12'b000111111111 : 12'b000111111111;
										assign node115 = (inp[6]) ? 12'b000011111111 : 12'b000111111111;
									assign node118 = (inp[5]) ? node122 : node119;
										assign node119 = (inp[2]) ? 12'b000011111111 : 12'b000111111111;
										assign node122 = (inp[10]) ? 12'b000000111111 : 12'b000011111111;
								assign node125 = (inp[11]) ? node133 : node126;
									assign node126 = (inp[6]) ? node130 : node127;
										assign node127 = (inp[2]) ? 12'b000011111111 : 12'b001111111111;
										assign node130 = (inp[5]) ? 12'b000001111111 : 12'b000001111111;
									assign node133 = (inp[5]) ? node135 : 12'b000001111111;
										assign node135 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
							assign node138 = (inp[6]) ? node150 : node139;
								assign node139 = (inp[5]) ? node145 : node140;
									assign node140 = (inp[2]) ? node142 : 12'b001111111111;
										assign node142 = (inp[4]) ? 12'b000001111111 : 12'b000011111111;
									assign node145 = (inp[11]) ? node147 : 12'b000001111111;
										assign node147 = (inp[4]) ? 12'b000001111111 : 12'b000001111111;
								assign node150 = (inp[11]) ? node152 : 12'b000001111111;
									assign node152 = (inp[5]) ? 12'b000000111111 : node153;
										assign node153 = (inp[10]) ? 12'b000000111111 : 12'b000001111111;
						assign node157 = (inp[2]) ? node179 : node158;
							assign node158 = (inp[6]) ? node170 : node159;
								assign node159 = (inp[4]) ? node163 : node160;
									assign node160 = (inp[10]) ? 12'b000011111111 : 12'b001111111111;
									assign node163 = (inp[10]) ? node167 : node164;
										assign node164 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
										assign node167 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
								assign node170 = (inp[11]) ? 12'b000000111111 : node171;
									assign node171 = (inp[5]) ? node175 : node172;
										assign node172 = (inp[10]) ? 12'b000001111111 : 12'b000111111111;
										assign node175 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
							assign node179 = (inp[8]) ? node191 : node180;
								assign node180 = (inp[4]) ? node184 : node181;
									assign node181 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
									assign node184 = (inp[11]) ? node188 : node185;
										assign node185 = (inp[5]) ? 12'b000000111111 : 12'b000011111111;
										assign node188 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
								assign node191 = (inp[5]) ? node199 : node192;
									assign node192 = (inp[6]) ? node196 : node193;
										assign node193 = (inp[4]) ? 12'b000000111111 : 12'b000000111111;
										assign node196 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
									assign node199 = (inp[6]) ? 12'b000000001111 : node200;
										assign node200 = (inp[4]) ? 12'b000000011111 : 12'b000000011111;
				assign node204 = (inp[4]) ? node310 : node205;
					assign node205 = (inp[10]) ? node259 : node206;
						assign node206 = (inp[6]) ? node234 : node207;
							assign node207 = (inp[2]) ? node221 : node208;
								assign node208 = (inp[9]) ? node216 : node209;
									assign node209 = (inp[11]) ? node213 : node210;
										assign node210 = (inp[5]) ? 12'b000111111111 : 12'b001111111111;
										assign node213 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
									assign node216 = (inp[8]) ? 12'b000011111111 : node217;
										assign node217 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
								assign node221 = (inp[8]) ? node229 : node222;
									assign node222 = (inp[11]) ? node226 : node223;
										assign node223 = (inp[9]) ? 12'b000011111111 : 12'b000111111111;
										assign node226 = (inp[9]) ? 12'b000011111111 : 12'b000001111111;
									assign node229 = (inp[3]) ? 12'b000001111111 : node230;
										assign node230 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
							assign node234 = (inp[11]) ? node246 : node235;
								assign node235 = (inp[9]) ? node241 : node236;
									assign node236 = (inp[8]) ? node238 : 12'b000111111111;
										assign node238 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
									assign node241 = (inp[5]) ? 12'b000000111111 : node242;
										assign node242 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
								assign node246 = (inp[3]) ? node252 : node247;
									assign node247 = (inp[8]) ? 12'b000001111111 : node248;
										assign node248 = (inp[2]) ? 12'b000001111111 : 12'b000001111111;
									assign node252 = (inp[2]) ? node256 : node253;
										assign node253 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
										assign node256 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
						assign node259 = (inp[6]) ? node285 : node260;
							assign node260 = (inp[11]) ? node274 : node261;
								assign node261 = (inp[5]) ? node269 : node262;
									assign node262 = (inp[8]) ? node266 : node263;
										assign node263 = (inp[9]) ? 12'b000011111111 : 12'b000111111111;
										assign node266 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
									assign node269 = (inp[2]) ? node271 : 12'b000001111111;
										assign node271 = (inp[3]) ? 12'b000001111111 : 12'b000011111111;
								assign node274 = (inp[3]) ? node280 : node275;
									assign node275 = (inp[9]) ? node277 : 12'b000011111111;
										assign node277 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
									assign node280 = (inp[5]) ? node282 : 12'b000000111111;
										assign node282 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
							assign node285 = (inp[2]) ? node299 : node286;
								assign node286 = (inp[8]) ? node292 : node287;
									assign node287 = (inp[9]) ? node289 : 12'b000011111111;
										assign node289 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node292 = (inp[5]) ? node296 : node293;
										assign node293 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
										assign node296 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
								assign node299 = (inp[3]) ? node305 : node300;
									assign node300 = (inp[8]) ? 12'b000000011111 : node301;
										assign node301 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node305 = (inp[9]) ? 12'b000000011111 : node306;
										assign node306 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
					assign node310 = (inp[8]) ? node360 : node311;
						assign node311 = (inp[5]) ? node337 : node312;
							assign node312 = (inp[9]) ? node326 : node313;
								assign node313 = (inp[6]) ? node321 : node314;
									assign node314 = (inp[10]) ? node318 : node315;
										assign node315 = (inp[2]) ? 12'b000011111111 : 12'b000111111111;
										assign node318 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
									assign node321 = (inp[11]) ? 12'b000001111111 : node322;
										assign node322 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
								assign node326 = (inp[2]) ? node332 : node327;
									assign node327 = (inp[6]) ? 12'b000001111111 : node328;
										assign node328 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
									assign node332 = (inp[3]) ? node334 : 12'b000001111111;
										assign node334 = (inp[11]) ? 12'b000000001111 : 12'b000000111111;
							assign node337 = (inp[6]) ? node351 : node338;
								assign node338 = (inp[11]) ? node346 : node339;
									assign node339 = (inp[3]) ? node343 : node340;
										assign node340 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
										assign node343 = (inp[10]) ? 12'b000000011111 : 12'b000001111111;
									assign node346 = (inp[2]) ? node348 : 12'b000000111111;
										assign node348 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
								assign node351 = (inp[9]) ? node355 : node352;
									assign node352 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
									assign node355 = (inp[10]) ? node357 : 12'b000000011111;
										assign node357 = (inp[2]) ? 12'b000000000111 : 12'b000000011111;
						assign node360 = (inp[10]) ? node384 : node361;
							assign node361 = (inp[3]) ? node369 : node362;
								assign node362 = (inp[11]) ? 12'b000000111111 : node363;
									assign node363 = (inp[6]) ? 12'b000000111111 : node364;
										assign node364 = (inp[5]) ? 12'b000000111111 : 12'b000011111111;
								assign node369 = (inp[2]) ? node377 : node370;
									assign node370 = (inp[11]) ? node374 : node371;
										assign node371 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
										assign node374 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
									assign node377 = (inp[11]) ? node381 : node378;
										assign node378 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
										assign node381 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
							assign node384 = (inp[3]) ? node400 : node385;
								assign node385 = (inp[2]) ? node393 : node386;
									assign node386 = (inp[11]) ? node390 : node387;
										assign node387 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
										assign node390 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
									assign node393 = (inp[11]) ? node397 : node394;
										assign node394 = (inp[9]) ? 12'b000000011111 : 12'b000000011111;
										assign node397 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
								assign node400 = (inp[6]) ? node406 : node401;
									assign node401 = (inp[11]) ? 12'b000000001111 : node402;
										assign node402 = (inp[2]) ? 12'b000000001111 : 12'b000000111111;
									assign node406 = (inp[9]) ? node408 : 12'b000000001111;
										assign node408 = (inp[11]) ? 12'b000000000111 : 12'b000000000111;
			assign node411 = (inp[4]) ? node617 : node412;
				assign node412 = (inp[9]) ? node514 : node413;
					assign node413 = (inp[6]) ? node467 : node414;
						assign node414 = (inp[2]) ? node440 : node415;
							assign node415 = (inp[3]) ? node429 : node416;
								assign node416 = (inp[11]) ? node424 : node417;
									assign node417 = (inp[10]) ? node421 : node418;
										assign node418 = (inp[1]) ? 12'b000111111111 : 12'b001111111111;
										assign node421 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
									assign node424 = (inp[5]) ? 12'b000011111111 : node425;
										assign node425 = (inp[8]) ? 12'b000111111111 : 12'b000011111111;
								assign node429 = (inp[1]) ? node435 : node430;
									assign node430 = (inp[8]) ? node432 : 12'b000011111111;
										assign node432 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
									assign node435 = (inp[10]) ? 12'b000000111111 : node436;
										assign node436 = (inp[8]) ? 12'b000001111111 : 12'b000111111111;
							assign node440 = (inp[11]) ? node454 : node441;
								assign node441 = (inp[1]) ? node449 : node442;
									assign node442 = (inp[5]) ? node446 : node443;
										assign node443 = (inp[8]) ? 12'b000011111111 : 12'b000111111111;
										assign node446 = (inp[3]) ? 12'b000001111111 : 12'b000011111111;
									assign node449 = (inp[10]) ? node451 : 12'b000011111111;
										assign node451 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
								assign node454 = (inp[10]) ? node460 : node455;
									assign node455 = (inp[8]) ? 12'b000001111111 : node456;
										assign node456 = (inp[3]) ? 12'b000001111111 : 12'b000011111111;
									assign node460 = (inp[3]) ? node464 : node461;
										assign node461 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node464 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
						assign node467 = (inp[5]) ? node485 : node468;
							assign node468 = (inp[3]) ? node472 : node469;
								assign node469 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
								assign node472 = (inp[10]) ? node480 : node473;
									assign node473 = (inp[1]) ? node477 : node474;
										assign node474 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
										assign node477 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
									assign node480 = (inp[11]) ? node482 : 12'b000000111111;
										assign node482 = (inp[1]) ? 12'b000000111111 : 12'b000000111111;
							assign node485 = (inp[3]) ? node501 : node486;
								assign node486 = (inp[11]) ? node494 : node487;
									assign node487 = (inp[8]) ? node491 : node488;
										assign node488 = (inp[2]) ? 12'b000001111111 : 12'b000011111111;
										assign node491 = (inp[2]) ? 12'b000000111111 : 12'b000001111111;
									assign node494 = (inp[2]) ? node498 : node495;
										assign node495 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node498 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
								assign node501 = (inp[10]) ? node509 : node502;
									assign node502 = (inp[8]) ? node506 : node503;
										assign node503 = (inp[2]) ? 12'b000000111111 : 12'b000000111111;
										assign node506 = (inp[2]) ? 12'b000000001111 : 12'b000000111111;
									assign node509 = (inp[2]) ? node511 : 12'b000000011111;
										assign node511 = (inp[1]) ? 12'b000000001111 : 12'b000000001111;
					assign node514 = (inp[8]) ? node570 : node515;
						assign node515 = (inp[11]) ? node543 : node516;
							assign node516 = (inp[1]) ? node530 : node517;
								assign node517 = (inp[6]) ? node523 : node518;
									assign node518 = (inp[5]) ? 12'b000001111111 : node519;
										assign node519 = (inp[10]) ? 12'b000011111111 : 12'b000111111111;
									assign node523 = (inp[10]) ? node527 : node524;
										assign node524 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
										assign node527 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
								assign node530 = (inp[3]) ? node538 : node531;
									assign node531 = (inp[10]) ? node535 : node532;
										assign node532 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
										assign node535 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
									assign node538 = (inp[10]) ? node540 : 12'b000000111111;
										assign node540 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
							assign node543 = (inp[5]) ? node557 : node544;
								assign node544 = (inp[2]) ? node550 : node545;
									assign node545 = (inp[3]) ? node547 : 12'b000011111111;
										assign node547 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
									assign node550 = (inp[10]) ? node554 : node551;
										assign node551 = (inp[3]) ? 12'b000000111111 : 12'b000000111111;
										assign node554 = (inp[6]) ? 12'b000000111111 : 12'b000000011111;
								assign node557 = (inp[1]) ? node565 : node558;
									assign node558 = (inp[10]) ? node562 : node559;
										assign node559 = (inp[2]) ? 12'b000000111111 : 12'b000000111111;
										assign node562 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
									assign node565 = (inp[6]) ? node567 : 12'b000000111111;
										assign node567 = (inp[10]) ? 12'b000000001111 : 12'b000000011111;
						assign node570 = (inp[6]) ? node596 : node571;
							assign node571 = (inp[2]) ? node585 : node572;
								assign node572 = (inp[1]) ? node580 : node573;
									assign node573 = (inp[11]) ? node577 : node574;
										assign node574 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
										assign node577 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
									assign node580 = (inp[10]) ? 12'b000000111111 : node581;
										assign node581 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
								assign node585 = (inp[11]) ? node591 : node586;
									assign node586 = (inp[3]) ? 12'b000001111111 : node587;
										assign node587 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
									assign node591 = (inp[10]) ? node593 : 12'b000000011111;
										assign node593 = (inp[1]) ? 12'b000000000111 : 12'b000000001111;
							assign node596 = (inp[1]) ? node606 : node597;
								assign node597 = (inp[3]) ? 12'b000000011111 : node598;
									assign node598 = (inp[2]) ? node602 : node599;
										assign node599 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
										assign node602 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
								assign node606 = (inp[5]) ? node612 : node607;
									assign node607 = (inp[11]) ? node609 : 12'b000000011111;
										assign node609 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
									assign node612 = (inp[2]) ? 12'b000000001111 : node613;
										assign node613 = (inp[10]) ? 12'b000000001111 : 12'b000000011111;
				assign node617 = (inp[10]) ? node731 : node618;
					assign node618 = (inp[5]) ? node672 : node619;
						assign node619 = (inp[1]) ? node647 : node620;
							assign node620 = (inp[6]) ? node632 : node621;
								assign node621 = (inp[9]) ? node627 : node622;
									assign node622 = (inp[11]) ? 12'b000011111111 : node623;
										assign node623 = (inp[2]) ? 12'b000011111111 : 12'b000111111111;
									assign node627 = (inp[3]) ? node629 : 12'b000011111111;
										assign node629 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
								assign node632 = (inp[8]) ? node640 : node633;
									assign node633 = (inp[3]) ? node637 : node634;
										assign node634 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
										assign node637 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node640 = (inp[9]) ? node644 : node641;
										assign node641 = (inp[2]) ? 12'b000000111111 : 12'b000000111111;
										assign node644 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
							assign node647 = (inp[11]) ? node657 : node648;
								assign node648 = (inp[6]) ? node654 : node649;
									assign node649 = (inp[2]) ? node651 : 12'b000001111111;
										assign node651 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
									assign node654 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
								assign node657 = (inp[2]) ? node665 : node658;
									assign node658 = (inp[8]) ? node662 : node659;
										assign node659 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
										assign node662 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
									assign node665 = (inp[9]) ? node669 : node666;
										assign node666 = (inp[6]) ? 12'b000000011111 : 12'b000000011111;
										assign node669 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
						assign node672 = (inp[6]) ? node702 : node673;
							assign node673 = (inp[3]) ? node689 : node674;
								assign node674 = (inp[2]) ? node682 : node675;
									assign node675 = (inp[8]) ? node679 : node676;
										assign node676 = (inp[1]) ? 12'b000001111111 : 12'b000001111111;
										assign node679 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
									assign node682 = (inp[9]) ? node686 : node683;
										assign node683 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node686 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
								assign node689 = (inp[11]) ? node697 : node690;
									assign node690 = (inp[8]) ? node694 : node691;
										assign node691 = (inp[1]) ? 12'b000000111111 : 12'b000001111111;
										assign node694 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
									assign node697 = (inp[1]) ? 12'b000000011111 : node698;
										assign node698 = (inp[2]) ? 12'b000000011111 : 12'b000000111111;
							assign node702 = (inp[9]) ? node718 : node703;
								assign node703 = (inp[11]) ? node711 : node704;
									assign node704 = (inp[8]) ? node708 : node705;
										assign node705 = (inp[3]) ? 12'b000001111111 : 12'b000000111111;
										assign node708 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
									assign node711 = (inp[2]) ? node715 : node712;
										assign node712 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
										assign node715 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
								assign node718 = (inp[1]) ? node726 : node719;
									assign node719 = (inp[11]) ? node723 : node720;
										assign node720 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
										assign node723 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
									assign node726 = (inp[2]) ? node728 : 12'b000000001111;
										assign node728 = (inp[11]) ? 12'b000000000011 : 12'b000000000111;
					assign node731 = (inp[8]) ? node791 : node732;
						assign node732 = (inp[9]) ? node762 : node733;
							assign node733 = (inp[3]) ? node747 : node734;
								assign node734 = (inp[1]) ? node742 : node735;
									assign node735 = (inp[6]) ? node739 : node736;
										assign node736 = (inp[11]) ? 12'b000001111111 : 12'b000011111111;
										assign node739 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
									assign node742 = (inp[11]) ? 12'b000000111111 : node743;
										assign node743 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
								assign node747 = (inp[2]) ? node755 : node748;
									assign node748 = (inp[11]) ? node752 : node749;
										assign node749 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
										assign node752 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
									assign node755 = (inp[11]) ? node759 : node756;
										assign node756 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
										assign node759 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
							assign node762 = (inp[3]) ? node778 : node763;
								assign node763 = (inp[5]) ? node771 : node764;
									assign node764 = (inp[2]) ? node768 : node765;
										assign node765 = (inp[6]) ? 12'b000000111111 : 12'b000000111111;
										assign node768 = (inp[11]) ? 12'b000000111111 : 12'b000000111111;
									assign node771 = (inp[2]) ? node775 : node772;
										assign node772 = (inp[1]) ? 12'b000000011111 : 12'b000000111111;
										assign node775 = (inp[11]) ? 12'b000000001111 : 12'b000000001111;
								assign node778 = (inp[6]) ? node784 : node779;
									assign node779 = (inp[2]) ? 12'b000000001111 : node780;
										assign node780 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
									assign node784 = (inp[1]) ? node788 : node785;
										assign node785 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
										assign node788 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
						assign node791 = (inp[5]) ? node815 : node792;
							assign node792 = (inp[11]) ? node802 : node793;
								assign node793 = (inp[3]) ? node799 : node794;
									assign node794 = (inp[6]) ? node796 : 12'b000000111111;
										assign node796 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
									assign node799 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
								assign node802 = (inp[6]) ? node808 : node803;
									assign node803 = (inp[9]) ? node805 : 12'b000000111111;
										assign node805 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
									assign node808 = (inp[2]) ? node812 : node809;
										assign node809 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
										assign node812 = (inp[3]) ? 12'b000000000111 : 12'b000000001111;
							assign node815 = (inp[9]) ? node825 : node816;
								assign node816 = (inp[3]) ? node820 : node817;
									assign node817 = (inp[11]) ? 12'b000000001111 : 12'b000000111111;
									assign node820 = (inp[6]) ? 12'b000000001111 : node821;
										assign node821 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
								assign node825 = (inp[2]) ? node831 : node826;
									assign node826 = (inp[6]) ? 12'b000000000111 : node827;
										assign node827 = (inp[1]) ? 12'b000000001111 : 12'b000000011111;
									assign node831 = (inp[11]) ? node835 : node832;
										assign node832 = (inp[1]) ? 12'b000000000111 : 12'b000000000111;
										assign node835 = (inp[3]) ? 12'b000000000011 : 12'b000000000111;
		assign node838 = (inp[1]) ? node1258 : node839;
			assign node839 = (inp[2]) ? node1045 : node840;
				assign node840 = (inp[4]) ? node946 : node841;
					assign node841 = (inp[11]) ? node897 : node842;
						assign node842 = (inp[10]) ? node870 : node843;
							assign node843 = (inp[9]) ? node857 : node844;
								assign node844 = (inp[3]) ? node850 : node845;
									assign node845 = (inp[8]) ? node847 : 12'b001111111111;
										assign node847 = (inp[5]) ? 12'b000111111111 : 12'b000111111111;
									assign node850 = (inp[8]) ? node854 : node851;
										assign node851 = (inp[0]) ? 12'b000111111111 : 12'b001111111111;
										assign node854 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
								assign node857 = (inp[5]) ? node863 : node858;
									assign node858 = (inp[8]) ? 12'b000011111111 : node859;
										assign node859 = (inp[3]) ? 12'b000011111111 : 12'b000111111111;
									assign node863 = (inp[6]) ? node867 : node864;
										assign node864 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
										assign node867 = (inp[3]) ? 12'b000001111111 : 12'b000000111111;
							assign node870 = (inp[8]) ? node884 : node871;
								assign node871 = (inp[0]) ? node877 : node872;
									assign node872 = (inp[9]) ? 12'b000011111111 : node873;
										assign node873 = (inp[5]) ? 12'b000011111111 : 12'b000111111111;
									assign node877 = (inp[3]) ? node881 : node878;
										assign node878 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
										assign node881 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
								assign node884 = (inp[6]) ? node892 : node885;
									assign node885 = (inp[9]) ? node889 : node886;
										assign node886 = (inp[5]) ? 12'b000001111111 : 12'b000001111111;
										assign node889 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
									assign node892 = (inp[0]) ? 12'b000000111111 : node893;
										assign node893 = (inp[3]) ? 12'b000000111111 : 12'b000011111111;
						assign node897 = (inp[3]) ? node923 : node898;
							assign node898 = (inp[9]) ? node910 : node899;
								assign node899 = (inp[6]) ? node905 : node900;
									assign node900 = (inp[0]) ? 12'b000011111111 : node901;
										assign node901 = (inp[10]) ? 12'b000011111111 : 12'b000111111111;
									assign node905 = (inp[8]) ? 12'b000001111111 : node906;
										assign node906 = (inp[10]) ? 12'b000001111111 : 12'b000111111111;
								assign node910 = (inp[0]) ? node918 : node911;
									assign node911 = (inp[8]) ? node915 : node912;
										assign node912 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
										assign node915 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
									assign node918 = (inp[8]) ? 12'b000000001111 : node919;
										assign node919 = (inp[5]) ? 12'b000000111111 : 12'b000001111111;
							assign node923 = (inp[9]) ? node937 : node924;
								assign node924 = (inp[8]) ? node930 : node925;
									assign node925 = (inp[5]) ? 12'b000001111111 : node926;
										assign node926 = (inp[0]) ? 12'b000011111111 : 12'b000011111111;
									assign node930 = (inp[0]) ? node934 : node931;
										assign node931 = (inp[10]) ? 12'b000000111111 : 12'b000000111111;
										assign node934 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
								assign node937 = (inp[10]) ? node939 : 12'b000000111111;
									assign node939 = (inp[5]) ? node943 : node940;
										assign node940 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
										assign node943 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
					assign node946 = (inp[5]) ? node996 : node947;
						assign node947 = (inp[10]) ? node975 : node948;
							assign node948 = (inp[6]) ? node960 : node949;
								assign node949 = (inp[11]) ? node955 : node950;
									assign node950 = (inp[9]) ? 12'b000001111111 : node951;
										assign node951 = (inp[3]) ? 12'b000011111111 : 12'b000111111111;
									assign node955 = (inp[0]) ? 12'b000001111111 : node956;
										assign node956 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
								assign node960 = (inp[3]) ? node968 : node961;
									assign node961 = (inp[0]) ? node965 : node962;
										assign node962 = (inp[9]) ? 12'b000001111111 : 12'b000001111111;
										assign node965 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
									assign node968 = (inp[0]) ? node972 : node969;
										assign node969 = (inp[9]) ? 12'b000000111111 : 12'b000000111111;
										assign node972 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
							assign node975 = (inp[8]) ? node987 : node976;
								assign node976 = (inp[0]) ? node982 : node977;
									assign node977 = (inp[11]) ? node979 : 12'b000001111111;
										assign node979 = (inp[6]) ? 12'b000001111111 : 12'b000000111111;
									assign node982 = (inp[11]) ? 12'b000000111111 : node983;
										assign node983 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
								assign node987 = (inp[0]) ? 12'b000000011111 : node988;
									assign node988 = (inp[3]) ? node992 : node989;
										assign node989 = (inp[9]) ? 12'b000000111111 : 12'b000000111111;
										assign node992 = (inp[11]) ? 12'b000000011111 : 12'b000001111111;
						assign node996 = (inp[9]) ? node1022 : node997;
							assign node997 = (inp[10]) ? node1011 : node998;
								assign node998 = (inp[0]) ? node1004 : node999;
									assign node999 = (inp[3]) ? node1001 : 12'b000111111111;
										assign node1001 = (inp[8]) ? 12'b000000111111 : 12'b000001111111;
									assign node1004 = (inp[11]) ? node1008 : node1005;
										assign node1005 = (inp[6]) ? 12'b000000111111 : 12'b000000111111;
										assign node1008 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
								assign node1011 = (inp[8]) ? node1017 : node1012;
									assign node1012 = (inp[6]) ? node1014 : 12'b000000111111;
										assign node1014 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
									assign node1017 = (inp[0]) ? 12'b000000011111 : node1018;
										assign node1018 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
							assign node1022 = (inp[3]) ? node1034 : node1023;
								assign node1023 = (inp[11]) ? node1027 : node1024;
									assign node1024 = (inp[8]) ? 12'b000000011111 : 12'b000001111111;
									assign node1027 = (inp[0]) ? node1031 : node1028;
										assign node1028 = (inp[8]) ? 12'b000000011111 : 12'b000000011111;
										assign node1031 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
								assign node1034 = (inp[6]) ? node1038 : node1035;
									assign node1035 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
									assign node1038 = (inp[8]) ? node1042 : node1039;
										assign node1039 = (inp[10]) ? 12'b000000000111 : 12'b000000001111;
										assign node1042 = (inp[11]) ? 12'b000000000011 : 12'b000000000111;
				assign node1045 = (inp[0]) ? node1143 : node1046;
					assign node1046 = (inp[10]) ? node1096 : node1047;
						assign node1047 = (inp[5]) ? node1075 : node1048;
							assign node1048 = (inp[4]) ? node1062 : node1049;
								assign node1049 = (inp[11]) ? node1057 : node1050;
									assign node1050 = (inp[9]) ? node1054 : node1051;
										assign node1051 = (inp[6]) ? 12'b000111111111 : 12'b000111111111;
										assign node1054 = (inp[8]) ? 12'b000011111111 : 12'b000011111111;
									assign node1057 = (inp[8]) ? node1059 : 12'b000011111111;
										assign node1059 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
								assign node1062 = (inp[8]) ? node1068 : node1063;
									assign node1063 = (inp[6]) ? 12'b000001111111 : node1064;
										assign node1064 = (inp[3]) ? 12'b000001111111 : 12'b000011111111;
									assign node1068 = (inp[6]) ? node1072 : node1069;
										assign node1069 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node1072 = (inp[3]) ? 12'b000000001111 : 12'b000000111111;
							assign node1075 = (inp[3]) ? node1087 : node1076;
								assign node1076 = (inp[11]) ? node1082 : node1077;
									assign node1077 = (inp[9]) ? 12'b000000111111 : node1078;
										assign node1078 = (inp[8]) ? 12'b000001111111 : 12'b000011111111;
									assign node1082 = (inp[9]) ? 12'b000000111111 : node1083;
										assign node1083 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
								assign node1087 = (inp[6]) ? node1093 : node1088;
									assign node1088 = (inp[11]) ? node1090 : 12'b000001111111;
										assign node1090 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
									assign node1093 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
						assign node1096 = (inp[6]) ? node1122 : node1097;
							assign node1097 = (inp[8]) ? node1109 : node1098;
								assign node1098 = (inp[9]) ? node1102 : node1099;
									assign node1099 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
									assign node1102 = (inp[3]) ? node1106 : node1103;
										assign node1103 = (inp[5]) ? 12'b000000111111 : 12'b000011111111;
										assign node1106 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
								assign node1109 = (inp[3]) ? node1117 : node1110;
									assign node1110 = (inp[5]) ? node1114 : node1111;
										assign node1111 = (inp[11]) ? 12'b000000111111 : 12'b000001111111;
										assign node1114 = (inp[11]) ? 12'b000000001111 : 12'b000000111111;
									assign node1117 = (inp[5]) ? node1119 : 12'b000000011111;
										assign node1119 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
							assign node1122 = (inp[3]) ? node1134 : node1123;
								assign node1123 = (inp[4]) ? node1129 : node1124;
									assign node1124 = (inp[9]) ? node1126 : 12'b000000111111;
										assign node1126 = (inp[8]) ? 12'b000000011111 : 12'b000000111111;
									assign node1129 = (inp[9]) ? node1131 : 12'b000000011111;
										assign node1131 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
								assign node1134 = (inp[11]) ? 12'b000000001111 : node1135;
									assign node1135 = (inp[4]) ? node1139 : node1136;
										assign node1136 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
										assign node1139 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
					assign node1143 = (inp[4]) ? node1203 : node1144;
						assign node1144 = (inp[11]) ? node1174 : node1145;
							assign node1145 = (inp[5]) ? node1161 : node1146;
								assign node1146 = (inp[3]) ? node1154 : node1147;
									assign node1147 = (inp[8]) ? node1151 : node1148;
										assign node1148 = (inp[10]) ? 12'b000001111111 : 12'b000011111111;
										assign node1151 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
									assign node1154 = (inp[10]) ? node1158 : node1155;
										assign node1155 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
										assign node1158 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
								assign node1161 = (inp[9]) ? node1169 : node1162;
									assign node1162 = (inp[3]) ? node1166 : node1163;
										assign node1163 = (inp[6]) ? 12'b000000111111 : 12'b000001111111;
										assign node1166 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
									assign node1169 = (inp[6]) ? node1171 : 12'b000000011111;
										assign node1171 = (inp[10]) ? 12'b000000001111 : 12'b000000111111;
							assign node1174 = (inp[8]) ? node1188 : node1175;
								assign node1175 = (inp[9]) ? node1183 : node1176;
									assign node1176 = (inp[3]) ? node1180 : node1177;
										assign node1177 = (inp[10]) ? 12'b000000111111 : 12'b000000111111;
										assign node1180 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
									assign node1183 = (inp[3]) ? 12'b000000011111 : node1184;
										assign node1184 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
								assign node1188 = (inp[6]) ? node1196 : node1189;
									assign node1189 = (inp[5]) ? node1193 : node1190;
										assign node1190 = (inp[10]) ? 12'b000000011111 : 12'b000000111111;
										assign node1193 = (inp[3]) ? 12'b000000000111 : 12'b000000001111;
									assign node1196 = (inp[9]) ? node1200 : node1197;
										assign node1197 = (inp[10]) ? 12'b000000001111 : 12'b000000001111;
										assign node1200 = (inp[10]) ? 12'b000000001111 : 12'b000000000111;
						assign node1203 = (inp[10]) ? node1233 : node1204;
							assign node1204 = (inp[3]) ? node1218 : node1205;
								assign node1205 = (inp[8]) ? node1211 : node1206;
									assign node1206 = (inp[5]) ? node1208 : 12'b000001111111;
										assign node1208 = (inp[6]) ? 12'b000000011111 : 12'b000000011111;
									assign node1211 = (inp[9]) ? node1215 : node1212;
										assign node1212 = (inp[11]) ? 12'b000000011111 : 12'b000000011111;
										assign node1215 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
								assign node1218 = (inp[8]) ? node1226 : node1219;
									assign node1219 = (inp[9]) ? node1223 : node1220;
										assign node1220 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
										assign node1223 = (inp[5]) ? 12'b000000001111 : 12'b000000001111;
									assign node1226 = (inp[11]) ? node1230 : node1227;
										assign node1227 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
										assign node1230 = (inp[5]) ? 12'b000000000111 : 12'b000000001111;
							assign node1233 = (inp[5]) ? node1245 : node1234;
								assign node1234 = (inp[11]) ? node1242 : node1235;
									assign node1235 = (inp[8]) ? node1239 : node1236;
										assign node1236 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
										assign node1239 = (inp[6]) ? 12'b000000000111 : 12'b000000011111;
									assign node1242 = (inp[6]) ? 12'b000000000111 : 12'b000000001111;
								assign node1245 = (inp[6]) ? node1251 : node1246;
									assign node1246 = (inp[8]) ? node1248 : 12'b000000001111;
										assign node1248 = (inp[9]) ? 12'b000000000111 : 12'b000000001111;
									assign node1251 = (inp[8]) ? node1255 : node1252;
										assign node1252 = (inp[3]) ? 12'b000000000111 : 12'b000000001111;
										assign node1255 = (inp[9]) ? 12'b000000000011 : 12'b000000001111;
			assign node1258 = (inp[10]) ? node1450 : node1259;
				assign node1259 = (inp[8]) ? node1351 : node1260;
					assign node1260 = (inp[11]) ? node1304 : node1261;
						assign node1261 = (inp[5]) ? node1285 : node1262;
							assign node1262 = (inp[4]) ? node1276 : node1263;
								assign node1263 = (inp[0]) ? node1269 : node1264;
									assign node1264 = (inp[6]) ? 12'b000011111111 : node1265;
										assign node1265 = (inp[3]) ? 12'b000011111111 : 12'b000111111111;
									assign node1269 = (inp[6]) ? node1273 : node1270;
										assign node1270 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
										assign node1273 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
								assign node1276 = (inp[2]) ? node1278 : 12'b000001111111;
									assign node1278 = (inp[6]) ? node1282 : node1279;
										assign node1279 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
										assign node1282 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
							assign node1285 = (inp[0]) ? node1293 : node1286;
								assign node1286 = (inp[4]) ? 12'b000000111111 : node1287;
									assign node1287 = (inp[3]) ? 12'b000001111111 : node1288;
										assign node1288 = (inp[9]) ? 12'b000001111111 : 12'b000011111111;
								assign node1293 = (inp[6]) ? node1297 : node1294;
									assign node1294 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
									assign node1297 = (inp[2]) ? node1301 : node1298;
										assign node1298 = (inp[3]) ? 12'b000000011111 : 12'b000001111111;
										assign node1301 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
						assign node1304 = (inp[2]) ? node1332 : node1305;
							assign node1305 = (inp[0]) ? node1319 : node1306;
								assign node1306 = (inp[6]) ? node1312 : node1307;
									assign node1307 = (inp[4]) ? 12'b000000111111 : node1308;
										assign node1308 = (inp[5]) ? 12'b000001111111 : 12'b000011111111;
									assign node1312 = (inp[9]) ? node1316 : node1313;
										assign node1313 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
										assign node1316 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
								assign node1319 = (inp[4]) ? node1327 : node1320;
									assign node1320 = (inp[3]) ? node1324 : node1321;
										assign node1321 = (inp[6]) ? 12'b000000111111 : 12'b000000111111;
										assign node1324 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
									assign node1327 = (inp[3]) ? node1329 : 12'b000000011111;
										assign node1329 = (inp[9]) ? 12'b000000001111 : 12'b000000011111;
							assign node1332 = (inp[5]) ? node1338 : node1333;
								assign node1333 = (inp[0]) ? 12'b000000011111 : node1334;
									assign node1334 = (inp[4]) ? 12'b000000111111 : 12'b000001111111;
								assign node1338 = (inp[4]) ? node1344 : node1339;
									assign node1339 = (inp[3]) ? node1341 : 12'b000000111111;
										assign node1341 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
									assign node1344 = (inp[9]) ? node1348 : node1345;
										assign node1345 = (inp[0]) ? 12'b000000001111 : 12'b000000001111;
										assign node1348 = (inp[0]) ? 12'b000000000111 : 12'b000000000111;
					assign node1351 = (inp[5]) ? node1399 : node1352;
						assign node1352 = (inp[0]) ? node1372 : node1353;
							assign node1353 = (inp[3]) ? node1365 : node1354;
								assign node1354 = (inp[4]) ? node1362 : node1355;
									assign node1355 = (inp[11]) ? node1359 : node1356;
										assign node1356 = (inp[2]) ? 12'b000001111111 : 12'b000001111111;
										assign node1359 = (inp[9]) ? 12'b000000111111 : 12'b000001111111;
									assign node1362 = (inp[2]) ? 12'b000000001111 : 12'b000000111111;
								assign node1365 = (inp[11]) ? node1367 : 12'b000000111111;
									assign node1367 = (inp[6]) ? 12'b000000011111 : node1368;
										assign node1368 = (inp[4]) ? 12'b000000011111 : 12'b000000111111;
							assign node1372 = (inp[2]) ? node1386 : node1373;
								assign node1373 = (inp[4]) ? node1381 : node1374;
									assign node1374 = (inp[6]) ? node1378 : node1375;
										assign node1375 = (inp[9]) ? 12'b000000111111 : 12'b000011111111;
										assign node1378 = (inp[3]) ? 12'b000000011111 : 12'b000000111111;
									assign node1381 = (inp[11]) ? node1383 : 12'b000000011111;
										assign node1383 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
								assign node1386 = (inp[9]) ? node1392 : node1387;
									assign node1387 = (inp[3]) ? node1389 : 12'b000000011111;
										assign node1389 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
									assign node1392 = (inp[3]) ? node1396 : node1393;
										assign node1393 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
										assign node1396 = (inp[6]) ? 12'b000000000111 : 12'b000000001111;
						assign node1399 = (inp[9]) ? node1421 : node1400;
							assign node1400 = (inp[0]) ? node1414 : node1401;
								assign node1401 = (inp[6]) ? node1407 : node1402;
									assign node1402 = (inp[3]) ? node1404 : 12'b000000111111;
										assign node1404 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
									assign node1407 = (inp[3]) ? node1411 : node1408;
										assign node1408 = (inp[2]) ? 12'b000000011111 : 12'b000001111111;
										assign node1411 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
								assign node1414 = (inp[11]) ? node1416 : 12'b000000011111;
									assign node1416 = (inp[6]) ? 12'b000000001111 : node1417;
										assign node1417 = (inp[4]) ? 12'b000000001111 : 12'b000000011111;
							assign node1421 = (inp[4]) ? node1437 : node1422;
								assign node1422 = (inp[3]) ? node1430 : node1423;
									assign node1423 = (inp[6]) ? node1427 : node1424;
										assign node1424 = (inp[0]) ? 12'b000000011111 : 12'b000000111111;
										assign node1427 = (inp[2]) ? 12'b000000001111 : 12'b000000011111;
									assign node1430 = (inp[11]) ? node1434 : node1431;
										assign node1431 = (inp[6]) ? 12'b000000001111 : 12'b000000011111;
										assign node1434 = (inp[2]) ? 12'b000000000111 : 12'b000000001111;
								assign node1437 = (inp[2]) ? node1445 : node1438;
									assign node1438 = (inp[0]) ? node1442 : node1439;
										assign node1439 = (inp[6]) ? 12'b000000001111 : 12'b000000001111;
										assign node1442 = (inp[6]) ? 12'b000000000011 : 12'b000000001111;
									assign node1445 = (inp[6]) ? node1447 : 12'b000000000111;
										assign node1447 = (inp[0]) ? 12'b000000000001 : 12'b000000000111;
				assign node1450 = (inp[2]) ? node1544 : node1451;
					assign node1451 = (inp[4]) ? node1495 : node1452;
						assign node1452 = (inp[8]) ? node1470 : node1453;
							assign node1453 = (inp[3]) ? node1461 : node1454;
								assign node1454 = (inp[6]) ? 12'b000000111111 : node1455;
									assign node1455 = (inp[11]) ? 12'b000001111111 : node1456;
										assign node1456 = (inp[0]) ? 12'b000001111111 : 12'b000011111111;
								assign node1461 = (inp[9]) ? 12'b000000011111 : node1462;
									assign node1462 = (inp[0]) ? node1466 : node1463;
										assign node1463 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
										assign node1466 = (inp[11]) ? 12'b000000011111 : 12'b000000011111;
							assign node1470 = (inp[6]) ? node1482 : node1471;
								assign node1471 = (inp[0]) ? node1479 : node1472;
									assign node1472 = (inp[3]) ? node1476 : node1473;
										assign node1473 = (inp[11]) ? 12'b000000011111 : 12'b000000111111;
										assign node1476 = (inp[5]) ? 12'b000000011111 : 12'b000000011111;
									assign node1479 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
								assign node1482 = (inp[9]) ? node1488 : node1483;
									assign node1483 = (inp[0]) ? node1485 : 12'b000001111111;
										assign node1485 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
									assign node1488 = (inp[3]) ? node1492 : node1489;
										assign node1489 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
										assign node1492 = (inp[5]) ? 12'b000000000111 : 12'b000000001111;
						assign node1495 = (inp[3]) ? node1519 : node1496;
							assign node1496 = (inp[11]) ? node1508 : node1497;
								assign node1497 = (inp[0]) ? node1503 : node1498;
									assign node1498 = (inp[6]) ? node1500 : 12'b000000111111;
										assign node1500 = (inp[8]) ? 12'b000000011111 : 12'b000000011111;
									assign node1503 = (inp[5]) ? node1505 : 12'b000000111111;
										assign node1505 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
								assign node1508 = (inp[5]) ? node1516 : node1509;
									assign node1509 = (inp[0]) ? node1513 : node1510;
										assign node1510 = (inp[9]) ? 12'b000000011111 : 12'b000000111111;
										assign node1513 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
									assign node1516 = (inp[0]) ? 12'b000000011111 : 12'b000000001111;
							assign node1519 = (inp[9]) ? node1535 : node1520;
								assign node1520 = (inp[8]) ? node1528 : node1521;
									assign node1521 = (inp[11]) ? node1525 : node1522;
										assign node1522 = (inp[6]) ? 12'b000000011111 : 12'b000000111111;
										assign node1525 = (inp[0]) ? 12'b000000001111 : 12'b000000011111;
									assign node1528 = (inp[6]) ? node1532 : node1529;
										assign node1529 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
										assign node1532 = (inp[5]) ? 12'b000000000011 : 12'b000000000111;
								assign node1535 = (inp[8]) ? node1541 : node1536;
									assign node1536 = (inp[6]) ? node1538 : 12'b000000001111;
										assign node1538 = (inp[11]) ? 12'b000000000111 : 12'b000000001111;
									assign node1541 = (inp[0]) ? 12'b000000000001 : 12'b000000000111;
					assign node1544 = (inp[0]) ? node1596 : node1545;
						assign node1545 = (inp[9]) ? node1569 : node1546;
							assign node1546 = (inp[5]) ? node1558 : node1547;
								assign node1547 = (inp[6]) ? node1553 : node1548;
									assign node1548 = (inp[11]) ? 12'b000000011111 : node1549;
										assign node1549 = (inp[3]) ? 12'b000000111111 : 12'b000001111111;
									assign node1553 = (inp[3]) ? node1555 : 12'b000000111111;
										assign node1555 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
								assign node1558 = (inp[8]) ? node1564 : node1559;
									assign node1559 = (inp[6]) ? 12'b000000011111 : node1560;
										assign node1560 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
									assign node1564 = (inp[11]) ? 12'b000000001111 : node1565;
										assign node1565 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
							assign node1569 = (inp[6]) ? node1581 : node1570;
								assign node1570 = (inp[8]) ? node1576 : node1571;
									assign node1571 = (inp[3]) ? node1573 : 12'b000000111111;
										assign node1573 = (inp[11]) ? 12'b000000001111 : 12'b000000011111;
									assign node1576 = (inp[4]) ? 12'b000000001111 : node1577;
										assign node1577 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
								assign node1581 = (inp[11]) ? node1589 : node1582;
									assign node1582 = (inp[4]) ? node1586 : node1583;
										assign node1583 = (inp[3]) ? 12'b000000001111 : 12'b000000011111;
										assign node1586 = (inp[5]) ? 12'b000000000111 : 12'b000000001111;
									assign node1589 = (inp[3]) ? node1593 : node1590;
										assign node1590 = (inp[5]) ? 12'b000000000111 : 12'b000000000111;
										assign node1593 = (inp[8]) ? 12'b000000000011 : 12'b000000000111;
						assign node1596 = (inp[6]) ? node1620 : node1597;
							assign node1597 = (inp[11]) ? node1611 : node1598;
								assign node1598 = (inp[9]) ? node1606 : node1599;
									assign node1599 = (inp[3]) ? node1603 : node1600;
										assign node1600 = (inp[5]) ? 12'b000000011111 : 12'b000000111111;
										assign node1603 = (inp[8]) ? 12'b000000001111 : 12'b000000011111;
									assign node1606 = (inp[3]) ? 12'b000000001111 : node1607;
										assign node1607 = (inp[5]) ? 12'b000000001111 : 12'b000000011111;
								assign node1611 = (inp[4]) ? node1615 : node1612;
									assign node1612 = (inp[3]) ? 12'b000000000111 : 12'b000000001111;
									assign node1615 = (inp[5]) ? node1617 : 12'b000000000111;
										assign node1617 = (inp[3]) ? 12'b000000000011 : 12'b000000000111;
							assign node1620 = (inp[9]) ? node1634 : node1621;
								assign node1621 = (inp[3]) ? node1627 : node1622;
									assign node1622 = (inp[8]) ? node1624 : 12'b000000011111;
										assign node1624 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
									assign node1627 = (inp[5]) ? node1631 : node1628;
										assign node1628 = (inp[4]) ? 12'b000000000111 : 12'b000000001111;
										assign node1631 = (inp[8]) ? 12'b000000000011 : 12'b000000000111;
								assign node1634 = (inp[3]) ? node1640 : node1635;
									assign node1635 = (inp[5]) ? node1637 : 12'b000000000111;
										assign node1637 = (inp[4]) ? 12'b000000000011 : 12'b000000000111;
									assign node1640 = (inp[5]) ? node1644 : node1641;
										assign node1641 = (inp[11]) ? 12'b000000000011 : 12'b000000000011;
										assign node1644 = (inp[11]) ? 12'b000000000001 : 12'b000000000011;

endmodule