module dtc_split66_bm30 (
	input  wire [14-1:0] inp,
	output wire [8-1:0] outp
);

	wire [8-1:0] node1;
	wire [8-1:0] node2;
	wire [8-1:0] node3;
	wire [8-1:0] node4;
	wire [8-1:0] node5;
	wire [8-1:0] node6;
	wire [8-1:0] node7;
	wire [8-1:0] node9;
	wire [8-1:0] node11;
	wire [8-1:0] node14;
	wire [8-1:0] node15;
	wire [8-1:0] node17;
	wire [8-1:0] node20;
	wire [8-1:0] node22;
	wire [8-1:0] node23;
	wire [8-1:0] node26;
	wire [8-1:0] node29;
	wire [8-1:0] node30;
	wire [8-1:0] node31;
	wire [8-1:0] node33;
	wire [8-1:0] node36;
	wire [8-1:0] node38;
	wire [8-1:0] node39;
	wire [8-1:0] node42;
	wire [8-1:0] node45;
	wire [8-1:0] node46;
	wire [8-1:0] node48;
	wire [8-1:0] node49;
	wire [8-1:0] node52;
	wire [8-1:0] node55;
	wire [8-1:0] node57;
	wire [8-1:0] node58;
	wire [8-1:0] node59;
	wire [8-1:0] node62;
	wire [8-1:0] node65;
	wire [8-1:0] node66;
	wire [8-1:0] node70;
	wire [8-1:0] node71;
	wire [8-1:0] node72;
	wire [8-1:0] node73;
	wire [8-1:0] node75;
	wire [8-1:0] node78;
	wire [8-1:0] node79;
	wire [8-1:0] node81;
	wire [8-1:0] node84;
	wire [8-1:0] node86;
	wire [8-1:0] node89;
	wire [8-1:0] node90;
	wire [8-1:0] node91;
	wire [8-1:0] node93;
	wire [8-1:0] node96;
	wire [8-1:0] node97;
	wire [8-1:0] node99;
	wire [8-1:0] node102;
	wire [8-1:0] node104;
	wire [8-1:0] node107;
	wire [8-1:0] node108;
	wire [8-1:0] node110;
	wire [8-1:0] node113;
	wire [8-1:0] node114;
	wire [8-1:0] node116;
	wire [8-1:0] node119;
	wire [8-1:0] node121;
	wire [8-1:0] node125;
	wire [8-1:0] node126;
	wire [8-1:0] node127;
	wire [8-1:0] node128;
	wire [8-1:0] node131;
	wire [8-1:0] node132;
	wire [8-1:0] node133;
	wire [8-1:0] node134;
	wire [8-1:0] node138;
	wire [8-1:0] node139;
	wire [8-1:0] node143;
	wire [8-1:0] node144;
	wire [8-1:0] node145;
	wire [8-1:0] node149;
	wire [8-1:0] node150;
	wire [8-1:0] node154;
	wire [8-1:0] node155;
	wire [8-1:0] node156;
	wire [8-1:0] node157;
	wire [8-1:0] node159;
	wire [8-1:0] node162;
	wire [8-1:0] node163;
	wire [8-1:0] node167;
	wire [8-1:0] node168;
	wire [8-1:0] node169;
	wire [8-1:0] node171;
	wire [8-1:0] node174;
	wire [8-1:0] node176;
	wire [8-1:0] node179;
	wire [8-1:0] node180;
	wire [8-1:0] node181;
	wire [8-1:0] node184;
	wire [8-1:0] node188;
	wire [8-1:0] node189;
	wire [8-1:0] node190;
	wire [8-1:0] node192;
	wire [8-1:0] node195;
	wire [8-1:0] node197;
	wire [8-1:0] node198;
	wire [8-1:0] node201;
	wire [8-1:0] node204;
	wire [8-1:0] node205;
	wire [8-1:0] node207;
	wire [8-1:0] node210;
	wire [8-1:0] node211;
	wire [8-1:0] node212;
	wire [8-1:0] node215;
	wire [8-1:0] node219;
	wire [8-1:0] node220;
	wire [8-1:0] node221;
	wire [8-1:0] node222;
	wire [8-1:0] node223;
	wire [8-1:0] node225;
	wire [8-1:0] node228;
	wire [8-1:0] node230;
	wire [8-1:0] node231;
	wire [8-1:0] node234;
	wire [8-1:0] node237;
	wire [8-1:0] node238;
	wire [8-1:0] node239;
	wire [8-1:0] node243;
	wire [8-1:0] node244;
	wire [8-1:0] node245;
	wire [8-1:0] node248;
	wire [8-1:0] node252;
	wire [8-1:0] node253;
	wire [8-1:0] node254;
	wire [8-1:0] node256;
	wire [8-1:0] node257;
	wire [8-1:0] node260;
	wire [8-1:0] node263;
	wire [8-1:0] node264;
	wire [8-1:0] node265;
	wire [8-1:0] node268;
	wire [8-1:0] node272;
	wire [8-1:0] node273;
	wire [8-1:0] node275;
	wire [8-1:0] node276;
	wire [8-1:0] node277;
	wire [8-1:0] node280;
	wire [8-1:0] node283;
	wire [8-1:0] node284;
	wire [8-1:0] node287;
	wire [8-1:0] node290;
	wire [8-1:0] node291;
	wire [8-1:0] node293;
	wire [8-1:0] node294;
	wire [8-1:0] node299;
	wire [8-1:0] node300;
	wire [8-1:0] node301;
	wire [8-1:0] node302;
	wire [8-1:0] node305;
	wire [8-1:0] node306;
	wire [8-1:0] node308;
	wire [8-1:0] node311;
	wire [8-1:0] node312;
	wire [8-1:0] node315;
	wire [8-1:0] node318;
	wire [8-1:0] node319;
	wire [8-1:0] node322;
	wire [8-1:0] node323;
	wire [8-1:0] node324;
	wire [8-1:0] node327;
	wire [8-1:0] node328;
	wire [8-1:0] node332;
	wire [8-1:0] node333;
	wire [8-1:0] node334;
	wire [8-1:0] node337;
	wire [8-1:0] node340;
	wire [8-1:0] node342;
	wire [8-1:0] node345;
	wire [8-1:0] node346;
	wire [8-1:0] node347;
	wire [8-1:0] node348;
	wire [8-1:0] node352;
	wire [8-1:0] node353;
	wire [8-1:0] node354;
	wire [8-1:0] node357;
	wire [8-1:0] node361;
	wire [8-1:0] node362;
	wire [8-1:0] node363;
	wire [8-1:0] node364;
	wire [8-1:0] node367;
	wire [8-1:0] node369;
	wire [8-1:0] node372;
	wire [8-1:0] node373;
	wire [8-1:0] node376;
	wire [8-1:0] node377;
	wire [8-1:0] node380;
	wire [8-1:0] node383;
	wire [8-1:0] node386;
	wire [8-1:0] node387;
	wire [8-1:0] node388;
	wire [8-1:0] node389;
	wire [8-1:0] node390;
	wire [8-1:0] node391;
	wire [8-1:0] node392;
	wire [8-1:0] node393;
	wire [8-1:0] node394;
	wire [8-1:0] node398;
	wire [8-1:0] node399;
	wire [8-1:0] node403;
	wire [8-1:0] node404;
	wire [8-1:0] node405;
	wire [8-1:0] node407;
	wire [8-1:0] node408;
	wire [8-1:0] node411;
	wire [8-1:0] node414;
	wire [8-1:0] node415;
	wire [8-1:0] node416;
	wire [8-1:0] node419;
	wire [8-1:0] node422;
	wire [8-1:0] node423;
	wire [8-1:0] node427;
	wire [8-1:0] node428;
	wire [8-1:0] node429;
	wire [8-1:0] node430;
	wire [8-1:0] node433;
	wire [8-1:0] node436;
	wire [8-1:0] node437;
	wire [8-1:0] node440;
	wire [8-1:0] node443;
	wire [8-1:0] node445;
	wire [8-1:0] node446;
	wire [8-1:0] node449;
	wire [8-1:0] node452;
	wire [8-1:0] node453;
	wire [8-1:0] node454;
	wire [8-1:0] node455;
	wire [8-1:0] node458;
	wire [8-1:0] node459;
	wire [8-1:0] node463;
	wire [8-1:0] node464;
	wire [8-1:0] node468;
	wire [8-1:0] node469;
	wire [8-1:0] node470;
	wire [8-1:0] node472;
	wire [8-1:0] node475;
	wire [8-1:0] node476;
	wire [8-1:0] node477;
	wire [8-1:0] node481;
	wire [8-1:0] node482;
	wire [8-1:0] node485;
	wire [8-1:0] node488;
	wire [8-1:0] node489;
	wire [8-1:0] node490;
	wire [8-1:0] node494;
	wire [8-1:0] node495;
	wire [8-1:0] node498;
	wire [8-1:0] node501;
	wire [8-1:0] node502;
	wire [8-1:0] node504;
	wire [8-1:0] node506;
	wire [8-1:0] node509;
	wire [8-1:0] node510;
	wire [8-1:0] node512;
	wire [8-1:0] node515;
	wire [8-1:0] node516;
	wire [8-1:0] node518;
	wire [8-1:0] node521;
	wire [8-1:0] node523;
	wire [8-1:0] node526;
	wire [8-1:0] node527;
	wire [8-1:0] node528;
	wire [8-1:0] node529;
	wire [8-1:0] node530;
	wire [8-1:0] node531;
	wire [8-1:0] node534;
	wire [8-1:0] node538;
	wire [8-1:0] node540;
	wire [8-1:0] node543;
	wire [8-1:0] node544;
	wire [8-1:0] node545;
	wire [8-1:0] node550;
	wire [8-1:0] node551;
	wire [8-1:0] node552;
	wire [8-1:0] node553;
	wire [8-1:0] node554;
	wire [8-1:0] node556;
	wire [8-1:0] node559;
	wire [8-1:0] node560;
	wire [8-1:0] node561;
	wire [8-1:0] node564;
	wire [8-1:0] node567;
	wire [8-1:0] node568;
	wire [8-1:0] node571;
	wire [8-1:0] node574;
	wire [8-1:0] node575;
	wire [8-1:0] node576;
	wire [8-1:0] node577;
	wire [8-1:0] node581;
	wire [8-1:0] node582;
	wire [8-1:0] node585;
	wire [8-1:0] node588;
	wire [8-1:0] node589;
	wire [8-1:0] node593;
	wire [8-1:0] node594;
	wire [8-1:0] node596;
	wire [8-1:0] node599;
	wire [8-1:0] node600;
	wire [8-1:0] node602;
	wire [8-1:0] node605;
	wire [8-1:0] node606;
	wire [8-1:0] node607;
	wire [8-1:0] node612;
	wire [8-1:0] node613;
	wire [8-1:0] node614;
	wire [8-1:0] node615;
	wire [8-1:0] node616;
	wire [8-1:0] node619;
	wire [8-1:0] node622;
	wire [8-1:0] node624;
	wire [8-1:0] node627;
	wire [8-1:0] node628;
	wire [8-1:0] node629;
	wire [8-1:0] node630;
	wire [8-1:0] node633;
	wire [8-1:0] node636;
	wire [8-1:0] node637;
	wire [8-1:0] node641;
	wire [8-1:0] node642;
	wire [8-1:0] node646;
	wire [8-1:0] node647;
	wire [8-1:0] node648;
	wire [8-1:0] node649;
	wire [8-1:0] node653;
	wire [8-1:0] node654;
	wire [8-1:0] node658;
	wire [8-1:0] node660;
	wire [8-1:0] node663;
	wire [8-1:0] node664;
	wire [8-1:0] node665;
	wire [8-1:0] node666;
	wire [8-1:0] node667;
	wire [8-1:0] node668;
	wire [8-1:0] node669;
	wire [8-1:0] node672;
	wire [8-1:0] node675;
	wire [8-1:0] node676;
	wire [8-1:0] node678;
	wire [8-1:0] node680;
	wire [8-1:0] node683;
	wire [8-1:0] node684;
	wire [8-1:0] node688;
	wire [8-1:0] node689;
	wire [8-1:0] node690;
	wire [8-1:0] node692;
	wire [8-1:0] node694;
	wire [8-1:0] node697;
	wire [8-1:0] node698;
	wire [8-1:0] node702;
	wire [8-1:0] node703;
	wire [8-1:0] node705;
	wire [8-1:0] node709;
	wire [8-1:0] node710;
	wire [8-1:0] node711;
	wire [8-1:0] node712;
	wire [8-1:0] node713;
	wire [8-1:0] node715;
	wire [8-1:0] node719;
	wire [8-1:0] node720;
	wire [8-1:0] node724;
	wire [8-1:0] node725;
	wire [8-1:0] node727;
	wire [8-1:0] node729;
	wire [8-1:0] node732;
	wire [8-1:0] node734;
	wire [8-1:0] node735;
	wire [8-1:0] node739;
	wire [8-1:0] node740;
	wire [8-1:0] node741;
	wire [8-1:0] node742;
	wire [8-1:0] node745;
	wire [8-1:0] node747;
	wire [8-1:0] node750;
	wire [8-1:0] node751;
	wire [8-1:0] node755;
	wire [8-1:0] node756;
	wire [8-1:0] node757;
	wire [8-1:0] node758;
	wire [8-1:0] node761;
	wire [8-1:0] node764;
	wire [8-1:0] node767;
	wire [8-1:0] node768;
	wire [8-1:0] node771;
	wire [8-1:0] node772;
	wire [8-1:0] node776;
	wire [8-1:0] node777;
	wire [8-1:0] node778;
	wire [8-1:0] node779;
	wire [8-1:0] node780;
	wire [8-1:0] node782;
	wire [8-1:0] node785;
	wire [8-1:0] node787;
	wire [8-1:0] node789;
	wire [8-1:0] node792;
	wire [8-1:0] node794;
	wire [8-1:0] node795;
	wire [8-1:0] node798;
	wire [8-1:0] node801;
	wire [8-1:0] node802;
	wire [8-1:0] node803;
	wire [8-1:0] node805;
	wire [8-1:0] node808;
	wire [8-1:0] node811;
	wire [8-1:0] node812;
	wire [8-1:0] node815;
	wire [8-1:0] node817;
	wire [8-1:0] node820;
	wire [8-1:0] node821;
	wire [8-1:0] node822;
	wire [8-1:0] node823;
	wire [8-1:0] node824;
	wire [8-1:0] node827;
	wire [8-1:0] node830;
	wire [8-1:0] node833;
	wire [8-1:0] node834;
	wire [8-1:0] node836;
	wire [8-1:0] node839;
	wire [8-1:0] node842;
	wire [8-1:0] node843;
	wire [8-1:0] node844;
	wire [8-1:0] node847;
	wire [8-1:0] node848;
	wire [8-1:0] node851;
	wire [8-1:0] node852;
	wire [8-1:0] node856;
	wire [8-1:0] node857;
	wire [8-1:0] node858;
	wire [8-1:0] node859;
	wire [8-1:0] node862;
	wire [8-1:0] node865;
	wire [8-1:0] node866;
	wire [8-1:0] node870;
	wire [8-1:0] node871;
	wire [8-1:0] node874;
	wire [8-1:0] node875;
	wire [8-1:0] node879;
	wire [8-1:0] node880;
	wire [8-1:0] node881;
	wire [8-1:0] node882;
	wire [8-1:0] node883;
	wire [8-1:0] node884;
	wire [8-1:0] node885;
	wire [8-1:0] node889;
	wire [8-1:0] node890;
	wire [8-1:0] node894;
	wire [8-1:0] node895;
	wire [8-1:0] node899;
	wire [8-1:0] node900;
	wire [8-1:0] node901;
	wire [8-1:0] node903;
	wire [8-1:0] node906;
	wire [8-1:0] node909;
	wire [8-1:0] node910;
	wire [8-1:0] node914;
	wire [8-1:0] node915;
	wire [8-1:0] node916;
	wire [8-1:0] node917;
	wire [8-1:0] node920;
	wire [8-1:0] node921;
	wire [8-1:0] node922;
	wire [8-1:0] node925;
	wire [8-1:0] node929;
	wire [8-1:0] node930;
	wire [8-1:0] node931;
	wire [8-1:0] node932;
	wire [8-1:0] node935;
	wire [8-1:0] node938;
	wire [8-1:0] node939;
	wire [8-1:0] node943;
	wire [8-1:0] node944;
	wire [8-1:0] node947;
	wire [8-1:0] node948;
	wire [8-1:0] node952;
	wire [8-1:0] node953;
	wire [8-1:0] node954;
	wire [8-1:0] node955;
	wire [8-1:0] node956;
	wire [8-1:0] node959;
	wire [8-1:0] node962;
	wire [8-1:0] node963;
	wire [8-1:0] node967;
	wire [8-1:0] node969;
	wire [8-1:0] node972;
	wire [8-1:0] node973;
	wire [8-1:0] node975;
	wire [8-1:0] node978;
	wire [8-1:0] node981;
	wire [8-1:0] node982;
	wire [8-1:0] node983;
	wire [8-1:0] node984;
	wire [8-1:0] node985;
	wire [8-1:0] node986;
	wire [8-1:0] node987;
	wire [8-1:0] node990;
	wire [8-1:0] node993;
	wire [8-1:0] node994;
	wire [8-1:0] node998;
	wire [8-1:0] node999;
	wire [8-1:0] node1001;
	wire [8-1:0] node1004;
	wire [8-1:0] node1005;
	wire [8-1:0] node1009;
	wire [8-1:0] node1010;
	wire [8-1:0] node1011;
	wire [8-1:0] node1012;
	wire [8-1:0] node1016;
	wire [8-1:0] node1018;
	wire [8-1:0] node1021;
	wire [8-1:0] node1022;
	wire [8-1:0] node1025;
	wire [8-1:0] node1028;
	wire [8-1:0] node1029;
	wire [8-1:0] node1030;
	wire [8-1:0] node1031;
	wire [8-1:0] node1034;
	wire [8-1:0] node1037;
	wire [8-1:0] node1038;
	wire [8-1:0] node1041;
	wire [8-1:0] node1042;
	wire [8-1:0] node1046;
	wire [8-1:0] node1047;
	wire [8-1:0] node1048;
	wire [8-1:0] node1051;
	wire [8-1:0] node1054;
	wire [8-1:0] node1057;
	wire [8-1:0] node1058;
	wire [8-1:0] node1059;
	wire [8-1:0] node1060;
	wire [8-1:0] node1062;
	wire [8-1:0] node1063;
	wire [8-1:0] node1067;
	wire [8-1:0] node1069;
	wire [8-1:0] node1070;
	wire [8-1:0] node1074;
	wire [8-1:0] node1075;
	wire [8-1:0] node1076;
	wire [8-1:0] node1079;
	wire [8-1:0] node1082;
	wire [8-1:0] node1084;
	wire [8-1:0] node1087;
	wire [8-1:0] node1088;
	wire [8-1:0] node1089;
	wire [8-1:0] node1092;
	wire [8-1:0] node1095;
	wire [8-1:0] node1098;
	wire [8-1:0] node1099;
	wire [8-1:0] node1100;
	wire [8-1:0] node1101;
	wire [8-1:0] node1102;
	wire [8-1:0] node1103;
	wire [8-1:0] node1104;
	wire [8-1:0] node1105;
	wire [8-1:0] node1108;
	wire [8-1:0] node1112;
	wire [8-1:0] node1113;
	wire [8-1:0] node1115;
	wire [8-1:0] node1118;
	wire [8-1:0] node1119;
	wire [8-1:0] node1123;
	wire [8-1:0] node1124;
	wire [8-1:0] node1125;
	wire [8-1:0] node1126;
	wire [8-1:0] node1130;
	wire [8-1:0] node1133;
	wire [8-1:0] node1134;
	wire [8-1:0] node1137;
	wire [8-1:0] node1138;
	wire [8-1:0] node1140;
	wire [8-1:0] node1141;
	wire [8-1:0] node1144;
	wire [8-1:0] node1148;
	wire [8-1:0] node1149;
	wire [8-1:0] node1150;
	wire [8-1:0] node1151;
	wire [8-1:0] node1152;
	wire [8-1:0] node1155;
	wire [8-1:0] node1156;
	wire [8-1:0] node1160;
	wire [8-1:0] node1161;
	wire [8-1:0] node1163;
	wire [8-1:0] node1166;
	wire [8-1:0] node1168;
	wire [8-1:0] node1171;
	wire [8-1:0] node1172;
	wire [8-1:0] node1173;
	wire [8-1:0] node1175;
	wire [8-1:0] node1178;
	wire [8-1:0] node1180;
	wire [8-1:0] node1183;
	wire [8-1:0] node1184;
	wire [8-1:0] node1185;
	wire [8-1:0] node1189;
	wire [8-1:0] node1190;
	wire [8-1:0] node1194;
	wire [8-1:0] node1195;
	wire [8-1:0] node1196;
	wire [8-1:0] node1197;
	wire [8-1:0] node1198;
	wire [8-1:0] node1201;
	wire [8-1:0] node1204;
	wire [8-1:0] node1206;
	wire [8-1:0] node1207;
	wire [8-1:0] node1211;
	wire [8-1:0] node1212;
	wire [8-1:0] node1214;
	wire [8-1:0] node1216;
	wire [8-1:0] node1219;
	wire [8-1:0] node1220;
	wire [8-1:0] node1223;
	wire [8-1:0] node1225;
	wire [8-1:0] node1228;
	wire [8-1:0] node1229;
	wire [8-1:0] node1230;
	wire [8-1:0] node1232;
	wire [8-1:0] node1234;
	wire [8-1:0] node1237;
	wire [8-1:0] node1238;
	wire [8-1:0] node1241;
	wire [8-1:0] node1244;
	wire [8-1:0] node1245;
	wire [8-1:0] node1246;
	wire [8-1:0] node1249;
	wire [8-1:0] node1250;
	wire [8-1:0] node1254;
	wire [8-1:0] node1256;
	wire [8-1:0] node1259;
	wire [8-1:0] node1260;
	wire [8-1:0] node1261;
	wire [8-1:0] node1262;
	wire [8-1:0] node1263;
	wire [8-1:0] node1264;
	wire [8-1:0] node1268;
	wire [8-1:0] node1270;
	wire [8-1:0] node1273;
	wire [8-1:0] node1274;
	wire [8-1:0] node1275;
	wire [8-1:0] node1278;
	wire [8-1:0] node1281;
	wire [8-1:0] node1282;
	wire [8-1:0] node1283;
	wire [8-1:0] node1288;
	wire [8-1:0] node1289;
	wire [8-1:0] node1290;
	wire [8-1:0] node1291;
	wire [8-1:0] node1295;
	wire [8-1:0] node1296;
	wire [8-1:0] node1300;
	wire [8-1:0] node1301;
	wire [8-1:0] node1302;
	wire [8-1:0] node1306;
	wire [8-1:0] node1307;
	wire [8-1:0] node1309;
	wire [8-1:0] node1312;
	wire [8-1:0] node1315;
	wire [8-1:0] node1316;
	wire [8-1:0] node1317;
	wire [8-1:0] node1318;
	wire [8-1:0] node1319;
	wire [8-1:0] node1321;
	wire [8-1:0] node1324;
	wire [8-1:0] node1326;
	wire [8-1:0] node1329;
	wire [8-1:0] node1331;
	wire [8-1:0] node1333;
	wire [8-1:0] node1336;
	wire [8-1:0] node1337;
	wire [8-1:0] node1338;
	wire [8-1:0] node1339;
	wire [8-1:0] node1344;
	wire [8-1:0] node1345;
	wire [8-1:0] node1346;
	wire [8-1:0] node1347;
	wire [8-1:0] node1352;
	wire [8-1:0] node1353;
	wire [8-1:0] node1357;
	wire [8-1:0] node1358;
	wire [8-1:0] node1359;
	wire [8-1:0] node1360;
	wire [8-1:0] node1362;
	wire [8-1:0] node1365;
	wire [8-1:0] node1368;
	wire [8-1:0] node1369;
	wire [8-1:0] node1371;
	wire [8-1:0] node1372;
	wire [8-1:0] node1375;
	wire [8-1:0] node1378;
	wire [8-1:0] node1380;
	wire [8-1:0] node1381;
	wire [8-1:0] node1384;
	wire [8-1:0] node1387;
	wire [8-1:0] node1388;
	wire [8-1:0] node1389;
	wire [8-1:0] node1391;
	wire [8-1:0] node1394;
	wire [8-1:0] node1395;
	wire [8-1:0] node1397;
	wire [8-1:0] node1400;
	wire [8-1:0] node1403;
	wire [8-1:0] node1404;
	wire [8-1:0] node1406;
	wire [8-1:0] node1409;
	wire [8-1:0] node1412;
	wire [8-1:0] node1413;
	wire [8-1:0] node1414;
	wire [8-1:0] node1415;
	wire [8-1:0] node1416;
	wire [8-1:0] node1417;
	wire [8-1:0] node1419;
	wire [8-1:0] node1420;
	wire [8-1:0] node1424;
	wire [8-1:0] node1425;
	wire [8-1:0] node1429;
	wire [8-1:0] node1430;
	wire [8-1:0] node1431;
	wire [8-1:0] node1432;
	wire [8-1:0] node1436;
	wire [8-1:0] node1437;
	wire [8-1:0] node1441;
	wire [8-1:0] node1442;
	wire [8-1:0] node1446;
	wire [8-1:0] node1447;
	wire [8-1:0] node1448;
	wire [8-1:0] node1449;
	wire [8-1:0] node1453;
	wire [8-1:0] node1454;
	wire [8-1:0] node1458;
	wire [8-1:0] node1459;
	wire [8-1:0] node1463;
	wire [8-1:0] node1464;
	wire [8-1:0] node1465;
	wire [8-1:0] node1466;
	wire [8-1:0] node1467;
	wire [8-1:0] node1468;
	wire [8-1:0] node1471;
	wire [8-1:0] node1474;
	wire [8-1:0] node1475;
	wire [8-1:0] node1477;
	wire [8-1:0] node1480;
	wire [8-1:0] node1481;
	wire [8-1:0] node1485;
	wire [8-1:0] node1486;
	wire [8-1:0] node1489;
	wire [8-1:0] node1491;
	wire [8-1:0] node1494;
	wire [8-1:0] node1495;
	wire [8-1:0] node1496;
	wire [8-1:0] node1498;
	wire [8-1:0] node1501;
	wire [8-1:0] node1502;
	wire [8-1:0] node1505;
	wire [8-1:0] node1507;
	wire [8-1:0] node1510;
	wire [8-1:0] node1511;
	wire [8-1:0] node1512;
	wire [8-1:0] node1515;
	wire [8-1:0] node1518;
	wire [8-1:0] node1519;
	wire [8-1:0] node1522;
	wire [8-1:0] node1525;
	wire [8-1:0] node1526;
	wire [8-1:0] node1527;
	wire [8-1:0] node1528;
	wire [8-1:0] node1529;
	wire [8-1:0] node1532;
	wire [8-1:0] node1535;
	wire [8-1:0] node1536;
	wire [8-1:0] node1539;
	wire [8-1:0] node1542;
	wire [8-1:0] node1543;
	wire [8-1:0] node1544;
	wire [8-1:0] node1547;
	wire [8-1:0] node1550;
	wire [8-1:0] node1551;
	wire [8-1:0] node1554;
	wire [8-1:0] node1557;
	wire [8-1:0] node1558;
	wire [8-1:0] node1559;
	wire [8-1:0] node1561;
	wire [8-1:0] node1564;
	wire [8-1:0] node1565;
	wire [8-1:0] node1569;
	wire [8-1:0] node1570;
	wire [8-1:0] node1572;
	wire [8-1:0] node1573;
	wire [8-1:0] node1576;
	wire [8-1:0] node1579;
	wire [8-1:0] node1580;
	wire [8-1:0] node1583;
	wire [8-1:0] node1584;
	wire [8-1:0] node1587;
	wire [8-1:0] node1590;
	wire [8-1:0] node1591;
	wire [8-1:0] node1592;
	wire [8-1:0] node1593;
	wire [8-1:0] node1594;
	wire [8-1:0] node1596;
	wire [8-1:0] node1598;
	wire [8-1:0] node1601;
	wire [8-1:0] node1603;
	wire [8-1:0] node1606;
	wire [8-1:0] node1607;
	wire [8-1:0] node1608;
	wire [8-1:0] node1611;
	wire [8-1:0] node1614;
	wire [8-1:0] node1615;
	wire [8-1:0] node1618;
	wire [8-1:0] node1621;
	wire [8-1:0] node1622;
	wire [8-1:0] node1623;
	wire [8-1:0] node1624;
	wire [8-1:0] node1628;
	wire [8-1:0] node1629;
	wire [8-1:0] node1632;
	wire [8-1:0] node1635;
	wire [8-1:0] node1636;
	wire [8-1:0] node1637;
	wire [8-1:0] node1640;
	wire [8-1:0] node1643;
	wire [8-1:0] node1644;
	wire [8-1:0] node1648;
	wire [8-1:0] node1649;
	wire [8-1:0] node1650;
	wire [8-1:0] node1651;
	wire [8-1:0] node1652;
	wire [8-1:0] node1654;
	wire [8-1:0] node1655;
	wire [8-1:0] node1658;
	wire [8-1:0] node1661;
	wire [8-1:0] node1662;
	wire [8-1:0] node1664;
	wire [8-1:0] node1668;
	wire [8-1:0] node1669;
	wire [8-1:0] node1670;
	wire [8-1:0] node1673;
	wire [8-1:0] node1676;
	wire [8-1:0] node1679;
	wire [8-1:0] node1680;
	wire [8-1:0] node1681;
	wire [8-1:0] node1682;
	wire [8-1:0] node1686;
	wire [8-1:0] node1687;
	wire [8-1:0] node1689;
	wire [8-1:0] node1693;
	wire [8-1:0] node1694;
	wire [8-1:0] node1695;
	wire [8-1:0] node1697;
	wire [8-1:0] node1700;
	wire [8-1:0] node1701;
	wire [8-1:0] node1705;
	wire [8-1:0] node1708;
	wire [8-1:0] node1709;
	wire [8-1:0] node1710;
	wire [8-1:0] node1711;
	wire [8-1:0] node1712;
	wire [8-1:0] node1713;
	wire [8-1:0] node1718;
	wire [8-1:0] node1719;
	wire [8-1:0] node1720;
	wire [8-1:0] node1724;
	wire [8-1:0] node1725;
	wire [8-1:0] node1729;
	wire [8-1:0] node1730;
	wire [8-1:0] node1731;
	wire [8-1:0] node1734;
	wire [8-1:0] node1735;
	wire [8-1:0] node1739;
	wire [8-1:0] node1740;
	wire [8-1:0] node1741;
	wire [8-1:0] node1745;
	wire [8-1:0] node1746;
	wire [8-1:0] node1750;
	wire [8-1:0] node1751;
	wire [8-1:0] node1752;
	wire [8-1:0] node1755;
	wire [8-1:0] node1756;
	wire [8-1:0] node1759;
	wire [8-1:0] node1762;
	wire [8-1:0] node1765;
	wire [8-1:0] node1766;
	wire [8-1:0] node1767;
	wire [8-1:0] node1768;
	wire [8-1:0] node1769;
	wire [8-1:0] node1770;
	wire [8-1:0] node1771;
	wire [8-1:0] node1772;
	wire [8-1:0] node1776;
	wire [8-1:0] node1778;
	wire [8-1:0] node1781;
	wire [8-1:0] node1782;
	wire [8-1:0] node1784;
	wire [8-1:0] node1787;
	wire [8-1:0] node1789;
	wire [8-1:0] node1792;
	wire [8-1:0] node1793;
	wire [8-1:0] node1794;
	wire [8-1:0] node1795;
	wire [8-1:0] node1796;
	wire [8-1:0] node1797;
	wire [8-1:0] node1798;
	wire [8-1:0] node1802;
	wire [8-1:0] node1803;
	wire [8-1:0] node1807;
	wire [8-1:0] node1808;
	wire [8-1:0] node1812;
	wire [8-1:0] node1813;
	wire [8-1:0] node1814;
	wire [8-1:0] node1815;
	wire [8-1:0] node1819;
	wire [8-1:0] node1820;
	wire [8-1:0] node1825;
	wire [8-1:0] node1826;
	wire [8-1:0] node1827;
	wire [8-1:0] node1828;
	wire [8-1:0] node1832;
	wire [8-1:0] node1833;
	wire [8-1:0] node1837;
	wire [8-1:0] node1838;
	wire [8-1:0] node1842;
	wire [8-1:0] node1843;
	wire [8-1:0] node1844;
	wire [8-1:0] node1845;
	wire [8-1:0] node1846;
	wire [8-1:0] node1847;
	wire [8-1:0] node1851;
	wire [8-1:0] node1852;
	wire [8-1:0] node1856;
	wire [8-1:0] node1857;
	wire [8-1:0] node1861;
	wire [8-1:0] node1862;
	wire [8-1:0] node1863;
	wire [8-1:0] node1864;
	wire [8-1:0] node1868;
	wire [8-1:0] node1871;
	wire [8-1:0] node1872;
	wire [8-1:0] node1876;
	wire [8-1:0] node1877;
	wire [8-1:0] node1878;
	wire [8-1:0] node1879;
	wire [8-1:0] node1880;
	wire [8-1:0] node1885;
	wire [8-1:0] node1886;
	wire [8-1:0] node1890;
	wire [8-1:0] node1891;
	wire [8-1:0] node1895;
	wire [8-1:0] node1896;
	wire [8-1:0] node1897;
	wire [8-1:0] node1898;
	wire [8-1:0] node1900;
	wire [8-1:0] node1903;
	wire [8-1:0] node1904;
	wire [8-1:0] node1908;
	wire [8-1:0] node1909;
	wire [8-1:0] node1910;
	wire [8-1:0] node1911;
	wire [8-1:0] node1915;
	wire [8-1:0] node1916;
	wire [8-1:0] node1917;
	wire [8-1:0] node1921;
	wire [8-1:0] node1922;
	wire [8-1:0] node1926;
	wire [8-1:0] node1927;
	wire [8-1:0] node1928;
	wire [8-1:0] node1929;
	wire [8-1:0] node1933;
	wire [8-1:0] node1934;
	wire [8-1:0] node1938;
	wire [8-1:0] node1939;
	wire [8-1:0] node1943;
	wire [8-1:0] node1944;
	wire [8-1:0] node1945;
	wire [8-1:0] node1946;
	wire [8-1:0] node1950;
	wire [8-1:0] node1951;
	wire [8-1:0] node1953;
	wire [8-1:0] node1956;
	wire [8-1:0] node1957;
	wire [8-1:0] node1961;
	wire [8-1:0] node1962;
	wire [8-1:0] node1966;
	wire [8-1:0] node1967;
	wire [8-1:0] node1968;
	wire [8-1:0] node1969;
	wire [8-1:0] node1970;
	wire [8-1:0] node1971;
	wire [8-1:0] node1973;
	wire [8-1:0] node1975;
	wire [8-1:0] node1978;
	wire [8-1:0] node1979;
	wire [8-1:0] node1982;
	wire [8-1:0] node1984;
	wire [8-1:0] node1987;
	wire [8-1:0] node1988;
	wire [8-1:0] node1989;
	wire [8-1:0] node1991;
	wire [8-1:0] node1993;
	wire [8-1:0] node1996;
	wire [8-1:0] node1998;
	wire [8-1:0] node2001;
	wire [8-1:0] node2002;
	wire [8-1:0] node2003;
	wire [8-1:0] node2006;
	wire [8-1:0] node2008;
	wire [8-1:0] node2011;
	wire [8-1:0] node2014;
	wire [8-1:0] node2015;
	wire [8-1:0] node2016;
	wire [8-1:0] node2017;
	wire [8-1:0] node2019;
	wire [8-1:0] node2021;
	wire [8-1:0] node2024;
	wire [8-1:0] node2027;
	wire [8-1:0] node2028;
	wire [8-1:0] node2029;
	wire [8-1:0] node2032;
	wire [8-1:0] node2034;
	wire [8-1:0] node2037;
	wire [8-1:0] node2040;
	wire [8-1:0] node2041;
	wire [8-1:0] node2042;
	wire [8-1:0] node2043;
	wire [8-1:0] node2045;
	wire [8-1:0] node2048;
	wire [8-1:0] node2050;
	wire [8-1:0] node2053;
	wire [8-1:0] node2054;
	wire [8-1:0] node2056;
	wire [8-1:0] node2059;
	wire [8-1:0] node2060;
	wire [8-1:0] node2064;
	wire [8-1:0] node2065;
	wire [8-1:0] node2069;
	wire [8-1:0] node2070;
	wire [8-1:0] node2071;
	wire [8-1:0] node2072;
	wire [8-1:0] node2073;
	wire [8-1:0] node2076;
	wire [8-1:0] node2077;
	wire [8-1:0] node2080;
	wire [8-1:0] node2083;
	wire [8-1:0] node2084;
	wire [8-1:0] node2085;
	wire [8-1:0] node2087;
	wire [8-1:0] node2089;
	wire [8-1:0] node2092;
	wire [8-1:0] node2093;
	wire [8-1:0] node2096;
	wire [8-1:0] node2098;
	wire [8-1:0] node2101;
	wire [8-1:0] node2102;
	wire [8-1:0] node2104;
	wire [8-1:0] node2105;
	wire [8-1:0] node2108;
	wire [8-1:0] node2111;
	wire [8-1:0] node2113;
	wire [8-1:0] node2114;
	wire [8-1:0] node2117;
	wire [8-1:0] node2120;
	wire [8-1:0] node2121;
	wire [8-1:0] node2122;
	wire [8-1:0] node2123;
	wire [8-1:0] node2124;
	wire [8-1:0] node2128;
	wire [8-1:0] node2130;
	wire [8-1:0] node2133;
	wire [8-1:0] node2134;
	wire [8-1:0] node2136;
	wire [8-1:0] node2139;
	wire [8-1:0] node2140;
	wire [8-1:0] node2143;
	wire [8-1:0] node2146;
	wire [8-1:0] node2147;
	wire [8-1:0] node2148;
	wire [8-1:0] node2149;
	wire [8-1:0] node2153;
	wire [8-1:0] node2154;
	wire [8-1:0] node2155;
	wire [8-1:0] node2158;
	wire [8-1:0] node2161;
	wire [8-1:0] node2164;
	wire [8-1:0] node2165;
	wire [8-1:0] node2166;
	wire [8-1:0] node2167;
	wire [8-1:0] node2171;
	wire [8-1:0] node2172;
	wire [8-1:0] node2176;
	wire [8-1:0] node2177;
	wire [8-1:0] node2180;
	wire [8-1:0] node2183;
	wire [8-1:0] node2184;
	wire [8-1:0] node2185;
	wire [8-1:0] node2186;
	wire [8-1:0] node2187;
	wire [8-1:0] node2188;
	wire [8-1:0] node2190;
	wire [8-1:0] node2193;
	wire [8-1:0] node2195;
	wire [8-1:0] node2198;
	wire [8-1:0] node2200;
	wire [8-1:0] node2203;
	wire [8-1:0] node2204;
	wire [8-1:0] node2205;
	wire [8-1:0] node2208;
	wire [8-1:0] node2209;
	wire [8-1:0] node2213;
	wire [8-1:0] node2214;
	wire [8-1:0] node2215;
	wire [8-1:0] node2220;
	wire [8-1:0] node2221;
	wire [8-1:0] node2222;
	wire [8-1:0] node2223;
	wire [8-1:0] node2226;
	wire [8-1:0] node2229;
	wire [8-1:0] node2232;
	wire [8-1:0] node2233;
	wire [8-1:0] node2234;
	wire [8-1:0] node2237;
	wire [8-1:0] node2240;
	wire [8-1:0] node2241;
	wire [8-1:0] node2244;
	wire [8-1:0] node2247;
	wire [8-1:0] node2248;
	wire [8-1:0] node2249;
	wire [8-1:0] node2250;
	wire [8-1:0] node2251;
	wire [8-1:0] node2253;
	wire [8-1:0] node2256;
	wire [8-1:0] node2259;
	wire [8-1:0] node2260;
	wire [8-1:0] node2261;
	wire [8-1:0] node2266;
	wire [8-1:0] node2267;
	wire [8-1:0] node2269;
	wire [8-1:0] node2270;
	wire [8-1:0] node2273;
	wire [8-1:0] node2276;
	wire [8-1:0] node2277;
	wire [8-1:0] node2278;
	wire [8-1:0] node2282;
	wire [8-1:0] node2283;
	wire [8-1:0] node2287;
	wire [8-1:0] node2288;
	wire [8-1:0] node2289;
	wire [8-1:0] node2292;
	wire [8-1:0] node2294;
	wire [8-1:0] node2297;
	wire [8-1:0] node2298;
	wire [8-1:0] node2299;
	wire [8-1:0] node2303;
	wire [8-1:0] node2304;
	wire [8-1:0] node2307;
	wire [8-1:0] node2310;
	wire [8-1:0] node2311;
	wire [8-1:0] node2312;
	wire [8-1:0] node2313;
	wire [8-1:0] node2314;
	wire [8-1:0] node2315;
	wire [8-1:0] node2319;
	wire [8-1:0] node2320;
	wire [8-1:0] node2323;
	wire [8-1:0] node2324;
	wire [8-1:0] node2327;
	wire [8-1:0] node2330;
	wire [8-1:0] node2331;
	wire [8-1:0] node2332;
	wire [8-1:0] node2334;
	wire [8-1:0] node2337;
	wire [8-1:0] node2339;
	wire [8-1:0] node2342;
	wire [8-1:0] node2343;
	wire [8-1:0] node2344;
	wire [8-1:0] node2347;
	wire [8-1:0] node2348;
	wire [8-1:0] node2350;
	wire [8-1:0] node2353;
	wire [8-1:0] node2356;
	wire [8-1:0] node2357;
	wire [8-1:0] node2360;
	wire [8-1:0] node2361;
	wire [8-1:0] node2364;
	wire [8-1:0] node2367;
	wire [8-1:0] node2368;
	wire [8-1:0] node2369;
	wire [8-1:0] node2370;
	wire [8-1:0] node2373;
	wire [8-1:0] node2376;
	wire [8-1:0] node2377;
	wire [8-1:0] node2378;
	wire [8-1:0] node2379;
	wire [8-1:0] node2382;
	wire [8-1:0] node2385;
	wire [8-1:0] node2386;
	wire [8-1:0] node2390;
	wire [8-1:0] node2391;
	wire [8-1:0] node2392;
	wire [8-1:0] node2393;
	wire [8-1:0] node2398;
	wire [8-1:0] node2399;
	wire [8-1:0] node2400;
	wire [8-1:0] node2404;
	wire [8-1:0] node2407;
	wire [8-1:0] node2408;
	wire [8-1:0] node2409;
	wire [8-1:0] node2410;
	wire [8-1:0] node2412;
	wire [8-1:0] node2413;
	wire [8-1:0] node2417;
	wire [8-1:0] node2419;
	wire [8-1:0] node2422;
	wire [8-1:0] node2423;
	wire [8-1:0] node2424;
	wire [8-1:0] node2428;
	wire [8-1:0] node2429;
	wire [8-1:0] node2432;
	wire [8-1:0] node2433;
	wire [8-1:0] node2437;
	wire [8-1:0] node2438;
	wire [8-1:0] node2439;
	wire [8-1:0] node2441;
	wire [8-1:0] node2444;
	wire [8-1:0] node2447;
	wire [8-1:0] node2448;
	wire [8-1:0] node2450;
	wire [8-1:0] node2453;
	wire [8-1:0] node2454;
	wire [8-1:0] node2455;
	wire [8-1:0] node2459;
	wire [8-1:0] node2460;
	wire [8-1:0] node2463;
	wire [8-1:0] node2466;
	wire [8-1:0] node2467;
	wire [8-1:0] node2468;
	wire [8-1:0] node2469;
	wire [8-1:0] node2470;
	wire [8-1:0] node2472;
	wire [8-1:0] node2475;
	wire [8-1:0] node2476;
	wire [8-1:0] node2478;
	wire [8-1:0] node2481;
	wire [8-1:0] node2484;
	wire [8-1:0] node2485;
	wire [8-1:0] node2487;
	wire [8-1:0] node2490;
	wire [8-1:0] node2491;
	wire [8-1:0] node2495;
	wire [8-1:0] node2496;
	wire [8-1:0] node2497;
	wire [8-1:0] node2498;
	wire [8-1:0] node2501;
	wire [8-1:0] node2502;
	wire [8-1:0] node2505;
	wire [8-1:0] node2508;
	wire [8-1:0] node2509;
	wire [8-1:0] node2510;
	wire [8-1:0] node2511;
	wire [8-1:0] node2516;
	wire [8-1:0] node2518;
	wire [8-1:0] node2520;
	wire [8-1:0] node2523;
	wire [8-1:0] node2524;
	wire [8-1:0] node2525;
	wire [8-1:0] node2526;
	wire [8-1:0] node2529;
	wire [8-1:0] node2531;
	wire [8-1:0] node2534;
	wire [8-1:0] node2537;
	wire [8-1:0] node2538;
	wire [8-1:0] node2539;
	wire [8-1:0] node2542;
	wire [8-1:0] node2545;
	wire [8-1:0] node2546;
	wire [8-1:0] node2549;
	wire [8-1:0] node2552;
	wire [8-1:0] node2553;
	wire [8-1:0] node2554;
	wire [8-1:0] node2555;
	wire [8-1:0] node2556;
	wire [8-1:0] node2558;
	wire [8-1:0] node2561;
	wire [8-1:0] node2564;
	wire [8-1:0] node2565;
	wire [8-1:0] node2567;
	wire [8-1:0] node2570;
	wire [8-1:0] node2571;
	wire [8-1:0] node2574;
	wire [8-1:0] node2576;
	wire [8-1:0] node2579;
	wire [8-1:0] node2580;
	wire [8-1:0] node2581;
	wire [8-1:0] node2583;
	wire [8-1:0] node2586;
	wire [8-1:0] node2587;
	wire [8-1:0] node2589;
	wire [8-1:0] node2593;
	wire [8-1:0] node2594;
	wire [8-1:0] node2596;
	wire [8-1:0] node2599;
	wire [8-1:0] node2600;
	wire [8-1:0] node2604;
	wire [8-1:0] node2605;
	wire [8-1:0] node2606;
	wire [8-1:0] node2607;
	wire [8-1:0] node2609;
	wire [8-1:0] node2612;
	wire [8-1:0] node2615;
	wire [8-1:0] node2616;
	wire [8-1:0] node2617;
	wire [8-1:0] node2619;
	wire [8-1:0] node2623;
	wire [8-1:0] node2624;
	wire [8-1:0] node2625;
	wire [8-1:0] node2630;
	wire [8-1:0] node2631;
	wire [8-1:0] node2632;
	wire [8-1:0] node2634;
	wire [8-1:0] node2637;
	wire [8-1:0] node2638;
	wire [8-1:0] node2641;
	wire [8-1:0] node2644;
	wire [8-1:0] node2645;
	wire [8-1:0] node2647;
	wire [8-1:0] node2650;
	wire [8-1:0] node2653;
	wire [8-1:0] node2654;
	wire [8-1:0] node2655;
	wire [8-1:0] node2656;
	wire [8-1:0] node2657;
	wire [8-1:0] node2658;
	wire [8-1:0] node2659;
	wire [8-1:0] node2661;
	wire [8-1:0] node2664;
	wire [8-1:0] node2665;
	wire [8-1:0] node2667;
	wire [8-1:0] node2670;
	wire [8-1:0] node2672;
	wire [8-1:0] node2675;
	wire [8-1:0] node2676;
	wire [8-1:0] node2677;
	wire [8-1:0] node2678;
	wire [8-1:0] node2679;
	wire [8-1:0] node2682;
	wire [8-1:0] node2685;
	wire [8-1:0] node2686;
	wire [8-1:0] node2689;
	wire [8-1:0] node2692;
	wire [8-1:0] node2693;
	wire [8-1:0] node2694;
	wire [8-1:0] node2698;
	wire [8-1:0] node2699;
	wire [8-1:0] node2703;
	wire [8-1:0] node2704;
	wire [8-1:0] node2705;
	wire [8-1:0] node2707;
	wire [8-1:0] node2710;
	wire [8-1:0] node2712;
	wire [8-1:0] node2713;
	wire [8-1:0] node2717;
	wire [8-1:0] node2718;
	wire [8-1:0] node2719;
	wire [8-1:0] node2722;
	wire [8-1:0] node2723;
	wire [8-1:0] node2727;
	wire [8-1:0] node2728;
	wire [8-1:0] node2731;
	wire [8-1:0] node2734;
	wire [8-1:0] node2735;
	wire [8-1:0] node2736;
	wire [8-1:0] node2737;
	wire [8-1:0] node2739;
	wire [8-1:0] node2742;
	wire [8-1:0] node2743;
	wire [8-1:0] node2744;
	wire [8-1:0] node2746;
	wire [8-1:0] node2750;
	wire [8-1:0] node2752;
	wire [8-1:0] node2755;
	wire [8-1:0] node2756;
	wire [8-1:0] node2757;
	wire [8-1:0] node2759;
	wire [8-1:0] node2763;
	wire [8-1:0] node2764;
	wire [8-1:0] node2766;
	wire [8-1:0] node2769;
	wire [8-1:0] node2772;
	wire [8-1:0] node2773;
	wire [8-1:0] node2774;
	wire [8-1:0] node2775;
	wire [8-1:0] node2777;
	wire [8-1:0] node2780;
	wire [8-1:0] node2783;
	wire [8-1:0] node2784;
	wire [8-1:0] node2787;
	wire [8-1:0] node2788;
	wire [8-1:0] node2792;
	wire [8-1:0] node2793;
	wire [8-1:0] node2795;
	wire [8-1:0] node2796;
	wire [8-1:0] node2799;
	wire [8-1:0] node2802;
	wire [8-1:0] node2803;
	wire [8-1:0] node2805;
	wire [8-1:0] node2808;
	wire [8-1:0] node2811;
	wire [8-1:0] node2812;
	wire [8-1:0] node2813;
	wire [8-1:0] node2814;
	wire [8-1:0] node2816;
	wire [8-1:0] node2819;
	wire [8-1:0] node2820;
	wire [8-1:0] node2823;
	wire [8-1:0] node2825;
	wire [8-1:0] node2828;
	wire [8-1:0] node2829;
	wire [8-1:0] node2830;
	wire [8-1:0] node2831;
	wire [8-1:0] node2835;
	wire [8-1:0] node2836;
	wire [8-1:0] node2839;
	wire [8-1:0] node2840;
	wire [8-1:0] node2844;
	wire [8-1:0] node2845;
	wire [8-1:0] node2847;
	wire [8-1:0] node2848;
	wire [8-1:0] node2852;
	wire [8-1:0] node2853;
	wire [8-1:0] node2856;
	wire [8-1:0] node2857;
	wire [8-1:0] node2860;
	wire [8-1:0] node2863;
	wire [8-1:0] node2864;
	wire [8-1:0] node2865;
	wire [8-1:0] node2866;
	wire [8-1:0] node2867;
	wire [8-1:0] node2868;
	wire [8-1:0] node2870;
	wire [8-1:0] node2873;
	wire [8-1:0] node2874;
	wire [8-1:0] node2878;
	wire [8-1:0] node2880;
	wire [8-1:0] node2882;
	wire [8-1:0] node2885;
	wire [8-1:0] node2886;
	wire [8-1:0] node2887;
	wire [8-1:0] node2889;
	wire [8-1:0] node2892;
	wire [8-1:0] node2893;
	wire [8-1:0] node2896;
	wire [8-1:0] node2899;
	wire [8-1:0] node2900;
	wire [8-1:0] node2903;
	wire [8-1:0] node2906;
	wire [8-1:0] node2907;
	wire [8-1:0] node2908;
	wire [8-1:0] node2909;
	wire [8-1:0] node2913;
	wire [8-1:0] node2915;
	wire [8-1:0] node2918;
	wire [8-1:0] node2919;
	wire [8-1:0] node2921;
	wire [8-1:0] node2922;
	wire [8-1:0] node2925;
	wire [8-1:0] node2928;
	wire [8-1:0] node2930;
	wire [8-1:0] node2933;
	wire [8-1:0] node2934;
	wire [8-1:0] node2935;
	wire [8-1:0] node2936;
	wire [8-1:0] node2938;
	wire [8-1:0] node2939;
	wire [8-1:0] node2942;
	wire [8-1:0] node2945;
	wire [8-1:0] node2946;
	wire [8-1:0] node2949;
	wire [8-1:0] node2952;
	wire [8-1:0] node2953;
	wire [8-1:0] node2954;
	wire [8-1:0] node2956;
	wire [8-1:0] node2959;
	wire [8-1:0] node2961;
	wire [8-1:0] node2964;
	wire [8-1:0] node2965;
	wire [8-1:0] node2968;
	wire [8-1:0] node2971;
	wire [8-1:0] node2972;
	wire [8-1:0] node2973;
	wire [8-1:0] node2975;
	wire [8-1:0] node2979;
	wire [8-1:0] node2980;
	wire [8-1:0] node2981;
	wire [8-1:0] node2984;
	wire [8-1:0] node2987;
	wire [8-1:0] node2989;
	wire [8-1:0] node2992;
	wire [8-1:0] node2993;
	wire [8-1:0] node2995;
	wire [8-1:0] node2997;
	wire [8-1:0] node3000;
	wire [8-1:0] node3001;
	wire [8-1:0] node3002;
	wire [8-1:0] node3003;
	wire [8-1:0] node3004;
	wire [8-1:0] node3006;
	wire [8-1:0] node3009;
	wire [8-1:0] node3010;
	wire [8-1:0] node3014;
	wire [8-1:0] node3015;
	wire [8-1:0] node3019;
	wire [8-1:0] node3020;
	wire [8-1:0] node3021;
	wire [8-1:0] node3022;
	wire [8-1:0] node3026;
	wire [8-1:0] node3027;
	wire [8-1:0] node3030;
	wire [8-1:0] node3033;
	wire [8-1:0] node3034;
	wire [8-1:0] node3035;
	wire [8-1:0] node3038;
	wire [8-1:0] node3041;
	wire [8-1:0] node3042;
	wire [8-1:0] node3045;
	wire [8-1:0] node3048;
	wire [8-1:0] node3049;
	wire [8-1:0] node3050;
	wire [8-1:0] node3052;
	wire [8-1:0] node3055;
	wire [8-1:0] node3056;
	wire [8-1:0] node3059;
	wire [8-1:0] node3062;
	wire [8-1:0] node3063;
	wire [8-1:0] node3064;
	wire [8-1:0] node3068;
	wire [8-1:0] node3069;
	wire [8-1:0] node3073;
	wire [8-1:0] node3074;
	wire [8-1:0] node3075;
	wire [8-1:0] node3076;
	wire [8-1:0] node3077;
	wire [8-1:0] node3078;
	wire [8-1:0] node3079;
	wire [8-1:0] node3081;
	wire [8-1:0] node3084;
	wire [8-1:0] node3086;
	wire [8-1:0] node3089;
	wire [8-1:0] node3090;
	wire [8-1:0] node3091;
	wire [8-1:0] node3092;
	wire [8-1:0] node3093;
	wire [8-1:0] node3097;
	wire [8-1:0] node3098;
	wire [8-1:0] node3102;
	wire [8-1:0] node3103;
	wire [8-1:0] node3104;
	wire [8-1:0] node3107;
	wire [8-1:0] node3110;
	wire [8-1:0] node3111;
	wire [8-1:0] node3114;
	wire [8-1:0] node3117;
	wire [8-1:0] node3118;
	wire [8-1:0] node3119;
	wire [8-1:0] node3121;
	wire [8-1:0] node3124;
	wire [8-1:0] node3126;
	wire [8-1:0] node3129;
	wire [8-1:0] node3130;
	wire [8-1:0] node3132;
	wire [8-1:0] node3135;
	wire [8-1:0] node3136;
	wire [8-1:0] node3139;
	wire [8-1:0] node3142;
	wire [8-1:0] node3143;
	wire [8-1:0] node3144;
	wire [8-1:0] node3145;
	wire [8-1:0] node3146;
	wire [8-1:0] node3149;
	wire [8-1:0] node3151;
	wire [8-1:0] node3154;
	wire [8-1:0] node3155;
	wire [8-1:0] node3158;
	wire [8-1:0] node3160;
	wire [8-1:0] node3163;
	wire [8-1:0] node3164;
	wire [8-1:0] node3165;
	wire [8-1:0] node3169;
	wire [8-1:0] node3171;
	wire [8-1:0] node3173;
	wire [8-1:0] node3176;
	wire [8-1:0] node3177;
	wire [8-1:0] node3178;
	wire [8-1:0] node3181;
	wire [8-1:0] node3182;
	wire [8-1:0] node3183;
	wire [8-1:0] node3187;
	wire [8-1:0] node3188;
	wire [8-1:0] node3192;
	wire [8-1:0] node3193;
	wire [8-1:0] node3194;
	wire [8-1:0] node3197;
	wire [8-1:0] node3199;
	wire [8-1:0] node3202;
	wire [8-1:0] node3203;
	wire [8-1:0] node3206;
	wire [8-1:0] node3209;
	wire [8-1:0] node3210;
	wire [8-1:0] node3211;
	wire [8-1:0] node3212;
	wire [8-1:0] node3214;
	wire [8-1:0] node3217;
	wire [8-1:0] node3219;
	wire [8-1:0] node3222;
	wire [8-1:0] node3223;
	wire [8-1:0] node3224;
	wire [8-1:0] node3225;
	wire [8-1:0] node3228;
	wire [8-1:0] node3229;
	wire [8-1:0] node3233;
	wire [8-1:0] node3234;
	wire [8-1:0] node3235;
	wire [8-1:0] node3238;
	wire [8-1:0] node3241;
	wire [8-1:0] node3242;
	wire [8-1:0] node3245;
	wire [8-1:0] node3248;
	wire [8-1:0] node3249;
	wire [8-1:0] node3251;
	wire [8-1:0] node3254;
	wire [8-1:0] node3255;
	wire [8-1:0] node3257;
	wire [8-1:0] node3260;
	wire [8-1:0] node3261;
	wire [8-1:0] node3265;
	wire [8-1:0] node3266;
	wire [8-1:0] node3267;
	wire [8-1:0] node3268;
	wire [8-1:0] node3269;
	wire [8-1:0] node3272;
	wire [8-1:0] node3274;
	wire [8-1:0] node3277;
	wire [8-1:0] node3278;
	wire [8-1:0] node3280;
	wire [8-1:0] node3283;
	wire [8-1:0] node3285;
	wire [8-1:0] node3288;
	wire [8-1:0] node3289;
	wire [8-1:0] node3291;
	wire [8-1:0] node3294;
	wire [8-1:0] node3295;
	wire [8-1:0] node3298;
	wire [8-1:0] node3299;
	wire [8-1:0] node3302;
	wire [8-1:0] node3305;
	wire [8-1:0] node3306;
	wire [8-1:0] node3307;
	wire [8-1:0] node3309;
	wire [8-1:0] node3312;
	wire [8-1:0] node3314;
	wire [8-1:0] node3316;
	wire [8-1:0] node3319;
	wire [8-1:0] node3320;
	wire [8-1:0] node3321;
	wire [8-1:0] node3324;
	wire [8-1:0] node3327;
	wire [8-1:0] node3328;
	wire [8-1:0] node3332;
	wire [8-1:0] node3333;
	wire [8-1:0] node3334;
	wire [8-1:0] node3335;
	wire [8-1:0] node3338;
	wire [8-1:0] node3339;
	wire [8-1:0] node3340;
	wire [8-1:0] node3341;
	wire [8-1:0] node3344;
	wire [8-1:0] node3347;
	wire [8-1:0] node3348;
	wire [8-1:0] node3351;
	wire [8-1:0] node3354;
	wire [8-1:0] node3355;
	wire [8-1:0] node3357;
	wire [8-1:0] node3360;
	wire [8-1:0] node3361;
	wire [8-1:0] node3364;
	wire [8-1:0] node3367;
	wire [8-1:0] node3368;
	wire [8-1:0] node3371;
	wire [8-1:0] node3372;
	wire [8-1:0] node3373;
	wire [8-1:0] node3376;
	wire [8-1:0] node3379;
	wire [8-1:0] node3380;
	wire [8-1:0] node3383;
	wire [8-1:0] node3386;
	wire [8-1:0] node3387;
	wire [8-1:0] node3388;
	wire [8-1:0] node3391;
	wire [8-1:0] node3392;
	wire [8-1:0] node3393;
	wire [8-1:0] node3396;
	wire [8-1:0] node3399;
	wire [8-1:0] node3400;
	wire [8-1:0] node3403;
	wire [8-1:0] node3406;
	wire [8-1:0] node3407;
	wire [8-1:0] node3409;
	wire [8-1:0] node3412;
	wire [8-1:0] node3414;
	wire [8-1:0] node3417;
	wire [8-1:0] node3418;
	wire [8-1:0] node3419;
	wire [8-1:0] node3420;
	wire [8-1:0] node3421;
	wire [8-1:0] node3422;
	wire [8-1:0] node3423;
	wire [8-1:0] node3424;
	wire [8-1:0] node3427;
	wire [8-1:0] node3430;
	wire [8-1:0] node3431;
	wire [8-1:0] node3432;
	wire [8-1:0] node3436;
	wire [8-1:0] node3439;
	wire [8-1:0] node3440;
	wire [8-1:0] node3442;
	wire [8-1:0] node3445;
	wire [8-1:0] node3447;
	wire [8-1:0] node3450;
	wire [8-1:0] node3451;
	wire [8-1:0] node3452;
	wire [8-1:0] node3454;
	wire [8-1:0] node3456;
	wire [8-1:0] node3459;
	wire [8-1:0] node3460;
	wire [8-1:0] node3461;
	wire [8-1:0] node3464;
	wire [8-1:0] node3467;
	wire [8-1:0] node3469;
	wire [8-1:0] node3472;
	wire [8-1:0] node3473;
	wire [8-1:0] node3474;
	wire [8-1:0] node3475;
	wire [8-1:0] node3478;
	wire [8-1:0] node3481;
	wire [8-1:0] node3482;
	wire [8-1:0] node3486;
	wire [8-1:0] node3487;
	wire [8-1:0] node3488;
	wire [8-1:0] node3492;
	wire [8-1:0] node3493;
	wire [8-1:0] node3496;
	wire [8-1:0] node3499;
	wire [8-1:0] node3500;
	wire [8-1:0] node3501;
	wire [8-1:0] node3502;
	wire [8-1:0] node3505;
	wire [8-1:0] node3508;
	wire [8-1:0] node3509;
	wire [8-1:0] node3511;
	wire [8-1:0] node3512;
	wire [8-1:0] node3515;
	wire [8-1:0] node3518;
	wire [8-1:0] node3519;
	wire [8-1:0] node3520;
	wire [8-1:0] node3525;
	wire [8-1:0] node3526;
	wire [8-1:0] node3527;
	wire [8-1:0] node3528;
	wire [8-1:0] node3529;
	wire [8-1:0] node3532;
	wire [8-1:0] node3535;
	wire [8-1:0] node3538;
	wire [8-1:0] node3539;
	wire [8-1:0] node3543;
	wire [8-1:0] node3544;
	wire [8-1:0] node3545;
	wire [8-1:0] node3546;
	wire [8-1:0] node3550;
	wire [8-1:0] node3551;
	wire [8-1:0] node3555;
	wire [8-1:0] node3556;
	wire [8-1:0] node3557;
	wire [8-1:0] node3561;
	wire [8-1:0] node3563;
	wire [8-1:0] node3566;
	wire [8-1:0] node3567;
	wire [8-1:0] node3568;
	wire [8-1:0] node3569;
	wire [8-1:0] node3571;
	wire [8-1:0] node3575;
	wire [8-1:0] node3576;
	wire [8-1:0] node3579;
	wire [8-1:0] node3580;
	wire [8-1:0] node3584;
	wire [8-1:0] node3585;
	wire [8-1:0] node3586;
	wire [8-1:0] node3588;
	wire [8-1:0] node3592;
	wire [8-1:0] node3593;
	wire [8-1:0] node3596;
	wire [8-1:0] node3597;
	wire [8-1:0] node3601;
	wire [8-1:0] node3602;
	wire [8-1:0] node3603;
	wire [8-1:0] node3604;
	wire [8-1:0] node3605;
	wire [8-1:0] node3606;
	wire [8-1:0] node3607;
	wire [8-1:0] node3610;
	wire [8-1:0] node3613;
	wire [8-1:0] node3614;
	wire [8-1:0] node3615;
	wire [8-1:0] node3618;
	wire [8-1:0] node3621;
	wire [8-1:0] node3622;
	wire [8-1:0] node3626;
	wire [8-1:0] node3627;
	wire [8-1:0] node3628;
	wire [8-1:0] node3631;
	wire [8-1:0] node3634;
	wire [8-1:0] node3636;
	wire [8-1:0] node3638;
	wire [8-1:0] node3641;
	wire [8-1:0] node3642;
	wire [8-1:0] node3643;
	wire [8-1:0] node3645;
	wire [8-1:0] node3648;
	wire [8-1:0] node3649;
	wire [8-1:0] node3651;
	wire [8-1:0] node3654;
	wire [8-1:0] node3657;
	wire [8-1:0] node3658;
	wire [8-1:0] node3660;
	wire [8-1:0] node3661;
	wire [8-1:0] node3665;
	wire [8-1:0] node3666;
	wire [8-1:0] node3669;
	wire [8-1:0] node3670;
	wire [8-1:0] node3673;
	wire [8-1:0] node3676;
	wire [8-1:0] node3677;
	wire [8-1:0] node3679;
	wire [8-1:0] node3682;
	wire [8-1:0] node3684;
	wire [8-1:0] node3687;
	wire [8-1:0] node3688;
	wire [8-1:0] node3689;
	wire [8-1:0] node3690;
	wire [8-1:0] node3691;
	wire [8-1:0] node3694;
	wire [8-1:0] node3695;
	wire [8-1:0] node3698;
	wire [8-1:0] node3701;
	wire [8-1:0] node3702;
	wire [8-1:0] node3703;
	wire [8-1:0] node3706;
	wire [8-1:0] node3709;
	wire [8-1:0] node3710;
	wire [8-1:0] node3713;
	wire [8-1:0] node3716;
	wire [8-1:0] node3717;
	wire [8-1:0] node3718;
	wire [8-1:0] node3720;
	wire [8-1:0] node3723;
	wire [8-1:0] node3724;
	wire [8-1:0] node3728;
	wire [8-1:0] node3729;
	wire [8-1:0] node3730;
	wire [8-1:0] node3734;
	wire [8-1:0] node3735;
	wire [8-1:0] node3739;
	wire [8-1:0] node3742;
	wire [8-1:0] node3743;
	wire [8-1:0] node3744;
	wire [8-1:0] node3745;
	wire [8-1:0] node3746;
	wire [8-1:0] node3747;
	wire [8-1:0] node3748;
	wire [8-1:0] node3749;
	wire [8-1:0] node3750;
	wire [8-1:0] node3751;
	wire [8-1:0] node3752;
	wire [8-1:0] node3756;
	wire [8-1:0] node3757;
	wire [8-1:0] node3761;
	wire [8-1:0] node3762;
	wire [8-1:0] node3763;
	wire [8-1:0] node3766;
	wire [8-1:0] node3767;
	wire [8-1:0] node3771;
	wire [8-1:0] node3772;
	wire [8-1:0] node3773;
	wire [8-1:0] node3775;
	wire [8-1:0] node3778;
	wire [8-1:0] node3780;
	wire [8-1:0] node3783;
	wire [8-1:0] node3786;
	wire [8-1:0] node3787;
	wire [8-1:0] node3788;
	wire [8-1:0] node3790;
	wire [8-1:0] node3793;
	wire [8-1:0] node3794;
	wire [8-1:0] node3798;
	wire [8-1:0] node3799;
	wire [8-1:0] node3800;
	wire [8-1:0] node3803;
	wire [8-1:0] node3806;
	wire [8-1:0] node3807;
	wire [8-1:0] node3809;
	wire [8-1:0] node3812;
	wire [8-1:0] node3813;
	wire [8-1:0] node3815;
	wire [8-1:0] node3819;
	wire [8-1:0] node3820;
	wire [8-1:0] node3821;
	wire [8-1:0] node3822;
	wire [8-1:0] node3824;
	wire [8-1:0] node3827;
	wire [8-1:0] node3828;
	wire [8-1:0] node3829;
	wire [8-1:0] node3832;
	wire [8-1:0] node3835;
	wire [8-1:0] node3836;
	wire [8-1:0] node3837;
	wire [8-1:0] node3842;
	wire [8-1:0] node3843;
	wire [8-1:0] node3844;
	wire [8-1:0] node3845;
	wire [8-1:0] node3849;
	wire [8-1:0] node3852;
	wire [8-1:0] node3853;
	wire [8-1:0] node3854;
	wire [8-1:0] node3858;
	wire [8-1:0] node3859;
	wire [8-1:0] node3863;
	wire [8-1:0] node3864;
	wire [8-1:0] node3865;
	wire [8-1:0] node3867;
	wire [8-1:0] node3868;
	wire [8-1:0] node3871;
	wire [8-1:0] node3874;
	wire [8-1:0] node3875;
	wire [8-1:0] node3878;
	wire [8-1:0] node3880;
	wire [8-1:0] node3882;
	wire [8-1:0] node3885;
	wire [8-1:0] node3886;
	wire [8-1:0] node3887;
	wire [8-1:0] node3888;
	wire [8-1:0] node3891;
	wire [8-1:0] node3894;
	wire [8-1:0] node3895;
	wire [8-1:0] node3898;
	wire [8-1:0] node3901;
	wire [8-1:0] node3903;
	wire [8-1:0] node3904;
	wire [8-1:0] node3907;
	wire [8-1:0] node3910;
	wire [8-1:0] node3911;
	wire [8-1:0] node3912;
	wire [8-1:0] node3913;
	wire [8-1:0] node3915;
	wire [8-1:0] node3916;
	wire [8-1:0] node3920;
	wire [8-1:0] node3921;
	wire [8-1:0] node3922;
	wire [8-1:0] node3923;
	wire [8-1:0] node3926;
	wire [8-1:0] node3929;
	wire [8-1:0] node3930;
	wire [8-1:0] node3934;
	wire [8-1:0] node3935;
	wire [8-1:0] node3938;
	wire [8-1:0] node3940;
	wire [8-1:0] node3943;
	wire [8-1:0] node3944;
	wire [8-1:0] node3945;
	wire [8-1:0] node3947;
	wire [8-1:0] node3949;
	wire [8-1:0] node3950;
	wire [8-1:0] node3953;
	wire [8-1:0] node3956;
	wire [8-1:0] node3957;
	wire [8-1:0] node3959;
	wire [8-1:0] node3962;
	wire [8-1:0] node3965;
	wire [8-1:0] node3966;
	wire [8-1:0] node3968;
	wire [8-1:0] node3972;
	wire [8-1:0] node3973;
	wire [8-1:0] node3974;
	wire [8-1:0] node3975;
	wire [8-1:0] node3976;
	wire [8-1:0] node3978;
	wire [8-1:0] node3981;
	wire [8-1:0] node3983;
	wire [8-1:0] node3986;
	wire [8-1:0] node3987;
	wire [8-1:0] node3989;
	wire [8-1:0] node3992;
	wire [8-1:0] node3994;
	wire [8-1:0] node3997;
	wire [8-1:0] node3998;
	wire [8-1:0] node3999;
	wire [8-1:0] node4002;
	wire [8-1:0] node4005;
	wire [8-1:0] node4006;
	wire [8-1:0] node4008;
	wire [8-1:0] node4010;
	wire [8-1:0] node4013;
	wire [8-1:0] node4014;
	wire [8-1:0] node4015;
	wire [8-1:0] node4020;
	wire [8-1:0] node4021;
	wire [8-1:0] node4022;
	wire [8-1:0] node4023;
	wire [8-1:0] node4025;
	wire [8-1:0] node4028;
	wire [8-1:0] node4031;
	wire [8-1:0] node4032;
	wire [8-1:0] node4034;
	wire [8-1:0] node4035;
	wire [8-1:0] node4039;
	wire [8-1:0] node4040;
	wire [8-1:0] node4044;
	wire [8-1:0] node4045;
	wire [8-1:0] node4047;
	wire [8-1:0] node4048;
	wire [8-1:0] node4049;
	wire [8-1:0] node4053;
	wire [8-1:0] node4056;
	wire [8-1:0] node4057;
	wire [8-1:0] node4059;
	wire [8-1:0] node4062;
	wire [8-1:0] node4063;
	wire [8-1:0] node4064;
	wire [8-1:0] node4067;
	wire [8-1:0] node4071;
	wire [8-1:0] node4072;
	wire [8-1:0] node4073;
	wire [8-1:0] node4074;
	wire [8-1:0] node4075;
	wire [8-1:0] node4076;
	wire [8-1:0] node4078;
	wire [8-1:0] node4081;
	wire [8-1:0] node4082;
	wire [8-1:0] node4083;
	wire [8-1:0] node4087;
	wire [8-1:0] node4088;
	wire [8-1:0] node4092;
	wire [8-1:0] node4093;
	wire [8-1:0] node4094;
	wire [8-1:0] node4097;
	wire [8-1:0] node4098;
	wire [8-1:0] node4102;
	wire [8-1:0] node4103;
	wire [8-1:0] node4107;
	wire [8-1:0] node4108;
	wire [8-1:0] node4109;
	wire [8-1:0] node4110;
	wire [8-1:0] node4114;
	wire [8-1:0] node4115;
	wire [8-1:0] node4119;
	wire [8-1:0] node4121;
	wire [8-1:0] node4124;
	wire [8-1:0] node4125;
	wire [8-1:0] node4126;
	wire [8-1:0] node4127;
	wire [8-1:0] node4128;
	wire [8-1:0] node4131;
	wire [8-1:0] node4134;
	wire [8-1:0] node4135;
	wire [8-1:0] node4137;
	wire [8-1:0] node4140;
	wire [8-1:0] node4142;
	wire [8-1:0] node4145;
	wire [8-1:0] node4146;
	wire [8-1:0] node4147;
	wire [8-1:0] node4150;
	wire [8-1:0] node4151;
	wire [8-1:0] node4154;
	wire [8-1:0] node4157;
	wire [8-1:0] node4158;
	wire [8-1:0] node4159;
	wire [8-1:0] node4163;
	wire [8-1:0] node4164;
	wire [8-1:0] node4168;
	wire [8-1:0] node4169;
	wire [8-1:0] node4170;
	wire [8-1:0] node4172;
	wire [8-1:0] node4175;
	wire [8-1:0] node4176;
	wire [8-1:0] node4179;
	wire [8-1:0] node4181;
	wire [8-1:0] node4184;
	wire [8-1:0] node4185;
	wire [8-1:0] node4186;
	wire [8-1:0] node4187;
	wire [8-1:0] node4190;
	wire [8-1:0] node4193;
	wire [8-1:0] node4195;
	wire [8-1:0] node4198;
	wire [8-1:0] node4199;
	wire [8-1:0] node4201;
	wire [8-1:0] node4203;
	wire [8-1:0] node4206;
	wire [8-1:0] node4207;
	wire [8-1:0] node4209;
	wire [8-1:0] node4212;
	wire [8-1:0] node4215;
	wire [8-1:0] node4216;
	wire [8-1:0] node4217;
	wire [8-1:0] node4218;
	wire [8-1:0] node4219;
	wire [8-1:0] node4220;
	wire [8-1:0] node4221;
	wire [8-1:0] node4224;
	wire [8-1:0] node4227;
	wire [8-1:0] node4228;
	wire [8-1:0] node4231;
	wire [8-1:0] node4234;
	wire [8-1:0] node4235;
	wire [8-1:0] node4236;
	wire [8-1:0] node4240;
	wire [8-1:0] node4241;
	wire [8-1:0] node4243;
	wire [8-1:0] node4246;
	wire [8-1:0] node4247;
	wire [8-1:0] node4251;
	wire [8-1:0] node4252;
	wire [8-1:0] node4253;
	wire [8-1:0] node4254;
	wire [8-1:0] node4257;
	wire [8-1:0] node4260;
	wire [8-1:0] node4261;
	wire [8-1:0] node4264;
	wire [8-1:0] node4267;
	wire [8-1:0] node4268;
	wire [8-1:0] node4269;
	wire [8-1:0] node4272;
	wire [8-1:0] node4275;
	wire [8-1:0] node4276;
	wire [8-1:0] node4277;
	wire [8-1:0] node4281;
	wire [8-1:0] node4284;
	wire [8-1:0] node4285;
	wire [8-1:0] node4286;
	wire [8-1:0] node4287;
	wire [8-1:0] node4291;
	wire [8-1:0] node4292;
	wire [8-1:0] node4296;
	wire [8-1:0] node4297;
	wire [8-1:0] node4298;
	wire [8-1:0] node4302;
	wire [8-1:0] node4303;
	wire [8-1:0] node4307;
	wire [8-1:0] node4308;
	wire [8-1:0] node4309;
	wire [8-1:0] node4310;
	wire [8-1:0] node4311;
	wire [8-1:0] node4312;
	wire [8-1:0] node4315;
	wire [8-1:0] node4318;
	wire [8-1:0] node4319;
	wire [8-1:0] node4323;
	wire [8-1:0] node4324;
	wire [8-1:0] node4325;
	wire [8-1:0] node4326;
	wire [8-1:0] node4330;
	wire [8-1:0] node4331;
	wire [8-1:0] node4334;
	wire [8-1:0] node4337;
	wire [8-1:0] node4338;
	wire [8-1:0] node4339;
	wire [8-1:0] node4343;
	wire [8-1:0] node4346;
	wire [8-1:0] node4347;
	wire [8-1:0] node4348;
	wire [8-1:0] node4349;
	wire [8-1:0] node4350;
	wire [8-1:0] node4354;
	wire [8-1:0] node4355;
	wire [8-1:0] node4358;
	wire [8-1:0] node4361;
	wire [8-1:0] node4362;
	wire [8-1:0] node4363;
	wire [8-1:0] node4366;
	wire [8-1:0] node4370;
	wire [8-1:0] node4371;
	wire [8-1:0] node4372;
	wire [8-1:0] node4374;
	wire [8-1:0] node4377;
	wire [8-1:0] node4378;
	wire [8-1:0] node4381;
	wire [8-1:0] node4384;
	wire [8-1:0] node4385;
	wire [8-1:0] node4387;
	wire [8-1:0] node4391;
	wire [8-1:0] node4392;
	wire [8-1:0] node4393;
	wire [8-1:0] node4394;
	wire [8-1:0] node4395;
	wire [8-1:0] node4399;
	wire [8-1:0] node4400;
	wire [8-1:0] node4403;
	wire [8-1:0] node4406;
	wire [8-1:0] node4407;
	wire [8-1:0] node4410;
	wire [8-1:0] node4411;
	wire [8-1:0] node4415;
	wire [8-1:0] node4416;
	wire [8-1:0] node4417;
	wire [8-1:0] node4421;
	wire [8-1:0] node4422;
	wire [8-1:0] node4425;
	wire [8-1:0] node4428;
	wire [8-1:0] node4429;
	wire [8-1:0] node4430;
	wire [8-1:0] node4431;
	wire [8-1:0] node4432;
	wire [8-1:0] node4434;
	wire [8-1:0] node4435;
	wire [8-1:0] node4439;
	wire [8-1:0] node4440;
	wire [8-1:0] node4441;
	wire [8-1:0] node4445;
	wire [8-1:0] node4446;
	wire [8-1:0] node4447;
	wire [8-1:0] node4450;
	wire [8-1:0] node4454;
	wire [8-1:0] node4455;
	wire [8-1:0] node4456;
	wire [8-1:0] node4457;
	wire [8-1:0] node4458;
	wire [8-1:0] node4461;
	wire [8-1:0] node4463;
	wire [8-1:0] node4466;
	wire [8-1:0] node4467;
	wire [8-1:0] node4468;
	wire [8-1:0] node4471;
	wire [8-1:0] node4474;
	wire [8-1:0] node4475;
	wire [8-1:0] node4479;
	wire [8-1:0] node4480;
	wire [8-1:0] node4481;
	wire [8-1:0] node4482;
	wire [8-1:0] node4485;
	wire [8-1:0] node4488;
	wire [8-1:0] node4489;
	wire [8-1:0] node4493;
	wire [8-1:0] node4494;
	wire [8-1:0] node4496;
	wire [8-1:0] node4500;
	wire [8-1:0] node4501;
	wire [8-1:0] node4502;
	wire [8-1:0] node4503;
	wire [8-1:0] node4504;
	wire [8-1:0] node4507;
	wire [8-1:0] node4510;
	wire [8-1:0] node4511;
	wire [8-1:0] node4512;
	wire [8-1:0] node4516;
	wire [8-1:0] node4518;
	wire [8-1:0] node4521;
	wire [8-1:0] node4522;
	wire [8-1:0] node4523;
	wire [8-1:0] node4524;
	wire [8-1:0] node4527;
	wire [8-1:0] node4531;
	wire [8-1:0] node4532;
	wire [8-1:0] node4533;
	wire [8-1:0] node4536;
	wire [8-1:0] node4540;
	wire [8-1:0] node4541;
	wire [8-1:0] node4542;
	wire [8-1:0] node4543;
	wire [8-1:0] node4547;
	wire [8-1:0] node4548;
	wire [8-1:0] node4553;
	wire [8-1:0] node4554;
	wire [8-1:0] node4555;
	wire [8-1:0] node4556;
	wire [8-1:0] node4557;
	wire [8-1:0] node4558;
	wire [8-1:0] node4562;
	wire [8-1:0] node4563;
	wire [8-1:0] node4565;
	wire [8-1:0] node4568;
	wire [8-1:0] node4571;
	wire [8-1:0] node4572;
	wire [8-1:0] node4573;
	wire [8-1:0] node4574;
	wire [8-1:0] node4578;
	wire [8-1:0] node4579;
	wire [8-1:0] node4582;
	wire [8-1:0] node4585;
	wire [8-1:0] node4586;
	wire [8-1:0] node4589;
	wire [8-1:0] node4592;
	wire [8-1:0] node4593;
	wire [8-1:0] node4594;
	wire [8-1:0] node4595;
	wire [8-1:0] node4596;
	wire [8-1:0] node4598;
	wire [8-1:0] node4603;
	wire [8-1:0] node4604;
	wire [8-1:0] node4608;
	wire [8-1:0] node4609;
	wire [8-1:0] node4611;
	wire [8-1:0] node4612;
	wire [8-1:0] node4615;
	wire [8-1:0] node4618;
	wire [8-1:0] node4621;
	wire [8-1:0] node4622;
	wire [8-1:0] node4623;
	wire [8-1:0] node4625;
	wire [8-1:0] node4626;
	wire [8-1:0] node4629;
	wire [8-1:0] node4632;
	wire [8-1:0] node4634;
	wire [8-1:0] node4637;
	wire [8-1:0] node4638;
	wire [8-1:0] node4640;
	wire [8-1:0] node4644;
	wire [8-1:0] node4645;
	wire [8-1:0] node4646;
	wire [8-1:0] node4647;
	wire [8-1:0] node4648;
	wire [8-1:0] node4649;
	wire [8-1:0] node4650;
	wire [8-1:0] node4653;
	wire [8-1:0] node4656;
	wire [8-1:0] node4657;
	wire [8-1:0] node4660;
	wire [8-1:0] node4661;
	wire [8-1:0] node4665;
	wire [8-1:0] node4666;
	wire [8-1:0] node4667;
	wire [8-1:0] node4669;
	wire [8-1:0] node4672;
	wire [8-1:0] node4674;
	wire [8-1:0] node4677;
	wire [8-1:0] node4678;
	wire [8-1:0] node4680;
	wire [8-1:0] node4683;
	wire [8-1:0] node4685;
	wire [8-1:0] node4688;
	wire [8-1:0] node4689;
	wire [8-1:0] node4690;
	wire [8-1:0] node4691;
	wire [8-1:0] node4693;
	wire [8-1:0] node4694;
	wire [8-1:0] node4698;
	wire [8-1:0] node4699;
	wire [8-1:0] node4702;
	wire [8-1:0] node4705;
	wire [8-1:0] node4706;
	wire [8-1:0] node4709;
	wire [8-1:0] node4711;
	wire [8-1:0] node4713;
	wire [8-1:0] node4716;
	wire [8-1:0] node4717;
	wire [8-1:0] node4718;
	wire [8-1:0] node4719;
	wire [8-1:0] node4722;
	wire [8-1:0] node4725;
	wire [8-1:0] node4727;
	wire [8-1:0] node4730;
	wire [8-1:0] node4732;
	wire [8-1:0] node4734;
	wire [8-1:0] node4737;
	wire [8-1:0] node4738;
	wire [8-1:0] node4739;
	wire [8-1:0] node4740;
	wire [8-1:0] node4741;
	wire [8-1:0] node4744;
	wire [8-1:0] node4747;
	wire [8-1:0] node4748;
	wire [8-1:0] node4749;
	wire [8-1:0] node4752;
	wire [8-1:0] node4754;
	wire [8-1:0] node4757;
	wire [8-1:0] node4760;
	wire [8-1:0] node4761;
	wire [8-1:0] node4762;
	wire [8-1:0] node4764;
	wire [8-1:0] node4767;
	wire [8-1:0] node4769;
	wire [8-1:0] node4772;
	wire [8-1:0] node4773;
	wire [8-1:0] node4775;
	wire [8-1:0] node4778;
	wire [8-1:0] node4780;
	wire [8-1:0] node4783;
	wire [8-1:0] node4784;
	wire [8-1:0] node4785;
	wire [8-1:0] node4787;
	wire [8-1:0] node4790;
	wire [8-1:0] node4791;
	wire [8-1:0] node4792;
	wire [8-1:0] node4794;
	wire [8-1:0] node4797;
	wire [8-1:0] node4798;
	wire [8-1:0] node4802;
	wire [8-1:0] node4804;
	wire [8-1:0] node4807;
	wire [8-1:0] node4808;
	wire [8-1:0] node4809;
	wire [8-1:0] node4810;
	wire [8-1:0] node4814;
	wire [8-1:0] node4815;
	wire [8-1:0] node4816;
	wire [8-1:0] node4819;
	wire [8-1:0] node4822;
	wire [8-1:0] node4825;
	wire [8-1:0] node4826;
	wire [8-1:0] node4827;
	wire [8-1:0] node4830;
	wire [8-1:0] node4832;
	wire [8-1:0] node4835;
	wire [8-1:0] node4837;
	wire [8-1:0] node4838;
	wire [8-1:0] node4842;
	wire [8-1:0] node4843;
	wire [8-1:0] node4844;
	wire [8-1:0] node4845;
	wire [8-1:0] node4846;
	wire [8-1:0] node4848;
	wire [8-1:0] node4851;
	wire [8-1:0] node4852;
	wire [8-1:0] node4854;
	wire [8-1:0] node4857;
	wire [8-1:0] node4859;
	wire [8-1:0] node4862;
	wire [8-1:0] node4863;
	wire [8-1:0] node4864;
	wire [8-1:0] node4866;
	wire [8-1:0] node4869;
	wire [8-1:0] node4871;
	wire [8-1:0] node4874;
	wire [8-1:0] node4875;
	wire [8-1:0] node4877;
	wire [8-1:0] node4880;
	wire [8-1:0] node4882;
	wire [8-1:0] node4885;
	wire [8-1:0] node4886;
	wire [8-1:0] node4887;
	wire [8-1:0] node4888;
	wire [8-1:0] node4892;
	wire [8-1:0] node4893;
	wire [8-1:0] node4894;
	wire [8-1:0] node4899;
	wire [8-1:0] node4900;
	wire [8-1:0] node4901;
	wire [8-1:0] node4904;
	wire [8-1:0] node4906;
	wire [8-1:0] node4909;
	wire [8-1:0] node4910;
	wire [8-1:0] node4911;
	wire [8-1:0] node4912;
	wire [8-1:0] node4915;
	wire [8-1:0] node4918;
	wire [8-1:0] node4920;
	wire [8-1:0] node4923;
	wire [8-1:0] node4924;
	wire [8-1:0] node4927;
	wire [8-1:0] node4929;
	wire [8-1:0] node4932;
	wire [8-1:0] node4933;
	wire [8-1:0] node4934;
	wire [8-1:0] node4935;
	wire [8-1:0] node4936;
	wire [8-1:0] node4937;
	wire [8-1:0] node4939;
	wire [8-1:0] node4943;
	wire [8-1:0] node4944;
	wire [8-1:0] node4945;
	wire [8-1:0] node4949;
	wire [8-1:0] node4952;
	wire [8-1:0] node4953;
	wire [8-1:0] node4954;
	wire [8-1:0] node4955;
	wire [8-1:0] node4958;
	wire [8-1:0] node4961;
	wire [8-1:0] node4962;
	wire [8-1:0] node4966;
	wire [8-1:0] node4967;
	wire [8-1:0] node4969;
	wire [8-1:0] node4972;
	wire [8-1:0] node4974;
	wire [8-1:0] node4977;
	wire [8-1:0] node4978;
	wire [8-1:0] node4979;
	wire [8-1:0] node4980;
	wire [8-1:0] node4984;
	wire [8-1:0] node4987;
	wire [8-1:0] node4988;
	wire [8-1:0] node4990;
	wire [8-1:0] node4993;
	wire [8-1:0] node4996;
	wire [8-1:0] node4997;
	wire [8-1:0] node4998;
	wire [8-1:0] node4999;
	wire [8-1:0] node5000;
	wire [8-1:0] node5003;
	wire [8-1:0] node5006;
	wire [8-1:0] node5007;
	wire [8-1:0] node5009;
	wire [8-1:0] node5012;
	wire [8-1:0] node5013;
	wire [8-1:0] node5017;
	wire [8-1:0] node5018;
	wire [8-1:0] node5019;
	wire [8-1:0] node5021;
	wire [8-1:0] node5024;
	wire [8-1:0] node5025;
	wire [8-1:0] node5029;
	wire [8-1:0] node5030;
	wire [8-1:0] node5033;
	wire [8-1:0] node5035;
	wire [8-1:0] node5038;
	wire [8-1:0] node5039;
	wire [8-1:0] node5040;
	wire [8-1:0] node5043;
	wire [8-1:0] node5046;
	wire [8-1:0] node5049;
	wire [8-1:0] node5050;
	wire [8-1:0] node5051;
	wire [8-1:0] node5052;
	wire [8-1:0] node5053;
	wire [8-1:0] node5054;
	wire [8-1:0] node5055;
	wire [8-1:0] node5056;
	wire [8-1:0] node5058;
	wire [8-1:0] node5061;
	wire [8-1:0] node5062;
	wire [8-1:0] node5063;
	wire [8-1:0] node5068;
	wire [8-1:0] node5069;
	wire [8-1:0] node5073;
	wire [8-1:0] node5074;
	wire [8-1:0] node5075;
	wire [8-1:0] node5076;
	wire [8-1:0] node5077;
	wire [8-1:0] node5082;
	wire [8-1:0] node5083;
	wire [8-1:0] node5087;
	wire [8-1:0] node5088;
	wire [8-1:0] node5090;
	wire [8-1:0] node5093;
	wire [8-1:0] node5095;
	wire [8-1:0] node5096;
	wire [8-1:0] node5100;
	wire [8-1:0] node5101;
	wire [8-1:0] node5102;
	wire [8-1:0] node5103;
	wire [8-1:0] node5104;
	wire [8-1:0] node5108;
	wire [8-1:0] node5109;
	wire [8-1:0] node5113;
	wire [8-1:0] node5115;
	wire [8-1:0] node5118;
	wire [8-1:0] node5119;
	wire [8-1:0] node5120;
	wire [8-1:0] node5121;
	wire [8-1:0] node5125;
	wire [8-1:0] node5126;
	wire [8-1:0] node5129;
	wire [8-1:0] node5132;
	wire [8-1:0] node5133;
	wire [8-1:0] node5134;
	wire [8-1:0] node5138;
	wire [8-1:0] node5139;
	wire [8-1:0] node5141;
	wire [8-1:0] node5144;
	wire [8-1:0] node5147;
	wire [8-1:0] node5148;
	wire [8-1:0] node5149;
	wire [8-1:0] node5150;
	wire [8-1:0] node5151;
	wire [8-1:0] node5155;
	wire [8-1:0] node5156;
	wire [8-1:0] node5157;
	wire [8-1:0] node5161;
	wire [8-1:0] node5163;
	wire [8-1:0] node5166;
	wire [8-1:0] node5167;
	wire [8-1:0] node5168;
	wire [8-1:0] node5172;
	wire [8-1:0] node5173;
	wire [8-1:0] node5175;
	wire [8-1:0] node5178;
	wire [8-1:0] node5180;
	wire [8-1:0] node5183;
	wire [8-1:0] node5184;
	wire [8-1:0] node5185;
	wire [8-1:0] node5189;
	wire [8-1:0] node5190;
	wire [8-1:0] node5191;
	wire [8-1:0] node5195;
	wire [8-1:0] node5197;
	wire [8-1:0] node5200;
	wire [8-1:0] node5201;
	wire [8-1:0] node5202;
	wire [8-1:0] node5203;
	wire [8-1:0] node5204;
	wire [8-1:0] node5205;
	wire [8-1:0] node5206;
	wire [8-1:0] node5209;
	wire [8-1:0] node5212;
	wire [8-1:0] node5213;
	wire [8-1:0] node5216;
	wire [8-1:0] node5219;
	wire [8-1:0] node5220;
	wire [8-1:0] node5221;
	wire [8-1:0] node5222;
	wire [8-1:0] node5225;
	wire [8-1:0] node5228;
	wire [8-1:0] node5230;
	wire [8-1:0] node5231;
	wire [8-1:0] node5234;
	wire [8-1:0] node5237;
	wire [8-1:0] node5238;
	wire [8-1:0] node5239;
	wire [8-1:0] node5240;
	wire [8-1:0] node5243;
	wire [8-1:0] node5246;
	wire [8-1:0] node5249;
	wire [8-1:0] node5250;
	wire [8-1:0] node5252;
	wire [8-1:0] node5255;
	wire [8-1:0] node5256;
	wire [8-1:0] node5259;
	wire [8-1:0] node5262;
	wire [8-1:0] node5263;
	wire [8-1:0] node5264;
	wire [8-1:0] node5265;
	wire [8-1:0] node5268;
	wire [8-1:0] node5271;
	wire [8-1:0] node5273;
	wire [8-1:0] node5275;
	wire [8-1:0] node5278;
	wire [8-1:0] node5279;
	wire [8-1:0] node5282;
	wire [8-1:0] node5283;
	wire [8-1:0] node5284;
	wire [8-1:0] node5286;
	wire [8-1:0] node5290;
	wire [8-1:0] node5292;
	wire [8-1:0] node5294;
	wire [8-1:0] node5297;
	wire [8-1:0] node5298;
	wire [8-1:0] node5299;
	wire [8-1:0] node5300;
	wire [8-1:0] node5301;
	wire [8-1:0] node5302;
	wire [8-1:0] node5305;
	wire [8-1:0] node5308;
	wire [8-1:0] node5309;
	wire [8-1:0] node5312;
	wire [8-1:0] node5315;
	wire [8-1:0] node5316;
	wire [8-1:0] node5318;
	wire [8-1:0] node5319;
	wire [8-1:0] node5322;
	wire [8-1:0] node5325;
	wire [8-1:0] node5327;
	wire [8-1:0] node5329;
	wire [8-1:0] node5332;
	wire [8-1:0] node5333;
	wire [8-1:0] node5334;
	wire [8-1:0] node5335;
	wire [8-1:0] node5339;
	wire [8-1:0] node5342;
	wire [8-1:0] node5343;
	wire [8-1:0] node5345;
	wire [8-1:0] node5347;
	wire [8-1:0] node5350;
	wire [8-1:0] node5351;
	wire [8-1:0] node5354;
	wire [8-1:0] node5355;
	wire [8-1:0] node5358;
	wire [8-1:0] node5361;
	wire [8-1:0] node5362;
	wire [8-1:0] node5363;
	wire [8-1:0] node5365;
	wire [8-1:0] node5368;
	wire [8-1:0] node5369;
	wire [8-1:0] node5372;
	wire [8-1:0] node5374;
	wire [8-1:0] node5377;
	wire [8-1:0] node5378;
	wire [8-1:0] node5379;
	wire [8-1:0] node5380;
	wire [8-1:0] node5383;
	wire [8-1:0] node5384;
	wire [8-1:0] node5388;
	wire [8-1:0] node5389;
	wire [8-1:0] node5391;
	wire [8-1:0] node5394;
	wire [8-1:0] node5395;
	wire [8-1:0] node5399;
	wire [8-1:0] node5400;
	wire [8-1:0] node5401;
	wire [8-1:0] node5404;
	wire [8-1:0] node5407;
	wire [8-1:0] node5408;
	wire [8-1:0] node5409;
	wire [8-1:0] node5412;
	wire [8-1:0] node5415;
	wire [8-1:0] node5417;
	wire [8-1:0] node5420;
	wire [8-1:0] node5421;
	wire [8-1:0] node5422;
	wire [8-1:0] node5423;
	wire [8-1:0] node5425;
	wire [8-1:0] node5428;
	wire [8-1:0] node5429;
	wire [8-1:0] node5431;
	wire [8-1:0] node5434;
	wire [8-1:0] node5436;
	wire [8-1:0] node5439;
	wire [8-1:0] node5440;
	wire [8-1:0] node5441;
	wire [8-1:0] node5442;
	wire [8-1:0] node5446;
	wire [8-1:0] node5449;
	wire [8-1:0] node5450;
	wire [8-1:0] node5452;
	wire [8-1:0] node5455;
	wire [8-1:0] node5456;
	wire [8-1:0] node5459;
	wire [8-1:0] node5461;
	wire [8-1:0] node5464;
	wire [8-1:0] node5465;
	wire [8-1:0] node5466;
	wire [8-1:0] node5467;
	wire [8-1:0] node5470;
	wire [8-1:0] node5472;
	wire [8-1:0] node5475;
	wire [8-1:0] node5476;
	wire [8-1:0] node5478;
	wire [8-1:0] node5481;
	wire [8-1:0] node5483;
	wire [8-1:0] node5485;
	wire [8-1:0] node5488;
	wire [8-1:0] node5489;
	wire [8-1:0] node5490;
	wire [8-1:0] node5491;
	wire [8-1:0] node5492;
	wire [8-1:0] node5493;
	wire [8-1:0] node5496;
	wire [8-1:0] node5500;
	wire [8-1:0] node5501;
	wire [8-1:0] node5504;
	wire [8-1:0] node5506;
	wire [8-1:0] node5509;
	wire [8-1:0] node5510;
	wire [8-1:0] node5511;
	wire [8-1:0] node5514;
	wire [8-1:0] node5515;
	wire [8-1:0] node5519;
	wire [8-1:0] node5521;
	wire [8-1:0] node5523;
	wire [8-1:0] node5526;
	wire [8-1:0] node5527;
	wire [8-1:0] node5528;
	wire [8-1:0] node5530;
	wire [8-1:0] node5533;
	wire [8-1:0] node5534;
	wire [8-1:0] node5537;
	wire [8-1:0] node5540;
	wire [8-1:0] node5541;
	wire [8-1:0] node5543;
	wire [8-1:0] node5546;
	wire [8-1:0] node5548;
	wire [8-1:0] node5549;
	wire [8-1:0] node5553;
	wire [8-1:0] node5554;
	wire [8-1:0] node5555;
	wire [8-1:0] node5556;
	wire [8-1:0] node5557;
	wire [8-1:0] node5558;
	wire [8-1:0] node5559;
	wire [8-1:0] node5560;
	wire [8-1:0] node5561;
	wire [8-1:0] node5564;
	wire [8-1:0] node5567;
	wire [8-1:0] node5568;
	wire [8-1:0] node5572;
	wire [8-1:0] node5573;
	wire [8-1:0] node5574;
	wire [8-1:0] node5577;
	wire [8-1:0] node5580;
	wire [8-1:0] node5582;
	wire [8-1:0] node5585;
	wire [8-1:0] node5586;
	wire [8-1:0] node5587;
	wire [8-1:0] node5588;
	wire [8-1:0] node5589;
	wire [8-1:0] node5592;
	wire [8-1:0] node5595;
	wire [8-1:0] node5596;
	wire [8-1:0] node5599;
	wire [8-1:0] node5602;
	wire [8-1:0] node5604;
	wire [8-1:0] node5607;
	wire [8-1:0] node5608;
	wire [8-1:0] node5609;
	wire [8-1:0] node5612;
	wire [8-1:0] node5613;
	wire [8-1:0] node5616;
	wire [8-1:0] node5619;
	wire [8-1:0] node5620;
	wire [8-1:0] node5621;
	wire [8-1:0] node5624;
	wire [8-1:0] node5627;
	wire [8-1:0] node5629;
	wire [8-1:0] node5632;
	wire [8-1:0] node5633;
	wire [8-1:0] node5634;
	wire [8-1:0] node5635;
	wire [8-1:0] node5637;
	wire [8-1:0] node5638;
	wire [8-1:0] node5641;
	wire [8-1:0] node5644;
	wire [8-1:0] node5645;
	wire [8-1:0] node5648;
	wire [8-1:0] node5651;
	wire [8-1:0] node5652;
	wire [8-1:0] node5653;
	wire [8-1:0] node5654;
	wire [8-1:0] node5657;
	wire [8-1:0] node5660;
	wire [8-1:0] node5662;
	wire [8-1:0] node5665;
	wire [8-1:0] node5666;
	wire [8-1:0] node5669;
	wire [8-1:0] node5672;
	wire [8-1:0] node5673;
	wire [8-1:0] node5674;
	wire [8-1:0] node5675;
	wire [8-1:0] node5678;
	wire [8-1:0] node5681;
	wire [8-1:0] node5682;
	wire [8-1:0] node5685;
	wire [8-1:0] node5688;
	wire [8-1:0] node5689;
	wire [8-1:0] node5690;
	wire [8-1:0] node5693;
	wire [8-1:0] node5696;
	wire [8-1:0] node5697;
	wire [8-1:0] node5701;
	wire [8-1:0] node5702;
	wire [8-1:0] node5703;
	wire [8-1:0] node5704;
	wire [8-1:0] node5705;
	wire [8-1:0] node5706;
	wire [8-1:0] node5708;
	wire [8-1:0] node5711;
	wire [8-1:0] node5712;
	wire [8-1:0] node5715;
	wire [8-1:0] node5718;
	wire [8-1:0] node5720;
	wire [8-1:0] node5721;
	wire [8-1:0] node5724;
	wire [8-1:0] node5727;
	wire [8-1:0] node5728;
	wire [8-1:0] node5729;
	wire [8-1:0] node5733;
	wire [8-1:0] node5734;
	wire [8-1:0] node5737;
	wire [8-1:0] node5739;
	wire [8-1:0] node5742;
	wire [8-1:0] node5743;
	wire [8-1:0] node5744;
	wire [8-1:0] node5745;
	wire [8-1:0] node5749;
	wire [8-1:0] node5750;
	wire [8-1:0] node5751;
	wire [8-1:0] node5755;
	wire [8-1:0] node5756;
	wire [8-1:0] node5760;
	wire [8-1:0] node5761;
	wire [8-1:0] node5762;
	wire [8-1:0] node5766;
	wire [8-1:0] node5767;
	wire [8-1:0] node5770;
	wire [8-1:0] node5772;
	wire [8-1:0] node5775;
	wire [8-1:0] node5776;
	wire [8-1:0] node5777;
	wire [8-1:0] node5778;
	wire [8-1:0] node5779;
	wire [8-1:0] node5782;
	wire [8-1:0] node5785;
	wire [8-1:0] node5786;
	wire [8-1:0] node5789;
	wire [8-1:0] node5792;
	wire [8-1:0] node5793;
	wire [8-1:0] node5794;
	wire [8-1:0] node5796;
	wire [8-1:0] node5799;
	wire [8-1:0] node5800;
	wire [8-1:0] node5803;
	wire [8-1:0] node5806;
	wire [8-1:0] node5808;
	wire [8-1:0] node5811;
	wire [8-1:0] node5812;
	wire [8-1:0] node5813;
	wire [8-1:0] node5814;
	wire [8-1:0] node5817;
	wire [8-1:0] node5820;
	wire [8-1:0] node5822;
	wire [8-1:0] node5825;
	wire [8-1:0] node5826;
	wire [8-1:0] node5827;
	wire [8-1:0] node5830;
	wire [8-1:0] node5833;
	wire [8-1:0] node5834;
	wire [8-1:0] node5837;
	wire [8-1:0] node5840;
	wire [8-1:0] node5841;
	wire [8-1:0] node5842;
	wire [8-1:0] node5843;
	wire [8-1:0] node5844;
	wire [8-1:0] node5845;
	wire [8-1:0] node5848;
	wire [8-1:0] node5851;
	wire [8-1:0] node5852;
	wire [8-1:0] node5856;
	wire [8-1:0] node5857;
	wire [8-1:0] node5858;
	wire [8-1:0] node5862;
	wire [8-1:0] node5863;
	wire [8-1:0] node5866;
	wire [8-1:0] node5869;
	wire [8-1:0] node5870;
	wire [8-1:0] node5871;
	wire [8-1:0] node5872;
	wire [8-1:0] node5875;
	wire [8-1:0] node5878;
	wire [8-1:0] node5879;
	wire [8-1:0] node5883;
	wire [8-1:0] node5884;
	wire [8-1:0] node5888;
	wire [8-1:0] node5889;
	wire [8-1:0] node5890;
	wire [8-1:0] node5892;
	wire [8-1:0] node5895;
	wire [8-1:0] node5897;
	wire [8-1:0] node5898;
	wire [8-1:0] node5902;
	wire [8-1:0] node5903;
	wire [8-1:0] node5904;
	wire [8-1:0] node5906;
	wire [8-1:0] node5910;
	wire [8-1:0] node5912;
	wire [8-1:0] node5914;
	wire [8-1:0] node5917;
	wire [8-1:0] node5918;
	wire [8-1:0] node5919;
	wire [8-1:0] node5920;
	wire [8-1:0] node5921;
	wire [8-1:0] node5922;
	wire [8-1:0] node5923;
	wire [8-1:0] node5924;
	wire [8-1:0] node5926;
	wire [8-1:0] node5930;
	wire [8-1:0] node5932;
	wire [8-1:0] node5934;
	wire [8-1:0] node5937;
	wire [8-1:0] node5938;
	wire [8-1:0] node5939;
	wire [8-1:0] node5940;
	wire [8-1:0] node5943;
	wire [8-1:0] node5947;
	wire [8-1:0] node5948;
	wire [8-1:0] node5951;
	wire [8-1:0] node5952;
	wire [8-1:0] node5955;
	wire [8-1:0] node5958;
	wire [8-1:0] node5959;
	wire [8-1:0] node5960;
	wire [8-1:0] node5963;
	wire [8-1:0] node5964;
	wire [8-1:0] node5967;
	wire [8-1:0] node5968;
	wire [8-1:0] node5971;
	wire [8-1:0] node5974;
	wire [8-1:0] node5975;
	wire [8-1:0] node5976;
	wire [8-1:0] node5977;
	wire [8-1:0] node5980;
	wire [8-1:0] node5983;
	wire [8-1:0] node5984;
	wire [8-1:0] node5988;
	wire [8-1:0] node5989;
	wire [8-1:0] node5990;
	wire [8-1:0] node5993;
	wire [8-1:0] node5997;
	wire [8-1:0] node5998;
	wire [8-1:0] node5999;
	wire [8-1:0] node6000;
	wire [8-1:0] node6001;
	wire [8-1:0] node6002;
	wire [8-1:0] node6007;
	wire [8-1:0] node6009;
	wire [8-1:0] node6010;
	wire [8-1:0] node6013;
	wire [8-1:0] node6016;
	wire [8-1:0] node6017;
	wire [8-1:0] node6018;
	wire [8-1:0] node6019;
	wire [8-1:0] node6023;
	wire [8-1:0] node6026;
	wire [8-1:0] node6027;
	wire [8-1:0] node6030;
	wire [8-1:0] node6031;
	wire [8-1:0] node6034;
	wire [8-1:0] node6037;
	wire [8-1:0] node6038;
	wire [8-1:0] node6039;
	wire [8-1:0] node6040;
	wire [8-1:0] node6041;
	wire [8-1:0] node6046;
	wire [8-1:0] node6047;
	wire [8-1:0] node6048;
	wire [8-1:0] node6052;
	wire [8-1:0] node6053;
	wire [8-1:0] node6057;
	wire [8-1:0] node6058;
	wire [8-1:0] node6059;
	wire [8-1:0] node6062;
	wire [8-1:0] node6064;
	wire [8-1:0] node6067;
	wire [8-1:0] node6068;
	wire [8-1:0] node6071;
	wire [8-1:0] node6074;
	wire [8-1:0] node6075;
	wire [8-1:0] node6076;
	wire [8-1:0] node6077;
	wire [8-1:0] node6078;
	wire [8-1:0] node6079;
	wire [8-1:0] node6082;
	wire [8-1:0] node6083;
	wire [8-1:0] node6087;
	wire [8-1:0] node6088;
	wire [8-1:0] node6089;
	wire [8-1:0] node6093;
	wire [8-1:0] node6096;
	wire [8-1:0] node6097;
	wire [8-1:0] node6098;
	wire [8-1:0] node6100;
	wire [8-1:0] node6103;
	wire [8-1:0] node6106;
	wire [8-1:0] node6107;
	wire [8-1:0] node6108;
	wire [8-1:0] node6111;
	wire [8-1:0] node6114;
	wire [8-1:0] node6116;
	wire [8-1:0] node6119;
	wire [8-1:0] node6120;
	wire [8-1:0] node6121;
	wire [8-1:0] node6122;
	wire [8-1:0] node6123;
	wire [8-1:0] node6126;
	wire [8-1:0] node6129;
	wire [8-1:0] node6132;
	wire [8-1:0] node6133;
	wire [8-1:0] node6135;
	wire [8-1:0] node6138;
	wire [8-1:0] node6139;
	wire [8-1:0] node6143;
	wire [8-1:0] node6144;
	wire [8-1:0] node6145;
	wire [8-1:0] node6147;
	wire [8-1:0] node6150;
	wire [8-1:0] node6153;
	wire [8-1:0] node6154;
	wire [8-1:0] node6155;
	wire [8-1:0] node6158;
	wire [8-1:0] node6162;
	wire [8-1:0] node6163;
	wire [8-1:0] node6164;
	wire [8-1:0] node6165;
	wire [8-1:0] node6166;
	wire [8-1:0] node6168;
	wire [8-1:0] node6171;
	wire [8-1:0] node6172;
	wire [8-1:0] node6176;
	wire [8-1:0] node6178;
	wire [8-1:0] node6179;
	wire [8-1:0] node6182;
	wire [8-1:0] node6185;
	wire [8-1:0] node6186;
	wire [8-1:0] node6187;
	wire [8-1:0] node6190;
	wire [8-1:0] node6191;
	wire [8-1:0] node6194;
	wire [8-1:0] node6197;
	wire [8-1:0] node6198;
	wire [8-1:0] node6199;
	wire [8-1:0] node6203;
	wire [8-1:0] node6204;
	wire [8-1:0] node6207;
	wire [8-1:0] node6210;
	wire [8-1:0] node6211;
	wire [8-1:0] node6212;
	wire [8-1:0] node6213;
	wire [8-1:0] node6214;
	wire [8-1:0] node6217;
	wire [8-1:0] node6220;
	wire [8-1:0] node6221;
	wire [8-1:0] node6224;
	wire [8-1:0] node6227;
	wire [8-1:0] node6228;
	wire [8-1:0] node6229;
	wire [8-1:0] node6232;
	wire [8-1:0] node6235;
	wire [8-1:0] node6236;
	wire [8-1:0] node6240;
	wire [8-1:0] node6241;
	wire [8-1:0] node6243;
	wire [8-1:0] node6246;
	wire [8-1:0] node6247;
	wire [8-1:0] node6249;
	wire [8-1:0] node6252;
	wire [8-1:0] node6255;
	wire [8-1:0] node6256;
	wire [8-1:0] node6257;
	wire [8-1:0] node6258;
	wire [8-1:0] node6259;
	wire [8-1:0] node6260;
	wire [8-1:0] node6262;
	wire [8-1:0] node6265;
	wire [8-1:0] node6268;
	wire [8-1:0] node6269;
	wire [8-1:0] node6270;
	wire [8-1:0] node6271;
	wire [8-1:0] node6274;
	wire [8-1:0] node6278;
	wire [8-1:0] node6281;
	wire [8-1:0] node6282;
	wire [8-1:0] node6283;
	wire [8-1:0] node6286;
	wire [8-1:0] node6289;
	wire [8-1:0] node6292;
	wire [8-1:0] node6293;
	wire [8-1:0] node6294;
	wire [8-1:0] node6295;
	wire [8-1:0] node6296;
	wire [8-1:0] node6299;
	wire [8-1:0] node6302;
	wire [8-1:0] node6305;
	wire [8-1:0] node6306;
	wire [8-1:0] node6309;
	wire [8-1:0] node6312;
	wire [8-1:0] node6313;
	wire [8-1:0] node6314;
	wire [8-1:0] node6317;
	wire [8-1:0] node6320;
	wire [8-1:0] node6323;
	wire [8-1:0] node6324;
	wire [8-1:0] node6325;
	wire [8-1:0] node6326;
	wire [8-1:0] node6327;
	wire [8-1:0] node6330;
	wire [8-1:0] node6333;
	wire [8-1:0] node6336;
	wire [8-1:0] node6337;
	wire [8-1:0] node6338;
	wire [8-1:0] node6341;
	wire [8-1:0] node6344;
	wire [8-1:0] node6347;
	wire [8-1:0] node6348;
	wire [8-1:0] node6349;
	wire [8-1:0] node6352;
	wire [8-1:0] node6355;
	wire [8-1:0] node6358;
	wire [8-1:0] node6359;
	wire [8-1:0] node6360;
	wire [8-1:0] node6361;
	wire [8-1:0] node6363;
	wire [8-1:0] node6364;
	wire [8-1:0] node6365;
	wire [8-1:0] node6366;
	wire [8-1:0] node6367;
	wire [8-1:0] node6368;
	wire [8-1:0] node6372;
	wire [8-1:0] node6373;
	wire [8-1:0] node6375;
	wire [8-1:0] node6378;
	wire [8-1:0] node6381;
	wire [8-1:0] node6382;
	wire [8-1:0] node6383;
	wire [8-1:0] node6387;
	wire [8-1:0] node6388;
	wire [8-1:0] node6389;
	wire [8-1:0] node6393;
	wire [8-1:0] node6396;
	wire [8-1:0] node6397;
	wire [8-1:0] node6398;
	wire [8-1:0] node6400;
	wire [8-1:0] node6403;
	wire [8-1:0] node6404;
	wire [8-1:0] node6408;
	wire [8-1:0] node6409;
	wire [8-1:0] node6413;
	wire [8-1:0] node6414;
	wire [8-1:0] node6415;
	wire [8-1:0] node6416;
	wire [8-1:0] node6417;
	wire [8-1:0] node6418;
	wire [8-1:0] node6423;
	wire [8-1:0] node6424;
	wire [8-1:0] node6426;
	wire [8-1:0] node6429;
	wire [8-1:0] node6430;
	wire [8-1:0] node6433;
	wire [8-1:0] node6436;
	wire [8-1:0] node6437;
	wire [8-1:0] node6438;
	wire [8-1:0] node6442;
	wire [8-1:0] node6443;
	wire [8-1:0] node6444;
	wire [8-1:0] node6449;
	wire [8-1:0] node6450;
	wire [8-1:0] node6451;
	wire [8-1:0] node6454;
	wire [8-1:0] node6455;
	wire [8-1:0] node6459;
	wire [8-1:0] node6460;
	wire [8-1:0] node6461;
	wire [8-1:0] node6463;
	wire [8-1:0] node6466;
	wire [8-1:0] node6469;
	wire [8-1:0] node6470;
	wire [8-1:0] node6472;
	wire [8-1:0] node6475;
	wire [8-1:0] node6476;
	wire [8-1:0] node6478;
	wire [8-1:0] node6482;
	wire [8-1:0] node6483;
	wire [8-1:0] node6484;
	wire [8-1:0] node6485;
	wire [8-1:0] node6487;
	wire [8-1:0] node6488;
	wire [8-1:0] node6492;
	wire [8-1:0] node6493;
	wire [8-1:0] node6494;
	wire [8-1:0] node6498;
	wire [8-1:0] node6499;
	wire [8-1:0] node6500;
	wire [8-1:0] node6503;
	wire [8-1:0] node6507;
	wire [8-1:0] node6508;
	wire [8-1:0] node6509;
	wire [8-1:0] node6510;
	wire [8-1:0] node6514;
	wire [8-1:0] node6515;
	wire [8-1:0] node6516;
	wire [8-1:0] node6519;
	wire [8-1:0] node6523;
	wire [8-1:0] node6524;
	wire [8-1:0] node6525;
	wire [8-1:0] node6526;
	wire [8-1:0] node6528;
	wire [8-1:0] node6532;
	wire [8-1:0] node6533;
	wire [8-1:0] node6535;
	wire [8-1:0] node6538;
	wire [8-1:0] node6540;
	wire [8-1:0] node6543;
	wire [8-1:0] node6546;
	wire [8-1:0] node6547;
	wire [8-1:0] node6548;
	wire [8-1:0] node6549;
	wire [8-1:0] node6550;
	wire [8-1:0] node6554;
	wire [8-1:0] node6555;
	wire [8-1:0] node6556;
	wire [8-1:0] node6559;
	wire [8-1:0] node6563;
	wire [8-1:0] node6564;
	wire [8-1:0] node6565;
	wire [8-1:0] node6566;
	wire [8-1:0] node6568;
	wire [8-1:0] node6571;
	wire [8-1:0] node6574;
	wire [8-1:0] node6575;
	wire [8-1:0] node6577;
	wire [8-1:0] node6580;
	wire [8-1:0] node6583;
	wire [8-1:0] node6586;
	wire [8-1:0] node6587;
	wire [8-1:0] node6588;
	wire [8-1:0] node6589;
	wire [8-1:0] node6590;
	wire [8-1:0] node6591;
	wire [8-1:0] node6595;
	wire [8-1:0] node6597;
	wire [8-1:0] node6600;
	wire [8-1:0] node6601;
	wire [8-1:0] node6603;
	wire [8-1:0] node6606;
	wire [8-1:0] node6609;
	wire [8-1:0] node6612;
	wire [8-1:0] node6613;
	wire [8-1:0] node6614;
	wire [8-1:0] node6615;
	wire [8-1:0] node6618;
	wire [8-1:0] node6619;
	wire [8-1:0] node6622;
	wire [8-1:0] node6624;
	wire [8-1:0] node6627;
	wire [8-1:0] node6628;
	wire [8-1:0] node6630;
	wire [8-1:0] node6633;
	wire [8-1:0] node6634;
	wire [8-1:0] node6638;
	wire [8-1:0] node6641;
	wire [8-1:0] node6642;
	wire [8-1:0] node6644;
	wire [8-1:0] node6645;
	wire [8-1:0] node6646;
	wire [8-1:0] node6647;
	wire [8-1:0] node6649;
	wire [8-1:0] node6652;
	wire [8-1:0] node6653;
	wire [8-1:0] node6655;
	wire [8-1:0] node6658;
	wire [8-1:0] node6660;
	wire [8-1:0] node6663;
	wire [8-1:0] node6664;
	wire [8-1:0] node6665;
	wire [8-1:0] node6667;
	wire [8-1:0] node6670;
	wire [8-1:0] node6671;
	wire [8-1:0] node6673;
	wire [8-1:0] node6676;
	wire [8-1:0] node6678;
	wire [8-1:0] node6681;
	wire [8-1:0] node6682;
	wire [8-1:0] node6684;
	wire [8-1:0] node6687;
	wire [8-1:0] node6688;
	wire [8-1:0] node6690;
	wire [8-1:0] node6692;
	wire [8-1:0] node6695;
	wire [8-1:0] node6697;
	wire [8-1:0] node6700;
	wire [8-1:0] node6701;
	wire [8-1:0] node6702;
	wire [8-1:0] node6703;
	wire [8-1:0] node6705;
	wire [8-1:0] node6708;
	wire [8-1:0] node6710;
	wire [8-1:0] node6713;
	wire [8-1:0] node6714;
	wire [8-1:0] node6715;
	wire [8-1:0] node6717;
	wire [8-1:0] node6720;
	wire [8-1:0] node6721;
	wire [8-1:0] node6724;
	wire [8-1:0] node6726;
	wire [8-1:0] node6729;
	wire [8-1:0] node6730;
	wire [8-1:0] node6732;
	wire [8-1:0] node6735;
	wire [8-1:0] node6737;
	wire [8-1:0] node6739;
	wire [8-1:0] node6742;
	wire [8-1:0] node6743;
	wire [8-1:0] node6744;
	wire [8-1:0] node6746;
	wire [8-1:0] node6749;
	wire [8-1:0] node6750;
	wire [8-1:0] node6752;
	wire [8-1:0] node6755;
	wire [8-1:0] node6756;
	wire [8-1:0] node6758;
	wire [8-1:0] node6762;
	wire [8-1:0] node6763;
	wire [8-1:0] node6764;
	wire [8-1:0] node6766;
	wire [8-1:0] node6769;
	wire [8-1:0] node6772;
	wire [8-1:0] node6773;
	wire [8-1:0] node6775;
	wire [8-1:0] node6778;
	wire [8-1:0] node6780;
	wire [8-1:0] node6782;
	wire [8-1:0] node6785;
	wire [8-1:0] node6786;
	wire [8-1:0] node6787;
	wire [8-1:0] node6788;
	wire [8-1:0] node6790;
	wire [8-1:0] node6792;
	wire [8-1:0] node6795;
	wire [8-1:0] node6796;
	wire [8-1:0] node6798;
	wire [8-1:0] node6799;
	wire [8-1:0] node6803;
	wire [8-1:0] node6804;
	wire [8-1:0] node6805;
	wire [8-1:0] node6809;
	wire [8-1:0] node6812;
	wire [8-1:0] node6813;
	wire [8-1:0] node6814;
	wire [8-1:0] node6816;
	wire [8-1:0] node6818;
	wire [8-1:0] node6821;
	wire [8-1:0] node6822;
	wire [8-1:0] node6824;
	wire [8-1:0] node6827;
	wire [8-1:0] node6830;
	wire [8-1:0] node6831;
	wire [8-1:0] node6832;
	wire [8-1:0] node6833;
	wire [8-1:0] node6836;
	wire [8-1:0] node6837;
	wire [8-1:0] node6841;
	wire [8-1:0] node6844;
	wire [8-1:0] node6847;
	wire [8-1:0] node6848;
	wire [8-1:0] node6849;
	wire [8-1:0] node6850;
	wire [8-1:0] node6852;
	wire [8-1:0] node6855;
	wire [8-1:0] node6856;
	wire [8-1:0] node6857;
	wire [8-1:0] node6860;
	wire [8-1:0] node6864;
	wire [8-1:0] node6865;
	wire [8-1:0] node6866;
	wire [8-1:0] node6867;
	wire [8-1:0] node6870;
	wire [8-1:0] node6874;
	wire [8-1:0] node6875;
	wire [8-1:0] node6876;
	wire [8-1:0] node6878;
	wire [8-1:0] node6881;
	wire [8-1:0] node6882;
	wire [8-1:0] node6887;
	wire [8-1:0] node6888;
	wire [8-1:0] node6889;
	wire [8-1:0] node6890;
	wire [8-1:0] node6891;
	wire [8-1:0] node6894;
	wire [8-1:0] node6898;
	wire [8-1:0] node6899;
	wire [8-1:0] node6900;
	wire [8-1:0] node6901;
	wire [8-1:0] node6904;
	wire [8-1:0] node6907;
	wire [8-1:0] node6911;
	wire [8-1:0] node6912;
	wire [8-1:0] node6913;
	wire [8-1:0] node6914;
	wire [8-1:0] node6915;
	wire [8-1:0] node6916;
	wire [8-1:0] node6921;
	wire [8-1:0] node6922;
	wire [8-1:0] node6925;
	wire [8-1:0] node6928;
	wire [8-1:0] node6929;
	wire [8-1:0] node6932;
	wire [8-1:0] node6935;
	wire [8-1:0] node6938;
	wire [8-1:0] node6939;
	wire [8-1:0] node6941;
	wire [8-1:0] node6942;
	wire [8-1:0] node6943;
	wire [8-1:0] node6944;
	wire [8-1:0] node6946;
	wire [8-1:0] node6949;
	wire [8-1:0] node6950;
	wire [8-1:0] node6952;
	wire [8-1:0] node6955;
	wire [8-1:0] node6956;
	wire [8-1:0] node6958;
	wire [8-1:0] node6961;
	wire [8-1:0] node6963;
	wire [8-1:0] node6966;
	wire [8-1:0] node6967;
	wire [8-1:0] node6968;
	wire [8-1:0] node6970;
	wire [8-1:0] node6973;
	wire [8-1:0] node6974;
	wire [8-1:0] node6976;
	wire [8-1:0] node6979;
	wire [8-1:0] node6980;
	wire [8-1:0] node6982;
	wire [8-1:0] node6985;
	wire [8-1:0] node6988;
	wire [8-1:0] node6989;
	wire [8-1:0] node6990;
	wire [8-1:0] node6992;
	wire [8-1:0] node6995;
	wire [8-1:0] node6996;
	wire [8-1:0] node6999;
	wire [8-1:0] node7001;
	wire [8-1:0] node7004;
	wire [8-1:0] node7005;
	wire [8-1:0] node7007;
	wire [8-1:0] node7010;
	wire [8-1:0] node7011;
	wire [8-1:0] node7015;
	wire [8-1:0] node7016;
	wire [8-1:0] node7017;
	wire [8-1:0] node7018;
	wire [8-1:0] node7020;
	wire [8-1:0] node7023;
	wire [8-1:0] node7024;
	wire [8-1:0] node7026;
	wire [8-1:0] node7029;
	wire [8-1:0] node7030;
	wire [8-1:0] node7032;
	wire [8-1:0] node7035;
	wire [8-1:0] node7037;
	wire [8-1:0] node7040;
	wire [8-1:0] node7041;
	wire [8-1:0] node7042;
	wire [8-1:0] node7044;
	wire [8-1:0] node7047;
	wire [8-1:0] node7048;
	wire [8-1:0] node7051;
	wire [8-1:0] node7054;
	wire [8-1:0] node7055;
	wire [8-1:0] node7057;
	wire [8-1:0] node7058;
	wire [8-1:0] node7062;
	wire [8-1:0] node7063;
	wire [8-1:0] node7065;
	wire [8-1:0] node7068;
	wire [8-1:0] node7069;
	wire [8-1:0] node7072;
	wire [8-1:0] node7075;
	wire [8-1:0] node7076;
	wire [8-1:0] node7077;
	wire [8-1:0] node7078;
	wire [8-1:0] node7080;
	wire [8-1:0] node7083;
	wire [8-1:0] node7085;
	wire [8-1:0] node7087;
	wire [8-1:0] node7090;
	wire [8-1:0] node7091;
	wire [8-1:0] node7092;
	wire [8-1:0] node7094;
	wire [8-1:0] node7097;
	wire [8-1:0] node7098;
	wire [8-1:0] node7101;
	wire [8-1:0] node7103;
	wire [8-1:0] node7106;
	wire [8-1:0] node7107;
	wire [8-1:0] node7109;
	wire [8-1:0] node7112;
	wire [8-1:0] node7114;
	wire [8-1:0] node7116;
	wire [8-1:0] node7119;
	wire [8-1:0] node7120;
	wire [8-1:0] node7121;
	wire [8-1:0] node7123;
	wire [8-1:0] node7126;
	wire [8-1:0] node7127;
	wire [8-1:0] node7131;
	wire [8-1:0] node7132;
	wire [8-1:0] node7134;
	wire [8-1:0] node7136;
	wire [8-1:0] node7139;
	wire [8-1:0] node7140;
	wire [8-1:0] node7142;
	wire [8-1:0] node7145;
	wire [8-1:0] node7148;
	wire [8-1:0] node7149;
	wire [8-1:0] node7150;
	wire [8-1:0] node7151;
	wire [8-1:0] node7153;
	wire [8-1:0] node7154;
	wire [8-1:0] node7158;
	wire [8-1:0] node7159;
	wire [8-1:0] node7160;
	wire [8-1:0] node7161;
	wire [8-1:0] node7163;
	wire [8-1:0] node7166;
	wire [8-1:0] node7168;
	wire [8-1:0] node7171;
	wire [8-1:0] node7173;
	wire [8-1:0] node7176;
	wire [8-1:0] node7177;
	wire [8-1:0] node7180;
	wire [8-1:0] node7183;
	wire [8-1:0] node7184;
	wire [8-1:0] node7185;
	wire [8-1:0] node7186;
	wire [8-1:0] node7187;
	wire [8-1:0] node7189;
	wire [8-1:0] node7190;
	wire [8-1:0] node7194;
	wire [8-1:0] node7195;
	wire [8-1:0] node7199;
	wire [8-1:0] node7200;
	wire [8-1:0] node7201;
	wire [8-1:0] node7204;
	wire [8-1:0] node7206;
	wire [8-1:0] node7209;
	wire [8-1:0] node7210;
	wire [8-1:0] node7214;
	wire [8-1:0] node7215;
	wire [8-1:0] node7216;
	wire [8-1:0] node7220;
	wire [8-1:0] node7221;
	wire [8-1:0] node7222;
	wire [8-1:0] node7225;
	wire [8-1:0] node7226;
	wire [8-1:0] node7230;
	wire [8-1:0] node7231;
	wire [8-1:0] node7235;
	wire [8-1:0] node7236;
	wire [8-1:0] node7237;
	wire [8-1:0] node7240;
	wire [8-1:0] node7243;
	wire [8-1:0] node7244;
	wire [8-1:0] node7247;
	wire [8-1:0] node7250;
	wire [8-1:0] node7251;
	wire [8-1:0] node7252;
	wire [8-1:0] node7253;
	wire [8-1:0] node7254;
	wire [8-1:0] node7255;
	wire [8-1:0] node7256;
	wire [8-1:0] node7257;
	wire [8-1:0] node7260;
	wire [8-1:0] node7264;
	wire [8-1:0] node7265;
	wire [8-1:0] node7268;
	wire [8-1:0] node7270;
	wire [8-1:0] node7273;
	wire [8-1:0] node7274;
	wire [8-1:0] node7276;
	wire [8-1:0] node7279;
	wire [8-1:0] node7281;
	wire [8-1:0] node7282;
	wire [8-1:0] node7286;
	wire [8-1:0] node7287;
	wire [8-1:0] node7288;
	wire [8-1:0] node7289;
	wire [8-1:0] node7290;
	wire [8-1:0] node7294;
	wire [8-1:0] node7295;
	wire [8-1:0] node7299;
	wire [8-1:0] node7301;
	wire [8-1:0] node7304;
	wire [8-1:0] node7305;
	wire [8-1:0] node7306;
	wire [8-1:0] node7307;
	wire [8-1:0] node7311;
	wire [8-1:0] node7314;
	wire [8-1:0] node7315;
	wire [8-1:0] node7318;
	wire [8-1:0] node7319;
	wire [8-1:0] node7323;
	wire [8-1:0] node7324;
	wire [8-1:0] node7325;
	wire [8-1:0] node7326;
	wire [8-1:0] node7330;
	wire [8-1:0] node7331;
	wire [8-1:0] node7332;
	wire [8-1:0] node7333;
	wire [8-1:0] node7337;
	wire [8-1:0] node7339;
	wire [8-1:0] node7342;
	wire [8-1:0] node7343;
	wire [8-1:0] node7347;
	wire [8-1:0] node7348;
	wire [8-1:0] node7349;
	wire [8-1:0] node7350;
	wire [8-1:0] node7352;
	wire [8-1:0] node7355;
	wire [8-1:0] node7356;
	wire [8-1:0] node7360;
	wire [8-1:0] node7361;
	wire [8-1:0] node7362;
	wire [8-1:0] node7363;
	wire [8-1:0] node7367;
	wire [8-1:0] node7370;
	wire [8-1:0] node7371;
	wire [8-1:0] node7375;
	wire [8-1:0] node7376;
	wire [8-1:0] node7377;
	wire [8-1:0] node7378;
	wire [8-1:0] node7382;
	wire [8-1:0] node7384;
	wire [8-1:0] node7387;
	wire [8-1:0] node7389;
	wire [8-1:0] node7390;
	wire [8-1:0] node7394;
	wire [8-1:0] node7395;
	wire [8-1:0] node7396;
	wire [8-1:0] node7397;
	wire [8-1:0] node7398;
	wire [8-1:0] node7401;
	wire [8-1:0] node7404;
	wire [8-1:0] node7405;
	wire [8-1:0] node7408;
	wire [8-1:0] node7411;
	wire [8-1:0] node7412;
	wire [8-1:0] node7413;
	wire [8-1:0] node7416;
	wire [8-1:0] node7419;
	wire [8-1:0] node7420;
	wire [8-1:0] node7423;
	wire [8-1:0] node7426;
	wire [8-1:0] node7427;
	wire [8-1:0] node7428;
	wire [8-1:0] node7429;
	wire [8-1:0] node7430;
	wire [8-1:0] node7433;
	wire [8-1:0] node7436;
	wire [8-1:0] node7437;
	wire [8-1:0] node7440;
	wire [8-1:0] node7443;
	wire [8-1:0] node7444;
	wire [8-1:0] node7445;
	wire [8-1:0] node7448;
	wire [8-1:0] node7451;
	wire [8-1:0] node7452;
	wire [8-1:0] node7455;
	wire [8-1:0] node7458;
	wire [8-1:0] node7459;
	wire [8-1:0] node7460;
	wire [8-1:0] node7461;
	wire [8-1:0] node7464;
	wire [8-1:0] node7467;
	wire [8-1:0] node7468;
	wire [8-1:0] node7471;
	wire [8-1:0] node7474;
	wire [8-1:0] node7475;
	wire [8-1:0] node7476;
	wire [8-1:0] node7479;
	wire [8-1:0] node7482;
	wire [8-1:0] node7483;
	wire [8-1:0] node7486;

	assign outp = (inp[4]) ? node3742 : node1;
		assign node1 = (inp[13]) ? node1765 : node2;
			assign node2 = (inp[7]) ? node386 : node3;
				assign node3 = (inp[11]) ? node125 : node4;
					assign node4 = (inp[0]) ? node70 : node5;
						assign node5 = (inp[1]) ? node29 : node6;
							assign node6 = (inp[8]) ? node14 : node7;
								assign node7 = (inp[2]) ? node9 : 8'b01111111;
									assign node9 = (inp[5]) ? node11 : 8'b00101111;
										assign node11 = (inp[6]) ? 8'b01111111 : 8'b00101111;
								assign node14 = (inp[2]) ? node20 : node15;
									assign node15 = (inp[5]) ? node17 : 8'b00111011;
										assign node17 = (inp[10]) ? 8'b01111111 : 8'b00111011;
									assign node20 = (inp[5]) ? node22 : 8'b00101011;
										assign node22 = (inp[10]) ? node26 : node23;
											assign node23 = (inp[6]) ? 8'b00111011 : 8'b00101011;
											assign node26 = (inp[6]) ? 8'b01111111 : 8'b00101111;
							assign node29 = (inp[2]) ? node45 : node30;
								assign node30 = (inp[8]) ? node36 : node31;
									assign node31 = (inp[5]) ? node33 : 8'b00111110;
										assign node33 = (inp[3]) ? 8'b01111111 : 8'b00111110;
									assign node36 = (inp[5]) ? node38 : 8'b00111010;
										assign node38 = (inp[10]) ? node42 : node39;
											assign node39 = (inp[3]) ? 8'b00111011 : 8'b00111010;
											assign node42 = (inp[3]) ? 8'b01111111 : 8'b00111110;
								assign node45 = (inp[8]) ? node55 : node46;
									assign node46 = (inp[5]) ? node48 : 8'b00101110;
										assign node48 = (inp[6]) ? node52 : node49;
											assign node49 = (inp[3]) ? 8'b00101111 : 8'b00101110;
											assign node52 = (inp[3]) ? 8'b01111111 : 8'b00111110;
									assign node55 = (inp[5]) ? node57 : 8'b00101010;
										assign node57 = (inp[6]) ? node65 : node58;
											assign node58 = (inp[10]) ? node62 : node59;
												assign node59 = (inp[3]) ? 8'b00101011 : 8'b00101010;
												assign node62 = (inp[3]) ? 8'b00101111 : 8'b00101110;
											assign node65 = (inp[10]) ? 8'b00111110 : node66;
												assign node66 = (inp[3]) ? 8'b00111011 : 8'b00111010;
						assign node70 = (inp[5]) ? 8'b01111111 : node71;
							assign node71 = (inp[3]) ? node89 : node72;
								assign node72 = (inp[2]) ? node78 : node73;
									assign node73 = (inp[8]) ? node75 : 8'b01111111;
										assign node75 = (inp[10]) ? 8'b00111011 : 8'b01111111;
									assign node78 = (inp[6]) ? node84 : node79;
										assign node79 = (inp[10]) ? node81 : 8'b01111111;
											assign node81 = (inp[8]) ? 8'b00111011 : 8'b01111111;
										assign node84 = (inp[8]) ? node86 : 8'b00101111;
											assign node86 = (inp[10]) ? 8'b00101011 : 8'b00101111;
								assign node89 = (inp[1]) ? node107 : node90;
									assign node90 = (inp[8]) ? node96 : node91;
										assign node91 = (inp[6]) ? node93 : 8'b01111111;
											assign node93 = (inp[2]) ? 8'b00101111 : 8'b01111111;
										assign node96 = (inp[10]) ? node102 : node97;
											assign node97 = (inp[2]) ? node99 : 8'b01111111;
												assign node99 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node102 = (inp[6]) ? node104 : 8'b00111011;
												assign node104 = (inp[2]) ? 8'b00101011 : 8'b00111011;
									assign node107 = (inp[10]) ? node113 : node108;
										assign node108 = (inp[6]) ? node110 : 8'b00111110;
											assign node110 = (inp[2]) ? 8'b00101110 : 8'b00111110;
										assign node113 = (inp[8]) ? node119 : node114;
											assign node114 = (inp[6]) ? node116 : 8'b00111110;
												assign node116 = (inp[2]) ? 8'b00101110 : 8'b00111110;
											assign node119 = (inp[2]) ? node121 : 8'b00111010;
												assign node121 = (inp[6]) ? 8'b00101010 : 8'b00111010;
					assign node125 = (inp[8]) ? node219 : node126;
						assign node126 = (inp[1]) ? node154 : node127;
							assign node127 = (inp[2]) ? node131 : node128;
								assign node128 = (inp[12]) ? 8'b01111111 : 8'b00101111;
								assign node131 = (inp[12]) ? node143 : node132;
									assign node132 = (inp[5]) ? node138 : node133;
										assign node133 = (inp[6]) ? 8'b00111110 : node134;
											assign node134 = (inp[0]) ? 8'b00101110 : 8'b00111110;
										assign node138 = (inp[0]) ? 8'b00101110 : node139;
											assign node139 = (inp[6]) ? 8'b00101110 : 8'b00111110;
									assign node143 = (inp[5]) ? node149 : node144;
										assign node144 = (inp[6]) ? 8'b00101111 : node145;
											assign node145 = (inp[0]) ? 8'b00111110 : 8'b00101111;
										assign node149 = (inp[0]) ? 8'b00111110 : node150;
											assign node150 = (inp[6]) ? 8'b00111110 : 8'b00101111;
							assign node154 = (inp[12]) ? node188 : node155;
								assign node155 = (inp[2]) ? node167 : node156;
									assign node156 = (inp[5]) ? node162 : node157;
										assign node157 = (inp[0]) ? node159 : 8'b00101110;
											assign node159 = (inp[3]) ? 8'b00101110 : 8'b00101011;
										assign node162 = (inp[0]) ? 8'b00101011 : node163;
											assign node163 = (inp[3]) ? 8'b00101011 : 8'b00101110;
									assign node167 = (inp[5]) ? node179 : node168;
										assign node168 = (inp[3]) ? node174 : node169;
											assign node169 = (inp[0]) ? node171 : 8'b00111011;
												assign node171 = (inp[6]) ? 8'b00111010 : 8'b00101010;
											assign node174 = (inp[0]) ? node176 : 8'b00111011;
												assign node176 = (inp[6]) ? 8'b00111011 : 8'b00101011;
										assign node179 = (inp[0]) ? 8'b00101010 : node180;
											assign node180 = (inp[6]) ? node184 : node181;
												assign node181 = (inp[3]) ? 8'b00111010 : 8'b00111011;
												assign node184 = (inp[3]) ? 8'b00101010 : 8'b00101011;
								assign node188 = (inp[0]) ? node204 : node189;
									assign node189 = (inp[2]) ? node195 : node190;
										assign node190 = (inp[5]) ? node192 : 8'b00111110;
											assign node192 = (inp[3]) ? 8'b00111011 : 8'b00111110;
										assign node195 = (inp[5]) ? node197 : 8'b00101110;
											assign node197 = (inp[6]) ? node201 : node198;
												assign node198 = (inp[3]) ? 8'b00101011 : 8'b00101110;
												assign node201 = (inp[3]) ? 8'b00111010 : 8'b00111011;
									assign node204 = (inp[2]) ? node210 : node205;
										assign node205 = (inp[3]) ? node207 : 8'b00111011;
											assign node207 = (inp[5]) ? 8'b00111011 : 8'b00111110;
										assign node210 = (inp[5]) ? 8'b00111010 : node211;
											assign node211 = (inp[6]) ? node215 : node212;
												assign node212 = (inp[3]) ? 8'b00111011 : 8'b00111010;
												assign node215 = (inp[3]) ? 8'b00101110 : 8'b00101011;
						assign node219 = (inp[12]) ? node299 : node220;
							assign node220 = (inp[2]) ? node252 : node221;
								assign node221 = (inp[0]) ? node237 : node222;
									assign node222 = (inp[1]) ? node228 : node223;
										assign node223 = (inp[10]) ? node225 : 8'b00101011;
											assign node225 = (inp[5]) ? 8'b00001111 : 8'b00101011;
										assign node228 = (inp[5]) ? node230 : 8'b00101010;
											assign node230 = (inp[3]) ? node234 : node231;
												assign node231 = (inp[10]) ? 8'b00001110 : 8'b00101010;
												assign node234 = (inp[10]) ? 8'b00001011 : 8'b00001111;
									assign node237 = (inp[1]) ? node243 : node238;
										assign node238 = (inp[5]) ? 8'b00001111 : node239;
											assign node239 = (inp[10]) ? 8'b00101011 : 8'b00001111;
										assign node243 = (inp[5]) ? 8'b00001011 : node244;
											assign node244 = (inp[3]) ? node248 : node245;
												assign node245 = (inp[10]) ? 8'b00001111 : 8'b00001011;
												assign node248 = (inp[10]) ? 8'b00101010 : 8'b00001110;
								assign node252 = (inp[1]) ? node272 : node253;
									assign node253 = (inp[0]) ? node263 : node254;
										assign node254 = (inp[5]) ? node256 : 8'b00111010;
											assign node256 = (inp[10]) ? node260 : node257;
												assign node257 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node260 = (inp[6]) ? 8'b00001110 : 8'b00011110;
										assign node263 = (inp[5]) ? 8'b00001110 : node264;
											assign node264 = (inp[10]) ? node268 : node265;
												assign node265 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node268 = (inp[6]) ? 8'b00111010 : 8'b00101010;
									assign node272 = (inp[0]) ? node290 : node273;
										assign node273 = (inp[5]) ? node275 : 8'b00011111;
											assign node275 = (inp[6]) ? node283 : node276;
												assign node276 = (inp[3]) ? node280 : node277;
													assign node277 = (inp[10]) ? 8'b00011011 : 8'b00011111;
													assign node280 = (inp[10]) ? 8'b00011010 : 8'b00011110;
												assign node283 = (inp[10]) ? node287 : node284;
													assign node284 = (inp[3]) ? 8'b00001110 : 8'b00001111;
													assign node287 = (inp[3]) ? 8'b00001010 : 8'b00001011;
										assign node290 = (inp[5]) ? 8'b00001010 : node291;
											assign node291 = (inp[10]) ? node293 : 8'b00011010;
												assign node293 = (inp[6]) ? 8'b00011111 : node294;
													assign node294 = (inp[3]) ? 8'b00001111 : 8'b00001110;
							assign node299 = (inp[5]) ? node345 : node300;
								assign node300 = (inp[2]) ? node318 : node301;
									assign node301 = (inp[0]) ? node305 : node302;
										assign node302 = (inp[1]) ? 8'b00111010 : 8'b00111011;
										assign node305 = (inp[10]) ? node311 : node306;
											assign node306 = (inp[1]) ? node308 : 8'b00011111;
												assign node308 = (inp[3]) ? 8'b00011110 : 8'b00011011;
											assign node311 = (inp[3]) ? node315 : node312;
												assign node312 = (inp[1]) ? 8'b00011111 : 8'b00111011;
												assign node315 = (inp[1]) ? 8'b00111010 : 8'b00111011;
									assign node318 = (inp[0]) ? node322 : node319;
										assign node319 = (inp[1]) ? 8'b00101010 : 8'b00101011;
										assign node322 = (inp[6]) ? node332 : node323;
											assign node323 = (inp[1]) ? node327 : node324;
												assign node324 = (inp[10]) ? 8'b00111010 : 8'b00011110;
												assign node327 = (inp[10]) ? 8'b00011110 : node328;
													assign node328 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node332 = (inp[10]) ? node340 : node333;
												assign node333 = (inp[3]) ? node337 : node334;
													assign node334 = (inp[1]) ? 8'b00001011 : 8'b00001111;
													assign node337 = (inp[1]) ? 8'b00001110 : 8'b00001111;
												assign node340 = (inp[1]) ? node342 : 8'b00101011;
													assign node342 = (inp[9]) ? 8'b00101010 : 8'b00001111;
								assign node345 = (inp[2]) ? node361 : node346;
									assign node346 = (inp[1]) ? node352 : node347;
										assign node347 = (inp[10]) ? 8'b00011111 : node348;
											assign node348 = (inp[0]) ? 8'b00011111 : 8'b00111011;
										assign node352 = (inp[0]) ? 8'b00011011 : node353;
											assign node353 = (inp[3]) ? node357 : node354;
												assign node354 = (inp[10]) ? 8'b00011110 : 8'b00111010;
												assign node357 = (inp[6]) ? 8'b00011011 : 8'b00011111;
									assign node361 = (inp[0]) ? node383 : node362;
										assign node362 = (inp[6]) ? node372 : node363;
											assign node363 = (inp[10]) ? node367 : node364;
												assign node364 = (inp[1]) ? 8'b00101010 : 8'b00101011;
												assign node367 = (inp[1]) ? node369 : 8'b00001111;
													assign node369 = (inp[3]) ? 8'b00001011 : 8'b00001110;
											assign node372 = (inp[1]) ? node376 : node373;
												assign node373 = (inp[10]) ? 8'b00011110 : 8'b00111010;
												assign node376 = (inp[3]) ? node380 : node377;
													assign node377 = (inp[10]) ? 8'b00011011 : 8'b00011111;
													assign node380 = (inp[10]) ? 8'b00011010 : 8'b00011110;
										assign node383 = (inp[1]) ? 8'b00011010 : 8'b00011110;
				assign node386 = (inp[9]) ? node1098 : node387;
					assign node387 = (inp[11]) ? node663 : node388;
						assign node388 = (inp[3]) ? node526 : node389;
							assign node389 = (inp[0]) ? node501 : node390;
								assign node390 = (inp[1]) ? node452 : node391;
									assign node391 = (inp[5]) ? node403 : node392;
										assign node392 = (inp[10]) ? node398 : node393;
											assign node393 = (inp[8]) ? 8'b00101011 : node394;
												assign node394 = (inp[2]) ? 8'b00101111 : 8'b01111111;
											assign node398 = (inp[6]) ? 8'b00101011 : node399;
												assign node399 = (inp[2]) ? 8'b00101011 : 8'b00111011;
										assign node403 = (inp[12]) ? node427 : node404;
											assign node404 = (inp[8]) ? node414 : node405;
												assign node405 = (inp[10]) ? node407 : 8'b00101111;
													assign node407 = (inp[2]) ? node411 : node408;
														assign node408 = (inp[6]) ? 8'b00101011 : 8'b00111011;
														assign node411 = (inp[6]) ? 8'b00111011 : 8'b00101011;
												assign node414 = (inp[10]) ? node422 : node415;
													assign node415 = (inp[6]) ? node419 : node416;
														assign node416 = (inp[2]) ? 8'b00101011 : 8'b00111011;
														assign node419 = (inp[2]) ? 8'b00111011 : 8'b00101011;
													assign node422 = (inp[2]) ? 8'b01111111 : node423;
														assign node423 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node427 = (inp[2]) ? node443 : node428;
												assign node428 = (inp[6]) ? node436 : node429;
													assign node429 = (inp[8]) ? node433 : node430;
														assign node430 = (inp[10]) ? 8'b00111011 : 8'b01111111;
														assign node433 = (inp[10]) ? 8'b01111111 : 8'b00111011;
													assign node436 = (inp[10]) ? node440 : node437;
														assign node437 = (inp[8]) ? 8'b00101011 : 8'b00101111;
														assign node440 = (inp[8]) ? 8'b00101111 : 8'b00101011;
												assign node443 = (inp[6]) ? node445 : 8'b00101111;
													assign node445 = (inp[10]) ? node449 : node446;
														assign node446 = (inp[8]) ? 8'b00111011 : 8'b01111111;
														assign node449 = (inp[8]) ? 8'b01111111 : 8'b00111011;
									assign node452 = (inp[5]) ? node468 : node453;
										assign node453 = (inp[10]) ? node463 : node454;
											assign node454 = (inp[8]) ? node458 : node455;
												assign node455 = (inp[2]) ? 8'b00101110 : 8'b00111110;
												assign node458 = (inp[2]) ? 8'b00101010 : node459;
													assign node459 = (inp[12]) ? 8'b00101010 : 8'b00111010;
											assign node463 = (inp[2]) ? 8'b00101010 : node464;
												assign node464 = (inp[6]) ? 8'b00101010 : 8'b00111010;
										assign node468 = (inp[8]) ? node488 : node469;
											assign node469 = (inp[10]) ? node475 : node470;
												assign node470 = (inp[2]) ? node472 : 8'b00101110;
													assign node472 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node475 = (inp[12]) ? node481 : node476;
													assign node476 = (inp[6]) ? 8'b00101010 : node477;
														assign node477 = (inp[2]) ? 8'b00101010 : 8'b00111010;
													assign node481 = (inp[6]) ? node485 : node482;
														assign node482 = (inp[2]) ? 8'b00101010 : 8'b00111010;
														assign node485 = (inp[2]) ? 8'b00111010 : 8'b00101010;
											assign node488 = (inp[10]) ? node494 : node489;
												assign node489 = (inp[2]) ? 8'b00111010 : node490;
													assign node490 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node494 = (inp[6]) ? node498 : node495;
													assign node495 = (inp[2]) ? 8'b00101110 : 8'b00111110;
													assign node498 = (inp[2]) ? 8'b00111110 : 8'b00101110;
								assign node501 = (inp[10]) ? node509 : node502;
									assign node502 = (inp[6]) ? node504 : 8'b01111111;
										assign node504 = (inp[5]) ? node506 : 8'b00101111;
											assign node506 = (inp[2]) ? 8'b01111111 : 8'b00101111;
									assign node509 = (inp[6]) ? node515 : node510;
										assign node510 = (inp[5]) ? node512 : 8'b00111011;
											assign node512 = (inp[8]) ? 8'b01111111 : 8'b00111011;
										assign node515 = (inp[2]) ? node521 : node516;
											assign node516 = (inp[5]) ? node518 : 8'b00101011;
												assign node518 = (inp[8]) ? 8'b00101111 : 8'b00101011;
											assign node521 = (inp[5]) ? node523 : 8'b00101011;
												assign node523 = (inp[8]) ? 8'b01111111 : 8'b00111011;
							assign node526 = (inp[5]) ? node550 : node527;
								assign node527 = (inp[10]) ? node543 : node528;
									assign node528 = (inp[6]) ? node538 : node529;
										assign node529 = (inp[0]) ? 8'b00111110 : node530;
											assign node530 = (inp[8]) ? node534 : node531;
												assign node531 = (inp[2]) ? 8'b00101110 : 8'b00111110;
												assign node534 = (inp[2]) ? 8'b00101010 : 8'b00111010;
										assign node538 = (inp[8]) ? node540 : 8'b00101110;
											assign node540 = (inp[0]) ? 8'b00101110 : 8'b00101010;
									assign node543 = (inp[6]) ? 8'b00101010 : node544;
										assign node544 = (inp[0]) ? 8'b00111010 : node545;
											assign node545 = (inp[2]) ? 8'b00101010 : 8'b00111010;
								assign node550 = (inp[1]) ? node612 : node551;
									assign node551 = (inp[0]) ? node593 : node552;
										assign node552 = (inp[8]) ? node574 : node553;
											assign node553 = (inp[10]) ? node559 : node554;
												assign node554 = (inp[2]) ? node556 : 8'b00111110;
													assign node556 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node559 = (inp[12]) ? node567 : node560;
													assign node560 = (inp[2]) ? node564 : node561;
														assign node561 = (inp[6]) ? 8'b00101010 : 8'b00111010;
														assign node564 = (inp[6]) ? 8'b00111010 : 8'b00101010;
													assign node567 = (inp[6]) ? node571 : node568;
														assign node568 = (inp[2]) ? 8'b00101010 : 8'b00111010;
														assign node571 = (inp[2]) ? 8'b00111010 : 8'b00101010;
											assign node574 = (inp[10]) ? node588 : node575;
												assign node575 = (inp[12]) ? node581 : node576;
													assign node576 = (inp[6]) ? 8'b00111010 : node577;
														assign node577 = (inp[2]) ? 8'b00101010 : 8'b00111010;
													assign node581 = (inp[2]) ? node585 : node582;
														assign node582 = (inp[6]) ? 8'b00101010 : 8'b00111010;
														assign node585 = (inp[6]) ? 8'b00111010 : 8'b00101010;
												assign node588 = (inp[2]) ? 8'b00111110 : node589;
													assign node589 = (inp[6]) ? 8'b00101110 : 8'b00111110;
										assign node593 = (inp[10]) ? node599 : node594;
											assign node594 = (inp[6]) ? node596 : 8'b00111110;
												assign node596 = (inp[2]) ? 8'b00111110 : 8'b00101110;
											assign node599 = (inp[8]) ? node605 : node600;
												assign node600 = (inp[6]) ? node602 : 8'b00111010;
													assign node602 = (inp[2]) ? 8'b00111010 : 8'b00101010;
												assign node605 = (inp[12]) ? 8'b00111110 : node606;
													assign node606 = (inp[2]) ? 8'b00111110 : node607;
														assign node607 = (inp[6]) ? 8'b00101110 : 8'b00111110;
									assign node612 = (inp[0]) ? node646 : node613;
										assign node613 = (inp[8]) ? node627 : node614;
											assign node614 = (inp[10]) ? node622 : node615;
												assign node615 = (inp[2]) ? node619 : node616;
													assign node616 = (inp[6]) ? 8'b00101111 : 8'b01111111;
													assign node619 = (inp[6]) ? 8'b01111111 : 8'b00101111;
												assign node622 = (inp[6]) ? node624 : 8'b00111011;
													assign node624 = (inp[2]) ? 8'b00111011 : 8'b00101011;
											assign node627 = (inp[10]) ? node641 : node628;
												assign node628 = (inp[12]) ? node636 : node629;
													assign node629 = (inp[6]) ? node633 : node630;
														assign node630 = (inp[2]) ? 8'b00101011 : 8'b00111011;
														assign node633 = (inp[2]) ? 8'b00111011 : 8'b00101011;
													assign node636 = (inp[6]) ? 8'b00111011 : node637;
														assign node637 = (inp[2]) ? 8'b00101011 : 8'b00111011;
												assign node641 = (inp[2]) ? 8'b00101111 : node642;
													assign node642 = (inp[6]) ? 8'b00101111 : 8'b01111111;
										assign node646 = (inp[8]) ? node658 : node647;
											assign node647 = (inp[10]) ? node653 : node648;
												assign node648 = (inp[2]) ? 8'b01111111 : node649;
													assign node649 = (inp[6]) ? 8'b00101111 : 8'b01111111;
												assign node653 = (inp[2]) ? 8'b00111011 : node654;
													assign node654 = (inp[6]) ? 8'b00101011 : 8'b00111011;
											assign node658 = (inp[6]) ? node660 : 8'b01111111;
												assign node660 = (inp[2]) ? 8'b01111111 : 8'b00101111;
						assign node663 = (inp[8]) ? node879 : node664;
							assign node664 = (inp[10]) ? node776 : node665;
								assign node665 = (inp[1]) ? node709 : node666;
									assign node666 = (inp[3]) ? node688 : node667;
										assign node667 = (inp[2]) ? node675 : node668;
											assign node668 = (inp[12]) ? node672 : node669;
												assign node669 = (inp[6]) ? 8'b00111110 : 8'b00101111;
												assign node672 = (inp[6]) ? 8'b00101111 : 8'b01111111;
											assign node675 = (inp[0]) ? node683 : node676;
												assign node676 = (inp[5]) ? node678 : 8'b00101111;
													assign node678 = (inp[6]) ? node680 : 8'b00101111;
														assign node680 = (inp[12]) ? 8'b00111110 : 8'b00101110;
												assign node683 = (inp[12]) ? 8'b00111110 : node684;
													assign node684 = (inp[6]) ? 8'b00111110 : 8'b00101110;
										assign node688 = (inp[12]) ? node702 : node689;
											assign node689 = (inp[0]) ? node697 : node690;
												assign node690 = (inp[2]) ? node692 : 8'b00111011;
													assign node692 = (inp[6]) ? node694 : 8'b00111011;
														assign node694 = (inp[5]) ? 8'b00101011 : 8'b00111011;
												assign node697 = (inp[2]) ? 8'b00101011 : node698;
													assign node698 = (inp[6]) ? 8'b00111011 : 8'b00101110;
											assign node702 = (inp[6]) ? 8'b00101110 : node703;
												assign node703 = (inp[2]) ? node705 : 8'b00111110;
													assign node705 = (inp[5]) ? 8'b00111011 : 8'b00101110;
									assign node709 = (inp[12]) ? node739 : node710;
										assign node710 = (inp[6]) ? node724 : node711;
											assign node711 = (inp[2]) ? node719 : node712;
												assign node712 = (inp[0]) ? 8'b00101011 : node713;
													assign node713 = (inp[3]) ? node715 : 8'b00101110;
														assign node715 = (inp[5]) ? 8'b00101011 : 8'b00101110;
												assign node719 = (inp[0]) ? 8'b00101010 : node720;
													assign node720 = (inp[3]) ? 8'b00111010 : 8'b00111011;
											assign node724 = (inp[2]) ? node732 : node725;
												assign node725 = (inp[0]) ? node727 : 8'b00111011;
													assign node727 = (inp[3]) ? node729 : 8'b00111010;
														assign node729 = (inp[5]) ? 8'b00111010 : 8'b00111011;
												assign node732 = (inp[5]) ? node734 : 8'b00111011;
													assign node734 = (inp[3]) ? 8'b00101010 : node735;
														assign node735 = (inp[0]) ? 8'b00101010 : 8'b00101011;
										assign node739 = (inp[5]) ? node755 : node740;
											assign node740 = (inp[6]) ? node750 : node741;
												assign node741 = (inp[0]) ? node745 : node742;
													assign node742 = (inp[2]) ? 8'b00101110 : 8'b00111110;
													assign node745 = (inp[2]) ? node747 : 8'b00111110;
														assign node747 = (inp[3]) ? 8'b00111011 : 8'b00111010;
												assign node750 = (inp[3]) ? 8'b00101110 : node751;
													assign node751 = (inp[0]) ? 8'b00101011 : 8'b00101110;
											assign node755 = (inp[3]) ? node767 : node756;
												assign node756 = (inp[0]) ? node764 : node757;
													assign node757 = (inp[6]) ? node761 : node758;
														assign node758 = (inp[2]) ? 8'b00101110 : 8'b00111110;
														assign node761 = (inp[2]) ? 8'b00111011 : 8'b00101110;
													assign node764 = (inp[2]) ? 8'b00111010 : 8'b00101011;
												assign node767 = (inp[2]) ? node771 : node768;
													assign node768 = (inp[6]) ? 8'b00101011 : 8'b00111011;
													assign node771 = (inp[0]) ? 8'b00111010 : node772;
														assign node772 = (inp[6]) ? 8'b00111010 : 8'b00101011;
								assign node776 = (inp[1]) ? node820 : node777;
									assign node777 = (inp[3]) ? node801 : node778;
										assign node778 = (inp[0]) ? node792 : node779;
											assign node779 = (inp[2]) ? node785 : node780;
												assign node780 = (inp[12]) ? node782 : 8'b00101011;
													assign node782 = (inp[6]) ? 8'b00101011 : 8'b00111011;
												assign node785 = (inp[12]) ? node787 : 8'b00111010;
													assign node787 = (inp[5]) ? node789 : 8'b00101011;
														assign node789 = (inp[6]) ? 8'b00111010 : 8'b00101011;
											assign node792 = (inp[5]) ? node794 : 8'b00111010;
												assign node794 = (inp[2]) ? node798 : node795;
													assign node795 = (inp[6]) ? 8'b00101011 : 8'b00111011;
													assign node798 = (inp[12]) ? 8'b00111010 : 8'b00101010;
										assign node801 = (inp[12]) ? node811 : node802;
											assign node802 = (inp[6]) ? node808 : node803;
												assign node803 = (inp[2]) ? node805 : 8'b00101010;
													assign node805 = (inp[0]) ? 8'b00001111 : 8'b00011111;
												assign node808 = (inp[5]) ? 8'b00001111 : 8'b00011111;
											assign node811 = (inp[2]) ? node815 : node812;
												assign node812 = (inp[6]) ? 8'b00101010 : 8'b00111010;
												assign node815 = (inp[0]) ? node817 : 8'b00101010;
													assign node817 = (inp[5]) ? 8'b00011111 : 8'b00101010;
									assign node820 = (inp[12]) ? node842 : node821;
										assign node821 = (inp[6]) ? node833 : node822;
											assign node822 = (inp[2]) ? node830 : node823;
												assign node823 = (inp[3]) ? node827 : node824;
													assign node824 = (inp[0]) ? 8'b00001111 : 8'b00101010;
													assign node827 = (inp[5]) ? 8'b00001111 : 8'b00101010;
												assign node830 = (inp[0]) ? 8'b00001110 : 8'b00011111;
											assign node833 = (inp[5]) ? node839 : node834;
												assign node834 = (inp[0]) ? node836 : 8'b00011111;
													assign node836 = (inp[3]) ? 8'b00011111 : 8'b00011110;
												assign node839 = (inp[0]) ? 8'b00011110 : 8'b00001110;
										assign node842 = (inp[5]) ? node856 : node843;
											assign node843 = (inp[0]) ? node847 : node844;
												assign node844 = (inp[2]) ? 8'b00101010 : 8'b00111010;
												assign node847 = (inp[3]) ? node851 : node848;
													assign node848 = (inp[6]) ? 8'b00001111 : 8'b00011111;
													assign node851 = (inp[6]) ? 8'b00101010 : node852;
														assign node852 = (inp[2]) ? 8'b00011111 : 8'b00111010;
											assign node856 = (inp[3]) ? node870 : node857;
												assign node857 = (inp[0]) ? node865 : node858;
													assign node858 = (inp[6]) ? node862 : node859;
														assign node859 = (inp[2]) ? 8'b00101010 : 8'b00111010;
														assign node862 = (inp[2]) ? 8'b00011111 : 8'b00101010;
													assign node865 = (inp[6]) ? 8'b00001111 : node866;
														assign node866 = (inp[2]) ? 8'b00011110 : 8'b00011111;
												assign node870 = (inp[2]) ? node874 : node871;
													assign node871 = (inp[6]) ? 8'b00001111 : 8'b00011111;
													assign node874 = (inp[0]) ? 8'b00011110 : node875;
														assign node875 = (inp[6]) ? 8'b00011110 : 8'b00001111;
							assign node879 = (inp[5]) ? node981 : node880;
								assign node880 = (inp[0]) ? node914 : node881;
									assign node881 = (inp[12]) ? node899 : node882;
										assign node882 = (inp[6]) ? node894 : node883;
											assign node883 = (inp[2]) ? node889 : node884;
												assign node884 = (inp[1]) ? 8'b00101010 : node885;
													assign node885 = (inp[3]) ? 8'b00101010 : 8'b00101011;
												assign node889 = (inp[3]) ? 8'b00011111 : node890;
													assign node890 = (inp[1]) ? 8'b00011111 : 8'b00111010;
											assign node894 = (inp[3]) ? 8'b00011111 : node895;
												assign node895 = (inp[1]) ? 8'b00011111 : 8'b00111010;
										assign node899 = (inp[2]) ? node909 : node900;
											assign node900 = (inp[6]) ? node906 : node901;
												assign node901 = (inp[10]) ? node903 : 8'b00111010;
													assign node903 = (inp[1]) ? 8'b00111010 : 8'b00111011;
												assign node906 = (inp[1]) ? 8'b00101010 : 8'b00101011;
											assign node909 = (inp[1]) ? 8'b00101010 : node910;
												assign node910 = (inp[3]) ? 8'b00101010 : 8'b00101011;
									assign node914 = (inp[10]) ? node952 : node915;
										assign node915 = (inp[1]) ? node929 : node916;
											assign node916 = (inp[2]) ? node920 : node917;
												assign node917 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node920 = (inp[3]) ? 8'b00001011 : node921;
													assign node921 = (inp[12]) ? node925 : node922;
														assign node922 = (inp[6]) ? 8'b00011110 : 8'b00001110;
														assign node925 = (inp[6]) ? 8'b00001111 : 8'b00011110;
											assign node929 = (inp[3]) ? node943 : node930;
												assign node930 = (inp[2]) ? node938 : node931;
													assign node931 = (inp[12]) ? node935 : node932;
														assign node932 = (inp[6]) ? 8'b00011010 : 8'b00001011;
														assign node935 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node938 = (inp[12]) ? 8'b00011010 : node939;
														assign node939 = (inp[6]) ? 8'b00011010 : 8'b00001010;
												assign node943 = (inp[12]) ? node947 : node944;
													assign node944 = (inp[6]) ? 8'b00011011 : 8'b00001011;
													assign node947 = (inp[2]) ? 8'b00011011 : node948;
														assign node948 = (inp[6]) ? 8'b00001110 : 8'b00011110;
										assign node952 = (inp[12]) ? node972 : node953;
											assign node953 = (inp[6]) ? node967 : node954;
												assign node954 = (inp[1]) ? node962 : node955;
													assign node955 = (inp[2]) ? node959 : node956;
														assign node956 = (inp[3]) ? 8'b00101010 : 8'b00101011;
														assign node959 = (inp[3]) ? 8'b00001111 : 8'b00101010;
													assign node962 = (inp[3]) ? 8'b00101010 : node963;
														assign node963 = (inp[2]) ? 8'b00001110 : 8'b00001111;
												assign node967 = (inp[2]) ? node969 : 8'b00011111;
													assign node969 = (inp[1]) ? 8'b00011110 : 8'b00111010;
											assign node972 = (inp[6]) ? node978 : node973;
												assign node973 = (inp[3]) ? node975 : 8'b00111010;
													assign node975 = (inp[2]) ? 8'b00011111 : 8'b00111010;
												assign node978 = (inp[3]) ? 8'b00101010 : 8'b00101011;
								assign node981 = (inp[1]) ? node1057 : node982;
									assign node982 = (inp[10]) ? node1028 : node983;
										assign node983 = (inp[0]) ? node1009 : node984;
											assign node984 = (inp[3]) ? node998 : node985;
												assign node985 = (inp[6]) ? node993 : node986;
													assign node986 = (inp[12]) ? node990 : node987;
														assign node987 = (inp[2]) ? 8'b00111010 : 8'b00101011;
														assign node990 = (inp[2]) ? 8'b00101011 : 8'b00111011;
													assign node993 = (inp[12]) ? 8'b00111010 : node994;
														assign node994 = (inp[2]) ? 8'b00101010 : 8'b00111010;
												assign node998 = (inp[12]) ? node1004 : node999;
													assign node999 = (inp[6]) ? node1001 : 8'b00011111;
														assign node1001 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node1004 = (inp[2]) ? 8'b00101010 : node1005;
														assign node1005 = (inp[6]) ? 8'b00101010 : 8'b00111010;
											assign node1009 = (inp[12]) ? node1021 : node1010;
												assign node1010 = (inp[6]) ? node1016 : node1011;
													assign node1011 = (inp[2]) ? 8'b00001110 : node1012;
														assign node1012 = (inp[3]) ? 8'b00001110 : 8'b00001111;
													assign node1016 = (inp[3]) ? node1018 : 8'b00001110;
														assign node1018 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node1021 = (inp[3]) ? node1025 : node1022;
													assign node1022 = (inp[2]) ? 8'b00011110 : 8'b00011111;
													assign node1025 = (inp[2]) ? 8'b00011011 : 8'b00011110;
										assign node1028 = (inp[3]) ? node1046 : node1029;
											assign node1029 = (inp[2]) ? node1037 : node1030;
												assign node1030 = (inp[6]) ? node1034 : node1031;
													assign node1031 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node1034 = (inp[12]) ? 8'b00001111 : 8'b00011110;
												assign node1037 = (inp[12]) ? node1041 : node1038;
													assign node1038 = (inp[6]) ? 8'b00001110 : 8'b00011110;
													assign node1041 = (inp[6]) ? 8'b00011110 : node1042;
														assign node1042 = (inp[0]) ? 8'b00011110 : 8'b00001111;
											assign node1046 = (inp[2]) ? node1054 : node1047;
												assign node1047 = (inp[6]) ? node1051 : node1048;
													assign node1048 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node1051 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node1054 = (inp[0]) ? 8'b00001011 : 8'b00011011;
									assign node1057 = (inp[0]) ? node1087 : node1058;
										assign node1058 = (inp[10]) ? node1074 : node1059;
											assign node1059 = (inp[3]) ? node1067 : node1060;
												assign node1060 = (inp[6]) ? node1062 : 8'b00101010;
													assign node1062 = (inp[2]) ? 8'b00011111 : node1063;
														assign node1063 = (inp[12]) ? 8'b00101010 : 8'b00011111;
												assign node1067 = (inp[12]) ? node1069 : 8'b00011110;
													assign node1069 = (inp[6]) ? 8'b00001111 : node1070;
														assign node1070 = (inp[2]) ? 8'b00001111 : 8'b00011111;
											assign node1074 = (inp[3]) ? node1082 : node1075;
												assign node1075 = (inp[12]) ? node1079 : node1076;
													assign node1076 = (inp[2]) ? 8'b00001011 : 8'b00011011;
													assign node1079 = (inp[2]) ? 8'b00011011 : 8'b00001110;
												assign node1082 = (inp[12]) ? node1084 : 8'b00011010;
													assign node1084 = (inp[6]) ? 8'b00011010 : 8'b00001011;
										assign node1087 = (inp[2]) ? node1095 : node1088;
											assign node1088 = (inp[6]) ? node1092 : node1089;
												assign node1089 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node1092 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node1095 = (inp[12]) ? 8'b00011010 : 8'b00001010;
					assign node1098 = (inp[8]) ? node1412 : node1099;
						assign node1099 = (inp[10]) ? node1259 : node1100;
							assign node1100 = (inp[11]) ? node1148 : node1101;
								assign node1101 = (inp[3]) ? node1123 : node1102;
									assign node1102 = (inp[6]) ? node1112 : node1103;
										assign node1103 = (inp[0]) ? 8'b00011111 : node1104;
											assign node1104 = (inp[1]) ? node1108 : node1105;
												assign node1105 = (inp[2]) ? 8'b00001111 : 8'b00011111;
												assign node1108 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node1112 = (inp[2]) ? node1118 : node1113;
											assign node1113 = (inp[1]) ? node1115 : 8'b00001111;
												assign node1115 = (inp[0]) ? 8'b00001111 : 8'b00001110;
											assign node1118 = (inp[5]) ? 8'b00011111 : node1119;
												assign node1119 = (inp[0]) ? 8'b00001111 : 8'b00001110;
									assign node1123 = (inp[1]) ? node1133 : node1124;
										assign node1124 = (inp[6]) ? node1130 : node1125;
											assign node1125 = (inp[0]) ? 8'b00011110 : node1126;
												assign node1126 = (inp[2]) ? 8'b00001110 : 8'b00011110;
											assign node1130 = (inp[2]) ? 8'b00011110 : 8'b00001110;
										assign node1133 = (inp[5]) ? node1137 : node1134;
											assign node1134 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node1137 = (inp[0]) ? 8'b00011111 : node1138;
												assign node1138 = (inp[12]) ? node1140 : 8'b00001111;
													assign node1140 = (inp[2]) ? node1144 : node1141;
														assign node1141 = (inp[6]) ? 8'b00001111 : 8'b00011111;
														assign node1144 = (inp[6]) ? 8'b00011111 : 8'b00001111;
								assign node1148 = (inp[1]) ? node1194 : node1149;
									assign node1149 = (inp[3]) ? node1171 : node1150;
										assign node1150 = (inp[12]) ? node1160 : node1151;
											assign node1151 = (inp[2]) ? node1155 : node1152;
												assign node1152 = (inp[6]) ? 8'b00011110 : 8'b00001111;
												assign node1155 = (inp[0]) ? 8'b00001110 : node1156;
													assign node1156 = (inp[6]) ? 8'b00001110 : 8'b00011110;
											assign node1160 = (inp[6]) ? node1166 : node1161;
												assign node1161 = (inp[2]) ? node1163 : 8'b00011111;
													assign node1163 = (inp[0]) ? 8'b00011110 : 8'b00001111;
												assign node1166 = (inp[5]) ? node1168 : 8'b00001111;
													assign node1168 = (inp[2]) ? 8'b00011110 : 8'b00001111;
										assign node1171 = (inp[12]) ? node1183 : node1172;
											assign node1172 = (inp[6]) ? node1178 : node1173;
												assign node1173 = (inp[2]) ? node1175 : 8'b00001110;
													assign node1175 = (inp[0]) ? 8'b00001011 : 8'b00011011;
												assign node1178 = (inp[2]) ? node1180 : 8'b00011011;
													assign node1180 = (inp[5]) ? 8'b00001011 : 8'b00011011;
											assign node1183 = (inp[5]) ? node1189 : node1184;
												assign node1184 = (inp[2]) ? 8'b00001110 : node1185;
													assign node1185 = (inp[6]) ? 8'b00001110 : 8'b00011110;
												assign node1189 = (inp[2]) ? 8'b00011011 : node1190;
													assign node1190 = (inp[6]) ? 8'b00001110 : 8'b00011110;
									assign node1194 = (inp[0]) ? node1228 : node1195;
										assign node1195 = (inp[2]) ? node1211 : node1196;
											assign node1196 = (inp[5]) ? node1204 : node1197;
												assign node1197 = (inp[6]) ? node1201 : node1198;
													assign node1198 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node1201 = (inp[3]) ? 8'b00001110 : 8'b00011011;
												assign node1204 = (inp[3]) ? node1206 : 8'b00001110;
													assign node1206 = (inp[6]) ? 8'b00011010 : node1207;
														assign node1207 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node1211 = (inp[3]) ? node1219 : node1212;
												assign node1212 = (inp[5]) ? node1214 : 8'b00011011;
													assign node1214 = (inp[6]) ? node1216 : 8'b00011011;
														assign node1216 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node1219 = (inp[12]) ? node1223 : node1220;
													assign node1220 = (inp[5]) ? 8'b00001010 : 8'b00011011;
													assign node1223 = (inp[5]) ? node1225 : 8'b00001110;
														assign node1225 = (inp[6]) ? 8'b00011010 : 8'b00001011;
										assign node1228 = (inp[12]) ? node1244 : node1229;
											assign node1229 = (inp[6]) ? node1237 : node1230;
												assign node1230 = (inp[2]) ? node1232 : 8'b00001011;
													assign node1232 = (inp[3]) ? node1234 : 8'b00001010;
														assign node1234 = (inp[5]) ? 8'b00001010 : 8'b00001011;
												assign node1237 = (inp[5]) ? node1241 : node1238;
													assign node1238 = (inp[3]) ? 8'b00011011 : 8'b00011010;
													assign node1241 = (inp[2]) ? 8'b00001010 : 8'b00011010;
											assign node1244 = (inp[6]) ? node1254 : node1245;
												assign node1245 = (inp[2]) ? node1249 : node1246;
													assign node1246 = (inp[5]) ? 8'b00011011 : 8'b00011110;
													assign node1249 = (inp[5]) ? 8'b00011010 : node1250;
														assign node1250 = (inp[3]) ? 8'b00011011 : 8'b00011010;
												assign node1254 = (inp[2]) ? node1256 : 8'b00001011;
													assign node1256 = (inp[5]) ? 8'b00011010 : 8'b00001011;
							assign node1259 = (inp[1]) ? node1315 : node1260;
								assign node1260 = (inp[3]) ? node1288 : node1261;
									assign node1261 = (inp[11]) ? node1273 : node1262;
										assign node1262 = (inp[6]) ? node1268 : node1263;
											assign node1263 = (inp[0]) ? 8'b00011011 : node1264;
												assign node1264 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node1268 = (inp[2]) ? node1270 : 8'b00001011;
												assign node1270 = (inp[5]) ? 8'b00011011 : 8'b00001011;
										assign node1273 = (inp[2]) ? node1281 : node1274;
											assign node1274 = (inp[6]) ? node1278 : node1275;
												assign node1275 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node1278 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node1281 = (inp[12]) ? 8'b00011010 : node1282;
												assign node1282 = (inp[6]) ? 8'b00011010 : node1283;
													assign node1283 = (inp[0]) ? 8'b00001010 : 8'b00011010;
									assign node1288 = (inp[2]) ? node1300 : node1289;
										assign node1289 = (inp[6]) ? node1295 : node1290;
											assign node1290 = (inp[12]) ? 8'b00011010 : node1291;
												assign node1291 = (inp[11]) ? 8'b00001010 : 8'b00011010;
											assign node1295 = (inp[12]) ? 8'b00000010 : node1296;
												assign node1296 = (inp[11]) ? 8'b11110111 : 8'b10000010;
										assign node1300 = (inp[11]) ? node1306 : node1301;
											assign node1301 = (inp[0]) ? 8'b10010000 : node1302;
												assign node1302 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node1306 = (inp[0]) ? node1312 : node1307;
												assign node1307 = (inp[12]) ? node1309 : 8'b11110111;
													assign node1309 = (inp[6]) ? 8'b11110101 : 8'b00000010;
												assign node1312 = (inp[12]) ? 8'b11110101 : 8'b10100101;
								assign node1315 = (inp[11]) ? node1357 : node1316;
									assign node1316 = (inp[5]) ? node1336 : node1317;
										assign node1317 = (inp[6]) ? node1329 : node1318;
											assign node1318 = (inp[2]) ? node1324 : node1319;
												assign node1319 = (inp[0]) ? node1321 : 8'b00011010;
													assign node1321 = (inp[3]) ? 8'b00011010 : 8'b10011001;
												assign node1324 = (inp[0]) ? node1326 : 8'b10000010;
													assign node1326 = (inp[3]) ? 8'b10010000 : 8'b10010001;
											assign node1329 = (inp[12]) ? node1331 : 8'b10000010;
												assign node1331 = (inp[0]) ? node1333 : 8'b00000010;
													assign node1333 = (inp[3]) ? 8'b00000010 : 8'b10000001;
										assign node1336 = (inp[2]) ? node1344 : node1337;
											assign node1337 = (inp[6]) ? 8'b10000001 : node1338;
												assign node1338 = (inp[0]) ? 8'b10011001 : node1339;
													assign node1339 = (inp[3]) ? 8'b10011001 : 8'b00011010;
											assign node1344 = (inp[3]) ? node1352 : node1345;
												assign node1345 = (inp[0]) ? 8'b10010001 : node1346;
													assign node1346 = (inp[6]) ? 8'b10010000 : node1347;
														assign node1347 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node1352 = (inp[0]) ? 8'b10010001 : node1353;
													assign node1353 = (inp[6]) ? 8'b10010001 : 8'b10000001;
									assign node1357 = (inp[0]) ? node1387 : node1358;
										assign node1358 = (inp[6]) ? node1368 : node1359;
											assign node1359 = (inp[2]) ? node1365 : node1360;
												assign node1360 = (inp[12]) ? node1362 : 8'b00001010;
													assign node1362 = (inp[5]) ? 8'b11111101 : 8'b00011010;
												assign node1365 = (inp[5]) ? 8'b00000010 : 8'b11110111;
											assign node1368 = (inp[12]) ? node1378 : node1369;
												assign node1369 = (inp[5]) ? node1371 : 8'b11110111;
													assign node1371 = (inp[3]) ? node1375 : node1372;
														assign node1372 = (inp[2]) ? 8'b10100101 : 8'b11110111;
														assign node1375 = (inp[2]) ? 8'b10100100 : 8'b10110100;
												assign node1378 = (inp[5]) ? node1380 : 8'b00000010;
													assign node1380 = (inp[2]) ? node1384 : node1381;
														assign node1381 = (inp[3]) ? 8'b10100101 : 8'b00000010;
														assign node1384 = (inp[3]) ? 8'b10110100 : 8'b11110101;
										assign node1387 = (inp[5]) ? node1403 : node1388;
											assign node1388 = (inp[3]) ? node1394 : node1389;
												assign node1389 = (inp[6]) ? node1391 : 8'b10101101;
													assign node1391 = (inp[12]) ? 8'b10100101 : 8'b10110100;
												assign node1394 = (inp[6]) ? node1400 : node1395;
													assign node1395 = (inp[2]) ? node1397 : 8'b00001010;
														assign node1397 = (inp[12]) ? 8'b11110101 : 8'b10100101;
													assign node1400 = (inp[12]) ? 8'b00000010 : 8'b11110111;
											assign node1403 = (inp[2]) ? node1409 : node1404;
												assign node1404 = (inp[6]) ? node1406 : 8'b10101101;
													assign node1406 = (inp[12]) ? 8'b10100101 : 8'b10110100;
												assign node1409 = (inp[12]) ? 8'b10110100 : 8'b10100100;
						assign node1412 = (inp[0]) ? node1590 : node1413;
							assign node1413 = (inp[5]) ? node1463 : node1414;
								assign node1414 = (inp[12]) ? node1446 : node1415;
									assign node1415 = (inp[11]) ? node1429 : node1416;
										assign node1416 = (inp[3]) ? node1424 : node1417;
											assign node1417 = (inp[1]) ? node1419 : 8'b00001011;
												assign node1419 = (inp[6]) ? 8'b10000010 : node1420;
													assign node1420 = (inp[2]) ? 8'b10000010 : 8'b00011010;
											assign node1424 = (inp[2]) ? 8'b10000010 : node1425;
												assign node1425 = (inp[6]) ? 8'b10000010 : 8'b00011010;
										assign node1429 = (inp[2]) ? node1441 : node1430;
											assign node1430 = (inp[6]) ? node1436 : node1431;
												assign node1431 = (inp[1]) ? 8'b00001010 : node1432;
													assign node1432 = (inp[3]) ? 8'b00001010 : 8'b00001011;
												assign node1436 = (inp[3]) ? 8'b11110111 : node1437;
													assign node1437 = (inp[10]) ? 8'b11110111 : 8'b00011010;
											assign node1441 = (inp[1]) ? 8'b11110111 : node1442;
												assign node1442 = (inp[3]) ? 8'b11110111 : 8'b00011010;
									assign node1446 = (inp[3]) ? node1458 : node1447;
										assign node1447 = (inp[1]) ? node1453 : node1448;
											assign node1448 = (inp[6]) ? 8'b00001011 : node1449;
												assign node1449 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node1453 = (inp[6]) ? 8'b00000010 : node1454;
												assign node1454 = (inp[2]) ? 8'b00000010 : 8'b00011010;
										assign node1458 = (inp[2]) ? 8'b00000010 : node1459;
											assign node1459 = (inp[6]) ? 8'b00000010 : 8'b00011010;
								assign node1463 = (inp[10]) ? node1525 : node1464;
									assign node1464 = (inp[3]) ? node1494 : node1465;
										assign node1465 = (inp[1]) ? node1485 : node1466;
											assign node1466 = (inp[11]) ? node1474 : node1467;
												assign node1467 = (inp[2]) ? node1471 : node1468;
													assign node1468 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node1471 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node1474 = (inp[2]) ? node1480 : node1475;
													assign node1475 = (inp[12]) ? node1477 : 8'b00001011;
														assign node1477 = (inp[6]) ? 8'b00001011 : 8'b00011011;
													assign node1480 = (inp[6]) ? 8'b00011010 : node1481;
														assign node1481 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node1485 = (inp[6]) ? node1489 : node1486;
												assign node1486 = (inp[12]) ? 8'b00000010 : 8'b00001010;
												assign node1489 = (inp[2]) ? node1491 : 8'b00000010;
													assign node1491 = (inp[12]) ? 8'b11110101 : 8'b10010000;
										assign node1494 = (inp[1]) ? node1510 : node1495;
											assign node1495 = (inp[6]) ? node1501 : node1496;
												assign node1496 = (inp[2]) ? node1498 : 8'b00011010;
													assign node1498 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node1501 = (inp[2]) ? node1505 : node1502;
													assign node1502 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node1505 = (inp[11]) ? node1507 : 8'b10010000;
														assign node1507 = (inp[12]) ? 8'b11110101 : 8'b10100101;
											assign node1510 = (inp[11]) ? node1518 : node1511;
												assign node1511 = (inp[6]) ? node1515 : node1512;
													assign node1512 = (inp[2]) ? 8'b10000001 : 8'b10011001;
													assign node1515 = (inp[2]) ? 8'b10010001 : 8'b10000001;
												assign node1518 = (inp[2]) ? node1522 : node1519;
													assign node1519 = (inp[12]) ? 8'b10100101 : 8'b10101101;
													assign node1522 = (inp[12]) ? 8'b10110100 : 8'b10100100;
									assign node1525 = (inp[11]) ? node1557 : node1526;
										assign node1526 = (inp[1]) ? node1542 : node1527;
											assign node1527 = (inp[3]) ? node1535 : node1528;
												assign node1528 = (inp[6]) ? node1532 : node1529;
													assign node1529 = (inp[2]) ? 8'b10001101 : 8'b10011101;
													assign node1532 = (inp[2]) ? 8'b10011101 : 8'b10001101;
												assign node1535 = (inp[6]) ? node1539 : node1536;
													assign node1536 = (inp[2]) ? 8'b10000100 : 8'b10011100;
													assign node1539 = (inp[2]) ? 8'b10010100 : 8'b10000100;
											assign node1542 = (inp[3]) ? node1550 : node1543;
												assign node1543 = (inp[6]) ? node1547 : node1544;
													assign node1544 = (inp[2]) ? 8'b10000100 : 8'b10011100;
													assign node1547 = (inp[12]) ? 8'b10000100 : 8'b10010100;
												assign node1550 = (inp[6]) ? node1554 : node1551;
													assign node1551 = (inp[2]) ? 8'b10000101 : 8'b10011101;
													assign node1554 = (inp[2]) ? 8'b10010101 : 8'b10000101;
										assign node1557 = (inp[3]) ? node1569 : node1558;
											assign node1558 = (inp[6]) ? node1564 : node1559;
												assign node1559 = (inp[1]) ? node1561 : 8'b10111100;
													assign node1561 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node1564 = (inp[1]) ? 8'b10100001 : node1565;
													assign node1565 = (inp[12]) ? 8'b10101101 : 8'b10111100;
											assign node1569 = (inp[6]) ? node1579 : node1570;
												assign node1570 = (inp[1]) ? node1572 : 8'b10111100;
													assign node1572 = (inp[2]) ? node1576 : node1573;
														assign node1573 = (inp[12]) ? 8'b10111001 : 8'b10101001;
														assign node1576 = (inp[12]) ? 8'b10100001 : 8'b10110000;
												assign node1579 = (inp[1]) ? node1583 : node1580;
													assign node1580 = (inp[2]) ? 8'b10100001 : 8'b10110001;
													assign node1583 = (inp[12]) ? node1587 : node1584;
														assign node1584 = (inp[2]) ? 8'b10100000 : 8'b10110000;
														assign node1587 = (inp[2]) ? 8'b10110000 : 8'b10100001;
							assign node1590 = (inp[11]) ? node1648 : node1591;
								assign node1591 = (inp[6]) ? node1621 : node1592;
									assign node1592 = (inp[3]) ? node1606 : node1593;
										assign node1593 = (inp[5]) ? node1601 : node1594;
											assign node1594 = (inp[10]) ? node1596 : 8'b10011101;
												assign node1596 = (inp[1]) ? node1598 : 8'b00011011;
													assign node1598 = (inp[2]) ? 8'b10010001 : 8'b10011001;
											assign node1601 = (inp[1]) ? node1603 : 8'b10011101;
												assign node1603 = (inp[2]) ? 8'b10010101 : 8'b10011101;
										assign node1606 = (inp[2]) ? node1614 : node1607;
											assign node1607 = (inp[5]) ? node1611 : node1608;
												assign node1608 = (inp[10]) ? 8'b00011010 : 8'b10011100;
												assign node1611 = (inp[1]) ? 8'b10011101 : 8'b10011100;
											assign node1614 = (inp[5]) ? node1618 : node1615;
												assign node1615 = (inp[10]) ? 8'b10010000 : 8'b10010100;
												assign node1618 = (inp[1]) ? 8'b10010101 : 8'b10010100;
									assign node1621 = (inp[5]) ? node1635 : node1622;
										assign node1622 = (inp[10]) ? node1628 : node1623;
											assign node1623 = (inp[3]) ? 8'b10000100 : node1624;
												assign node1624 = (inp[1]) ? 8'b10000101 : 8'b10001101;
											assign node1628 = (inp[3]) ? node1632 : node1629;
												assign node1629 = (inp[1]) ? 8'b10000001 : 8'b00001011;
												assign node1632 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node1635 = (inp[2]) ? node1643 : node1636;
											assign node1636 = (inp[3]) ? node1640 : node1637;
												assign node1637 = (inp[1]) ? 8'b10000101 : 8'b10001101;
												assign node1640 = (inp[1]) ? 8'b10000101 : 8'b10000100;
											assign node1643 = (inp[1]) ? 8'b10010101 : node1644;
												assign node1644 = (inp[3]) ? 8'b10010100 : 8'b10011101;
								assign node1648 = (inp[1]) ? node1708 : node1649;
									assign node1649 = (inp[3]) ? node1679 : node1650;
										assign node1650 = (inp[5]) ? node1668 : node1651;
											assign node1651 = (inp[10]) ? node1661 : node1652;
												assign node1652 = (inp[2]) ? node1654 : 8'b10101101;
													assign node1654 = (inp[6]) ? node1658 : node1655;
														assign node1655 = (inp[12]) ? 8'b10111100 : 8'b10101100;
														assign node1658 = (inp[12]) ? 8'b10101101 : 8'b10111100;
												assign node1661 = (inp[6]) ? 8'b00001011 : node1662;
													assign node1662 = (inp[12]) ? node1664 : 8'b00001011;
														assign node1664 = (inp[2]) ? 8'b00011010 : 8'b00011011;
											assign node1668 = (inp[2]) ? node1676 : node1669;
												assign node1669 = (inp[12]) ? node1673 : node1670;
													assign node1670 = (inp[6]) ? 8'b10111100 : 8'b10101101;
													assign node1673 = (inp[6]) ? 8'b10101101 : 8'b11111101;
												assign node1676 = (inp[12]) ? 8'b10111100 : 8'b10101100;
										assign node1679 = (inp[2]) ? node1693 : node1680;
											assign node1680 = (inp[6]) ? node1686 : node1681;
												assign node1681 = (inp[12]) ? 8'b10111100 : node1682;
													assign node1682 = (inp[5]) ? 8'b10101100 : 8'b00001010;
												assign node1686 = (inp[12]) ? 8'b10100100 : node1687;
													assign node1687 = (inp[10]) ? node1689 : 8'b10110001;
														assign node1689 = (inp[5]) ? 8'b10110001 : 8'b11110111;
											assign node1693 = (inp[5]) ? node1705 : node1694;
												assign node1694 = (inp[6]) ? node1700 : node1695;
													assign node1695 = (inp[12]) ? node1697 : 8'b10100101;
														assign node1697 = (inp[10]) ? 8'b11110101 : 8'b10110001;
													assign node1700 = (inp[10]) ? 8'b00000010 : node1701;
														assign node1701 = (inp[12]) ? 8'b10100100 : 8'b10110001;
												assign node1705 = (inp[12]) ? 8'b10110001 : 8'b10100001;
									assign node1708 = (inp[2]) ? node1750 : node1709;
										assign node1709 = (inp[6]) ? node1729 : node1710;
											assign node1710 = (inp[12]) ? node1718 : node1711;
												assign node1711 = (inp[5]) ? 8'b10101001 : node1712;
													assign node1712 = (inp[3]) ? 8'b10101100 : node1713;
														assign node1713 = (inp[10]) ? 8'b10101101 : 8'b10101001;
												assign node1718 = (inp[3]) ? node1724 : node1719;
													assign node1719 = (inp[5]) ? 8'b10111001 : node1720;
														assign node1720 = (inp[10]) ? 8'b11111101 : 8'b10111001;
													assign node1724 = (inp[10]) ? 8'b00011010 : node1725;
														assign node1725 = (inp[5]) ? 8'b10111001 : 8'b10111100;
											assign node1729 = (inp[12]) ? node1739 : node1730;
												assign node1730 = (inp[3]) ? node1734 : node1731;
													assign node1731 = (inp[10]) ? 8'b10110100 : 8'b10110000;
													assign node1734 = (inp[5]) ? 8'b10110000 : node1735;
														assign node1735 = (inp[10]) ? 8'b11110111 : 8'b10110001;
												assign node1739 = (inp[3]) ? node1745 : node1740;
													assign node1740 = (inp[5]) ? 8'b10100001 : node1741;
														assign node1741 = (inp[10]) ? 8'b10100101 : 8'b10100001;
													assign node1745 = (inp[10]) ? 8'b00000010 : node1746;
														assign node1746 = (inp[5]) ? 8'b10100001 : 8'b10100100;
										assign node1750 = (inp[5]) ? node1762 : node1751;
											assign node1751 = (inp[10]) ? node1755 : node1752;
												assign node1752 = (inp[3]) ? 8'b10110001 : 8'b10110000;
												assign node1755 = (inp[3]) ? node1759 : node1756;
													assign node1756 = (inp[6]) ? 8'b10100101 : 8'b10100100;
													assign node1759 = (inp[12]) ? 8'b00000010 : 8'b11110111;
											assign node1762 = (inp[12]) ? 8'b10110000 : 8'b10100000;
			assign node1765 = (inp[5]) ? node2653 : node1766;
				assign node1766 = (inp[0]) ? node1966 : node1767;
					assign node1767 = (inp[8]) ? node1895 : node1768;
						assign node1768 = (inp[7]) ? node1792 : node1769;
							assign node1769 = (inp[1]) ? node1781 : node1770;
								assign node1770 = (inp[2]) ? node1776 : node1771;
									assign node1771 = (inp[12]) ? 8'b00011111 : node1772;
										assign node1772 = (inp[11]) ? 8'b00001111 : 8'b00011111;
									assign node1776 = (inp[11]) ? node1778 : 8'b00001111;
										assign node1778 = (inp[12]) ? 8'b00001111 : 8'b00011110;
								assign node1781 = (inp[2]) ? node1787 : node1782;
									assign node1782 = (inp[11]) ? node1784 : 8'b00011110;
										assign node1784 = (inp[12]) ? 8'b00011110 : 8'b00001110;
									assign node1787 = (inp[11]) ? node1789 : 8'b00001110;
										assign node1789 = (inp[12]) ? 8'b00001110 : 8'b00011011;
							assign node1792 = (inp[10]) ? node1842 : node1793;
								assign node1793 = (inp[12]) ? node1825 : node1794;
									assign node1794 = (inp[11]) ? node1812 : node1795;
										assign node1795 = (inp[6]) ? node1807 : node1796;
											assign node1796 = (inp[2]) ? node1802 : node1797;
												assign node1797 = (inp[3]) ? 8'b00011110 : node1798;
													assign node1798 = (inp[1]) ? 8'b00011110 : 8'b00011111;
												assign node1802 = (inp[3]) ? 8'b00001110 : node1803;
													assign node1803 = (inp[9]) ? 8'b00001110 : 8'b00001111;
											assign node1807 = (inp[1]) ? 8'b00001110 : node1808;
												assign node1808 = (inp[3]) ? 8'b00001110 : 8'b00001111;
										assign node1812 = (inp[3]) ? 8'b00011011 : node1813;
											assign node1813 = (inp[1]) ? node1819 : node1814;
												assign node1814 = (inp[6]) ? 8'b00011110 : node1815;
													assign node1815 = (inp[2]) ? 8'b00011110 : 8'b00001111;
												assign node1819 = (inp[6]) ? 8'b00011011 : node1820;
													assign node1820 = (inp[2]) ? 8'b00011011 : 8'b00001110;
									assign node1825 = (inp[3]) ? node1837 : node1826;
										assign node1826 = (inp[1]) ? node1832 : node1827;
											assign node1827 = (inp[2]) ? 8'b00001111 : node1828;
												assign node1828 = (inp[6]) ? 8'b00001111 : 8'b00011111;
											assign node1832 = (inp[6]) ? 8'b00001110 : node1833;
												assign node1833 = (inp[9]) ? 8'b00011110 : 8'b00001110;
										assign node1837 = (inp[6]) ? 8'b00001110 : node1838;
											assign node1838 = (inp[2]) ? 8'b00001110 : 8'b00011110;
								assign node1842 = (inp[12]) ? node1876 : node1843;
									assign node1843 = (inp[11]) ? node1861 : node1844;
										assign node1844 = (inp[1]) ? node1856 : node1845;
											assign node1845 = (inp[3]) ? node1851 : node1846;
												assign node1846 = (inp[6]) ? 8'b00001011 : node1847;
													assign node1847 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node1851 = (inp[2]) ? 8'b10000010 : node1852;
													assign node1852 = (inp[6]) ? 8'b10000010 : 8'b00011010;
											assign node1856 = (inp[2]) ? 8'b10000010 : node1857;
												assign node1857 = (inp[6]) ? 8'b10000010 : 8'b00011010;
										assign node1861 = (inp[6]) ? node1871 : node1862;
											assign node1862 = (inp[2]) ? node1868 : node1863;
												assign node1863 = (inp[1]) ? 8'b00001010 : node1864;
													assign node1864 = (inp[3]) ? 8'b00001010 : 8'b00001011;
												assign node1868 = (inp[3]) ? 8'b11110111 : 8'b00011010;
											assign node1871 = (inp[3]) ? 8'b11110111 : node1872;
												assign node1872 = (inp[1]) ? 8'b11110111 : 8'b00011010;
									assign node1876 = (inp[2]) ? node1890 : node1877;
										assign node1877 = (inp[6]) ? node1885 : node1878;
											assign node1878 = (inp[11]) ? 8'b00011010 : node1879;
												assign node1879 = (inp[3]) ? 8'b00011010 : node1880;
													assign node1880 = (inp[1]) ? 8'b00011010 : 8'b00011011;
											assign node1885 = (inp[1]) ? 8'b00000010 : node1886;
												assign node1886 = (inp[3]) ? 8'b00000010 : 8'b00001011;
										assign node1890 = (inp[1]) ? 8'b00000010 : node1891;
											assign node1891 = (inp[3]) ? 8'b00000010 : 8'b00001011;
						assign node1895 = (inp[1]) ? node1943 : node1896;
							assign node1896 = (inp[7]) ? node1908 : node1897;
								assign node1897 = (inp[2]) ? node1903 : node1898;
									assign node1898 = (inp[11]) ? node1900 : 8'b00011011;
										assign node1900 = (inp[12]) ? 8'b00011011 : 8'b00001011;
									assign node1903 = (inp[12]) ? 8'b00001011 : node1904;
										assign node1904 = (inp[11]) ? 8'b00011010 : 8'b00001011;
								assign node1908 = (inp[3]) ? node1926 : node1909;
									assign node1909 = (inp[11]) ? node1915 : node1910;
										assign node1910 = (inp[6]) ? 8'b00001011 : node1911;
											assign node1911 = (inp[2]) ? 8'b00001011 : 8'b00011011;
										assign node1915 = (inp[12]) ? node1921 : node1916;
											assign node1916 = (inp[6]) ? 8'b00011010 : node1917;
												assign node1917 = (inp[2]) ? 8'b00011010 : 8'b00001011;
											assign node1921 = (inp[2]) ? 8'b00001011 : node1922;
												assign node1922 = (inp[6]) ? 8'b00001011 : 8'b00011011;
									assign node1926 = (inp[12]) ? node1938 : node1927;
										assign node1927 = (inp[11]) ? node1933 : node1928;
											assign node1928 = (inp[2]) ? 8'b10000010 : node1929;
												assign node1929 = (inp[6]) ? 8'b10000010 : 8'b00011010;
											assign node1933 = (inp[6]) ? 8'b11110111 : node1934;
												assign node1934 = (inp[2]) ? 8'b11110111 : 8'b00001010;
										assign node1938 = (inp[2]) ? 8'b00000010 : node1939;
											assign node1939 = (inp[6]) ? 8'b00000010 : 8'b00011010;
							assign node1943 = (inp[2]) ? node1961 : node1944;
								assign node1944 = (inp[7]) ? node1950 : node1945;
									assign node1945 = (inp[12]) ? 8'b00011010 : node1946;
										assign node1946 = (inp[11]) ? 8'b00001010 : 8'b00011010;
									assign node1950 = (inp[6]) ? node1956 : node1951;
										assign node1951 = (inp[11]) ? node1953 : 8'b00011010;
											assign node1953 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node1956 = (inp[12]) ? 8'b00000010 : node1957;
											assign node1957 = (inp[11]) ? 8'b11110111 : 8'b10000010;
								assign node1961 = (inp[12]) ? 8'b00000010 : node1962;
									assign node1962 = (inp[11]) ? 8'b11110111 : 8'b10000010;
					assign node1966 = (inp[9]) ? node2310 : node1967;
						assign node1967 = (inp[11]) ? node2069 : node1968;
							assign node1968 = (inp[3]) ? node2014 : node1969;
								assign node1969 = (inp[10]) ? node1987 : node1970;
									assign node1970 = (inp[6]) ? node1978 : node1971;
										assign node1971 = (inp[8]) ? node1973 : 8'b11111101;
											assign node1973 = (inp[1]) ? node1975 : 8'b11111101;
												assign node1975 = (inp[2]) ? 8'b11110101 : 8'b11111101;
										assign node1978 = (inp[7]) ? node1982 : node1979;
											assign node1979 = (inp[2]) ? 8'b10101101 : 8'b11111101;
											assign node1982 = (inp[8]) ? node1984 : 8'b10101101;
												assign node1984 = (inp[1]) ? 8'b10100101 : 8'b10101101;
									assign node1987 = (inp[6]) ? node2001 : node1988;
										assign node1988 = (inp[7]) ? node1996 : node1989;
											assign node1989 = (inp[8]) ? node1991 : 8'b11111101;
												assign node1991 = (inp[1]) ? node1993 : 8'b10111001;
													assign node1993 = (inp[2]) ? 8'b10110001 : 8'b10111001;
											assign node1996 = (inp[2]) ? node1998 : 8'b10111001;
												assign node1998 = (inp[1]) ? 8'b10110001 : 8'b10111001;
										assign node2001 = (inp[7]) ? node2011 : node2002;
											assign node2002 = (inp[8]) ? node2006 : node2003;
												assign node2003 = (inp[2]) ? 8'b10101101 : 8'b11111101;
												assign node2006 = (inp[2]) ? node2008 : 8'b10111001;
													assign node2008 = (inp[1]) ? 8'b10100001 : 8'b10101001;
											assign node2011 = (inp[1]) ? 8'b10100001 : 8'b10101001;
								assign node2014 = (inp[10]) ? node2040 : node2015;
									assign node2015 = (inp[6]) ? node2027 : node2016;
										assign node2016 = (inp[1]) ? node2024 : node2017;
											assign node2017 = (inp[7]) ? node2019 : 8'b11111101;
												assign node2019 = (inp[2]) ? node2021 : 8'b10111100;
													assign node2021 = (inp[8]) ? 8'b10110100 : 8'b10111100;
											assign node2024 = (inp[2]) ? 8'b10110100 : 8'b10111100;
										assign node2027 = (inp[7]) ? node2037 : node2028;
											assign node2028 = (inp[2]) ? node2032 : node2029;
												assign node2029 = (inp[1]) ? 8'b10111100 : 8'b11111101;
												assign node2032 = (inp[1]) ? node2034 : 8'b10101101;
													assign node2034 = (inp[8]) ? 8'b10100100 : 8'b10101100;
											assign node2037 = (inp[8]) ? 8'b10100100 : 8'b10101100;
									assign node2040 = (inp[7]) ? node2064 : node2041;
										assign node2041 = (inp[8]) ? node2053 : node2042;
											assign node2042 = (inp[1]) ? node2048 : node2043;
												assign node2043 = (inp[12]) ? node2045 : 8'b11111101;
													assign node2045 = (inp[6]) ? 8'b10101101 : 8'b11111101;
												assign node2048 = (inp[6]) ? node2050 : 8'b10111100;
													assign node2050 = (inp[2]) ? 8'b10101100 : 8'b10111100;
											assign node2053 = (inp[1]) ? node2059 : node2054;
												assign node2054 = (inp[6]) ? node2056 : 8'b10111001;
													assign node2056 = (inp[2]) ? 8'b10101001 : 8'b10111001;
												assign node2059 = (inp[6]) ? 8'b10100000 : node2060;
													assign node2060 = (inp[2]) ? 8'b10110000 : 8'b10111000;
										assign node2064 = (inp[6]) ? 8'b10100000 : node2065;
											assign node2065 = (inp[2]) ? 8'b10110000 : 8'b10111000;
							assign node2069 = (inp[8]) ? node2183 : node2070;
								assign node2070 = (inp[1]) ? node2120 : node2071;
									assign node2071 = (inp[7]) ? node2083 : node2072;
										assign node2072 = (inp[2]) ? node2076 : node2073;
											assign node2073 = (inp[12]) ? 8'b11111101 : 8'b10101101;
											assign node2076 = (inp[6]) ? node2080 : node2077;
												assign node2077 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node2080 = (inp[12]) ? 8'b10101101 : 8'b10111100;
										assign node2083 = (inp[10]) ? node2101 : node2084;
											assign node2084 = (inp[2]) ? node2092 : node2085;
												assign node2085 = (inp[3]) ? node2087 : 8'b10111100;
													assign node2087 = (inp[12]) ? node2089 : 8'b10101100;
														assign node2089 = (inp[6]) ? 8'b10101100 : 8'b10111100;
												assign node2092 = (inp[6]) ? node2096 : node2093;
													assign node2093 = (inp[3]) ? 8'b10111001 : 8'b10111100;
													assign node2096 = (inp[12]) ? node2098 : 8'b10111100;
														assign node2098 = (inp[3]) ? 8'b10101100 : 8'b10101101;
											assign node2101 = (inp[3]) ? node2111 : node2102;
												assign node2102 = (inp[2]) ? node2104 : 8'b10101001;
													assign node2104 = (inp[6]) ? node2108 : node2105;
														assign node2105 = (inp[12]) ? 8'b10111000 : 8'b10101000;
														assign node2108 = (inp[12]) ? 8'b10101001 : 8'b10111000;
												assign node2111 = (inp[2]) ? node2113 : 8'b10111000;
													assign node2113 = (inp[6]) ? node2117 : node2114;
														assign node2114 = (inp[12]) ? 8'b10010101 : 8'b10000101;
														assign node2117 = (inp[12]) ? 8'b10100000 : 8'b10010101;
									assign node2120 = (inp[7]) ? node2146 : node2121;
										assign node2121 = (inp[6]) ? node2133 : node2122;
											assign node2122 = (inp[12]) ? node2128 : node2123;
												assign node2123 = (inp[3]) ? 8'b10101001 : node2124;
													assign node2124 = (inp[2]) ? 8'b10101000 : 8'b10101001;
												assign node2128 = (inp[2]) ? node2130 : 8'b10111001;
													assign node2130 = (inp[3]) ? 8'b10111001 : 8'b10111000;
											assign node2133 = (inp[3]) ? node2139 : node2134;
												assign node2134 = (inp[12]) ? node2136 : 8'b10111000;
													assign node2136 = (inp[2]) ? 8'b10101001 : 8'b10111001;
												assign node2139 = (inp[12]) ? node2143 : node2140;
													assign node2140 = (inp[2]) ? 8'b10111001 : 8'b10101100;
													assign node2143 = (inp[2]) ? 8'b10101100 : 8'b10111100;
										assign node2146 = (inp[10]) ? node2164 : node2147;
											assign node2147 = (inp[2]) ? node2153 : node2148;
												assign node2148 = (inp[3]) ? 8'b10111001 : node2149;
													assign node2149 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node2153 = (inp[6]) ? node2161 : node2154;
													assign node2154 = (inp[3]) ? node2158 : node2155;
														assign node2155 = (inp[12]) ? 8'b10111000 : 8'b10101000;
														assign node2158 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node2161 = (inp[3]) ? 8'b10101100 : 8'b10101001;
											assign node2164 = (inp[3]) ? node2176 : node2165;
												assign node2165 = (inp[2]) ? node2171 : node2166;
													assign node2166 = (inp[6]) ? 8'b10010100 : node2167;
														assign node2167 = (inp[12]) ? 8'b10011101 : 8'b10001101;
													assign node2171 = (inp[12]) ? 8'b10000101 : node2172;
														assign node2172 = (inp[6]) ? 8'b10010100 : 8'b10000100;
												assign node2176 = (inp[6]) ? node2180 : node2177;
													assign node2177 = (inp[12]) ? 8'b10111000 : 8'b10101000;
													assign node2180 = (inp[12]) ? 8'b10100000 : 8'b10010101;
								assign node2183 = (inp[10]) ? node2247 : node2184;
									assign node2184 = (inp[1]) ? node2220 : node2185;
										assign node2185 = (inp[3]) ? node2203 : node2186;
											assign node2186 = (inp[2]) ? node2198 : node2187;
												assign node2187 = (inp[12]) ? node2193 : node2188;
													assign node2188 = (inp[6]) ? node2190 : 8'b10001101;
														assign node2190 = (inp[7]) ? 8'b10011100 : 8'b10001101;
													assign node2193 = (inp[7]) ? node2195 : 8'b10011101;
														assign node2195 = (inp[6]) ? 8'b10001101 : 8'b10011101;
												assign node2198 = (inp[12]) ? node2200 : 8'b10011100;
													assign node2200 = (inp[6]) ? 8'b10001101 : 8'b10011100;
											assign node2203 = (inp[7]) ? node2213 : node2204;
												assign node2204 = (inp[2]) ? node2208 : node2205;
													assign node2205 = (inp[12]) ? 8'b10011101 : 8'b10001101;
													assign node2208 = (inp[6]) ? 8'b10001101 : node2209;
														assign node2209 = (inp[12]) ? 8'b10011100 : 8'b10001100;
												assign node2213 = (inp[12]) ? 8'b10000100 : node2214;
													assign node2214 = (inp[6]) ? 8'b10010001 : node2215;
														assign node2215 = (inp[2]) ? 8'b10000001 : 8'b10001100;
										assign node2220 = (inp[2]) ? node2232 : node2221;
											assign node2221 = (inp[3]) ? node2229 : node2222;
												assign node2222 = (inp[7]) ? node2226 : node2223;
													assign node2223 = (inp[12]) ? 8'b10011001 : 8'b10001001;
													assign node2226 = (inp[6]) ? 8'b10010000 : 8'b10011001;
												assign node2229 = (inp[12]) ? 8'b10011100 : 8'b10001100;
											assign node2232 = (inp[3]) ? node2240 : node2233;
												assign node2233 = (inp[6]) ? node2237 : node2234;
													assign node2234 = (inp[12]) ? 8'b10010000 : 8'b10000000;
													assign node2237 = (inp[12]) ? 8'b10000001 : 8'b10010000;
												assign node2240 = (inp[12]) ? node2244 : node2241;
													assign node2241 = (inp[6]) ? 8'b10010001 : 8'b10000001;
													assign node2244 = (inp[7]) ? 8'b10000100 : 8'b10010001;
									assign node2247 = (inp[1]) ? node2287 : node2248;
										assign node2248 = (inp[3]) ? node2266 : node2249;
											assign node2249 = (inp[2]) ? node2259 : node2250;
												assign node2250 = (inp[12]) ? node2256 : node2251;
													assign node2251 = (inp[6]) ? node2253 : 8'b10101001;
														assign node2253 = (inp[7]) ? 8'b10111000 : 8'b10101001;
													assign node2256 = (inp[6]) ? 8'b10101001 : 8'b10111001;
												assign node2259 = (inp[7]) ? 8'b10111000 : node2260;
													assign node2260 = (inp[12]) ? 8'b10101001 : node2261;
														assign node2261 = (inp[6]) ? 8'b10111000 : 8'b10101000;
											assign node2266 = (inp[7]) ? node2276 : node2267;
												assign node2267 = (inp[6]) ? node2269 : 8'b10101000;
													assign node2269 = (inp[12]) ? node2273 : node2270;
														assign node2270 = (inp[2]) ? 8'b10111000 : 8'b10101001;
														assign node2273 = (inp[2]) ? 8'b10101001 : 8'b10111001;
												assign node2276 = (inp[2]) ? node2282 : node2277;
													assign node2277 = (inp[6]) ? 8'b10100000 : node2278;
														assign node2278 = (inp[12]) ? 8'b10111000 : 8'b10101000;
													assign node2282 = (inp[6]) ? 8'b10100000 : node2283;
														assign node2283 = (inp[12]) ? 8'b10010101 : 8'b10000101;
										assign node2287 = (inp[2]) ? node2297 : node2288;
											assign node2288 = (inp[3]) ? node2292 : node2289;
												assign node2289 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node2292 = (inp[7]) ? node2294 : 8'b10111000;
													assign node2294 = (inp[6]) ? 8'b10100000 : 8'b10101000;
											assign node2297 = (inp[3]) ? node2303 : node2298;
												assign node2298 = (inp[6]) ? 8'b10010100 : node2299;
													assign node2299 = (inp[12]) ? 8'b10010100 : 8'b10000100;
												assign node2303 = (inp[12]) ? node2307 : node2304;
													assign node2304 = (inp[6]) ? 8'b10010101 : 8'b10000101;
													assign node2307 = (inp[6]) ? 8'b10100000 : 8'b10010101;
						assign node2310 = (inp[8]) ? node2466 : node2311;
							assign node2311 = (inp[7]) ? node2367 : node2312;
								assign node2312 = (inp[1]) ? node2330 : node2313;
									assign node2313 = (inp[2]) ? node2319 : node2314;
										assign node2314 = (inp[12]) ? 8'b00011111 : node2315;
											assign node2315 = (inp[11]) ? 8'b00001111 : 8'b00011111;
										assign node2319 = (inp[11]) ? node2323 : node2320;
											assign node2320 = (inp[6]) ? 8'b00001111 : 8'b00011111;
											assign node2323 = (inp[6]) ? node2327 : node2324;
												assign node2324 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node2327 = (inp[12]) ? 8'b00001111 : 8'b00011110;
									assign node2330 = (inp[11]) ? node2342 : node2331;
										assign node2331 = (inp[3]) ? node2337 : node2332;
											assign node2332 = (inp[6]) ? node2334 : 8'b00011111;
												assign node2334 = (inp[2]) ? 8'b00001111 : 8'b00011111;
											assign node2337 = (inp[6]) ? node2339 : 8'b00011110;
												assign node2339 = (inp[2]) ? 8'b00001110 : 8'b00011110;
										assign node2342 = (inp[3]) ? node2356 : node2343;
											assign node2343 = (inp[2]) ? node2347 : node2344;
												assign node2344 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node2347 = (inp[10]) ? node2353 : node2348;
													assign node2348 = (inp[6]) ? node2350 : 8'b00011010;
														assign node2350 = (inp[12]) ? 8'b00001011 : 8'b00011010;
													assign node2353 = (inp[6]) ? 8'b00001011 : 8'b00001010;
											assign node2356 = (inp[2]) ? node2360 : node2357;
												assign node2357 = (inp[10]) ? 8'b00001110 : 8'b00011110;
												assign node2360 = (inp[6]) ? node2364 : node2361;
													assign node2361 = (inp[12]) ? 8'b00011011 : 8'b00001011;
													assign node2364 = (inp[12]) ? 8'b00001110 : 8'b00011011;
								assign node2367 = (inp[10]) ? node2407 : node2368;
									assign node2368 = (inp[11]) ? node2376 : node2369;
										assign node2369 = (inp[6]) ? node2373 : node2370;
											assign node2370 = (inp[3]) ? 8'b00011110 : 8'b00011111;
											assign node2373 = (inp[3]) ? 8'b00001110 : 8'b00001111;
										assign node2376 = (inp[1]) ? node2390 : node2377;
											assign node2377 = (inp[12]) ? node2385 : node2378;
												assign node2378 = (inp[3]) ? node2382 : node2379;
													assign node2379 = (inp[6]) ? 8'b00011110 : 8'b00001110;
													assign node2382 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node2385 = (inp[3]) ? 8'b00001110 : node2386;
													assign node2386 = (inp[6]) ? 8'b00001111 : 8'b00011111;
											assign node2390 = (inp[3]) ? node2398 : node2391;
												assign node2391 = (inp[6]) ? 8'b00011010 : node2392;
													assign node2392 = (inp[12]) ? 8'b00011010 : node2393;
														assign node2393 = (inp[2]) ? 8'b00001010 : 8'b00001011;
												assign node2398 = (inp[12]) ? node2404 : node2399;
													assign node2399 = (inp[6]) ? 8'b00011011 : node2400;
														assign node2400 = (inp[2]) ? 8'b00001011 : 8'b00001110;
													assign node2404 = (inp[6]) ? 8'b00001110 : 8'b00011011;
									assign node2407 = (inp[1]) ? node2437 : node2408;
										assign node2408 = (inp[3]) ? node2422 : node2409;
											assign node2409 = (inp[6]) ? node2417 : node2410;
												assign node2410 = (inp[11]) ? node2412 : 8'b00011011;
													assign node2412 = (inp[2]) ? 8'b00001010 : node2413;
														assign node2413 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node2417 = (inp[11]) ? node2419 : 8'b00001011;
													assign node2419 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node2422 = (inp[2]) ? node2428 : node2423;
												assign node2423 = (inp[6]) ? 8'b00000010 : node2424;
													assign node2424 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node2428 = (inp[6]) ? node2432 : node2429;
													assign node2429 = (inp[11]) ? 8'b10100101 : 8'b10010000;
													assign node2432 = (inp[12]) ? 8'b00000010 : node2433;
														assign node2433 = (inp[11]) ? 8'b11110111 : 8'b10000010;
										assign node2437 = (inp[11]) ? node2447 : node2438;
											assign node2438 = (inp[6]) ? node2444 : node2439;
												assign node2439 = (inp[3]) ? node2441 : 8'b10011001;
													assign node2441 = (inp[2]) ? 8'b10010000 : 8'b00011010;
												assign node2444 = (inp[3]) ? 8'b10000010 : 8'b10000001;
											assign node2447 = (inp[3]) ? node2453 : node2448;
												assign node2448 = (inp[2]) ? node2450 : 8'b10110100;
													assign node2450 = (inp[12]) ? 8'b10100101 : 8'b10100100;
												assign node2453 = (inp[2]) ? node2459 : node2454;
													assign node2454 = (inp[6]) ? 8'b11110111 : node2455;
														assign node2455 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node2459 = (inp[6]) ? node2463 : node2460;
														assign node2460 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node2463 = (inp[12]) ? 8'b00000010 : 8'b11110111;
							assign node2466 = (inp[10]) ? node2552 : node2467;
								assign node2467 = (inp[11]) ? node2495 : node2468;
									assign node2468 = (inp[3]) ? node2484 : node2469;
										assign node2469 = (inp[6]) ? node2475 : node2470;
											assign node2470 = (inp[1]) ? node2472 : 8'b10011101;
												assign node2472 = (inp[2]) ? 8'b10010101 : 8'b10011101;
											assign node2475 = (inp[7]) ? node2481 : node2476;
												assign node2476 = (inp[2]) ? node2478 : 8'b10011101;
													assign node2478 = (inp[12]) ? 8'b10000101 : 8'b10001101;
												assign node2481 = (inp[1]) ? 8'b10000101 : 8'b10001101;
										assign node2484 = (inp[7]) ? node2490 : node2485;
											assign node2485 = (inp[1]) ? node2487 : 8'b10011101;
												assign node2487 = (inp[2]) ? 8'b10000100 : 8'b10011100;
											assign node2490 = (inp[6]) ? 8'b10000100 : node2491;
												assign node2491 = (inp[2]) ? 8'b10010100 : 8'b10011100;
									assign node2495 = (inp[1]) ? node2523 : node2496;
										assign node2496 = (inp[7]) ? node2508 : node2497;
											assign node2497 = (inp[2]) ? node2501 : node2498;
												assign node2498 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node2501 = (inp[6]) ? node2505 : node2502;
													assign node2502 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node2505 = (inp[12]) ? 8'b10101101 : 8'b10111100;
											assign node2508 = (inp[2]) ? node2516 : node2509;
												assign node2509 = (inp[12]) ? 8'b10111100 : node2510;
													assign node2510 = (inp[6]) ? 8'b10111100 : node2511;
														assign node2511 = (inp[3]) ? 8'b10101100 : 8'b10101101;
												assign node2516 = (inp[3]) ? node2518 : 8'b10111100;
													assign node2518 = (inp[6]) ? node2520 : 8'b10110001;
														assign node2520 = (inp[12]) ? 8'b10100100 : 8'b10110001;
										assign node2523 = (inp[2]) ? node2537 : node2524;
											assign node2524 = (inp[3]) ? node2534 : node2525;
												assign node2525 = (inp[6]) ? node2529 : node2526;
													assign node2526 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node2529 = (inp[12]) ? node2531 : 8'b10110000;
														assign node2531 = (inp[7]) ? 8'b10100001 : 8'b10111001;
												assign node2534 = (inp[7]) ? 8'b10100100 : 8'b10101100;
											assign node2537 = (inp[3]) ? node2545 : node2538;
												assign node2538 = (inp[6]) ? node2542 : node2539;
													assign node2539 = (inp[12]) ? 8'b10110000 : 8'b10100000;
													assign node2542 = (inp[12]) ? 8'b10100001 : 8'b10110000;
												assign node2545 = (inp[7]) ? node2549 : node2546;
													assign node2546 = (inp[6]) ? 8'b10110001 : 8'b10100001;
													assign node2549 = (inp[6]) ? 8'b10100100 : 8'b10110001;
								assign node2552 = (inp[1]) ? node2604 : node2553;
									assign node2553 = (inp[6]) ? node2579 : node2554;
										assign node2554 = (inp[12]) ? node2564 : node2555;
											assign node2555 = (inp[11]) ? node2561 : node2556;
												assign node2556 = (inp[7]) ? node2558 : 8'b00011011;
													assign node2558 = (inp[3]) ? 8'b00011010 : 8'b00011011;
												assign node2561 = (inp[2]) ? 8'b00001010 : 8'b00001011;
											assign node2564 = (inp[7]) ? node2570 : node2565;
												assign node2565 = (inp[11]) ? node2567 : 8'b00011011;
													assign node2567 = (inp[2]) ? 8'b00011010 : 8'b00011011;
												assign node2570 = (inp[3]) ? node2574 : node2571;
													assign node2571 = (inp[11]) ? 8'b00011010 : 8'b00011011;
													assign node2574 = (inp[2]) ? node2576 : 8'b00011010;
														assign node2576 = (inp[11]) ? 8'b11110101 : 8'b10010000;
										assign node2579 = (inp[7]) ? node2593 : node2580;
											assign node2580 = (inp[2]) ? node2586 : node2581;
												assign node2581 = (inp[11]) ? node2583 : 8'b00011011;
													assign node2583 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node2586 = (inp[3]) ? 8'b00001011 : node2587;
													assign node2587 = (inp[11]) ? node2589 : 8'b00001011;
														assign node2589 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node2593 = (inp[3]) ? node2599 : node2594;
												assign node2594 = (inp[11]) ? node2596 : 8'b00001011;
													assign node2596 = (inp[12]) ? 8'b00001011 : 8'b00011010;
												assign node2599 = (inp[12]) ? 8'b00000010 : node2600;
													assign node2600 = (inp[11]) ? 8'b11110111 : 8'b10000010;
									assign node2604 = (inp[3]) ? node2630 : node2605;
										assign node2605 = (inp[11]) ? node2615 : node2606;
											assign node2606 = (inp[2]) ? node2612 : node2607;
												assign node2607 = (inp[7]) ? node2609 : 8'b10011001;
													assign node2609 = (inp[6]) ? 8'b10000001 : 8'b10011001;
												assign node2612 = (inp[6]) ? 8'b10000001 : 8'b10010001;
											assign node2615 = (inp[2]) ? node2623 : node2616;
												assign node2616 = (inp[12]) ? 8'b11111101 : node2617;
													assign node2617 = (inp[7]) ? node2619 : 8'b10101101;
														assign node2619 = (inp[6]) ? 8'b10110100 : 8'b10101101;
												assign node2623 = (inp[7]) ? 8'b10110100 : node2624;
													assign node2624 = (inp[6]) ? 8'b10100101 : node2625;
														assign node2625 = (inp[12]) ? 8'b10110100 : 8'b10100100;
										assign node2630 = (inp[2]) ? node2644 : node2631;
											assign node2631 = (inp[7]) ? node2637 : node2632;
												assign node2632 = (inp[11]) ? node2634 : 8'b00011010;
													assign node2634 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node2637 = (inp[6]) ? node2641 : node2638;
													assign node2638 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node2641 = (inp[12]) ? 8'b00000010 : 8'b10000010;
											assign node2644 = (inp[6]) ? node2650 : node2645;
												assign node2645 = (inp[11]) ? node2647 : 8'b10010000;
													assign node2647 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node2650 = (inp[12]) ? 8'b00000010 : 8'b10000010;
				assign node2653 = (inp[11]) ? node3073 : node2654;
					assign node2654 = (inp[0]) ? node2992 : node2655;
						assign node2655 = (inp[9]) ? node2811 : node2656;
							assign node2656 = (inp[8]) ? node2734 : node2657;
								assign node2657 = (inp[7]) ? node2675 : node2658;
									assign node2658 = (inp[2]) ? node2664 : node2659;
										assign node2659 = (inp[1]) ? node2661 : 8'b00011111;
											assign node2661 = (inp[3]) ? 8'b00011111 : 8'b00011110;
										assign node2664 = (inp[6]) ? node2670 : node2665;
											assign node2665 = (inp[1]) ? node2667 : 8'b00001111;
												assign node2667 = (inp[3]) ? 8'b00001111 : 8'b00001110;
											assign node2670 = (inp[1]) ? node2672 : 8'b00011111;
												assign node2672 = (inp[3]) ? 8'b00011111 : 8'b00011110;
									assign node2675 = (inp[10]) ? node2703 : node2676;
										assign node2676 = (inp[2]) ? node2692 : node2677;
											assign node2677 = (inp[6]) ? node2685 : node2678;
												assign node2678 = (inp[3]) ? node2682 : node2679;
													assign node2679 = (inp[1]) ? 8'b00011110 : 8'b00011111;
													assign node2682 = (inp[1]) ? 8'b00011111 : 8'b00011110;
												assign node2685 = (inp[3]) ? node2689 : node2686;
													assign node2686 = (inp[1]) ? 8'b00001110 : 8'b00001111;
													assign node2689 = (inp[1]) ? 8'b00001111 : 8'b00001110;
											assign node2692 = (inp[6]) ? node2698 : node2693;
												assign node2693 = (inp[1]) ? 8'b00001111 : node2694;
													assign node2694 = (inp[3]) ? 8'b00001110 : 8'b00001111;
												assign node2698 = (inp[1]) ? 8'b00011111 : node2699;
													assign node2699 = (inp[3]) ? 8'b00011110 : 8'b00011111;
										assign node2703 = (inp[1]) ? node2717 : node2704;
											assign node2704 = (inp[3]) ? node2710 : node2705;
												assign node2705 = (inp[2]) ? node2707 : 8'b00001011;
													assign node2707 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node2710 = (inp[12]) ? node2712 : 8'b10000010;
													assign node2712 = (inp[2]) ? 8'b10010000 : node2713;
														assign node2713 = (inp[6]) ? 8'b00000010 : 8'b00011010;
											assign node2717 = (inp[3]) ? node2727 : node2718;
												assign node2718 = (inp[6]) ? node2722 : node2719;
													assign node2719 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node2722 = (inp[2]) ? 8'b10010000 : node2723;
														assign node2723 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node2727 = (inp[2]) ? node2731 : node2728;
													assign node2728 = (inp[6]) ? 8'b10000001 : 8'b10011001;
													assign node2731 = (inp[6]) ? 8'b10010001 : 8'b10000001;
								assign node2734 = (inp[10]) ? node2772 : node2735;
									assign node2735 = (inp[1]) ? node2755 : node2736;
										assign node2736 = (inp[7]) ? node2742 : node2737;
											assign node2737 = (inp[2]) ? node2739 : 8'b00011011;
												assign node2739 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node2742 = (inp[3]) ? node2750 : node2743;
												assign node2743 = (inp[12]) ? 8'b00011011 : node2744;
													assign node2744 = (inp[2]) ? node2746 : 8'b00001011;
														assign node2746 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node2750 = (inp[2]) ? node2752 : 8'b00011010;
													assign node2752 = (inp[6]) ? 8'b10010000 : 8'b10000010;
										assign node2755 = (inp[3]) ? node2763 : node2756;
											assign node2756 = (inp[2]) ? 8'b10010000 : node2757;
												assign node2757 = (inp[7]) ? node2759 : 8'b00011010;
													assign node2759 = (inp[6]) ? 8'b00000010 : 8'b00011010;
											assign node2763 = (inp[2]) ? node2769 : node2764;
												assign node2764 = (inp[7]) ? node2766 : 8'b10011001;
													assign node2766 = (inp[6]) ? 8'b10000001 : 8'b10011001;
												assign node2769 = (inp[6]) ? 8'b10010001 : 8'b10000001;
									assign node2772 = (inp[1]) ? node2792 : node2773;
										assign node2773 = (inp[3]) ? node2783 : node2774;
											assign node2774 = (inp[2]) ? node2780 : node2775;
												assign node2775 = (inp[7]) ? node2777 : 8'b10011101;
													assign node2777 = (inp[6]) ? 8'b10001101 : 8'b10011101;
												assign node2780 = (inp[6]) ? 8'b10011101 : 8'b10001101;
											assign node2783 = (inp[7]) ? node2787 : node2784;
												assign node2784 = (inp[2]) ? 8'b10001101 : 8'b10011101;
												assign node2787 = (inp[2]) ? 8'b10000100 : node2788;
													assign node2788 = (inp[6]) ? 8'b10000100 : 8'b10011100;
										assign node2792 = (inp[3]) ? node2802 : node2793;
											assign node2793 = (inp[6]) ? node2795 : 8'b10000100;
												assign node2795 = (inp[7]) ? node2799 : node2796;
													assign node2796 = (inp[2]) ? 8'b10010100 : 8'b10011100;
													assign node2799 = (inp[2]) ? 8'b10010100 : 8'b10000100;
											assign node2802 = (inp[2]) ? node2808 : node2803;
												assign node2803 = (inp[6]) ? node2805 : 8'b10011101;
													assign node2805 = (inp[7]) ? 8'b10000101 : 8'b10011101;
												assign node2808 = (inp[7]) ? 8'b10000101 : 8'b10010101;
							assign node2811 = (inp[7]) ? node2863 : node2812;
								assign node2812 = (inp[1]) ? node2828 : node2813;
									assign node2813 = (inp[8]) ? node2819 : node2814;
										assign node2814 = (inp[2]) ? node2816 : 8'b11111101;
											assign node2816 = (inp[6]) ? 8'b11111101 : 8'b10101101;
										assign node2819 = (inp[10]) ? node2823 : node2820;
											assign node2820 = (inp[2]) ? 8'b10101001 : 8'b10111001;
											assign node2823 = (inp[2]) ? node2825 : 8'b11111101;
												assign node2825 = (inp[6]) ? 8'b11111101 : 8'b10101101;
									assign node2828 = (inp[3]) ? node2844 : node2829;
										assign node2829 = (inp[8]) ? node2835 : node2830;
											assign node2830 = (inp[6]) ? 8'b10111100 : node2831;
												assign node2831 = (inp[2]) ? 8'b10101100 : 8'b10111100;
											assign node2835 = (inp[2]) ? node2839 : node2836;
												assign node2836 = (inp[10]) ? 8'b10111100 : 8'b10111000;
												assign node2839 = (inp[10]) ? 8'b10110100 : node2840;
													assign node2840 = (inp[6]) ? 8'b10110000 : 8'b10100000;
										assign node2844 = (inp[8]) ? node2852 : node2845;
											assign node2845 = (inp[12]) ? node2847 : 8'b11111101;
												assign node2847 = (inp[10]) ? 8'b11111101 : node2848;
													assign node2848 = (inp[6]) ? 8'b11111101 : 8'b10101101;
											assign node2852 = (inp[2]) ? node2856 : node2853;
												assign node2853 = (inp[10]) ? 8'b11111101 : 8'b10111001;
												assign node2856 = (inp[6]) ? node2860 : node2857;
													assign node2857 = (inp[10]) ? 8'b10100101 : 8'b10100001;
													assign node2860 = (inp[10]) ? 8'b11110101 : 8'b10110001;
								assign node2863 = (inp[6]) ? node2933 : node2864;
									assign node2864 = (inp[2]) ? node2906 : node2865;
										assign node2865 = (inp[3]) ? node2885 : node2866;
											assign node2866 = (inp[1]) ? node2878 : node2867;
												assign node2867 = (inp[12]) ? node2873 : node2868;
													assign node2868 = (inp[8]) ? node2870 : 8'b11111101;
														assign node2870 = (inp[10]) ? 8'b11111101 : 8'b10111001;
													assign node2873 = (inp[8]) ? 8'b11111101 : node2874;
														assign node2874 = (inp[10]) ? 8'b10111001 : 8'b11111101;
												assign node2878 = (inp[12]) ? node2880 : 8'b10111100;
													assign node2880 = (inp[8]) ? node2882 : 8'b10111100;
														assign node2882 = (inp[10]) ? 8'b10111100 : 8'b10111000;
											assign node2885 = (inp[1]) ? node2899 : node2886;
												assign node2886 = (inp[12]) ? node2892 : node2887;
													assign node2887 = (inp[10]) ? node2889 : 8'b10111100;
														assign node2889 = (inp[8]) ? 8'b10111100 : 8'b10111000;
													assign node2892 = (inp[8]) ? node2896 : node2893;
														assign node2893 = (inp[10]) ? 8'b10111000 : 8'b10111100;
														assign node2896 = (inp[10]) ? 8'b10111100 : 8'b10111000;
												assign node2899 = (inp[10]) ? node2903 : node2900;
													assign node2900 = (inp[8]) ? 8'b10111001 : 8'b11111101;
													assign node2903 = (inp[8]) ? 8'b11111101 : 8'b10111001;
										assign node2906 = (inp[1]) ? node2918 : node2907;
											assign node2907 = (inp[3]) ? node2913 : node2908;
												assign node2908 = (inp[10]) ? 8'b10101101 : node2909;
													assign node2909 = (inp[8]) ? 8'b10101001 : 8'b10101101;
												assign node2913 = (inp[10]) ? node2915 : 8'b10101100;
													assign node2915 = (inp[8]) ? 8'b10100100 : 8'b10100000;
											assign node2918 = (inp[3]) ? node2928 : node2919;
												assign node2919 = (inp[12]) ? node2921 : 8'b10100000;
													assign node2921 = (inp[10]) ? node2925 : node2922;
														assign node2922 = (inp[8]) ? 8'b10100000 : 8'b10101100;
														assign node2925 = (inp[8]) ? 8'b10100100 : 8'b10100000;
												assign node2928 = (inp[8]) ? node2930 : 8'b10101101;
													assign node2930 = (inp[10]) ? 8'b10100101 : 8'b10100001;
									assign node2933 = (inp[2]) ? node2971 : node2934;
										assign node2934 = (inp[8]) ? node2952 : node2935;
											assign node2935 = (inp[10]) ? node2945 : node2936;
												assign node2936 = (inp[12]) ? node2938 : 8'b10101101;
													assign node2938 = (inp[1]) ? node2942 : node2939;
														assign node2939 = (inp[3]) ? 8'b10101100 : 8'b10101101;
														assign node2942 = (inp[3]) ? 8'b10101101 : 8'b10101100;
												assign node2945 = (inp[3]) ? node2949 : node2946;
													assign node2946 = (inp[1]) ? 8'b10100000 : 8'b10101001;
													assign node2949 = (inp[1]) ? 8'b10100001 : 8'b10100000;
											assign node2952 = (inp[10]) ? node2964 : node2953;
												assign node2953 = (inp[12]) ? node2959 : node2954;
													assign node2954 = (inp[1]) ? node2956 : 8'b10100000;
														assign node2956 = (inp[3]) ? 8'b10100001 : 8'b10100000;
													assign node2959 = (inp[1]) ? node2961 : 8'b10101001;
														assign node2961 = (inp[3]) ? 8'b10100001 : 8'b10100000;
												assign node2964 = (inp[3]) ? node2968 : node2965;
													assign node2965 = (inp[1]) ? 8'b10100100 : 8'b10101101;
													assign node2968 = (inp[1]) ? 8'b10100101 : 8'b10100100;
										assign node2971 = (inp[8]) ? node2979 : node2972;
											assign node2972 = (inp[10]) ? 8'b10111001 : node2973;
												assign node2973 = (inp[1]) ? node2975 : 8'b11111101;
													assign node2975 = (inp[3]) ? 8'b11111101 : 8'b10111100;
											assign node2979 = (inp[10]) ? node2987 : node2980;
												assign node2980 = (inp[1]) ? node2984 : node2981;
													assign node2981 = (inp[3]) ? 8'b10110000 : 8'b10111001;
													assign node2984 = (inp[3]) ? 8'b10110001 : 8'b10110000;
												assign node2987 = (inp[1]) ? node2989 : 8'b11111101;
													assign node2989 = (inp[3]) ? 8'b11110101 : 8'b10110100;
						assign node2992 = (inp[7]) ? node3000 : node2993;
							assign node2993 = (inp[1]) ? node2995 : 8'b11111101;
								assign node2995 = (inp[2]) ? node2997 : 8'b11111101;
									assign node2997 = (inp[8]) ? 8'b11110101 : 8'b11111101;
							assign node3000 = (inp[2]) ? node3048 : node3001;
								assign node3001 = (inp[6]) ? node3019 : node3002;
									assign node3002 = (inp[8]) ? node3014 : node3003;
										assign node3003 = (inp[10]) ? node3009 : node3004;
											assign node3004 = (inp[3]) ? node3006 : 8'b11111101;
												assign node3006 = (inp[1]) ? 8'b11111101 : 8'b10111100;
											assign node3009 = (inp[1]) ? 8'b10111001 : node3010;
												assign node3010 = (inp[3]) ? 8'b10111000 : 8'b10111001;
										assign node3014 = (inp[1]) ? 8'b11111101 : node3015;
											assign node3015 = (inp[3]) ? 8'b10111100 : 8'b11111101;
									assign node3019 = (inp[3]) ? node3033 : node3020;
										assign node3020 = (inp[1]) ? node3026 : node3021;
											assign node3021 = (inp[8]) ? 8'b10101101 : node3022;
												assign node3022 = (inp[10]) ? 8'b10101001 : 8'b10101101;
											assign node3026 = (inp[10]) ? node3030 : node3027;
												assign node3027 = (inp[8]) ? 8'b10100101 : 8'b10101101;
												assign node3030 = (inp[8]) ? 8'b10100101 : 8'b10100001;
										assign node3033 = (inp[1]) ? node3041 : node3034;
											assign node3034 = (inp[10]) ? node3038 : node3035;
												assign node3035 = (inp[8]) ? 8'b10100100 : 8'b10101100;
												assign node3038 = (inp[8]) ? 8'b10100100 : 8'b10100000;
											assign node3041 = (inp[10]) ? node3045 : node3042;
												assign node3042 = (inp[8]) ? 8'b10100101 : 8'b10101101;
												assign node3045 = (inp[8]) ? 8'b10100101 : 8'b10100001;
								assign node3048 = (inp[3]) ? node3062 : node3049;
									assign node3049 = (inp[10]) ? node3055 : node3050;
										assign node3050 = (inp[8]) ? node3052 : 8'b11111101;
											assign node3052 = (inp[1]) ? 8'b11110101 : 8'b11111101;
										assign node3055 = (inp[8]) ? node3059 : node3056;
											assign node3056 = (inp[1]) ? 8'b10110001 : 8'b10111001;
											assign node3059 = (inp[1]) ? 8'b11110101 : 8'b11111101;
									assign node3062 = (inp[1]) ? node3068 : node3063;
										assign node3063 = (inp[8]) ? 8'b10110100 : node3064;
											assign node3064 = (inp[10]) ? 8'b10110000 : 8'b10111100;
										assign node3068 = (inp[8]) ? 8'b11110101 : node3069;
											assign node3069 = (inp[10]) ? 8'b10110001 : 8'b11111101;
					assign node3073 = (inp[2]) ? node3417 : node3074;
						assign node3074 = (inp[0]) ? node3332 : node3075;
							assign node3075 = (inp[9]) ? node3209 : node3076;
								assign node3076 = (inp[8]) ? node3142 : node3077;
									assign node3077 = (inp[7]) ? node3089 : node3078;
										assign node3078 = (inp[12]) ? node3084 : node3079;
											assign node3079 = (inp[1]) ? node3081 : 8'b00001111;
												assign node3081 = (inp[3]) ? 8'b00001011 : 8'b00001110;
											assign node3084 = (inp[1]) ? node3086 : 8'b00011111;
												assign node3086 = (inp[3]) ? 8'b00011011 : 8'b00011110;
										assign node3089 = (inp[10]) ? node3117 : node3090;
											assign node3090 = (inp[1]) ? node3102 : node3091;
												assign node3091 = (inp[3]) ? node3097 : node3092;
													assign node3092 = (inp[6]) ? 8'b00001111 : node3093;
														assign node3093 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node3097 = (inp[6]) ? 8'b00001110 : node3098;
														assign node3098 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node3102 = (inp[3]) ? node3110 : node3103;
													assign node3103 = (inp[6]) ? node3107 : node3104;
														assign node3104 = (inp[12]) ? 8'b00011110 : 8'b00001110;
														assign node3107 = (inp[12]) ? 8'b00001110 : 8'b00011011;
													assign node3110 = (inp[6]) ? node3114 : node3111;
														assign node3111 = (inp[12]) ? 8'b00011011 : 8'b00001011;
														assign node3114 = (inp[12]) ? 8'b00001011 : 8'b00011010;
											assign node3117 = (inp[3]) ? node3129 : node3118;
												assign node3118 = (inp[6]) ? node3124 : node3119;
													assign node3119 = (inp[12]) ? node3121 : 8'b00001011;
														assign node3121 = (inp[1]) ? 8'b00011010 : 8'b00011011;
													assign node3124 = (inp[1]) ? node3126 : 8'b00011010;
														assign node3126 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node3129 = (inp[1]) ? node3135 : node3130;
													assign node3130 = (inp[6]) ? node3132 : 8'b00001010;
														assign node3132 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node3135 = (inp[6]) ? node3139 : node3136;
														assign node3136 = (inp[12]) ? 8'b11111101 : 8'b10101101;
														assign node3139 = (inp[12]) ? 8'b10100101 : 8'b10110100;
									assign node3142 = (inp[10]) ? node3176 : node3143;
										assign node3143 = (inp[3]) ? node3163 : node3144;
											assign node3144 = (inp[1]) ? node3154 : node3145;
												assign node3145 = (inp[12]) ? node3149 : node3146;
													assign node3146 = (inp[7]) ? 8'b00011010 : 8'b00001011;
													assign node3149 = (inp[6]) ? node3151 : 8'b00011011;
														assign node3151 = (inp[7]) ? 8'b00001011 : 8'b00011011;
												assign node3154 = (inp[12]) ? node3158 : node3155;
													assign node3155 = (inp[7]) ? 8'b11110111 : 8'b00001010;
													assign node3158 = (inp[6]) ? node3160 : 8'b00011010;
														assign node3160 = (inp[7]) ? 8'b00000010 : 8'b00011010;
											assign node3163 = (inp[1]) ? node3169 : node3164;
												assign node3164 = (inp[7]) ? 8'b11110111 : node3165;
													assign node3165 = (inp[12]) ? 8'b00011011 : 8'b00001011;
												assign node3169 = (inp[12]) ? node3171 : 8'b10101101;
													assign node3171 = (inp[7]) ? node3173 : 8'b11111101;
														assign node3173 = (inp[6]) ? 8'b10100101 : 8'b11111101;
										assign node3176 = (inp[1]) ? node3192 : node3177;
											assign node3177 = (inp[7]) ? node3181 : node3178;
												assign node3178 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node3181 = (inp[3]) ? node3187 : node3182;
													assign node3182 = (inp[6]) ? 8'b10111100 : node3183;
														assign node3183 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node3187 = (inp[6]) ? 8'b10100100 : node3188;
														assign node3188 = (inp[12]) ? 8'b10111100 : 8'b10101100;
											assign node3192 = (inp[3]) ? node3202 : node3193;
												assign node3193 = (inp[7]) ? node3197 : node3194;
													assign node3194 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node3197 = (inp[6]) ? node3199 : 8'b10101100;
														assign node3199 = (inp[12]) ? 8'b10100100 : 8'b10110001;
												assign node3202 = (inp[6]) ? node3206 : node3203;
													assign node3203 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node3206 = (inp[12]) ? 8'b10100001 : 8'b10101001;
								assign node3209 = (inp[8]) ? node3265 : node3210;
									assign node3210 = (inp[7]) ? node3222 : node3211;
										assign node3211 = (inp[12]) ? node3217 : node3212;
											assign node3212 = (inp[1]) ? node3214 : 8'b10101101;
												assign node3214 = (inp[3]) ? 8'b10101001 : 8'b10101100;
											assign node3217 = (inp[1]) ? node3219 : 8'b11111101;
												assign node3219 = (inp[3]) ? 8'b10111001 : 8'b10111100;
										assign node3222 = (inp[10]) ? node3248 : node3223;
											assign node3223 = (inp[6]) ? node3233 : node3224;
												assign node3224 = (inp[12]) ? node3228 : node3225;
													assign node3225 = (inp[3]) ? 8'b10101100 : 8'b10101101;
													assign node3228 = (inp[1]) ? 8'b10111100 : node3229;
														assign node3229 = (inp[3]) ? 8'b10111100 : 8'b11111101;
												assign node3233 = (inp[12]) ? node3241 : node3234;
													assign node3234 = (inp[3]) ? node3238 : node3235;
														assign node3235 = (inp[1]) ? 8'b10111001 : 8'b10111100;
														assign node3238 = (inp[1]) ? 8'b10111000 : 8'b10111001;
													assign node3241 = (inp[1]) ? node3245 : node3242;
														assign node3242 = (inp[3]) ? 8'b10101100 : 8'b10101101;
														assign node3245 = (inp[3]) ? 8'b10101001 : 8'b10101100;
											assign node3248 = (inp[6]) ? node3254 : node3249;
												assign node3249 = (inp[12]) ? node3251 : 8'b10101000;
													assign node3251 = (inp[1]) ? 8'b10011101 : 8'b10111000;
												assign node3254 = (inp[1]) ? node3260 : node3255;
													assign node3255 = (inp[3]) ? node3257 : 8'b10111000;
														assign node3257 = (inp[12]) ? 8'b10100000 : 8'b10010101;
													assign node3260 = (inp[12]) ? 8'b10000101 : node3261;
														assign node3261 = (inp[3]) ? 8'b10010100 : 8'b10010101;
									assign node3265 = (inp[10]) ? node3305 : node3266;
										assign node3266 = (inp[3]) ? node3288 : node3267;
											assign node3267 = (inp[1]) ? node3277 : node3268;
												assign node3268 = (inp[12]) ? node3272 : node3269;
													assign node3269 = (inp[6]) ? 8'b10111000 : 8'b10101001;
													assign node3272 = (inp[7]) ? node3274 : 8'b10111001;
														assign node3274 = (inp[6]) ? 8'b10101001 : 8'b10111001;
												assign node3277 = (inp[12]) ? node3283 : node3278;
													assign node3278 = (inp[7]) ? node3280 : 8'b10101000;
														assign node3280 = (inp[6]) ? 8'b10010101 : 8'b10101000;
													assign node3283 = (inp[7]) ? node3285 : 8'b10111000;
														assign node3285 = (inp[6]) ? 8'b10100000 : 8'b10111000;
											assign node3288 = (inp[1]) ? node3294 : node3289;
												assign node3289 = (inp[7]) ? node3291 : 8'b10101001;
													assign node3291 = (inp[6]) ? 8'b10010101 : 8'b10111000;
												assign node3294 = (inp[6]) ? node3298 : node3295;
													assign node3295 = (inp[12]) ? 8'b10011101 : 8'b10001101;
													assign node3298 = (inp[7]) ? node3302 : node3299;
														assign node3299 = (inp[12]) ? 8'b10011101 : 8'b10001101;
														assign node3302 = (inp[12]) ? 8'b10000101 : 8'b10010100;
										assign node3305 = (inp[1]) ? node3319 : node3306;
											assign node3306 = (inp[6]) ? node3312 : node3307;
												assign node3307 = (inp[3]) ? node3309 : 8'b10001101;
													assign node3309 = (inp[7]) ? 8'b10001100 : 8'b10001101;
												assign node3312 = (inp[12]) ? node3314 : 8'b10010001;
													assign node3314 = (inp[7]) ? node3316 : 8'b10011101;
														assign node3316 = (inp[3]) ? 8'b10000100 : 8'b10001101;
											assign node3319 = (inp[3]) ? node3327 : node3320;
												assign node3320 = (inp[7]) ? node3324 : node3321;
													assign node3321 = (inp[12]) ? 8'b10011100 : 8'b10001100;
													assign node3324 = (inp[12]) ? 8'b10000100 : 8'b10010001;
												assign node3327 = (inp[12]) ? 8'b10011001 : node3328;
													assign node3328 = (inp[6]) ? 8'b10010000 : 8'b10001001;
							assign node3332 = (inp[8]) ? node3386 : node3333;
								assign node3333 = (inp[1]) ? node3367 : node3334;
									assign node3334 = (inp[7]) ? node3338 : node3335;
										assign node3335 = (inp[12]) ? 8'b11111101 : 8'b10101101;
										assign node3338 = (inp[10]) ? node3354 : node3339;
											assign node3339 = (inp[3]) ? node3347 : node3340;
												assign node3340 = (inp[6]) ? node3344 : node3341;
													assign node3341 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node3344 = (inp[12]) ? 8'b10101101 : 8'b10111100;
												assign node3347 = (inp[12]) ? node3351 : node3348;
													assign node3348 = (inp[6]) ? 8'b10111001 : 8'b10101100;
													assign node3351 = (inp[6]) ? 8'b10101100 : 8'b10111100;
											assign node3354 = (inp[3]) ? node3360 : node3355;
												assign node3355 = (inp[12]) ? node3357 : 8'b10111000;
													assign node3357 = (inp[6]) ? 8'b10101001 : 8'b10111001;
												assign node3360 = (inp[6]) ? node3364 : node3361;
													assign node3361 = (inp[9]) ? 8'b10111000 : 8'b10101000;
													assign node3364 = (inp[12]) ? 8'b10100000 : 8'b10010101;
									assign node3367 = (inp[7]) ? node3371 : node3368;
										assign node3368 = (inp[12]) ? 8'b10111001 : 8'b10101001;
										assign node3371 = (inp[10]) ? node3379 : node3372;
											assign node3372 = (inp[6]) ? node3376 : node3373;
												assign node3373 = (inp[12]) ? 8'b10111001 : 8'b10101001;
												assign node3376 = (inp[12]) ? 8'b10101001 : 8'b10111000;
											assign node3379 = (inp[6]) ? node3383 : node3380;
												assign node3380 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node3383 = (inp[9]) ? 8'b10010100 : 8'b10000101;
								assign node3386 = (inp[1]) ? node3406 : node3387;
									assign node3387 = (inp[7]) ? node3391 : node3388;
										assign node3388 = (inp[12]) ? 8'b10011101 : 8'b10001101;
										assign node3391 = (inp[3]) ? node3399 : node3392;
											assign node3392 = (inp[6]) ? node3396 : node3393;
												assign node3393 = (inp[12]) ? 8'b10011101 : 8'b10001101;
												assign node3396 = (inp[12]) ? 8'b10001101 : 8'b10011100;
											assign node3399 = (inp[6]) ? node3403 : node3400;
												assign node3400 = (inp[12]) ? 8'b10011100 : 8'b10001100;
												assign node3403 = (inp[12]) ? 8'b10000100 : 8'b10010001;
									assign node3406 = (inp[12]) ? node3412 : node3407;
										assign node3407 = (inp[6]) ? node3409 : 8'b10001001;
											assign node3409 = (inp[7]) ? 8'b10010000 : 8'b10001001;
										assign node3412 = (inp[7]) ? node3414 : 8'b10011001;
											assign node3414 = (inp[6]) ? 8'b10000001 : 8'b10011001;
						assign node3417 = (inp[8]) ? node3601 : node3418;
							assign node3418 = (inp[0]) ? node3566 : node3419;
								assign node3419 = (inp[9]) ? node3499 : node3420;
									assign node3420 = (inp[10]) ? node3450 : node3421;
										assign node3421 = (inp[1]) ? node3439 : node3422;
											assign node3422 = (inp[3]) ? node3430 : node3423;
												assign node3423 = (inp[6]) ? node3427 : node3424;
													assign node3424 = (inp[12]) ? 8'b00001111 : 8'b00011110;
													assign node3427 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node3430 = (inp[6]) ? node3436 : node3431;
													assign node3431 = (inp[12]) ? 8'b00001110 : node3432;
														assign node3432 = (inp[7]) ? 8'b00011011 : 8'b00011110;
													assign node3436 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node3439 = (inp[6]) ? node3445 : node3440;
												assign node3440 = (inp[12]) ? node3442 : 8'b00011011;
													assign node3442 = (inp[3]) ? 8'b00001011 : 8'b00001110;
												assign node3445 = (inp[3]) ? node3447 : 8'b00011011;
													assign node3447 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node3450 = (inp[7]) ? node3472 : node3451;
											assign node3451 = (inp[1]) ? node3459 : node3452;
												assign node3452 = (inp[3]) ? node3454 : 8'b00001111;
													assign node3454 = (inp[6]) ? node3456 : 8'b00011110;
														assign node3456 = (inp[12]) ? 8'b00011110 : 8'b00001110;
												assign node3459 = (inp[3]) ? node3467 : node3460;
													assign node3460 = (inp[6]) ? node3464 : node3461;
														assign node3461 = (inp[12]) ? 8'b00001110 : 8'b00011011;
														assign node3464 = (inp[12]) ? 8'b00011011 : 8'b00001011;
													assign node3467 = (inp[12]) ? node3469 : 8'b00011010;
														assign node3469 = (inp[6]) ? 8'b00011010 : 8'b00001011;
											assign node3472 = (inp[1]) ? node3486 : node3473;
												assign node3473 = (inp[3]) ? node3481 : node3474;
													assign node3474 = (inp[12]) ? node3478 : node3475;
														assign node3475 = (inp[6]) ? 8'b00001010 : 8'b00011010;
														assign node3478 = (inp[6]) ? 8'b00011010 : 8'b00001011;
													assign node3481 = (inp[6]) ? 8'b11110101 : node3482;
														assign node3482 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node3486 = (inp[3]) ? node3492 : node3487;
													assign node3487 = (inp[12]) ? 8'b00000010 : node3488;
														assign node3488 = (inp[6]) ? 8'b10100101 : 8'b11110111;
													assign node3492 = (inp[6]) ? node3496 : node3493;
														assign node3493 = (inp[12]) ? 8'b10100101 : 8'b10110100;
														assign node3496 = (inp[12]) ? 8'b10110100 : 8'b10100100;
									assign node3499 = (inp[7]) ? node3525 : node3500;
										assign node3500 = (inp[1]) ? node3508 : node3501;
											assign node3501 = (inp[12]) ? node3505 : node3502;
												assign node3502 = (inp[6]) ? 8'b10101100 : 8'b10111100;
												assign node3505 = (inp[6]) ? 8'b10111100 : 8'b10101101;
											assign node3508 = (inp[3]) ? node3518 : node3509;
												assign node3509 = (inp[10]) ? node3511 : 8'b10111001;
													assign node3511 = (inp[12]) ? node3515 : node3512;
														assign node3512 = (inp[6]) ? 8'b10101001 : 8'b10111001;
														assign node3515 = (inp[6]) ? 8'b10111001 : 8'b10101100;
												assign node3518 = (inp[10]) ? 8'b10111000 : node3519;
													assign node3519 = (inp[12]) ? 8'b10101001 : node3520;
														assign node3520 = (inp[6]) ? 8'b10101000 : 8'b10111000;
										assign node3525 = (inp[10]) ? node3543 : node3526;
											assign node3526 = (inp[3]) ? node3538 : node3527;
												assign node3527 = (inp[1]) ? node3535 : node3528;
													assign node3528 = (inp[6]) ? node3532 : node3529;
														assign node3529 = (inp[12]) ? 8'b10101101 : 8'b10111100;
														assign node3532 = (inp[12]) ? 8'b10111100 : 8'b10101100;
													assign node3535 = (inp[12]) ? 8'b10101100 : 8'b10101001;
												assign node3538 = (inp[6]) ? 8'b10111000 : node3539;
													assign node3539 = (inp[1]) ? 8'b10101001 : 8'b10111001;
											assign node3543 = (inp[1]) ? node3555 : node3544;
												assign node3544 = (inp[3]) ? node3550 : node3545;
													assign node3545 = (inp[12]) ? 8'b10101001 : node3546;
														assign node3546 = (inp[6]) ? 8'b10101000 : 8'b10111000;
													assign node3550 = (inp[12]) ? 8'b10100000 : node3551;
														assign node3551 = (inp[6]) ? 8'b10000101 : 8'b10010101;
												assign node3555 = (inp[3]) ? node3561 : node3556;
													assign node3556 = (inp[12]) ? 8'b10010101 : node3557;
														assign node3557 = (inp[6]) ? 8'b10000101 : 8'b10010101;
													assign node3561 = (inp[12]) ? node3563 : 8'b10010100;
														assign node3563 = (inp[6]) ? 8'b10010100 : 8'b10000101;
								assign node3566 = (inp[12]) ? node3584 : node3567;
									assign node3567 = (inp[10]) ? node3575 : node3568;
										assign node3568 = (inp[1]) ? 8'b10101000 : node3569;
											assign node3569 = (inp[3]) ? node3571 : 8'b10101100;
												assign node3571 = (inp[7]) ? 8'b10101001 : 8'b10101100;
										assign node3575 = (inp[7]) ? node3579 : node3576;
											assign node3576 = (inp[1]) ? 8'b10101000 : 8'b10101100;
											assign node3579 = (inp[1]) ? 8'b10000100 : node3580;
												assign node3580 = (inp[3]) ? 8'b10000101 : 8'b10101000;
									assign node3584 = (inp[10]) ? node3592 : node3585;
										assign node3585 = (inp[1]) ? 8'b10111000 : node3586;
											assign node3586 = (inp[7]) ? node3588 : 8'b10111100;
												assign node3588 = (inp[3]) ? 8'b10111001 : 8'b10111100;
										assign node3592 = (inp[7]) ? node3596 : node3593;
											assign node3593 = (inp[1]) ? 8'b10111000 : 8'b10111100;
											assign node3596 = (inp[1]) ? 8'b10010100 : node3597;
												assign node3597 = (inp[3]) ? 8'b10010101 : 8'b10111000;
							assign node3601 = (inp[1]) ? node3687 : node3602;
								assign node3602 = (inp[0]) ? node3676 : node3603;
									assign node3603 = (inp[10]) ? node3641 : node3604;
										assign node3604 = (inp[9]) ? node3626 : node3605;
											assign node3605 = (inp[3]) ? node3613 : node3606;
												assign node3606 = (inp[6]) ? node3610 : node3607;
													assign node3607 = (inp[12]) ? 8'b00001011 : 8'b00011010;
													assign node3610 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node3613 = (inp[7]) ? node3621 : node3614;
													assign node3614 = (inp[6]) ? node3618 : node3615;
														assign node3615 = (inp[12]) ? 8'b00001011 : 8'b00011010;
														assign node3618 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node3621 = (inp[12]) ? 8'b00000010 : node3622;
														assign node3622 = (inp[6]) ? 8'b10100101 : 8'b11110111;
											assign node3626 = (inp[3]) ? node3634 : node3627;
												assign node3627 = (inp[12]) ? node3631 : node3628;
													assign node3628 = (inp[6]) ? 8'b10101000 : 8'b10111000;
													assign node3631 = (inp[6]) ? 8'b10111000 : 8'b10101001;
												assign node3634 = (inp[7]) ? node3636 : 8'b10101000;
													assign node3636 = (inp[6]) ? node3638 : 8'b10100000;
														assign node3638 = (inp[12]) ? 8'b10010101 : 8'b10000101;
										assign node3641 = (inp[9]) ? node3657 : node3642;
											assign node3642 = (inp[7]) ? node3648 : node3643;
												assign node3643 = (inp[6]) ? node3645 : 8'b10101101;
													assign node3645 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node3648 = (inp[3]) ? node3654 : node3649;
													assign node3649 = (inp[12]) ? node3651 : 8'b10111100;
														assign node3651 = (inp[6]) ? 8'b10111100 : 8'b10101101;
													assign node3654 = (inp[6]) ? 8'b10100001 : 8'b10110001;
											assign node3657 = (inp[7]) ? node3665 : node3658;
												assign node3658 = (inp[3]) ? node3660 : 8'b10011100;
													assign node3660 = (inp[12]) ? 8'b10001101 : node3661;
														assign node3661 = (inp[6]) ? 8'b10001100 : 8'b10011100;
												assign node3665 = (inp[3]) ? node3669 : node3666;
													assign node3666 = (inp[6]) ? 8'b10001100 : 8'b10001101;
													assign node3669 = (inp[6]) ? node3673 : node3670;
														assign node3670 = (inp[12]) ? 8'b10000100 : 8'b10010001;
														assign node3673 = (inp[12]) ? 8'b10010001 : 8'b10000001;
									assign node3676 = (inp[12]) ? node3682 : node3677;
										assign node3677 = (inp[7]) ? node3679 : 8'b10001100;
											assign node3679 = (inp[3]) ? 8'b10000001 : 8'b10001100;
										assign node3682 = (inp[3]) ? node3684 : 8'b10011100;
											assign node3684 = (inp[7]) ? 8'b10010001 : 8'b10011100;
								assign node3687 = (inp[0]) ? node3739 : node3688;
									assign node3688 = (inp[9]) ? node3716 : node3689;
										assign node3689 = (inp[10]) ? node3701 : node3690;
											assign node3690 = (inp[6]) ? node3694 : node3691;
												assign node3691 = (inp[3]) ? 8'b10100101 : 8'b00000010;
												assign node3694 = (inp[3]) ? node3698 : node3695;
													assign node3695 = (inp[12]) ? 8'b11110101 : 8'b10100101;
													assign node3698 = (inp[12]) ? 8'b10110100 : 8'b10100100;
											assign node3701 = (inp[3]) ? node3709 : node3702;
												assign node3702 = (inp[6]) ? node3706 : node3703;
													assign node3703 = (inp[7]) ? 8'b10100100 : 8'b10110001;
													assign node3706 = (inp[12]) ? 8'b10110001 : 8'b10100001;
												assign node3709 = (inp[6]) ? node3713 : node3710;
													assign node3710 = (inp[12]) ? 8'b10100001 : 8'b10110000;
													assign node3713 = (inp[12]) ? 8'b10110000 : 8'b10100000;
										assign node3716 = (inp[10]) ? node3728 : node3717;
											assign node3717 = (inp[3]) ? node3723 : node3718;
												assign node3718 = (inp[6]) ? node3720 : 8'b10100000;
													assign node3720 = (inp[12]) ? 8'b10010101 : 8'b10000101;
												assign node3723 = (inp[12]) ? 8'b10000101 : node3724;
													assign node3724 = (inp[6]) ? 8'b10000100 : 8'b10010100;
											assign node3728 = (inp[3]) ? node3734 : node3729;
												assign node3729 = (inp[12]) ? 8'b10000100 : node3730;
													assign node3730 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node3734 = (inp[12]) ? 8'b10010000 : node3735;
													assign node3735 = (inp[6]) ? 8'b10000000 : 8'b10010000;
									assign node3739 = (inp[12]) ? 8'b10010000 : 8'b10000000;
		assign node3742 = (inp[7]) ? node6358 : node3743;
			assign node3743 = (inp[13]) ? node5049 : node3744;
				assign node3744 = (inp[9]) ? node4428 : node3745;
					assign node3745 = (inp[8]) ? node4071 : node3746;
						assign node3746 = (inp[10]) ? node3910 : node3747;
							assign node3747 = (inp[1]) ? node3819 : node3748;
								assign node3748 = (inp[3]) ? node3786 : node3749;
									assign node3749 = (inp[2]) ? node3761 : node3750;
										assign node3750 = (inp[6]) ? node3756 : node3751;
											assign node3751 = (inp[12]) ? 8'b00000010 : node3752;
												assign node3752 = (inp[11]) ? 8'b11110111 : 8'b10000010;
											assign node3756 = (inp[12]) ? 8'b00011010 : node3757;
												assign node3757 = (inp[11]) ? 8'b00001010 : 8'b00011010;
										assign node3761 = (inp[11]) ? node3771 : node3762;
											assign node3762 = (inp[5]) ? node3766 : node3763;
												assign node3763 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node3766 = (inp[0]) ? 8'b10010000 : node3767;
													assign node3767 = (inp[6]) ? 8'b10010000 : 8'b10000010;
											assign node3771 = (inp[12]) ? node3783 : node3772;
												assign node3772 = (inp[0]) ? node3778 : node3773;
													assign node3773 = (inp[6]) ? node3775 : 8'b11110111;
														assign node3775 = (inp[5]) ? 8'b10100101 : 8'b11110111;
													assign node3778 = (inp[6]) ? node3780 : 8'b10100101;
														assign node3780 = (inp[5]) ? 8'b10100101 : 8'b11110111;
												assign node3783 = (inp[5]) ? 8'b11110101 : 8'b00000010;
									assign node3786 = (inp[11]) ? node3798 : node3787;
										assign node3787 = (inp[6]) ? node3793 : node3788;
											assign node3788 = (inp[2]) ? node3790 : 8'b00001011;
												assign node3790 = (inp[0]) ? 8'b00011011 : 8'b00001011;
											assign node3793 = (inp[5]) ? 8'b00011011 : node3794;
												assign node3794 = (inp[2]) ? 8'b00001011 : 8'b00011011;
										assign node3798 = (inp[2]) ? node3806 : node3799;
											assign node3799 = (inp[6]) ? node3803 : node3800;
												assign node3800 = (inp[12]) ? 8'b00001011 : 8'b00011010;
												assign node3803 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node3806 = (inp[12]) ? node3812 : node3807;
												assign node3807 = (inp[5]) ? node3809 : 8'b00011010;
													assign node3809 = (inp[0]) ? 8'b00001010 : 8'b00011010;
												assign node3812 = (inp[0]) ? 8'b00011010 : node3813;
													assign node3813 = (inp[6]) ? node3815 : 8'b00001011;
														assign node3815 = (inp[5]) ? 8'b00011010 : 8'b00001011;
								assign node3819 = (inp[11]) ? node3863 : node3820;
									assign node3820 = (inp[5]) ? node3842 : node3821;
										assign node3821 = (inp[0]) ? node3827 : node3822;
											assign node3822 = (inp[12]) ? node3824 : 8'b10000010;
												assign node3824 = (inp[2]) ? 8'b00000010 : 8'b00011010;
											assign node3827 = (inp[3]) ? node3835 : node3828;
												assign node3828 = (inp[6]) ? node3832 : node3829;
													assign node3829 = (inp[2]) ? 8'b10010001 : 8'b10000001;
													assign node3832 = (inp[2]) ? 8'b10000001 : 8'b10011001;
												assign node3835 = (inp[12]) ? 8'b00000010 : node3836;
													assign node3836 = (inp[6]) ? 8'b00011010 : node3837;
														assign node3837 = (inp[2]) ? 8'b10010000 : 8'b10000010;
										assign node3842 = (inp[6]) ? node3852 : node3843;
											assign node3843 = (inp[0]) ? node3849 : node3844;
												assign node3844 = (inp[3]) ? 8'b10000001 : node3845;
													assign node3845 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node3849 = (inp[2]) ? 8'b10010001 : 8'b10000001;
											assign node3852 = (inp[2]) ? node3858 : node3853;
												assign node3853 = (inp[3]) ? 8'b10011001 : node3854;
													assign node3854 = (inp[0]) ? 8'b10011001 : 8'b00011010;
												assign node3858 = (inp[0]) ? 8'b10010001 : node3859;
													assign node3859 = (inp[3]) ? 8'b10010001 : 8'b10010000;
									assign node3863 = (inp[0]) ? node3885 : node3864;
										assign node3864 = (inp[12]) ? node3874 : node3865;
											assign node3865 = (inp[5]) ? node3867 : 8'b11110111;
												assign node3867 = (inp[6]) ? node3871 : node3868;
													assign node3868 = (inp[3]) ? 8'b10110100 : 8'b11110111;
													assign node3871 = (inp[3]) ? 8'b10101101 : 8'b10100101;
											assign node3874 = (inp[3]) ? node3878 : node3875;
												assign node3875 = (inp[6]) ? 8'b00011010 : 8'b00000010;
												assign node3878 = (inp[5]) ? node3880 : 8'b00000010;
													assign node3880 = (inp[6]) ? node3882 : 8'b10100101;
														assign node3882 = (inp[2]) ? 8'b10110100 : 8'b11111101;
										assign node3885 = (inp[6]) ? node3901 : node3886;
											assign node3886 = (inp[5]) ? node3894 : node3887;
												assign node3887 = (inp[2]) ? node3891 : node3888;
													assign node3888 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node3891 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node3894 = (inp[2]) ? node3898 : node3895;
													assign node3895 = (inp[12]) ? 8'b10100101 : 8'b10110100;
													assign node3898 = (inp[12]) ? 8'b10110100 : 8'b10100100;
											assign node3901 = (inp[5]) ? node3903 : 8'b00001010;
												assign node3903 = (inp[2]) ? node3907 : node3904;
													assign node3904 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node3907 = (inp[12]) ? 8'b10110100 : 8'b10100100;
							assign node3910 = (inp[11]) ? node3972 : node3911;
								assign node3911 = (inp[6]) ? node3943 : node3912;
									assign node3912 = (inp[0]) ? node3920 : node3913;
										assign node3913 = (inp[3]) ? node3915 : 8'b00001110;
											assign node3915 = (inp[5]) ? 8'b00001111 : node3916;
												assign node3916 = (inp[1]) ? 8'b00001110 : 8'b00001111;
										assign node3920 = (inp[2]) ? node3934 : node3921;
											assign node3921 = (inp[5]) ? node3929 : node3922;
												assign node3922 = (inp[1]) ? node3926 : node3923;
													assign node3923 = (inp[3]) ? 8'b00001111 : 8'b00001110;
													assign node3926 = (inp[3]) ? 8'b00001110 : 8'b00001111;
												assign node3929 = (inp[3]) ? 8'b00001111 : node3930;
													assign node3930 = (inp[1]) ? 8'b00001111 : 8'b00001110;
											assign node3934 = (inp[1]) ? node3938 : node3935;
												assign node3935 = (inp[3]) ? 8'b00011111 : 8'b00011110;
												assign node3938 = (inp[3]) ? node3940 : 8'b00011111;
													assign node3940 = (inp[5]) ? 8'b00011111 : 8'b00011110;
									assign node3943 = (inp[5]) ? node3965 : node3944;
										assign node3944 = (inp[2]) ? node3956 : node3945;
											assign node3945 = (inp[0]) ? node3947 : 8'b00011110;
												assign node3947 = (inp[12]) ? node3949 : 8'b00011110;
													assign node3949 = (inp[1]) ? node3953 : node3950;
														assign node3950 = (inp[3]) ? 8'b00011111 : 8'b00011110;
														assign node3953 = (inp[3]) ? 8'b00011110 : 8'b00011111;
											assign node3956 = (inp[3]) ? node3962 : node3957;
												assign node3957 = (inp[0]) ? node3959 : 8'b00001110;
													assign node3959 = (inp[1]) ? 8'b00001111 : 8'b00001110;
												assign node3962 = (inp[1]) ? 8'b00001110 : 8'b00001111;
										assign node3965 = (inp[3]) ? 8'b00011111 : node3966;
											assign node3966 = (inp[1]) ? node3968 : 8'b00011110;
												assign node3968 = (inp[0]) ? 8'b00011111 : 8'b00011110;
								assign node3972 = (inp[1]) ? node4020 : node3973;
									assign node3973 = (inp[3]) ? node3997 : node3974;
										assign node3974 = (inp[12]) ? node3986 : node3975;
											assign node3975 = (inp[6]) ? node3981 : node3976;
												assign node3976 = (inp[2]) ? node3978 : 8'b00011011;
													assign node3978 = (inp[0]) ? 8'b00001011 : 8'b00011011;
												assign node3981 = (inp[2]) ? node3983 : 8'b00001110;
													assign node3983 = (inp[5]) ? 8'b00001011 : 8'b00011011;
											assign node3986 = (inp[6]) ? node3992 : node3987;
												assign node3987 = (inp[0]) ? node3989 : 8'b00001110;
													assign node3989 = (inp[2]) ? 8'b00011011 : 8'b00001110;
												assign node3992 = (inp[2]) ? node3994 : 8'b00011110;
													assign node3994 = (inp[5]) ? 8'b00011011 : 8'b00001110;
										assign node3997 = (inp[2]) ? node4005 : node3998;
											assign node3998 = (inp[6]) ? node4002 : node3999;
												assign node3999 = (inp[12]) ? 8'b00001111 : 8'b00011110;
												assign node4002 = (inp[12]) ? 8'b00011111 : 8'b00001111;
											assign node4005 = (inp[5]) ? node4013 : node4006;
												assign node4006 = (inp[0]) ? node4008 : 8'b00001111;
													assign node4008 = (inp[6]) ? node4010 : 8'b00011110;
														assign node4010 = (inp[12]) ? 8'b00001111 : 8'b00011110;
												assign node4013 = (inp[12]) ? 8'b00011110 : node4014;
													assign node4014 = (inp[6]) ? 8'b00001110 : node4015;
														assign node4015 = (inp[0]) ? 8'b00001110 : 8'b00011110;
									assign node4020 = (inp[12]) ? node4044 : node4021;
										assign node4021 = (inp[6]) ? node4031 : node4022;
											assign node4022 = (inp[0]) ? node4028 : node4023;
												assign node4023 = (inp[3]) ? node4025 : 8'b00011011;
													assign node4025 = (inp[5]) ? 8'b00011010 : 8'b00011011;
												assign node4028 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node4031 = (inp[2]) ? node4039 : node4032;
												assign node4032 = (inp[0]) ? node4034 : 8'b00001110;
													assign node4034 = (inp[5]) ? 8'b00001011 : node4035;
														assign node4035 = (inp[3]) ? 8'b00001110 : 8'b00001011;
												assign node4039 = (inp[0]) ? 8'b00001010 : node4040;
													assign node4040 = (inp[3]) ? 8'b00011011 : 8'b00001011;
										assign node4044 = (inp[6]) ? node4056 : node4045;
											assign node4045 = (inp[0]) ? node4047 : 8'b00001110;
												assign node4047 = (inp[2]) ? node4053 : node4048;
													assign node4048 = (inp[5]) ? 8'b00001011 : node4049;
														assign node4049 = (inp[3]) ? 8'b00001110 : 8'b00001011;
													assign node4053 = (inp[5]) ? 8'b00011010 : 8'b00011011;
											assign node4056 = (inp[5]) ? node4062 : node4057;
												assign node4057 = (inp[3]) ? node4059 : 8'b00011011;
													assign node4059 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node4062 = (inp[0]) ? 8'b00011011 : node4063;
													assign node4063 = (inp[3]) ? node4067 : node4064;
														assign node4064 = (inp[2]) ? 8'b00011011 : 8'b00011110;
														assign node4067 = (inp[2]) ? 8'b00011010 : 8'b00011011;
						assign node4071 = (inp[0]) ? node4215 : node4072;
							assign node4072 = (inp[5]) ? node4124 : node4073;
								assign node4073 = (inp[12]) ? node4107 : node4074;
									assign node4074 = (inp[11]) ? node4092 : node4075;
										assign node4075 = (inp[6]) ? node4081 : node4076;
											assign node4076 = (inp[3]) ? node4078 : 8'b10000010;
												assign node4078 = (inp[1]) ? 8'b10000010 : 8'b00001011;
											assign node4081 = (inp[2]) ? node4087 : node4082;
												assign node4082 = (inp[1]) ? 8'b00011010 : node4083;
													assign node4083 = (inp[3]) ? 8'b00011011 : 8'b00011010;
												assign node4087 = (inp[1]) ? 8'b10000010 : node4088;
													assign node4088 = (inp[3]) ? 8'b00001011 : 8'b10000010;
										assign node4092 = (inp[1]) ? node4102 : node4093;
											assign node4093 = (inp[6]) ? node4097 : node4094;
												assign node4094 = (inp[10]) ? 8'b11110111 : 8'b00011010;
												assign node4097 = (inp[2]) ? 8'b00011010 : node4098;
													assign node4098 = (inp[3]) ? 8'b00001011 : 8'b00001010;
											assign node4102 = (inp[2]) ? 8'b11110111 : node4103;
												assign node4103 = (inp[6]) ? 8'b00001010 : 8'b11110111;
									assign node4107 = (inp[2]) ? node4119 : node4108;
										assign node4108 = (inp[6]) ? node4114 : node4109;
											assign node4109 = (inp[1]) ? 8'b00000010 : node4110;
												assign node4110 = (inp[3]) ? 8'b00001011 : 8'b00000010;
											assign node4114 = (inp[1]) ? 8'b00011010 : node4115;
												assign node4115 = (inp[3]) ? 8'b00011011 : 8'b00011010;
										assign node4119 = (inp[3]) ? node4121 : 8'b00000010;
											assign node4121 = (inp[1]) ? 8'b00000010 : 8'b00001011;
								assign node4124 = (inp[10]) ? node4168 : node4125;
									assign node4125 = (inp[3]) ? node4145 : node4126;
										assign node4126 = (inp[11]) ? node4134 : node4127;
											assign node4127 = (inp[6]) ? node4131 : node4128;
												assign node4128 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node4131 = (inp[2]) ? 8'b10010000 : 8'b00011010;
											assign node4134 = (inp[12]) ? node4140 : node4135;
												assign node4135 = (inp[6]) ? node4137 : 8'b11110111;
													assign node4137 = (inp[1]) ? 8'b10100101 : 8'b00001010;
												assign node4140 = (inp[6]) ? node4142 : 8'b00000010;
													assign node4142 = (inp[2]) ? 8'b11110101 : 8'b00011010;
										assign node4145 = (inp[1]) ? node4157 : node4146;
											assign node4146 = (inp[11]) ? node4150 : node4147;
												assign node4147 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node4150 = (inp[12]) ? node4154 : node4151;
													assign node4151 = (inp[6]) ? 8'b00001011 : 8'b00011010;
													assign node4154 = (inp[6]) ? 8'b00011010 : 8'b00001011;
											assign node4157 = (inp[11]) ? node4163 : node4158;
												assign node4158 = (inp[12]) ? 8'b10000001 : node4159;
													assign node4159 = (inp[2]) ? 8'b10010001 : 8'b10011001;
												assign node4163 = (inp[6]) ? 8'b11111101 : node4164;
													assign node4164 = (inp[2]) ? 8'b10110100 : 8'b10100101;
									assign node4168 = (inp[11]) ? node4184 : node4169;
										assign node4169 = (inp[6]) ? node4175 : node4170;
											assign node4170 = (inp[3]) ? node4172 : 8'b10000100;
												assign node4172 = (inp[1]) ? 8'b10000101 : 8'b10001101;
											assign node4175 = (inp[3]) ? node4179 : node4176;
												assign node4176 = (inp[2]) ? 8'b10010100 : 8'b10011100;
												assign node4179 = (inp[2]) ? node4181 : 8'b10011101;
													assign node4181 = (inp[1]) ? 8'b10010101 : 8'b10011101;
										assign node4184 = (inp[1]) ? node4198 : node4185;
											assign node4185 = (inp[3]) ? node4193 : node4186;
												assign node4186 = (inp[6]) ? node4190 : node4187;
													assign node4187 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node4190 = (inp[12]) ? 8'b10110001 : 8'b10100001;
												assign node4193 = (inp[6]) ? node4195 : 8'b10101101;
													assign node4195 = (inp[2]) ? 8'b10101100 : 8'b10101101;
											assign node4198 = (inp[3]) ? node4206 : node4199;
												assign node4199 = (inp[12]) ? node4201 : 8'b10110001;
													assign node4201 = (inp[6]) ? node4203 : 8'b10100100;
														assign node4203 = (inp[2]) ? 8'b10110001 : 8'b10111100;
												assign node4206 = (inp[2]) ? node4212 : node4207;
													assign node4207 = (inp[12]) ? node4209 : 8'b10110000;
														assign node4209 = (inp[6]) ? 8'b10111001 : 8'b10100001;
													assign node4212 = (inp[12]) ? 8'b10110000 : 8'b10100000;
							assign node4215 = (inp[11]) ? node4307 : node4216;
								assign node4216 = (inp[5]) ? node4284 : node4217;
									assign node4217 = (inp[10]) ? node4251 : node4218;
										assign node4218 = (inp[1]) ? node4234 : node4219;
											assign node4219 = (inp[3]) ? node4227 : node4220;
												assign node4220 = (inp[6]) ? node4224 : node4221;
													assign node4221 = (inp[2]) ? 8'b10010100 : 8'b10000100;
													assign node4224 = (inp[2]) ? 8'b10000100 : 8'b10011100;
												assign node4227 = (inp[2]) ? node4231 : node4228;
													assign node4228 = (inp[6]) ? 8'b10011101 : 8'b10001101;
													assign node4231 = (inp[6]) ? 8'b10001101 : 8'b10011101;
											assign node4234 = (inp[3]) ? node4240 : node4235;
												assign node4235 = (inp[2]) ? 8'b10000101 : node4236;
													assign node4236 = (inp[6]) ? 8'b10011101 : 8'b10000101;
												assign node4240 = (inp[12]) ? node4246 : node4241;
													assign node4241 = (inp[2]) ? node4243 : 8'b10000100;
														assign node4243 = (inp[6]) ? 8'b10000100 : 8'b10010100;
													assign node4246 = (inp[2]) ? 8'b10000100 : node4247;
														assign node4247 = (inp[6]) ? 8'b10011100 : 8'b10000100;
										assign node4251 = (inp[1]) ? node4267 : node4252;
											assign node4252 = (inp[3]) ? node4260 : node4253;
												assign node4253 = (inp[2]) ? node4257 : node4254;
													assign node4254 = (inp[6]) ? 8'b00011010 : 8'b00000010;
													assign node4257 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node4260 = (inp[6]) ? node4264 : node4261;
													assign node4261 = (inp[2]) ? 8'b00011011 : 8'b00001011;
													assign node4264 = (inp[2]) ? 8'b00001011 : 8'b00011011;
											assign node4267 = (inp[3]) ? node4275 : node4268;
												assign node4268 = (inp[2]) ? node4272 : node4269;
													assign node4269 = (inp[6]) ? 8'b10011001 : 8'b10000001;
													assign node4272 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node4275 = (inp[2]) ? node4281 : node4276;
													assign node4276 = (inp[6]) ? 8'b00011010 : node4277;
														assign node4277 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node4281 = (inp[6]) ? 8'b10000010 : 8'b10010000;
									assign node4284 = (inp[3]) ? node4296 : node4285;
										assign node4285 = (inp[1]) ? node4291 : node4286;
											assign node4286 = (inp[2]) ? 8'b10010100 : node4287;
												assign node4287 = (inp[6]) ? 8'b10011100 : 8'b10000100;
											assign node4291 = (inp[2]) ? 8'b10010101 : node4292;
												assign node4292 = (inp[6]) ? 8'b10011101 : 8'b10000101;
										assign node4296 = (inp[1]) ? node4302 : node4297;
											assign node4297 = (inp[2]) ? 8'b10011101 : node4298;
												assign node4298 = (inp[6]) ? 8'b10011101 : 8'b10001101;
											assign node4302 = (inp[2]) ? 8'b10010101 : node4303;
												assign node4303 = (inp[6]) ? 8'b10011101 : 8'b10000101;
								assign node4307 = (inp[5]) ? node4391 : node4308;
									assign node4308 = (inp[10]) ? node4346 : node4309;
										assign node4309 = (inp[1]) ? node4323 : node4310;
											assign node4310 = (inp[3]) ? node4318 : node4311;
												assign node4311 = (inp[2]) ? node4315 : node4312;
													assign node4312 = (inp[6]) ? 8'b10101100 : 8'b10100100;
													assign node4315 = (inp[12]) ? 8'b10100100 : 8'b10110001;
												assign node4318 = (inp[12]) ? 8'b10111100 : node4319;
													assign node4319 = (inp[2]) ? 8'b10101100 : 8'b10101101;
											assign node4323 = (inp[6]) ? node4337 : node4324;
												assign node4324 = (inp[3]) ? node4330 : node4325;
													assign node4325 = (inp[2]) ? 8'b10110000 : node4326;
														assign node4326 = (inp[12]) ? 8'b10100001 : 8'b10110000;
													assign node4330 = (inp[2]) ? node4334 : node4331;
														assign node4331 = (inp[12]) ? 8'b10100100 : 8'b10110001;
														assign node4334 = (inp[12]) ? 8'b10110001 : 8'b10100001;
												assign node4337 = (inp[3]) ? node4343 : node4338;
													assign node4338 = (inp[2]) ? 8'b10100001 : node4339;
														assign node4339 = (inp[12]) ? 8'b10111001 : 8'b10101001;
													assign node4343 = (inp[12]) ? 8'b10111100 : 8'b10101100;
										assign node4346 = (inp[3]) ? node4370 : node4347;
											assign node4347 = (inp[1]) ? node4361 : node4348;
												assign node4348 = (inp[6]) ? node4354 : node4349;
													assign node4349 = (inp[2]) ? 8'b11110101 : node4350;
														assign node4350 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node4354 = (inp[2]) ? node4358 : node4355;
														assign node4355 = (inp[12]) ? 8'b00011010 : 8'b00001010;
														assign node4358 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node4361 = (inp[12]) ? 8'b10100101 : node4362;
													assign node4362 = (inp[2]) ? node4366 : node4363;
														assign node4363 = (inp[6]) ? 8'b10101101 : 8'b10110100;
														assign node4366 = (inp[6]) ? 8'b10110100 : 8'b10100100;
											assign node4370 = (inp[1]) ? node4384 : node4371;
												assign node4371 = (inp[12]) ? node4377 : node4372;
													assign node4372 = (inp[6]) ? node4374 : 8'b00011010;
														assign node4374 = (inp[2]) ? 8'b00011010 : 8'b00001011;
													assign node4377 = (inp[6]) ? node4381 : node4378;
														assign node4378 = (inp[2]) ? 8'b00011010 : 8'b00001011;
														assign node4381 = (inp[2]) ? 8'b00001011 : 8'b00011011;
												assign node4384 = (inp[12]) ? 8'b00011010 : node4385;
													assign node4385 = (inp[6]) ? node4387 : 8'b11110111;
														assign node4387 = (inp[2]) ? 8'b11110111 : 8'b00001010;
									assign node4391 = (inp[12]) ? node4415 : node4392;
										assign node4392 = (inp[6]) ? node4406 : node4393;
											assign node4393 = (inp[2]) ? node4399 : node4394;
												assign node4394 = (inp[1]) ? 8'b10110000 : node4395;
													assign node4395 = (inp[3]) ? 8'b10111100 : 8'b10110001;
												assign node4399 = (inp[3]) ? node4403 : node4400;
													assign node4400 = (inp[1]) ? 8'b10100000 : 8'b10100001;
													assign node4403 = (inp[1]) ? 8'b10100000 : 8'b10101100;
											assign node4406 = (inp[2]) ? node4410 : node4407;
												assign node4407 = (inp[1]) ? 8'b10101001 : 8'b10101100;
												assign node4410 = (inp[1]) ? 8'b10100000 : node4411;
													assign node4411 = (inp[10]) ? 8'b10100001 : 8'b10101100;
										assign node4415 = (inp[2]) ? node4421 : node4416;
											assign node4416 = (inp[6]) ? 8'b10111001 : node4417;
												assign node4417 = (inp[3]) ? 8'b10101101 : 8'b10100001;
											assign node4421 = (inp[3]) ? node4425 : node4422;
												assign node4422 = (inp[1]) ? 8'b10110000 : 8'b10110001;
												assign node4425 = (inp[1]) ? 8'b10110000 : 8'b10111100;
					assign node4428 = (inp[11]) ? node4644 : node4429;
						assign node4429 = (inp[3]) ? node4553 : node4430;
							assign node4430 = (inp[0]) ? node4454 : node4431;
								assign node4431 = (inp[10]) ? node4439 : node4432;
									assign node4432 = (inp[6]) ? node4434 : 8'b00101010;
										assign node4434 = (inp[5]) ? 8'b00111010 : node4435;
											assign node4435 = (inp[2]) ? 8'b00101010 : 8'b00111010;
									assign node4439 = (inp[6]) ? node4445 : node4440;
										assign node4440 = (inp[5]) ? 8'b00101110 : node4441;
											assign node4441 = (inp[8]) ? 8'b00101010 : 8'b00101110;
										assign node4445 = (inp[5]) ? 8'b00111110 : node4446;
											assign node4446 = (inp[2]) ? node4450 : node4447;
												assign node4447 = (inp[8]) ? 8'b00111010 : 8'b00111110;
												assign node4450 = (inp[8]) ? 8'b00101010 : 8'b00101110;
								assign node4454 = (inp[1]) ? node4500 : node4455;
									assign node4455 = (inp[8]) ? node4479 : node4456;
										assign node4456 = (inp[10]) ? node4466 : node4457;
											assign node4457 = (inp[2]) ? node4461 : node4458;
												assign node4458 = (inp[6]) ? 8'b00111010 : 8'b00101010;
												assign node4461 = (inp[6]) ? node4463 : 8'b00111010;
													assign node4463 = (inp[5]) ? 8'b00111010 : 8'b00101010;
											assign node4466 = (inp[5]) ? node4474 : node4467;
												assign node4467 = (inp[12]) ? node4471 : node4468;
													assign node4468 = (inp[6]) ? 8'b00101110 : 8'b00111110;
													assign node4471 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node4474 = (inp[2]) ? 8'b00111110 : node4475;
													assign node4475 = (inp[6]) ? 8'b00111110 : 8'b00101110;
										assign node4479 = (inp[10]) ? node4493 : node4480;
											assign node4480 = (inp[5]) ? node4488 : node4481;
												assign node4481 = (inp[2]) ? node4485 : node4482;
													assign node4482 = (inp[6]) ? 8'b00111110 : 8'b00101110;
													assign node4485 = (inp[6]) ? 8'b00101110 : 8'b00111110;
												assign node4488 = (inp[2]) ? 8'b00111110 : node4489;
													assign node4489 = (inp[6]) ? 8'b00111110 : 8'b00101110;
											assign node4493 = (inp[5]) ? 8'b00111110 : node4494;
												assign node4494 = (inp[6]) ? node4496 : 8'b00111010;
													assign node4496 = (inp[2]) ? 8'b00101010 : 8'b00111010;
									assign node4500 = (inp[5]) ? node4540 : node4501;
										assign node4501 = (inp[12]) ? node4521 : node4502;
											assign node4502 = (inp[6]) ? node4510 : node4503;
												assign node4503 = (inp[8]) ? node4507 : node4504;
													assign node4504 = (inp[10]) ? 8'b01111111 : 8'b00111011;
													assign node4507 = (inp[10]) ? 8'b00111011 : 8'b01111111;
												assign node4510 = (inp[2]) ? node4516 : node4511;
													assign node4511 = (inp[8]) ? 8'b00111011 : node4512;
														assign node4512 = (inp[10]) ? 8'b01111111 : 8'b00111011;
													assign node4516 = (inp[8]) ? node4518 : 8'b00101011;
														assign node4518 = (inp[10]) ? 8'b00101011 : 8'b00101111;
											assign node4521 = (inp[2]) ? node4531 : node4522;
												assign node4522 = (inp[6]) ? 8'b01111111 : node4523;
													assign node4523 = (inp[10]) ? node4527 : node4524;
														assign node4524 = (inp[8]) ? 8'b00101111 : 8'b00101011;
														assign node4527 = (inp[8]) ? 8'b00101011 : 8'b00101111;
												assign node4531 = (inp[6]) ? 8'b00101011 : node4532;
													assign node4532 = (inp[8]) ? node4536 : node4533;
														assign node4533 = (inp[10]) ? 8'b01111111 : 8'b00111011;
														assign node4536 = (inp[10]) ? 8'b00111011 : 8'b01111111;
										assign node4540 = (inp[6]) ? 8'b01111111 : node4541;
											assign node4541 = (inp[2]) ? node4547 : node4542;
												assign node4542 = (inp[8]) ? 8'b00101111 : node4543;
													assign node4543 = (inp[10]) ? 8'b00101111 : 8'b00101011;
												assign node4547 = (inp[8]) ? 8'b01111111 : node4548;
													assign node4548 = (inp[10]) ? 8'b01111111 : 8'b00111011;
							assign node4553 = (inp[5]) ? node4621 : node4554;
								assign node4554 = (inp[1]) ? node4592 : node4555;
									assign node4555 = (inp[2]) ? node4571 : node4556;
										assign node4556 = (inp[6]) ? node4562 : node4557;
											assign node4557 = (inp[8]) ? 8'b00101011 : node4558;
												assign node4558 = (inp[10]) ? 8'b00101111 : 8'b00101011;
											assign node4562 = (inp[10]) ? node4568 : node4563;
												assign node4563 = (inp[8]) ? node4565 : 8'b00111011;
													assign node4565 = (inp[0]) ? 8'b01111111 : 8'b00111011;
												assign node4568 = (inp[8]) ? 8'b00111011 : 8'b01111111;
										assign node4571 = (inp[6]) ? node4585 : node4572;
											assign node4572 = (inp[0]) ? node4578 : node4573;
												assign node4573 = (inp[8]) ? 8'b00101011 : node4574;
													assign node4574 = (inp[10]) ? 8'b00101111 : 8'b00101011;
												assign node4578 = (inp[8]) ? node4582 : node4579;
													assign node4579 = (inp[10]) ? 8'b01111111 : 8'b00111011;
													assign node4582 = (inp[10]) ? 8'b00111011 : 8'b01111111;
											assign node4585 = (inp[10]) ? node4589 : node4586;
												assign node4586 = (inp[8]) ? 8'b00101111 : 8'b00101011;
												assign node4589 = (inp[8]) ? 8'b00101011 : 8'b00101111;
									assign node4592 = (inp[0]) ? node4608 : node4593;
										assign node4593 = (inp[8]) ? node4603 : node4594;
											assign node4594 = (inp[10]) ? 8'b00101110 : node4595;
												assign node4595 = (inp[12]) ? 8'b00101010 : node4596;
													assign node4596 = (inp[6]) ? node4598 : 8'b00101010;
														assign node4598 = (inp[2]) ? 8'b00101010 : 8'b00111010;
											assign node4603 = (inp[2]) ? 8'b00101010 : node4604;
												assign node4604 = (inp[6]) ? 8'b00111010 : 8'b00101010;
										assign node4608 = (inp[10]) ? node4618 : node4609;
											assign node4609 = (inp[8]) ? node4611 : 8'b00101010;
												assign node4611 = (inp[6]) ? node4615 : node4612;
													assign node4612 = (inp[2]) ? 8'b00111110 : 8'b00101110;
													assign node4615 = (inp[2]) ? 8'b00101110 : 8'b00111110;
											assign node4618 = (inp[8]) ? 8'b00111010 : 8'b00111110;
								assign node4621 = (inp[6]) ? node4637 : node4622;
									assign node4622 = (inp[10]) ? node4632 : node4623;
										assign node4623 = (inp[0]) ? node4625 : 8'b00101011;
											assign node4625 = (inp[2]) ? node4629 : node4626;
												assign node4626 = (inp[8]) ? 8'b00101111 : 8'b00101011;
												assign node4629 = (inp[8]) ? 8'b01111111 : 8'b00111011;
										assign node4632 = (inp[2]) ? node4634 : 8'b00101111;
											assign node4634 = (inp[0]) ? 8'b01111111 : 8'b00101111;
									assign node4637 = (inp[10]) ? 8'b01111111 : node4638;
										assign node4638 = (inp[0]) ? node4640 : 8'b00111011;
											assign node4640 = (inp[8]) ? 8'b01111111 : 8'b00111011;
						assign node4644 = (inp[8]) ? node4842 : node4645;
							assign node4645 = (inp[10]) ? node4737 : node4646;
								assign node4646 = (inp[1]) ? node4688 : node4647;
									assign node4647 = (inp[3]) ? node4665 : node4648;
										assign node4648 = (inp[2]) ? node4656 : node4649;
											assign node4649 = (inp[6]) ? node4653 : node4650;
												assign node4650 = (inp[12]) ? 8'b00101010 : 8'b00011111;
												assign node4653 = (inp[12]) ? 8'b00111010 : 8'b00101010;
											assign node4656 = (inp[0]) ? node4660 : node4657;
												assign node4657 = (inp[6]) ? 8'b00011111 : 8'b00101010;
												assign node4660 = (inp[12]) ? 8'b00011111 : node4661;
													assign node4661 = (inp[5]) ? 8'b00001111 : 8'b00011111;
										assign node4665 = (inp[12]) ? node4677 : node4666;
											assign node4666 = (inp[6]) ? node4672 : node4667;
												assign node4667 = (inp[0]) ? node4669 : 8'b00111010;
													assign node4669 = (inp[2]) ? 8'b00101010 : 8'b00111010;
												assign node4672 = (inp[2]) ? node4674 : 8'b00101011;
													assign node4674 = (inp[5]) ? 8'b00101010 : 8'b00111010;
											assign node4677 = (inp[6]) ? node4683 : node4678;
												assign node4678 = (inp[2]) ? node4680 : 8'b00101011;
													assign node4680 = (inp[0]) ? 8'b00111010 : 8'b00101011;
												assign node4683 = (inp[2]) ? node4685 : 8'b00111011;
													assign node4685 = (inp[5]) ? 8'b00111010 : 8'b00101011;
									assign node4688 = (inp[5]) ? node4716 : node4689;
										assign node4689 = (inp[12]) ? node4705 : node4690;
											assign node4690 = (inp[6]) ? node4698 : node4691;
												assign node4691 = (inp[0]) ? node4693 : 8'b00011111;
													assign node4693 = (inp[3]) ? 8'b00011111 : node4694;
														assign node4694 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node4698 = (inp[2]) ? node4702 : node4699;
													assign node4699 = (inp[0]) ? 8'b00001111 : 8'b00101010;
													assign node4702 = (inp[0]) ? 8'b00011110 : 8'b00011111;
											assign node4705 = (inp[0]) ? node4709 : node4706;
												assign node4706 = (inp[2]) ? 8'b00101010 : 8'b00111010;
												assign node4709 = (inp[3]) ? node4711 : 8'b00001111;
													assign node4711 = (inp[6]) ? node4713 : 8'b00011111;
														assign node4713 = (inp[2]) ? 8'b00101010 : 8'b00111010;
										assign node4716 = (inp[12]) ? node4730 : node4717;
											assign node4717 = (inp[6]) ? node4725 : node4718;
												assign node4718 = (inp[0]) ? node4722 : node4719;
													assign node4719 = (inp[3]) ? 8'b00011110 : 8'b00011111;
													assign node4722 = (inp[2]) ? 8'b00001110 : 8'b00011110;
												assign node4725 = (inp[3]) ? node4727 : 8'b00101010;
													assign node4727 = (inp[2]) ? 8'b00001110 : 8'b00001111;
											assign node4730 = (inp[6]) ? node4732 : 8'b00001111;
												assign node4732 = (inp[2]) ? node4734 : 8'b00011111;
													assign node4734 = (inp[3]) ? 8'b00011110 : 8'b00011111;
								assign node4737 = (inp[1]) ? node4783 : node4738;
									assign node4738 = (inp[3]) ? node4760 : node4739;
										assign node4739 = (inp[2]) ? node4747 : node4740;
											assign node4740 = (inp[12]) ? node4744 : node4741;
												assign node4741 = (inp[6]) ? 8'b00101110 : 8'b00111011;
												assign node4744 = (inp[6]) ? 8'b00111110 : 8'b00101110;
											assign node4747 = (inp[12]) ? node4757 : node4748;
												assign node4748 = (inp[0]) ? node4752 : node4749;
													assign node4749 = (inp[6]) ? 8'b00101011 : 8'b00111011;
													assign node4752 = (inp[6]) ? node4754 : 8'b00101011;
														assign node4754 = (inp[5]) ? 8'b00101011 : 8'b00111011;
												assign node4757 = (inp[5]) ? 8'b00111011 : 8'b00101110;
										assign node4760 = (inp[12]) ? node4772 : node4761;
											assign node4761 = (inp[6]) ? node4767 : node4762;
												assign node4762 = (inp[0]) ? node4764 : 8'b00111110;
													assign node4764 = (inp[2]) ? 8'b00101110 : 8'b00111110;
												assign node4767 = (inp[2]) ? node4769 : 8'b00101111;
													assign node4769 = (inp[5]) ? 8'b00101110 : 8'b00111110;
											assign node4772 = (inp[6]) ? node4778 : node4773;
												assign node4773 = (inp[2]) ? node4775 : 8'b00101111;
													assign node4775 = (inp[0]) ? 8'b00111110 : 8'b00101111;
												assign node4778 = (inp[2]) ? node4780 : 8'b01111111;
													assign node4780 = (inp[5]) ? 8'b00111110 : 8'b00101111;
									assign node4783 = (inp[12]) ? node4807 : node4784;
										assign node4784 = (inp[0]) ? node4790 : node4785;
											assign node4785 = (inp[5]) ? node4787 : 8'b00111011;
												assign node4787 = (inp[3]) ? 8'b00101011 : 8'b00111011;
											assign node4790 = (inp[6]) ? node4802 : node4791;
												assign node4791 = (inp[2]) ? node4797 : node4792;
													assign node4792 = (inp[3]) ? node4794 : 8'b00111010;
														assign node4794 = (inp[5]) ? 8'b00111010 : 8'b00111011;
													assign node4797 = (inp[5]) ? 8'b00101010 : node4798;
														assign node4798 = (inp[3]) ? 8'b00101011 : 8'b00101010;
												assign node4802 = (inp[2]) ? node4804 : 8'b00101011;
													assign node4804 = (inp[3]) ? 8'b00111011 : 8'b00111010;
										assign node4807 = (inp[5]) ? node4825 : node4808;
											assign node4808 = (inp[0]) ? node4814 : node4809;
												assign node4809 = (inp[2]) ? 8'b00101110 : node4810;
													assign node4810 = (inp[6]) ? 8'b00111110 : 8'b00101110;
												assign node4814 = (inp[3]) ? node4822 : node4815;
													assign node4815 = (inp[2]) ? node4819 : node4816;
														assign node4816 = (inp[6]) ? 8'b00111011 : 8'b00101011;
														assign node4819 = (inp[6]) ? 8'b00101011 : 8'b00111010;
													assign node4822 = (inp[2]) ? 8'b00101110 : 8'b00111110;
											assign node4825 = (inp[6]) ? node4835 : node4826;
												assign node4826 = (inp[3]) ? node4830 : node4827;
													assign node4827 = (inp[0]) ? 8'b00111010 : 8'b00101110;
													assign node4830 = (inp[2]) ? node4832 : 8'b00101011;
														assign node4832 = (inp[0]) ? 8'b00111010 : 8'b00101011;
												assign node4835 = (inp[2]) ? node4837 : 8'b00111011;
													assign node4837 = (inp[0]) ? 8'b00111010 : node4838;
														assign node4838 = (inp[3]) ? 8'b00111010 : 8'b00111011;
							assign node4842 = (inp[0]) ? node4932 : node4843;
								assign node4843 = (inp[12]) ? node4885 : node4844;
									assign node4844 = (inp[6]) ? node4862 : node4845;
										assign node4845 = (inp[3]) ? node4851 : node4846;
											assign node4846 = (inp[5]) ? node4848 : 8'b00011111;
												assign node4848 = (inp[10]) ? 8'b00011011 : 8'b00011111;
											assign node4851 = (inp[1]) ? node4857 : node4852;
												assign node4852 = (inp[10]) ? node4854 : 8'b00111010;
													assign node4854 = (inp[5]) ? 8'b00011110 : 8'b00111010;
												assign node4857 = (inp[5]) ? node4859 : 8'b00011111;
													assign node4859 = (inp[10]) ? 8'b00011010 : 8'b00011110;
										assign node4862 = (inp[2]) ? node4874 : node4863;
											assign node4863 = (inp[3]) ? node4869 : node4864;
												assign node4864 = (inp[10]) ? node4866 : 8'b00101010;
													assign node4866 = (inp[5]) ? 8'b00001110 : 8'b00101010;
												assign node4869 = (inp[10]) ? node4871 : 8'b00101011;
													assign node4871 = (inp[5]) ? 8'b00001111 : 8'b00101011;
											assign node4874 = (inp[5]) ? node4880 : node4875;
												assign node4875 = (inp[3]) ? node4877 : 8'b00011111;
													assign node4877 = (inp[1]) ? 8'b00011111 : 8'b00111010;
												assign node4880 = (inp[1]) ? node4882 : 8'b00001011;
													assign node4882 = (inp[10]) ? 8'b00001010 : 8'b00001110;
									assign node4885 = (inp[5]) ? node4899 : node4886;
										assign node4886 = (inp[3]) ? node4892 : node4887;
											assign node4887 = (inp[2]) ? 8'b00101010 : node4888;
												assign node4888 = (inp[6]) ? 8'b00111010 : 8'b00101010;
											assign node4892 = (inp[1]) ? 8'b00101010 : node4893;
												assign node4893 = (inp[2]) ? 8'b00101011 : node4894;
													assign node4894 = (inp[6]) ? 8'b00111011 : 8'b00101011;
										assign node4899 = (inp[6]) ? node4909 : node4900;
											assign node4900 = (inp[3]) ? node4904 : node4901;
												assign node4901 = (inp[10]) ? 8'b00001110 : 8'b00101010;
												assign node4904 = (inp[1]) ? node4906 : 8'b00101011;
													assign node4906 = (inp[10]) ? 8'b00001011 : 8'b00001111;
											assign node4909 = (inp[10]) ? node4923 : node4910;
												assign node4910 = (inp[1]) ? node4918 : node4911;
													assign node4911 = (inp[2]) ? node4915 : node4912;
														assign node4912 = (inp[3]) ? 8'b00111011 : 8'b00111010;
														assign node4915 = (inp[3]) ? 8'b00111010 : 8'b00011111;
													assign node4918 = (inp[3]) ? node4920 : 8'b00011111;
														assign node4920 = (inp[2]) ? 8'b00011110 : 8'b00011111;
												assign node4923 = (inp[2]) ? node4927 : node4924;
													assign node4924 = (inp[3]) ? 8'b00011111 : 8'b00011110;
													assign node4927 = (inp[3]) ? node4929 : 8'b00011011;
														assign node4929 = (inp[1]) ? 8'b00011010 : 8'b00011110;
								assign node4932 = (inp[1]) ? node4996 : node4933;
									assign node4933 = (inp[5]) ? node4977 : node4934;
										assign node4934 = (inp[10]) ? node4952 : node4935;
											assign node4935 = (inp[12]) ? node4943 : node4936;
												assign node4936 = (inp[3]) ? 8'b00011110 : node4937;
													assign node4937 = (inp[2]) ? node4939 : 8'b00011011;
														assign node4939 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node4943 = (inp[6]) ? node4949 : node4944;
													assign node4944 = (inp[2]) ? 8'b00011110 : node4945;
														assign node4945 = (inp[3]) ? 8'b00001111 : 8'b00001110;
													assign node4949 = (inp[3]) ? 8'b00011111 : 8'b00011110;
											assign node4952 = (inp[3]) ? node4966 : node4953;
												assign node4953 = (inp[2]) ? node4961 : node4954;
													assign node4954 = (inp[12]) ? node4958 : node4955;
														assign node4955 = (inp[6]) ? 8'b00101010 : 8'b00011111;
														assign node4958 = (inp[6]) ? 8'b00111010 : 8'b00101010;
													assign node4961 = (inp[6]) ? 8'b00011111 : node4962;
														assign node4962 = (inp[12]) ? 8'b00011111 : 8'b00001111;
												assign node4966 = (inp[2]) ? node4972 : node4967;
													assign node4967 = (inp[6]) ? node4969 : 8'b00101011;
														assign node4969 = (inp[12]) ? 8'b00111011 : 8'b00101011;
													assign node4972 = (inp[6]) ? node4974 : 8'b00111010;
														assign node4974 = (inp[12]) ? 8'b00101011 : 8'b00111010;
										assign node4977 = (inp[3]) ? node4987 : node4978;
											assign node4978 = (inp[2]) ? node4984 : node4979;
												assign node4979 = (inp[10]) ? 8'b00001110 : node4980;
													assign node4980 = (inp[12]) ? 8'b00001110 : 8'b00011011;
												assign node4984 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node4987 = (inp[2]) ? node4993 : node4988;
												assign node4988 = (inp[12]) ? node4990 : 8'b00011110;
													assign node4990 = (inp[6]) ? 8'b00011111 : 8'b00001111;
												assign node4993 = (inp[12]) ? 8'b00011110 : 8'b00001110;
									assign node4996 = (inp[5]) ? node5038 : node4997;
										assign node4997 = (inp[10]) ? node5017 : node4998;
											assign node4998 = (inp[6]) ? node5006 : node4999;
												assign node4999 = (inp[12]) ? node5003 : node5000;
													assign node5000 = (inp[3]) ? 8'b00001011 : 8'b00001010;
													assign node5003 = (inp[3]) ? 8'b00011011 : 8'b00001011;
												assign node5006 = (inp[2]) ? node5012 : node5007;
													assign node5007 = (inp[3]) ? node5009 : 8'b00011011;
														assign node5009 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node5012 = (inp[12]) ? 8'b00001011 : node5013;
														assign node5013 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node5017 = (inp[3]) ? node5029 : node5018;
												assign node5018 = (inp[2]) ? node5024 : node5019;
													assign node5019 = (inp[6]) ? node5021 : 8'b00011110;
														assign node5021 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node5024 = (inp[12]) ? 8'b00011110 : node5025;
														assign node5025 = (inp[6]) ? 8'b00011110 : 8'b00001110;
												assign node5029 = (inp[12]) ? node5033 : node5030;
													assign node5030 = (inp[2]) ? 8'b00001111 : 8'b00011111;
													assign node5033 = (inp[2]) ? node5035 : 8'b00101010;
														assign node5035 = (inp[6]) ? 8'b00101010 : 8'b00011111;
										assign node5038 = (inp[2]) ? node5046 : node5039;
											assign node5039 = (inp[12]) ? node5043 : node5040;
												assign node5040 = (inp[6]) ? 8'b00001011 : 8'b00011010;
												assign node5043 = (inp[6]) ? 8'b00011011 : 8'b00001011;
											assign node5046 = (inp[12]) ? 8'b00011010 : 8'b00001010;
				assign node5049 = (inp[0]) ? node5553 : node5050;
					assign node5050 = (inp[5]) ? node5200 : node5051;
						assign node5051 = (inp[12]) ? node5147 : node5052;
							assign node5052 = (inp[11]) ? node5100 : node5053;
								assign node5053 = (inp[6]) ? node5073 : node5054;
									assign node5054 = (inp[8]) ? node5068 : node5055;
										assign node5055 = (inp[10]) ? node5061 : node5056;
											assign node5056 = (inp[3]) ? node5058 : 8'b10000010;
												assign node5058 = (inp[2]) ? 8'b00001011 : 8'b10000010;
											assign node5061 = (inp[9]) ? 8'b00001110 : node5062;
												assign node5062 = (inp[2]) ? 8'b00001110 : node5063;
													assign node5063 = (inp[1]) ? 8'b00001110 : 8'b00001111;
										assign node5068 = (inp[1]) ? 8'b10000010 : node5069;
											assign node5069 = (inp[3]) ? 8'b00001011 : 8'b10000010;
									assign node5073 = (inp[2]) ? node5087 : node5074;
										assign node5074 = (inp[8]) ? node5082 : node5075;
											assign node5075 = (inp[10]) ? 8'b00011110 : node5076;
												assign node5076 = (inp[1]) ? 8'b00011010 : node5077;
													assign node5077 = (inp[3]) ? 8'b00011011 : 8'b00011010;
											assign node5082 = (inp[1]) ? 8'b00011010 : node5083;
												assign node5083 = (inp[3]) ? 8'b00011011 : 8'b00011010;
										assign node5087 = (inp[3]) ? node5093 : node5088;
											assign node5088 = (inp[10]) ? node5090 : 8'b10000010;
												assign node5090 = (inp[8]) ? 8'b10000010 : 8'b00001110;
											assign node5093 = (inp[1]) ? node5095 : 8'b00001011;
												assign node5095 = (inp[8]) ? 8'b10000010 : node5096;
													assign node5096 = (inp[10]) ? 8'b00001110 : 8'b10000010;
								assign node5100 = (inp[6]) ? node5118 : node5101;
									assign node5101 = (inp[8]) ? node5113 : node5102;
										assign node5102 = (inp[10]) ? node5108 : node5103;
											assign node5103 = (inp[1]) ? 8'b11110111 : node5104;
												assign node5104 = (inp[3]) ? 8'b00011010 : 8'b11110111;
											assign node5108 = (inp[1]) ? 8'b00011011 : node5109;
												assign node5109 = (inp[3]) ? 8'b00011110 : 8'b00011011;
										assign node5113 = (inp[3]) ? node5115 : 8'b11110111;
											assign node5115 = (inp[1]) ? 8'b11110111 : 8'b00011010;
									assign node5118 = (inp[2]) ? node5132 : node5119;
										assign node5119 = (inp[3]) ? node5125 : node5120;
											assign node5120 = (inp[8]) ? 8'b00001010 : node5121;
												assign node5121 = (inp[10]) ? 8'b00001110 : 8'b00001010;
											assign node5125 = (inp[8]) ? node5129 : node5126;
												assign node5126 = (inp[1]) ? 8'b00001110 : 8'b00001111;
												assign node5129 = (inp[1]) ? 8'b00001010 : 8'b00001011;
										assign node5132 = (inp[3]) ? node5138 : node5133;
											assign node5133 = (inp[8]) ? 8'b11110111 : node5134;
												assign node5134 = (inp[10]) ? 8'b00011011 : 8'b11110111;
											assign node5138 = (inp[1]) ? node5144 : node5139;
												assign node5139 = (inp[10]) ? node5141 : 8'b00011010;
													assign node5141 = (inp[8]) ? 8'b00011010 : 8'b00011110;
												assign node5144 = (inp[10]) ? 8'b00011011 : 8'b11110111;
							assign node5147 = (inp[2]) ? node5183 : node5148;
								assign node5148 = (inp[6]) ? node5166 : node5149;
									assign node5149 = (inp[10]) ? node5155 : node5150;
										assign node5150 = (inp[1]) ? 8'b00000010 : node5151;
											assign node5151 = (inp[3]) ? 8'b00001011 : 8'b00000010;
										assign node5155 = (inp[8]) ? node5161 : node5156;
											assign node5156 = (inp[1]) ? 8'b00001110 : node5157;
												assign node5157 = (inp[3]) ? 8'b00001111 : 8'b00001110;
											assign node5161 = (inp[3]) ? node5163 : 8'b00000010;
												assign node5163 = (inp[1]) ? 8'b00000010 : 8'b00001011;
									assign node5166 = (inp[3]) ? node5172 : node5167;
										assign node5167 = (inp[8]) ? 8'b00011010 : node5168;
											assign node5168 = (inp[10]) ? 8'b00011110 : 8'b00011010;
										assign node5172 = (inp[1]) ? node5178 : node5173;
											assign node5173 = (inp[10]) ? node5175 : 8'b00011011;
												assign node5175 = (inp[8]) ? 8'b00011011 : 8'b00011111;
											assign node5178 = (inp[10]) ? node5180 : 8'b00011010;
												assign node5180 = (inp[8]) ? 8'b00011010 : 8'b00011110;
								assign node5183 = (inp[3]) ? node5189 : node5184;
									assign node5184 = (inp[8]) ? 8'b00000010 : node5185;
										assign node5185 = (inp[10]) ? 8'b00001110 : 8'b00000010;
									assign node5189 = (inp[1]) ? node5195 : node5190;
										assign node5190 = (inp[8]) ? 8'b00001011 : node5191;
											assign node5191 = (inp[10]) ? 8'b00001111 : 8'b00001011;
										assign node5195 = (inp[10]) ? node5197 : 8'b00000010;
											assign node5197 = (inp[8]) ? 8'b00000010 : 8'b00001110;
						assign node5200 = (inp[9]) ? node5420 : node5201;
							assign node5201 = (inp[8]) ? node5297 : node5202;
								assign node5202 = (inp[10]) ? node5262 : node5203;
									assign node5203 = (inp[11]) ? node5219 : node5204;
										assign node5204 = (inp[6]) ? node5212 : node5205;
											assign node5205 = (inp[3]) ? node5209 : node5206;
												assign node5206 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node5209 = (inp[1]) ? 8'b10000001 : 8'b00001011;
											assign node5212 = (inp[3]) ? node5216 : node5213;
												assign node5213 = (inp[2]) ? 8'b10010000 : 8'b00011010;
												assign node5216 = (inp[1]) ? 8'b10011001 : 8'b00011011;
										assign node5219 = (inp[1]) ? node5237 : node5220;
											assign node5220 = (inp[3]) ? node5228 : node5221;
												assign node5221 = (inp[6]) ? node5225 : node5222;
													assign node5222 = (inp[12]) ? 8'b00000010 : 8'b11110111;
													assign node5225 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node5228 = (inp[2]) ? node5230 : 8'b00001011;
													assign node5230 = (inp[6]) ? node5234 : node5231;
														assign node5231 = (inp[12]) ? 8'b00001011 : 8'b00011010;
														assign node5234 = (inp[12]) ? 8'b00011010 : 8'b00001010;
											assign node5237 = (inp[2]) ? node5249 : node5238;
												assign node5238 = (inp[3]) ? node5246 : node5239;
													assign node5239 = (inp[6]) ? node5243 : node5240;
														assign node5240 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node5243 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node5246 = (inp[12]) ? 8'b11111101 : 8'b10101101;
												assign node5249 = (inp[3]) ? node5255 : node5250;
													assign node5250 = (inp[6]) ? node5252 : 8'b11110111;
														assign node5252 = (inp[12]) ? 8'b11110101 : 8'b10100101;
													assign node5255 = (inp[6]) ? node5259 : node5256;
														assign node5256 = (inp[12]) ? 8'b10100101 : 8'b10110100;
														assign node5259 = (inp[12]) ? 8'b10110100 : 8'b10100100;
									assign node5262 = (inp[6]) ? node5278 : node5263;
										assign node5263 = (inp[12]) ? node5271 : node5264;
											assign node5264 = (inp[11]) ? node5268 : node5265;
												assign node5265 = (inp[3]) ? 8'b00001111 : 8'b00001110;
												assign node5268 = (inp[3]) ? 8'b00011110 : 8'b00011011;
											assign node5271 = (inp[3]) ? node5273 : 8'b00001110;
												assign node5273 = (inp[11]) ? node5275 : 8'b00001111;
													assign node5275 = (inp[1]) ? 8'b00001011 : 8'b00001111;
										assign node5278 = (inp[11]) ? node5282 : node5279;
											assign node5279 = (inp[3]) ? 8'b00011111 : 8'b00011110;
											assign node5282 = (inp[12]) ? node5290 : node5283;
												assign node5283 = (inp[1]) ? 8'b00001011 : node5284;
													assign node5284 = (inp[3]) ? node5286 : 8'b00001110;
														assign node5286 = (inp[2]) ? 8'b00001110 : 8'b00001111;
												assign node5290 = (inp[2]) ? node5292 : 8'b00011110;
													assign node5292 = (inp[3]) ? node5294 : 8'b00011011;
														assign node5294 = (inp[1]) ? 8'b00011010 : 8'b00011110;
								assign node5297 = (inp[10]) ? node5361 : node5298;
									assign node5298 = (inp[1]) ? node5332 : node5299;
										assign node5299 = (inp[3]) ? node5315 : node5300;
											assign node5300 = (inp[11]) ? node5308 : node5301;
												assign node5301 = (inp[6]) ? node5305 : node5302;
													assign node5302 = (inp[12]) ? 8'b00000010 : 8'b10000010;
													assign node5305 = (inp[2]) ? 8'b10010000 : 8'b00011010;
												assign node5308 = (inp[12]) ? node5312 : node5309;
													assign node5309 = (inp[6]) ? 8'b00001010 : 8'b11110111;
													assign node5312 = (inp[6]) ? 8'b11110101 : 8'b00000010;
											assign node5315 = (inp[2]) ? node5325 : node5316;
												assign node5316 = (inp[11]) ? node5318 : 8'b00001011;
													assign node5318 = (inp[12]) ? node5322 : node5319;
														assign node5319 = (inp[6]) ? 8'b00001011 : 8'b00011010;
														assign node5322 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node5325 = (inp[11]) ? node5327 : 8'b00011011;
													assign node5327 = (inp[6]) ? node5329 : 8'b00011010;
														assign node5329 = (inp[12]) ? 8'b00011010 : 8'b00001010;
										assign node5332 = (inp[11]) ? node5342 : node5333;
											assign node5333 = (inp[3]) ? node5339 : node5334;
												assign node5334 = (inp[6]) ? 8'b00011010 : node5335;
													assign node5335 = (inp[12]) ? 8'b00000010 : 8'b10000010;
												assign node5339 = (inp[2]) ? 8'b10010001 : 8'b10011001;
											assign node5342 = (inp[3]) ? node5350 : node5343;
												assign node5343 = (inp[6]) ? node5345 : 8'b11110111;
													assign node5345 = (inp[2]) ? node5347 : 8'b00001010;
														assign node5347 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node5350 = (inp[2]) ? node5354 : node5351;
													assign node5351 = (inp[6]) ? 8'b10101101 : 8'b10110100;
													assign node5354 = (inp[12]) ? node5358 : node5355;
														assign node5355 = (inp[6]) ? 8'b10100100 : 8'b10110100;
														assign node5358 = (inp[6]) ? 8'b10110100 : 8'b10100101;
									assign node5361 = (inp[11]) ? node5377 : node5362;
										assign node5362 = (inp[3]) ? node5368 : node5363;
											assign node5363 = (inp[6]) ? node5365 : 8'b10000100;
												assign node5365 = (inp[2]) ? 8'b10010100 : 8'b10011100;
											assign node5368 = (inp[6]) ? node5372 : node5369;
												assign node5369 = (inp[1]) ? 8'b10000101 : 8'b10001101;
												assign node5372 = (inp[1]) ? node5374 : 8'b10011101;
													assign node5374 = (inp[2]) ? 8'b10010101 : 8'b10011101;
										assign node5377 = (inp[1]) ? node5399 : node5378;
											assign node5378 = (inp[3]) ? node5388 : node5379;
												assign node5379 = (inp[6]) ? node5383 : node5380;
													assign node5380 = (inp[12]) ? 8'b10100100 : 8'b10110001;
													assign node5383 = (inp[2]) ? 8'b10110001 : node5384;
														assign node5384 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node5388 = (inp[2]) ? node5394 : node5389;
													assign node5389 = (inp[12]) ? node5391 : 8'b10111100;
														assign node5391 = (inp[6]) ? 8'b11111101 : 8'b10101101;
													assign node5394 = (inp[12]) ? 8'b10111100 : node5395;
														assign node5395 = (inp[6]) ? 8'b10101100 : 8'b10111100;
											assign node5399 = (inp[2]) ? node5407 : node5400;
												assign node5400 = (inp[3]) ? node5404 : node5401;
													assign node5401 = (inp[12]) ? 8'b10100100 : 8'b10101100;
													assign node5404 = (inp[6]) ? 8'b10101001 : 8'b10110000;
												assign node5407 = (inp[3]) ? node5415 : node5408;
													assign node5408 = (inp[6]) ? node5412 : node5409;
														assign node5409 = (inp[12]) ? 8'b10100100 : 8'b10110001;
														assign node5412 = (inp[12]) ? 8'b10110001 : 8'b10100001;
													assign node5415 = (inp[6]) ? node5417 : 8'b10100001;
														assign node5417 = (inp[12]) ? 8'b10110000 : 8'b10100000;
							assign node5420 = (inp[6]) ? node5464 : node5421;
								assign node5421 = (inp[3]) ? node5439 : node5422;
									assign node5422 = (inp[11]) ? node5428 : node5423;
										assign node5423 = (inp[10]) ? node5425 : 8'b10100000;
											assign node5425 = (inp[8]) ? 8'b10100100 : 8'b10101100;
										assign node5428 = (inp[12]) ? node5434 : node5429;
											assign node5429 = (inp[10]) ? node5431 : 8'b10010101;
												assign node5431 = (inp[8]) ? 8'b10010001 : 8'b10111001;
											assign node5434 = (inp[10]) ? node5436 : 8'b10100000;
												assign node5436 = (inp[8]) ? 8'b10000100 : 8'b10101100;
									assign node5439 = (inp[1]) ? node5449 : node5440;
										assign node5440 = (inp[10]) ? node5446 : node5441;
											assign node5441 = (inp[12]) ? 8'b10101001 : node5442;
												assign node5442 = (inp[11]) ? 8'b10111000 : 8'b10101001;
											assign node5446 = (inp[11]) ? 8'b10011100 : 8'b10101101;
										assign node5449 = (inp[11]) ? node5455 : node5450;
											assign node5450 = (inp[10]) ? node5452 : 8'b10100001;
												assign node5452 = (inp[8]) ? 8'b10100101 : 8'b10101101;
											assign node5455 = (inp[12]) ? node5459 : node5456;
												assign node5456 = (inp[10]) ? 8'b10111000 : 8'b10010100;
												assign node5459 = (inp[10]) ? node5461 : 8'b10000101;
													assign node5461 = (inp[8]) ? 8'b10000001 : 8'b10101001;
								assign node5464 = (inp[11]) ? node5488 : node5465;
									assign node5465 = (inp[10]) ? node5475 : node5466;
										assign node5466 = (inp[3]) ? node5470 : node5467;
											assign node5467 = (inp[2]) ? 8'b10110000 : 8'b10111000;
											assign node5470 = (inp[1]) ? node5472 : 8'b10111001;
												assign node5472 = (inp[2]) ? 8'b10110001 : 8'b10111001;
										assign node5475 = (inp[3]) ? node5481 : node5476;
											assign node5476 = (inp[8]) ? node5478 : 8'b10111100;
												assign node5478 = (inp[12]) ? 8'b10110100 : 8'b10111100;
											assign node5481 = (inp[1]) ? node5483 : 8'b11111101;
												assign node5483 = (inp[8]) ? node5485 : 8'b11111101;
													assign node5485 = (inp[2]) ? 8'b11110101 : 8'b11111101;
									assign node5488 = (inp[12]) ? node5526 : node5489;
										assign node5489 = (inp[8]) ? node5509 : node5490;
											assign node5490 = (inp[10]) ? node5500 : node5491;
												assign node5491 = (inp[1]) ? 8'b10001101 : node5492;
													assign node5492 = (inp[3]) ? node5496 : node5493;
														assign node5493 = (inp[2]) ? 8'b10000101 : 8'b10101000;
														assign node5496 = (inp[2]) ? 8'b10101000 : 8'b10101001;
												assign node5500 = (inp[2]) ? node5504 : node5501;
													assign node5501 = (inp[3]) ? 8'b10101101 : 8'b10101100;
													assign node5504 = (inp[3]) ? node5506 : 8'b10101001;
														assign node5506 = (inp[1]) ? 8'b10101000 : 8'b10101100;
											assign node5509 = (inp[2]) ? node5519 : node5510;
												assign node5510 = (inp[3]) ? node5514 : node5511;
													assign node5511 = (inp[10]) ? 8'b10001100 : 8'b10101000;
													assign node5514 = (inp[1]) ? 8'b10001101 : node5515;
														assign node5515 = (inp[10]) ? 8'b10001101 : 8'b10101001;
												assign node5519 = (inp[3]) ? node5521 : 8'b10000001;
													assign node5521 = (inp[1]) ? node5523 : 8'b10101000;
														assign node5523 = (inp[10]) ? 8'b10000000 : 8'b10000100;
										assign node5526 = (inp[2]) ? node5540 : node5527;
											assign node5527 = (inp[3]) ? node5533 : node5528;
												assign node5528 = (inp[10]) ? node5530 : 8'b10111000;
													assign node5530 = (inp[8]) ? 8'b10011100 : 8'b10111100;
												assign node5533 = (inp[1]) ? node5537 : node5534;
													assign node5534 = (inp[10]) ? 8'b11111101 : 8'b10111001;
													assign node5537 = (inp[10]) ? 8'b10011001 : 8'b10011101;
											assign node5540 = (inp[3]) ? node5546 : node5541;
												assign node5541 = (inp[10]) ? node5543 : 8'b10010101;
													assign node5543 = (inp[8]) ? 8'b10010001 : 8'b10111001;
												assign node5546 = (inp[10]) ? node5548 : 8'b10010100;
													assign node5548 = (inp[8]) ? 8'b10011100 : node5549;
														assign node5549 = (inp[1]) ? 8'b10111000 : 8'b10111100;
					assign node5553 = (inp[11]) ? node5917 : node5554;
						assign node5554 = (inp[5]) ? node5840 : node5555;
							assign node5555 = (inp[9]) ? node5701 : node5556;
								assign node5556 = (inp[1]) ? node5632 : node5557;
									assign node5557 = (inp[3]) ? node5585 : node5558;
										assign node5558 = (inp[10]) ? node5572 : node5559;
											assign node5559 = (inp[8]) ? node5567 : node5560;
												assign node5560 = (inp[2]) ? node5564 : node5561;
													assign node5561 = (inp[6]) ? 8'b10111000 : 8'b10100000;
													assign node5564 = (inp[6]) ? 8'b10100000 : 8'b10110000;
												assign node5567 = (inp[6]) ? 8'b10111100 : node5568;
													assign node5568 = (inp[2]) ? 8'b10110100 : 8'b10100100;
											assign node5572 = (inp[8]) ? node5580 : node5573;
												assign node5573 = (inp[6]) ? node5577 : node5574;
													assign node5574 = (inp[2]) ? 8'b10111100 : 8'b10101100;
													assign node5577 = (inp[2]) ? 8'b10101100 : 8'b10111100;
												assign node5580 = (inp[6]) ? node5582 : 8'b10100000;
													assign node5582 = (inp[2]) ? 8'b10100000 : 8'b10111000;
										assign node5585 = (inp[12]) ? node5607 : node5586;
											assign node5586 = (inp[6]) ? node5602 : node5587;
												assign node5587 = (inp[2]) ? node5595 : node5588;
													assign node5588 = (inp[10]) ? node5592 : node5589;
														assign node5589 = (inp[8]) ? 8'b10101101 : 8'b10101001;
														assign node5592 = (inp[8]) ? 8'b10101001 : 8'b10101101;
													assign node5595 = (inp[10]) ? node5599 : node5596;
														assign node5596 = (inp[8]) ? 8'b11111101 : 8'b10111001;
														assign node5599 = (inp[8]) ? 8'b10111001 : 8'b11111101;
												assign node5602 = (inp[10]) ? node5604 : 8'b11111101;
													assign node5604 = (inp[8]) ? 8'b10111001 : 8'b11111101;
											assign node5607 = (inp[8]) ? node5619 : node5608;
												assign node5608 = (inp[10]) ? node5612 : node5609;
													assign node5609 = (inp[2]) ? 8'b10101001 : 8'b10111001;
													assign node5612 = (inp[6]) ? node5616 : node5613;
														assign node5613 = (inp[2]) ? 8'b11111101 : 8'b10101101;
														assign node5616 = (inp[2]) ? 8'b10101101 : 8'b11111101;
												assign node5619 = (inp[10]) ? node5627 : node5620;
													assign node5620 = (inp[2]) ? node5624 : node5621;
														assign node5621 = (inp[6]) ? 8'b11111101 : 8'b10101101;
														assign node5624 = (inp[6]) ? 8'b10101101 : 8'b11111101;
													assign node5627 = (inp[2]) ? node5629 : 8'b10101001;
														assign node5629 = (inp[6]) ? 8'b10101001 : 8'b10111001;
									assign node5632 = (inp[3]) ? node5672 : node5633;
										assign node5633 = (inp[6]) ? node5651 : node5634;
											assign node5634 = (inp[2]) ? node5644 : node5635;
												assign node5635 = (inp[12]) ? node5637 : 8'b10100001;
													assign node5637 = (inp[8]) ? node5641 : node5638;
														assign node5638 = (inp[10]) ? 8'b10101101 : 8'b10100001;
														assign node5641 = (inp[10]) ? 8'b10100001 : 8'b10100101;
												assign node5644 = (inp[10]) ? node5648 : node5645;
													assign node5645 = (inp[8]) ? 8'b11110101 : 8'b10110001;
													assign node5648 = (inp[8]) ? 8'b10110001 : 8'b11111101;
											assign node5651 = (inp[2]) ? node5665 : node5652;
												assign node5652 = (inp[12]) ? node5660 : node5653;
													assign node5653 = (inp[10]) ? node5657 : node5654;
														assign node5654 = (inp[8]) ? 8'b11111101 : 8'b10111001;
														assign node5657 = (inp[8]) ? 8'b10111001 : 8'b11111101;
													assign node5660 = (inp[8]) ? node5662 : 8'b10111001;
														assign node5662 = (inp[10]) ? 8'b10111001 : 8'b11111101;
												assign node5665 = (inp[8]) ? node5669 : node5666;
													assign node5666 = (inp[10]) ? 8'b10101101 : 8'b10100001;
													assign node5669 = (inp[10]) ? 8'b10100001 : 8'b10100101;
										assign node5672 = (inp[2]) ? node5688 : node5673;
											assign node5673 = (inp[6]) ? node5681 : node5674;
												assign node5674 = (inp[8]) ? node5678 : node5675;
													assign node5675 = (inp[10]) ? 8'b10101100 : 8'b10100000;
													assign node5678 = (inp[10]) ? 8'b10100000 : 8'b10100100;
												assign node5681 = (inp[10]) ? node5685 : node5682;
													assign node5682 = (inp[8]) ? 8'b10111100 : 8'b10111000;
													assign node5685 = (inp[8]) ? 8'b10111000 : 8'b10111100;
											assign node5688 = (inp[6]) ? node5696 : node5689;
												assign node5689 = (inp[8]) ? node5693 : node5690;
													assign node5690 = (inp[10]) ? 8'b10111100 : 8'b10110000;
													assign node5693 = (inp[10]) ? 8'b10110000 : 8'b10110100;
												assign node5696 = (inp[10]) ? 8'b10100000 : node5697;
													assign node5697 = (inp[8]) ? 8'b10100100 : 8'b10100000;
								assign node5701 = (inp[8]) ? node5775 : node5702;
									assign node5702 = (inp[10]) ? node5742 : node5703;
										assign node5703 = (inp[1]) ? node5727 : node5704;
											assign node5704 = (inp[3]) ? node5718 : node5705;
												assign node5705 = (inp[12]) ? node5711 : node5706;
													assign node5706 = (inp[2]) ? node5708 : 8'b10000010;
														assign node5708 = (inp[6]) ? 8'b10000010 : 8'b10010000;
													assign node5711 = (inp[2]) ? node5715 : node5712;
														assign node5712 = (inp[6]) ? 8'b00011010 : 8'b00000010;
														assign node5715 = (inp[6]) ? 8'b00000010 : 8'b10010000;
												assign node5718 = (inp[12]) ? node5720 : 8'b00001011;
													assign node5720 = (inp[2]) ? node5724 : node5721;
														assign node5721 = (inp[6]) ? 8'b00011011 : 8'b00001011;
														assign node5724 = (inp[6]) ? 8'b00001011 : 8'b00011011;
											assign node5727 = (inp[3]) ? node5733 : node5728;
												assign node5728 = (inp[2]) ? 8'b10000001 : node5729;
													assign node5729 = (inp[6]) ? 8'b10011001 : 8'b10000001;
												assign node5733 = (inp[6]) ? node5737 : node5734;
													assign node5734 = (inp[2]) ? 8'b10010000 : 8'b10000010;
													assign node5737 = (inp[2]) ? node5739 : 8'b00011010;
														assign node5739 = (inp[12]) ? 8'b00000010 : 8'b10000010;
										assign node5742 = (inp[6]) ? node5760 : node5743;
											assign node5743 = (inp[2]) ? node5749 : node5744;
												assign node5744 = (inp[1]) ? 8'b00001111 : node5745;
													assign node5745 = (inp[3]) ? 8'b00001111 : 8'b00001110;
												assign node5749 = (inp[12]) ? node5755 : node5750;
													assign node5750 = (inp[3]) ? 8'b00011110 : node5751;
														assign node5751 = (inp[1]) ? 8'b00011111 : 8'b00011110;
													assign node5755 = (inp[1]) ? 8'b00011111 : node5756;
														assign node5756 = (inp[3]) ? 8'b00011111 : 8'b00011110;
											assign node5760 = (inp[2]) ? node5766 : node5761;
												assign node5761 = (inp[1]) ? 8'b00011110 : node5762;
													assign node5762 = (inp[3]) ? 8'b00011111 : 8'b00011110;
												assign node5766 = (inp[12]) ? node5770 : node5767;
													assign node5767 = (inp[1]) ? 8'b00001110 : 8'b00001111;
													assign node5770 = (inp[1]) ? node5772 : 8'b00001110;
														assign node5772 = (inp[3]) ? 8'b00001110 : 8'b00001111;
									assign node5775 = (inp[10]) ? node5811 : node5776;
										assign node5776 = (inp[3]) ? node5792 : node5777;
											assign node5777 = (inp[1]) ? node5785 : node5778;
												assign node5778 = (inp[6]) ? node5782 : node5779;
													assign node5779 = (inp[2]) ? 8'b10010100 : 8'b10000100;
													assign node5782 = (inp[2]) ? 8'b10000100 : 8'b10011100;
												assign node5785 = (inp[6]) ? node5789 : node5786;
													assign node5786 = (inp[2]) ? 8'b10010101 : 8'b10000101;
													assign node5789 = (inp[2]) ? 8'b10000101 : 8'b10011101;
											assign node5792 = (inp[1]) ? node5806 : node5793;
												assign node5793 = (inp[12]) ? node5799 : node5794;
													assign node5794 = (inp[6]) ? node5796 : 8'b10001101;
														assign node5796 = (inp[2]) ? 8'b10001101 : 8'b10011101;
													assign node5799 = (inp[2]) ? node5803 : node5800;
														assign node5800 = (inp[6]) ? 8'b10011101 : 8'b10001101;
														assign node5803 = (inp[6]) ? 8'b10001101 : 8'b10011101;
												assign node5806 = (inp[2]) ? node5808 : 8'b10011100;
													assign node5808 = (inp[6]) ? 8'b10000100 : 8'b10010100;
										assign node5811 = (inp[1]) ? node5825 : node5812;
											assign node5812 = (inp[3]) ? node5820 : node5813;
												assign node5813 = (inp[2]) ? node5817 : node5814;
													assign node5814 = (inp[6]) ? 8'b00011010 : 8'b00000010;
													assign node5817 = (inp[6]) ? 8'b10000010 : 8'b10010000;
												assign node5820 = (inp[2]) ? node5822 : 8'b00001011;
													assign node5822 = (inp[6]) ? 8'b00001011 : 8'b00011011;
											assign node5825 = (inp[3]) ? node5833 : node5826;
												assign node5826 = (inp[2]) ? node5830 : node5827;
													assign node5827 = (inp[6]) ? 8'b10011001 : 8'b10000001;
													assign node5830 = (inp[6]) ? 8'b10000001 : 8'b10010001;
												assign node5833 = (inp[6]) ? node5837 : node5834;
													assign node5834 = (inp[2]) ? 8'b10010000 : 8'b10000010;
													assign node5837 = (inp[2]) ? 8'b00000010 : 8'b00011010;
							assign node5840 = (inp[6]) ? node5888 : node5841;
								assign node5841 = (inp[2]) ? node5869 : node5842;
									assign node5842 = (inp[10]) ? node5856 : node5843;
										assign node5843 = (inp[8]) ? node5851 : node5844;
											assign node5844 = (inp[3]) ? node5848 : node5845;
												assign node5845 = (inp[1]) ? 8'b10100001 : 8'b10100000;
												assign node5848 = (inp[1]) ? 8'b10100001 : 8'b10101001;
											assign node5851 = (inp[1]) ? 8'b10100101 : node5852;
												assign node5852 = (inp[9]) ? 8'b10100100 : 8'b10101101;
										assign node5856 = (inp[8]) ? node5862 : node5857;
											assign node5857 = (inp[3]) ? 8'b10101101 : node5858;
												assign node5858 = (inp[1]) ? 8'b10101101 : 8'b10101100;
											assign node5862 = (inp[3]) ? node5866 : node5863;
												assign node5863 = (inp[1]) ? 8'b10100101 : 8'b10100100;
												assign node5866 = (inp[1]) ? 8'b10100101 : 8'b10101101;
									assign node5869 = (inp[1]) ? node5883 : node5870;
										assign node5870 = (inp[3]) ? node5878 : node5871;
											assign node5871 = (inp[10]) ? node5875 : node5872;
												assign node5872 = (inp[8]) ? 8'b10110100 : 8'b10110000;
												assign node5875 = (inp[8]) ? 8'b10110100 : 8'b10111100;
											assign node5878 = (inp[10]) ? 8'b11111101 : node5879;
												assign node5879 = (inp[8]) ? 8'b11111101 : 8'b10111001;
										assign node5883 = (inp[8]) ? 8'b11110101 : node5884;
											assign node5884 = (inp[10]) ? 8'b11111101 : 8'b10110001;
								assign node5888 = (inp[3]) ? node5902 : node5889;
									assign node5889 = (inp[1]) ? node5895 : node5890;
										assign node5890 = (inp[2]) ? node5892 : 8'b10111100;
											assign node5892 = (inp[8]) ? 8'b10110100 : 8'b10110000;
										assign node5895 = (inp[2]) ? node5897 : 8'b11111101;
											assign node5897 = (inp[8]) ? 8'b11110101 : node5898;
												assign node5898 = (inp[10]) ? 8'b11111101 : 8'b10110001;
									assign node5902 = (inp[10]) ? node5910 : node5903;
										assign node5903 = (inp[8]) ? 8'b11111101 : node5904;
											assign node5904 = (inp[2]) ? node5906 : 8'b10111001;
												assign node5906 = (inp[1]) ? 8'b10110001 : 8'b10111001;
										assign node5910 = (inp[8]) ? node5912 : 8'b11111101;
											assign node5912 = (inp[2]) ? node5914 : 8'b11111101;
												assign node5914 = (inp[1]) ? 8'b11110101 : 8'b11111101;
						assign node5917 = (inp[5]) ? node6255 : node5918;
							assign node5918 = (inp[9]) ? node6074 : node5919;
								assign node5919 = (inp[8]) ? node5997 : node5920;
									assign node5920 = (inp[10]) ? node5958 : node5921;
										assign node5921 = (inp[3]) ? node5937 : node5922;
											assign node5922 = (inp[1]) ? node5930 : node5923;
												assign node5923 = (inp[6]) ? 8'b10111000 : node5924;
													assign node5924 = (inp[12]) ? node5926 : 8'b10010101;
														assign node5926 = (inp[2]) ? 8'b10010101 : 8'b10100000;
												assign node5930 = (inp[12]) ? node5932 : 8'b10010100;
													assign node5932 = (inp[6]) ? node5934 : 8'b10010100;
														assign node5934 = (inp[2]) ? 8'b10000101 : 8'b10011101;
											assign node5937 = (inp[1]) ? node5947 : node5938;
												assign node5938 = (inp[6]) ? 8'b10101001 : node5939;
													assign node5939 = (inp[12]) ? node5943 : node5940;
														assign node5940 = (inp[2]) ? 8'b10101000 : 8'b10111000;
														assign node5943 = (inp[2]) ? 8'b10111000 : 8'b10101001;
												assign node5947 = (inp[6]) ? node5951 : node5948;
													assign node5948 = (inp[2]) ? 8'b10000101 : 8'b10010101;
													assign node5951 = (inp[2]) ? node5955 : node5952;
														assign node5952 = (inp[12]) ? 8'b10111000 : 8'b10101000;
														assign node5955 = (inp[12]) ? 8'b10100000 : 8'b10010101;
										assign node5958 = (inp[3]) ? node5974 : node5959;
											assign node5959 = (inp[12]) ? node5963 : node5960;
												assign node5960 = (inp[1]) ? 8'b10111000 : 8'b10111001;
												assign node5963 = (inp[1]) ? node5967 : node5964;
													assign node5964 = (inp[2]) ? 8'b10101100 : 8'b10111100;
													assign node5967 = (inp[6]) ? node5971 : node5968;
														assign node5968 = (inp[2]) ? 8'b10111000 : 8'b10101001;
														assign node5971 = (inp[2]) ? 8'b10101001 : 8'b10111001;
											assign node5974 = (inp[1]) ? node5988 : node5975;
												assign node5975 = (inp[2]) ? node5983 : node5976;
													assign node5976 = (inp[6]) ? node5980 : node5977;
														assign node5977 = (inp[12]) ? 8'b10101101 : 8'b10111100;
														assign node5980 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node5983 = (inp[6]) ? 8'b10111100 : node5984;
														assign node5984 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node5988 = (inp[2]) ? 8'b10101001 : node5989;
													assign node5989 = (inp[12]) ? node5993 : node5990;
														assign node5990 = (inp[6]) ? 8'b10101100 : 8'b10111001;
														assign node5993 = (inp[6]) ? 8'b10111100 : 8'b10101100;
									assign node5997 = (inp[3]) ? node6037 : node5998;
										assign node5998 = (inp[6]) ? node6016 : node5999;
											assign node5999 = (inp[10]) ? node6007 : node6000;
												assign node6000 = (inp[12]) ? 8'b10000100 : node6001;
													assign node6001 = (inp[1]) ? 8'b10010000 : node6002;
														assign node6002 = (inp[2]) ? 8'b10000001 : 8'b10010001;
												assign node6007 = (inp[1]) ? node6009 : 8'b10010101;
													assign node6009 = (inp[2]) ? node6013 : node6010;
														assign node6010 = (inp[12]) ? 8'b10000101 : 8'b10010100;
														assign node6013 = (inp[12]) ? 8'b10010100 : 8'b10000100;
											assign node6016 = (inp[2]) ? node6026 : node6017;
												assign node6017 = (inp[12]) ? node6023 : node6018;
													assign node6018 = (inp[1]) ? 8'b10001101 : node6019;
														assign node6019 = (inp[10]) ? 8'b10101000 : 8'b10001100;
													assign node6023 = (inp[1]) ? 8'b10011101 : 8'b10011100;
												assign node6026 = (inp[12]) ? node6030 : node6027;
													assign node6027 = (inp[1]) ? 8'b10010100 : 8'b10010101;
													assign node6030 = (inp[1]) ? node6034 : node6031;
														assign node6031 = (inp[10]) ? 8'b10100000 : 8'b10000100;
														assign node6034 = (inp[10]) ? 8'b10000101 : 8'b10000001;
										assign node6037 = (inp[10]) ? node6057 : node6038;
											assign node6038 = (inp[6]) ? node6046 : node6039;
												assign node6039 = (inp[1]) ? 8'b10000100 : node6040;
													assign node6040 = (inp[12]) ? 8'b10011100 : node6041;
														assign node6041 = (inp[2]) ? 8'b10001100 : 8'b10011100;
												assign node6046 = (inp[1]) ? node6052 : node6047;
													assign node6047 = (inp[2]) ? 8'b10001101 : node6048;
														assign node6048 = (inp[12]) ? 8'b10011101 : 8'b10001101;
													assign node6052 = (inp[2]) ? 8'b10010001 : node6053;
														assign node6053 = (inp[12]) ? 8'b10011100 : 8'b10001100;
											assign node6057 = (inp[1]) ? node6067 : node6058;
												assign node6058 = (inp[6]) ? node6062 : node6059;
													assign node6059 = (inp[2]) ? 8'b10101000 : 8'b10101001;
													assign node6062 = (inp[12]) ? node6064 : 8'b10101001;
														assign node6064 = (inp[2]) ? 8'b10101001 : 8'b10111001;
												assign node6067 = (inp[2]) ? node6071 : node6068;
													assign node6068 = (inp[12]) ? 8'b10111000 : 8'b10101000;
													assign node6071 = (inp[12]) ? 8'b10100000 : 8'b10010101;
								assign node6074 = (inp[8]) ? node6162 : node6075;
									assign node6075 = (inp[10]) ? node6119 : node6076;
										assign node6076 = (inp[1]) ? node6096 : node6077;
											assign node6077 = (inp[3]) ? node6087 : node6078;
												assign node6078 = (inp[6]) ? node6082 : node6079;
													assign node6079 = (inp[12]) ? 8'b11110101 : 8'b11110111;
													assign node6082 = (inp[2]) ? 8'b00000010 : node6083;
														assign node6083 = (inp[12]) ? 8'b00011010 : 8'b00001010;
												assign node6087 = (inp[6]) ? node6093 : node6088;
													assign node6088 = (inp[12]) ? 8'b00011010 : node6089;
														assign node6089 = (inp[2]) ? 8'b00001010 : 8'b00011010;
													assign node6093 = (inp[12]) ? 8'b00011011 : 8'b00001011;
											assign node6096 = (inp[3]) ? node6106 : node6097;
												assign node6097 = (inp[6]) ? node6103 : node6098;
													assign node6098 = (inp[12]) ? node6100 : 8'b10110100;
														assign node6100 = (inp[2]) ? 8'b10110100 : 8'b10100101;
													assign node6103 = (inp[2]) ? 8'b10100101 : 8'b11111101;
												assign node6106 = (inp[2]) ? node6114 : node6107;
													assign node6107 = (inp[6]) ? node6111 : node6108;
														assign node6108 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node6111 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node6114 = (inp[6]) ? node6116 : 8'b11110101;
														assign node6116 = (inp[12]) ? 8'b00000010 : 8'b11110111;
										assign node6119 = (inp[1]) ? node6143 : node6120;
											assign node6120 = (inp[3]) ? node6132 : node6121;
												assign node6121 = (inp[2]) ? node6129 : node6122;
													assign node6122 = (inp[6]) ? node6126 : node6123;
														assign node6123 = (inp[12]) ? 8'b00001110 : 8'b00011011;
														assign node6126 = (inp[12]) ? 8'b00011110 : 8'b00001110;
													assign node6129 = (inp[6]) ? 8'b00011011 : 8'b00001011;
												assign node6132 = (inp[2]) ? node6138 : node6133;
													assign node6133 = (inp[6]) ? node6135 : 8'b00001111;
														assign node6135 = (inp[12]) ? 8'b00011111 : 8'b00001111;
													assign node6138 = (inp[6]) ? 8'b00011110 : node6139;
														assign node6139 = (inp[12]) ? 8'b00011110 : 8'b00001110;
											assign node6143 = (inp[12]) ? node6153 : node6144;
												assign node6144 = (inp[6]) ? node6150 : node6145;
													assign node6145 = (inp[2]) ? node6147 : 8'b00011010;
														assign node6147 = (inp[3]) ? 8'b00001011 : 8'b00001010;
													assign node6150 = (inp[3]) ? 8'b00001110 : 8'b00001011;
												assign node6153 = (inp[3]) ? 8'b00011011 : node6154;
													assign node6154 = (inp[6]) ? node6158 : node6155;
														assign node6155 = (inp[2]) ? 8'b00011010 : 8'b00001011;
														assign node6158 = (inp[2]) ? 8'b00001011 : 8'b00011011;
									assign node6162 = (inp[10]) ? node6210 : node6163;
										assign node6163 = (inp[1]) ? node6185 : node6164;
											assign node6164 = (inp[3]) ? node6176 : node6165;
												assign node6165 = (inp[6]) ? node6171 : node6166;
													assign node6166 = (inp[2]) ? node6168 : 8'b10100100;
														assign node6168 = (inp[12]) ? 8'b10110001 : 8'b10100001;
													assign node6171 = (inp[2]) ? 8'b10100100 : node6172;
														assign node6172 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node6176 = (inp[6]) ? node6178 : 8'b10111100;
													assign node6178 = (inp[2]) ? node6182 : node6179;
														assign node6179 = (inp[12]) ? 8'b11111101 : 8'b10101101;
														assign node6182 = (inp[12]) ? 8'b10101101 : 8'b10111100;
											assign node6185 = (inp[2]) ? node6197 : node6186;
												assign node6186 = (inp[6]) ? node6190 : node6187;
													assign node6187 = (inp[3]) ? 8'b10110001 : 8'b10100001;
													assign node6190 = (inp[3]) ? node6194 : node6191;
														assign node6191 = (inp[12]) ? 8'b10111001 : 8'b10101001;
														assign node6194 = (inp[12]) ? 8'b10111100 : 8'b10101100;
												assign node6197 = (inp[3]) ? node6203 : node6198;
													assign node6198 = (inp[12]) ? 8'b10100001 : node6199;
														assign node6199 = (inp[6]) ? 8'b10110000 : 8'b10100000;
													assign node6203 = (inp[6]) ? node6207 : node6204;
														assign node6204 = (inp[12]) ? 8'b10110001 : 8'b10100001;
														assign node6207 = (inp[12]) ? 8'b10100100 : 8'b10110001;
										assign node6210 = (inp[3]) ? node6240 : node6211;
											assign node6211 = (inp[1]) ? node6227 : node6212;
												assign node6212 = (inp[2]) ? node6220 : node6213;
													assign node6213 = (inp[6]) ? node6217 : node6214;
														assign node6214 = (inp[12]) ? 8'b00000010 : 8'b11110111;
														assign node6217 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node6220 = (inp[6]) ? node6224 : node6221;
														assign node6221 = (inp[12]) ? 8'b11110101 : 8'b10100101;
														assign node6224 = (inp[12]) ? 8'b00000010 : 8'b11110111;
												assign node6227 = (inp[2]) ? node6235 : node6228;
													assign node6228 = (inp[6]) ? node6232 : node6229;
														assign node6229 = (inp[12]) ? 8'b10100101 : 8'b10110100;
														assign node6232 = (inp[12]) ? 8'b11111101 : 8'b10101101;
													assign node6235 = (inp[12]) ? 8'b10110100 : node6236;
														assign node6236 = (inp[6]) ? 8'b10110100 : 8'b10100100;
											assign node6240 = (inp[6]) ? node6246 : node6241;
												assign node6241 = (inp[1]) ? node6243 : 8'b00011010;
													assign node6243 = (inp[12]) ? 8'b11110101 : 8'b10100101;
												assign node6246 = (inp[2]) ? node6252 : node6247;
													assign node6247 = (inp[1]) ? node6249 : 8'b00001011;
														assign node6249 = (inp[12]) ? 8'b00011010 : 8'b00001010;
													assign node6252 = (inp[1]) ? 8'b00000010 : 8'b00011010;
							assign node6255 = (inp[8]) ? node6323 : node6256;
								assign node6256 = (inp[10]) ? node6292 : node6257;
									assign node6257 = (inp[1]) ? node6281 : node6258;
										assign node6258 = (inp[3]) ? node6268 : node6259;
											assign node6259 = (inp[2]) ? node6265 : node6260;
												assign node6260 = (inp[12]) ? node6262 : 8'b10010101;
													assign node6262 = (inp[6]) ? 8'b10111000 : 8'b10100000;
												assign node6265 = (inp[12]) ? 8'b10010101 : 8'b10000101;
											assign node6268 = (inp[2]) ? node6278 : node6269;
												assign node6269 = (inp[9]) ? 8'b10111000 : node6270;
													assign node6270 = (inp[12]) ? node6274 : node6271;
														assign node6271 = (inp[6]) ? 8'b10101001 : 8'b10111000;
														assign node6274 = (inp[6]) ? 8'b10111001 : 8'b10101001;
												assign node6278 = (inp[12]) ? 8'b10111000 : 8'b10101000;
										assign node6281 = (inp[2]) ? node6289 : node6282;
											assign node6282 = (inp[6]) ? node6286 : node6283;
												assign node6283 = (inp[12]) ? 8'b10000101 : 8'b10010100;
												assign node6286 = (inp[12]) ? 8'b10011101 : 8'b10001101;
											assign node6289 = (inp[12]) ? 8'b10010100 : 8'b10000100;
									assign node6292 = (inp[1]) ? node6312 : node6293;
										assign node6293 = (inp[12]) ? node6305 : node6294;
											assign node6294 = (inp[3]) ? node6302 : node6295;
												assign node6295 = (inp[6]) ? node6299 : node6296;
													assign node6296 = (inp[9]) ? 8'b10111001 : 8'b10101001;
													assign node6299 = (inp[2]) ? 8'b10101001 : 8'b10101100;
												assign node6302 = (inp[2]) ? 8'b10101100 : 8'b10101101;
											assign node6305 = (inp[3]) ? node6309 : node6306;
												assign node6306 = (inp[2]) ? 8'b10111001 : 8'b10101100;
												assign node6309 = (inp[2]) ? 8'b10111100 : 8'b11111101;
										assign node6312 = (inp[2]) ? node6320 : node6313;
											assign node6313 = (inp[6]) ? node6317 : node6314;
												assign node6314 = (inp[12]) ? 8'b10101001 : 8'b10111000;
												assign node6317 = (inp[12]) ? 8'b10111001 : 8'b10101001;
											assign node6320 = (inp[12]) ? 8'b10111000 : 8'b10101000;
								assign node6323 = (inp[1]) ? node6347 : node6324;
									assign node6324 = (inp[3]) ? node6336 : node6325;
										assign node6325 = (inp[2]) ? node6333 : node6326;
											assign node6326 = (inp[6]) ? node6330 : node6327;
												assign node6327 = (inp[12]) ? 8'b10000100 : 8'b10010001;
												assign node6330 = (inp[12]) ? 8'b10011100 : 8'b10001100;
											assign node6333 = (inp[12]) ? 8'b10010001 : 8'b10000001;
										assign node6336 = (inp[2]) ? node6344 : node6337;
											assign node6337 = (inp[6]) ? node6341 : node6338;
												assign node6338 = (inp[12]) ? 8'b10001101 : 8'b10011100;
												assign node6341 = (inp[12]) ? 8'b10011101 : 8'b10001101;
											assign node6344 = (inp[12]) ? 8'b10011100 : 8'b10001100;
									assign node6347 = (inp[2]) ? node6355 : node6348;
										assign node6348 = (inp[6]) ? node6352 : node6349;
											assign node6349 = (inp[12]) ? 8'b10000001 : 8'b10010000;
											assign node6352 = (inp[12]) ? 8'b10011001 : 8'b10001001;
										assign node6355 = (inp[12]) ? 8'b10010000 : 8'b10000000;
			assign node6358 = (inp[12]) ? node6938 : node6359;
				assign node6359 = (inp[11]) ? node6641 : node6360;
					assign node6360 = (inp[5]) ? node6482 : node6361;
						assign node6361 = (inp[0]) ? node6363 : 8'b10000010;
							assign node6363 = (inp[2]) ? node6413 : node6364;
								assign node6364 = (inp[3]) ? node6396 : node6365;
									assign node6365 = (inp[1]) ? node6381 : node6366;
										assign node6366 = (inp[13]) ? node6372 : node6367;
											assign node6367 = (inp[10]) ? 8'b10000010 : node6368;
												assign node6368 = (inp[8]) ? 8'b10000100 : 8'b10000010;
											assign node6372 = (inp[9]) ? node6378 : node6373;
												assign node6373 = (inp[8]) ? node6375 : 8'b10100000;
													assign node6375 = (inp[10]) ? 8'b10100000 : 8'b10100100;
												assign node6378 = (inp[8]) ? 8'b10000100 : 8'b10000010;
										assign node6381 = (inp[13]) ? node6387 : node6382;
											assign node6382 = (inp[10]) ? 8'b10000001 : node6383;
												assign node6383 = (inp[8]) ? 8'b10000101 : 8'b10000001;
											assign node6387 = (inp[9]) ? node6393 : node6388;
												assign node6388 = (inp[10]) ? 8'b10100001 : node6389;
													assign node6389 = (inp[8]) ? 8'b10100101 : 8'b10100001;
												assign node6393 = (inp[8]) ? 8'b10000101 : 8'b10000001;
									assign node6396 = (inp[9]) ? node6408 : node6397;
										assign node6397 = (inp[13]) ? node6403 : node6398;
											assign node6398 = (inp[8]) ? node6400 : 8'b10000010;
												assign node6400 = (inp[10]) ? 8'b10000010 : 8'b10000100;
											assign node6403 = (inp[10]) ? 8'b10100000 : node6404;
												assign node6404 = (inp[8]) ? 8'b10100100 : 8'b10100000;
										assign node6408 = (inp[10]) ? 8'b10000010 : node6409;
											assign node6409 = (inp[8]) ? 8'b10000100 : 8'b10000010;
								assign node6413 = (inp[6]) ? node6449 : node6414;
									assign node6414 = (inp[9]) ? node6436 : node6415;
										assign node6415 = (inp[13]) ? node6423 : node6416;
											assign node6416 = (inp[3]) ? 8'b10010000 : node6417;
												assign node6417 = (inp[1]) ? 8'b10010001 : node6418;
													assign node6418 = (inp[10]) ? 8'b10010000 : 8'b10010100;
											assign node6423 = (inp[8]) ? node6429 : node6424;
												assign node6424 = (inp[1]) ? node6426 : 8'b10110000;
													assign node6426 = (inp[3]) ? 8'b10110000 : 8'b10110001;
												assign node6429 = (inp[10]) ? node6433 : node6430;
													assign node6430 = (inp[1]) ? 8'b11110101 : 8'b10110100;
													assign node6433 = (inp[3]) ? 8'b10110000 : 8'b10110001;
										assign node6436 = (inp[8]) ? node6442 : node6437;
											assign node6437 = (inp[3]) ? 8'b10010000 : node6438;
												assign node6438 = (inp[1]) ? 8'b10010001 : 8'b10010000;
											assign node6442 = (inp[10]) ? 8'b10010000 : node6443;
												assign node6443 = (inp[3]) ? 8'b10010100 : node6444;
													assign node6444 = (inp[1]) ? 8'b10010101 : 8'b10010100;
									assign node6449 = (inp[1]) ? node6459 : node6450;
										assign node6450 = (inp[9]) ? node6454 : node6451;
											assign node6451 = (inp[13]) ? 8'b10100000 : 8'b10000010;
											assign node6454 = (inp[10]) ? 8'b10000010 : node6455;
												assign node6455 = (inp[8]) ? 8'b10000100 : 8'b10000010;
										assign node6459 = (inp[3]) ? node6469 : node6460;
											assign node6460 = (inp[13]) ? node6466 : node6461;
												assign node6461 = (inp[8]) ? node6463 : 8'b10000001;
													assign node6463 = (inp[10]) ? 8'b10000001 : 8'b10000101;
												assign node6466 = (inp[9]) ? 8'b10000001 : 8'b10100001;
											assign node6469 = (inp[8]) ? node6475 : node6470;
												assign node6470 = (inp[13]) ? node6472 : 8'b10000010;
													assign node6472 = (inp[9]) ? 8'b10000010 : 8'b10100000;
												assign node6475 = (inp[10]) ? 8'b10000010 : node6476;
													assign node6476 = (inp[13]) ? node6478 : 8'b10000100;
														assign node6478 = (inp[9]) ? 8'b10000100 : 8'b10100100;
						assign node6482 = (inp[13]) ? node6546 : node6483;
							assign node6483 = (inp[2]) ? node6507 : node6484;
								assign node6484 = (inp[1]) ? node6492 : node6485;
									assign node6485 = (inp[8]) ? node6487 : 8'b10000010;
										assign node6487 = (inp[10]) ? 8'b10000100 : node6488;
											assign node6488 = (inp[0]) ? 8'b10000100 : 8'b10000010;
									assign node6492 = (inp[8]) ? node6498 : node6493;
										assign node6493 = (inp[0]) ? 8'b10000001 : node6494;
											assign node6494 = (inp[3]) ? 8'b10000001 : 8'b10000010;
										assign node6498 = (inp[0]) ? 8'b10000101 : node6499;
											assign node6499 = (inp[10]) ? node6503 : node6500;
												assign node6500 = (inp[3]) ? 8'b10000001 : 8'b10000010;
												assign node6503 = (inp[3]) ? 8'b10000101 : 8'b10000100;
								assign node6507 = (inp[8]) ? node6523 : node6508;
									assign node6508 = (inp[1]) ? node6514 : node6509;
										assign node6509 = (inp[0]) ? 8'b10010000 : node6510;
											assign node6510 = (inp[6]) ? 8'b10010000 : 8'b10000010;
										assign node6514 = (inp[0]) ? 8'b10010001 : node6515;
											assign node6515 = (inp[3]) ? node6519 : node6516;
												assign node6516 = (inp[6]) ? 8'b10010000 : 8'b10000010;
												assign node6519 = (inp[6]) ? 8'b10010001 : 8'b10000001;
									assign node6523 = (inp[0]) ? node6543 : node6524;
										assign node6524 = (inp[10]) ? node6532 : node6525;
											assign node6525 = (inp[6]) ? 8'b10010000 : node6526;
												assign node6526 = (inp[3]) ? node6528 : 8'b10000010;
													assign node6528 = (inp[1]) ? 8'b10000001 : 8'b10000010;
											assign node6532 = (inp[6]) ? node6538 : node6533;
												assign node6533 = (inp[3]) ? node6535 : 8'b10000100;
													assign node6535 = (inp[1]) ? 8'b10000101 : 8'b10000100;
												assign node6538 = (inp[3]) ? node6540 : 8'b10010100;
													assign node6540 = (inp[1]) ? 8'b10010101 : 8'b10010100;
										assign node6543 = (inp[1]) ? 8'b10010101 : 8'b10010100;
							assign node6546 = (inp[8]) ? node6586 : node6547;
								assign node6547 = (inp[1]) ? node6563 : node6548;
									assign node6548 = (inp[2]) ? node6554 : node6549;
										assign node6549 = (inp[9]) ? 8'b10100000 : node6550;
											assign node6550 = (inp[0]) ? 8'b10100000 : 8'b10000010;
										assign node6554 = (inp[0]) ? 8'b10110000 : node6555;
											assign node6555 = (inp[6]) ? node6559 : node6556;
												assign node6556 = (inp[9]) ? 8'b10100000 : 8'b10000010;
												assign node6559 = (inp[9]) ? 8'b10110000 : 8'b10010000;
									assign node6563 = (inp[0]) ? node6583 : node6564;
										assign node6564 = (inp[9]) ? node6574 : node6565;
											assign node6565 = (inp[3]) ? node6571 : node6566;
												assign node6566 = (inp[2]) ? node6568 : 8'b10000010;
													assign node6568 = (inp[6]) ? 8'b10010000 : 8'b10000010;
												assign node6571 = (inp[2]) ? 8'b10010001 : 8'b10000001;
											assign node6574 = (inp[3]) ? node6580 : node6575;
												assign node6575 = (inp[6]) ? node6577 : 8'b10100000;
													assign node6577 = (inp[2]) ? 8'b10110000 : 8'b10100000;
												assign node6580 = (inp[6]) ? 8'b10110001 : 8'b10100001;
										assign node6583 = (inp[2]) ? 8'b10110001 : 8'b10100001;
								assign node6586 = (inp[1]) ? node6612 : node6587;
									assign node6587 = (inp[0]) ? node6609 : node6588;
										assign node6588 = (inp[10]) ? node6600 : node6589;
											assign node6589 = (inp[9]) ? node6595 : node6590;
												assign node6590 = (inp[3]) ? 8'b10000010 : node6591;
													assign node6591 = (inp[6]) ? 8'b10010000 : 8'b10000010;
												assign node6595 = (inp[2]) ? node6597 : 8'b10100000;
													assign node6597 = (inp[6]) ? 8'b10110000 : 8'b10100000;
											assign node6600 = (inp[9]) ? node6606 : node6601;
												assign node6601 = (inp[2]) ? node6603 : 8'b10000100;
													assign node6603 = (inp[6]) ? 8'b10010100 : 8'b10000100;
												assign node6606 = (inp[6]) ? 8'b10110100 : 8'b10100100;
										assign node6609 = (inp[2]) ? 8'b10110100 : 8'b10100100;
									assign node6612 = (inp[0]) ? node6638 : node6613;
										assign node6613 = (inp[10]) ? node6627 : node6614;
											assign node6614 = (inp[9]) ? node6618 : node6615;
												assign node6615 = (inp[2]) ? 8'b10010001 : 8'b10000001;
												assign node6618 = (inp[3]) ? node6622 : node6619;
													assign node6619 = (inp[6]) ? 8'b10110000 : 8'b10100000;
													assign node6622 = (inp[6]) ? node6624 : 8'b10100001;
														assign node6624 = (inp[2]) ? 8'b10110001 : 8'b10100001;
											assign node6627 = (inp[3]) ? node6633 : node6628;
												assign node6628 = (inp[9]) ? node6630 : 8'b10000100;
													assign node6630 = (inp[6]) ? 8'b10110100 : 8'b10100100;
												assign node6633 = (inp[9]) ? 8'b10100101 : node6634;
													assign node6634 = (inp[6]) ? 8'b10010101 : 8'b10000101;
										assign node6638 = (inp[2]) ? 8'b11110101 : 8'b10100101;
					assign node6641 = (inp[0]) ? node6785 : node6642;
						assign node6642 = (inp[5]) ? node6644 : 8'b11110111;
							assign node6644 = (inp[8]) ? node6700 : node6645;
								assign node6645 = (inp[1]) ? node6663 : node6646;
									assign node6646 = (inp[2]) ? node6652 : node6647;
										assign node6647 = (inp[9]) ? node6649 : 8'b11110111;
											assign node6649 = (inp[13]) ? 8'b10010101 : 8'b11110111;
										assign node6652 = (inp[6]) ? node6658 : node6653;
											assign node6653 = (inp[13]) ? node6655 : 8'b11110111;
												assign node6655 = (inp[9]) ? 8'b10010101 : 8'b11110111;
											assign node6658 = (inp[13]) ? node6660 : 8'b10100101;
												assign node6660 = (inp[9]) ? 8'b10000101 : 8'b10100101;
									assign node6663 = (inp[3]) ? node6681 : node6664;
										assign node6664 = (inp[13]) ? node6670 : node6665;
											assign node6665 = (inp[2]) ? node6667 : 8'b11110111;
												assign node6667 = (inp[6]) ? 8'b10100101 : 8'b11110111;
											assign node6670 = (inp[9]) ? node6676 : node6671;
												assign node6671 = (inp[6]) ? node6673 : 8'b11110111;
													assign node6673 = (inp[2]) ? 8'b10100101 : 8'b11110111;
												assign node6676 = (inp[2]) ? node6678 : 8'b10010101;
													assign node6678 = (inp[6]) ? 8'b10000101 : 8'b10010101;
										assign node6681 = (inp[9]) ? node6687 : node6682;
											assign node6682 = (inp[2]) ? node6684 : 8'b10110100;
												assign node6684 = (inp[6]) ? 8'b10100100 : 8'b10110100;
											assign node6687 = (inp[13]) ? node6695 : node6688;
												assign node6688 = (inp[10]) ? node6690 : 8'b10110100;
													assign node6690 = (inp[2]) ? node6692 : 8'b10110100;
														assign node6692 = (inp[6]) ? 8'b10100100 : 8'b10110100;
												assign node6695 = (inp[6]) ? node6697 : 8'b10010100;
													assign node6697 = (inp[2]) ? 8'b10000100 : 8'b10010100;
								assign node6700 = (inp[10]) ? node6742 : node6701;
									assign node6701 = (inp[9]) ? node6713 : node6702;
										assign node6702 = (inp[6]) ? node6708 : node6703;
											assign node6703 = (inp[1]) ? node6705 : 8'b11110111;
												assign node6705 = (inp[3]) ? 8'b10110100 : 8'b11110111;
											assign node6708 = (inp[2]) ? node6710 : 8'b11110111;
												assign node6710 = (inp[1]) ? 8'b10100100 : 8'b10100101;
										assign node6713 = (inp[13]) ? node6729 : node6714;
											assign node6714 = (inp[3]) ? node6720 : node6715;
												assign node6715 = (inp[6]) ? node6717 : 8'b11110111;
													assign node6717 = (inp[2]) ? 8'b10100101 : 8'b11110111;
												assign node6720 = (inp[1]) ? node6724 : node6721;
													assign node6721 = (inp[6]) ? 8'b10100101 : 8'b11110111;
													assign node6724 = (inp[2]) ? node6726 : 8'b10110100;
														assign node6726 = (inp[6]) ? 8'b10100100 : 8'b10110100;
											assign node6729 = (inp[1]) ? node6735 : node6730;
												assign node6730 = (inp[6]) ? node6732 : 8'b10010101;
													assign node6732 = (inp[2]) ? 8'b10000101 : 8'b10010101;
												assign node6735 = (inp[3]) ? node6737 : 8'b10000101;
													assign node6737 = (inp[6]) ? node6739 : 8'b10010100;
														assign node6739 = (inp[2]) ? 8'b10000100 : 8'b10010100;
									assign node6742 = (inp[1]) ? node6762 : node6743;
										assign node6743 = (inp[6]) ? node6749 : node6744;
											assign node6744 = (inp[13]) ? node6746 : 8'b10110001;
												assign node6746 = (inp[9]) ? 8'b10010001 : 8'b10110001;
											assign node6749 = (inp[2]) ? node6755 : node6750;
												assign node6750 = (inp[9]) ? node6752 : 8'b10110001;
													assign node6752 = (inp[13]) ? 8'b10010001 : 8'b10110001;
												assign node6755 = (inp[3]) ? 8'b10100001 : node6756;
													assign node6756 = (inp[13]) ? node6758 : 8'b10100001;
														assign node6758 = (inp[9]) ? 8'b10000001 : 8'b10100001;
										assign node6762 = (inp[3]) ? node6772 : node6763;
											assign node6763 = (inp[9]) ? node6769 : node6764;
												assign node6764 = (inp[6]) ? node6766 : 8'b10110001;
													assign node6766 = (inp[2]) ? 8'b10100001 : 8'b10110001;
												assign node6769 = (inp[13]) ? 8'b10010001 : 8'b10110001;
											assign node6772 = (inp[2]) ? node6778 : node6773;
												assign node6773 = (inp[9]) ? node6775 : 8'b10110000;
													assign node6775 = (inp[13]) ? 8'b10010000 : 8'b10110000;
												assign node6778 = (inp[6]) ? node6780 : 8'b10110000;
													assign node6780 = (inp[13]) ? node6782 : 8'b10100000;
														assign node6782 = (inp[9]) ? 8'b10000000 : 8'b10100000;
						assign node6785 = (inp[8]) ? node6847 : node6786;
							assign node6786 = (inp[13]) ? node6812 : node6787;
								assign node6787 = (inp[2]) ? node6795 : node6788;
									assign node6788 = (inp[1]) ? node6790 : 8'b11110111;
										assign node6790 = (inp[3]) ? node6792 : 8'b10110100;
											assign node6792 = (inp[5]) ? 8'b10110100 : 8'b11110111;
									assign node6795 = (inp[6]) ? node6803 : node6796;
										assign node6796 = (inp[1]) ? node6798 : 8'b10100101;
											assign node6798 = (inp[5]) ? 8'b10100100 : node6799;
												assign node6799 = (inp[3]) ? 8'b10100101 : 8'b10100100;
										assign node6803 = (inp[5]) ? node6809 : node6804;
											assign node6804 = (inp[3]) ? 8'b11110111 : node6805;
												assign node6805 = (inp[1]) ? 8'b10110100 : 8'b11110111;
											assign node6809 = (inp[1]) ? 8'b10100100 : 8'b10100101;
								assign node6812 = (inp[2]) ? node6830 : node6813;
									assign node6813 = (inp[9]) ? node6821 : node6814;
										assign node6814 = (inp[1]) ? node6816 : 8'b10010101;
											assign node6816 = (inp[3]) ? node6818 : 8'b10010100;
												assign node6818 = (inp[5]) ? 8'b10010100 : 8'b10010101;
										assign node6821 = (inp[5]) ? node6827 : node6822;
											assign node6822 = (inp[1]) ? node6824 : 8'b11110111;
												assign node6824 = (inp[3]) ? 8'b11110111 : 8'b10110100;
											assign node6827 = (inp[1]) ? 8'b10010100 : 8'b10010101;
									assign node6830 = (inp[5]) ? node6844 : node6831;
										assign node6831 = (inp[9]) ? node6841 : node6832;
											assign node6832 = (inp[6]) ? node6836 : node6833;
												assign node6833 = (inp[3]) ? 8'b10000101 : 8'b10000100;
												assign node6836 = (inp[3]) ? 8'b10010101 : node6837;
													assign node6837 = (inp[1]) ? 8'b10010100 : 8'b10010101;
											assign node6841 = (inp[6]) ? 8'b11110111 : 8'b10100101;
										assign node6844 = (inp[1]) ? 8'b10000100 : 8'b10000101;
							assign node6847 = (inp[2]) ? node6887 : node6848;
								assign node6848 = (inp[13]) ? node6864 : node6849;
									assign node6849 = (inp[1]) ? node6855 : node6850;
										assign node6850 = (inp[10]) ? node6852 : 8'b10110001;
											assign node6852 = (inp[5]) ? 8'b10110001 : 8'b11110111;
										assign node6855 = (inp[5]) ? 8'b10110000 : node6856;
											assign node6856 = (inp[3]) ? node6860 : node6857;
												assign node6857 = (inp[10]) ? 8'b10110100 : 8'b10110000;
												assign node6860 = (inp[10]) ? 8'b11110111 : 8'b10110001;
									assign node6864 = (inp[1]) ? node6874 : node6865;
										assign node6865 = (inp[5]) ? 8'b10010001 : node6866;
											assign node6866 = (inp[9]) ? node6870 : node6867;
												assign node6867 = (inp[10]) ? 8'b10010101 : 8'b10010001;
												assign node6870 = (inp[10]) ? 8'b11110111 : 8'b10110001;
										assign node6874 = (inp[5]) ? 8'b10010000 : node6875;
											assign node6875 = (inp[9]) ? node6881 : node6876;
												assign node6876 = (inp[3]) ? node6878 : 8'b10010000;
													assign node6878 = (inp[10]) ? 8'b10010101 : 8'b10010001;
												assign node6881 = (inp[3]) ? 8'b10110001 : node6882;
													assign node6882 = (inp[10]) ? 8'b10110100 : 8'b10110000;
								assign node6887 = (inp[13]) ? node6911 : node6888;
									assign node6888 = (inp[1]) ? node6898 : node6889;
										assign node6889 = (inp[5]) ? 8'b10100001 : node6890;
											assign node6890 = (inp[10]) ? node6894 : node6891;
												assign node6891 = (inp[6]) ? 8'b10110001 : 8'b10100001;
												assign node6894 = (inp[6]) ? 8'b11110111 : 8'b10100101;
										assign node6898 = (inp[5]) ? 8'b10100000 : node6899;
											assign node6899 = (inp[6]) ? node6907 : node6900;
												assign node6900 = (inp[3]) ? node6904 : node6901;
													assign node6901 = (inp[10]) ? 8'b10100100 : 8'b10100000;
													assign node6904 = (inp[10]) ? 8'b10100101 : 8'b10100001;
												assign node6907 = (inp[3]) ? 8'b10110001 : 8'b10110000;
									assign node6911 = (inp[5]) ? node6935 : node6912;
										assign node6912 = (inp[9]) ? node6928 : node6913;
											assign node6913 = (inp[6]) ? node6921 : node6914;
												assign node6914 = (inp[10]) ? 8'b10000101 : node6915;
													assign node6915 = (inp[3]) ? 8'b10000001 : node6916;
														assign node6916 = (inp[1]) ? 8'b10000000 : 8'b10000001;
												assign node6921 = (inp[10]) ? node6925 : node6922;
													assign node6922 = (inp[3]) ? 8'b10010001 : 8'b10010000;
													assign node6925 = (inp[1]) ? 8'b10010100 : 8'b10010101;
											assign node6928 = (inp[10]) ? node6932 : node6929;
												assign node6929 = (inp[6]) ? 8'b10110001 : 8'b10100001;
												assign node6932 = (inp[6]) ? 8'b11110111 : 8'b10100101;
										assign node6935 = (inp[1]) ? 8'b10000000 : 8'b10000001;
				assign node6938 = (inp[0]) ? node7148 : node6939;
					assign node6939 = (inp[5]) ? node6941 : 8'b00000010;
						assign node6941 = (inp[2]) ? node7015 : node6942;
							assign node6942 = (inp[3]) ? node6966 : node6943;
								assign node6943 = (inp[10]) ? node6949 : node6944;
									assign node6944 = (inp[13]) ? node6946 : 8'b00000010;
										assign node6946 = (inp[9]) ? 8'b10100000 : 8'b00000010;
									assign node6949 = (inp[8]) ? node6955 : node6950;
										assign node6950 = (inp[13]) ? node6952 : 8'b00000010;
											assign node6952 = (inp[9]) ? 8'b10100000 : 8'b00000010;
										assign node6955 = (inp[11]) ? node6961 : node6956;
											assign node6956 = (inp[13]) ? node6958 : 8'b10000100;
												assign node6958 = (inp[9]) ? 8'b10100100 : 8'b10000100;
											assign node6961 = (inp[13]) ? node6963 : 8'b10100100;
												assign node6963 = (inp[1]) ? 8'b10000100 : 8'b10100100;
								assign node6966 = (inp[1]) ? node6988 : node6967;
									assign node6967 = (inp[10]) ? node6973 : node6968;
										assign node6968 = (inp[13]) ? node6970 : 8'b00000010;
											assign node6970 = (inp[9]) ? 8'b10100000 : 8'b00000010;
										assign node6973 = (inp[8]) ? node6979 : node6974;
											assign node6974 = (inp[13]) ? node6976 : 8'b00000010;
												assign node6976 = (inp[9]) ? 8'b10100000 : 8'b00000010;
											assign node6979 = (inp[11]) ? node6985 : node6980;
												assign node6980 = (inp[9]) ? node6982 : 8'b10000100;
													assign node6982 = (inp[13]) ? 8'b10100100 : 8'b10000100;
												assign node6985 = (inp[13]) ? 8'b10000100 : 8'b10100100;
									assign node6988 = (inp[11]) ? node7004 : node6989;
										assign node6989 = (inp[13]) ? node6995 : node6990;
											assign node6990 = (inp[8]) ? node6992 : 8'b10000001;
												assign node6992 = (inp[10]) ? 8'b10000101 : 8'b10000001;
											assign node6995 = (inp[9]) ? node6999 : node6996;
												assign node6996 = (inp[8]) ? 8'b10000101 : 8'b10000001;
												assign node6999 = (inp[8]) ? node7001 : 8'b10100001;
													assign node7001 = (inp[10]) ? 8'b10100101 : 8'b10100001;
										assign node7004 = (inp[9]) ? node7010 : node7005;
											assign node7005 = (inp[8]) ? node7007 : 8'b10100101;
												assign node7007 = (inp[10]) ? 8'b10100001 : 8'b10100101;
											assign node7010 = (inp[13]) ? 8'b10000101 : node7011;
												assign node7011 = (inp[10]) ? 8'b10100001 : 8'b10100101;
							assign node7015 = (inp[6]) ? node7075 : node7016;
								assign node7016 = (inp[1]) ? node7040 : node7017;
									assign node7017 = (inp[8]) ? node7023 : node7018;
										assign node7018 = (inp[9]) ? node7020 : 8'b00000010;
											assign node7020 = (inp[13]) ? 8'b10100000 : 8'b00000010;
										assign node7023 = (inp[10]) ? node7029 : node7024;
											assign node7024 = (inp[13]) ? node7026 : 8'b00000010;
												assign node7026 = (inp[9]) ? 8'b10100000 : 8'b00000010;
											assign node7029 = (inp[11]) ? node7035 : node7030;
												assign node7030 = (inp[13]) ? node7032 : 8'b10000100;
													assign node7032 = (inp[9]) ? 8'b10100100 : 8'b10000100;
												assign node7035 = (inp[9]) ? node7037 : 8'b10100100;
													assign node7037 = (inp[13]) ? 8'b10000100 : 8'b10100100;
									assign node7040 = (inp[3]) ? node7054 : node7041;
										assign node7041 = (inp[8]) ? node7047 : node7042;
											assign node7042 = (inp[9]) ? node7044 : 8'b00000010;
												assign node7044 = (inp[13]) ? 8'b10100000 : 8'b00000010;
											assign node7047 = (inp[10]) ? node7051 : node7048;
												assign node7048 = (inp[13]) ? 8'b10100000 : 8'b00000010;
												assign node7051 = (inp[13]) ? 8'b10100100 : 8'b10000100;
										assign node7054 = (inp[11]) ? node7062 : node7055;
											assign node7055 = (inp[10]) ? node7057 : 8'b10000001;
												assign node7057 = (inp[8]) ? 8'b10100101 : node7058;
													assign node7058 = (inp[9]) ? 8'b10100001 : 8'b10000001;
											assign node7062 = (inp[13]) ? node7068 : node7063;
												assign node7063 = (inp[8]) ? node7065 : 8'b10100101;
													assign node7065 = (inp[10]) ? 8'b10100001 : 8'b10100101;
												assign node7068 = (inp[8]) ? node7072 : node7069;
													assign node7069 = (inp[9]) ? 8'b10000101 : 8'b10100101;
													assign node7072 = (inp[9]) ? 8'b10000001 : 8'b10100001;
								assign node7075 = (inp[11]) ? node7119 : node7076;
									assign node7076 = (inp[3]) ? node7090 : node7077;
										assign node7077 = (inp[13]) ? node7083 : node7078;
											assign node7078 = (inp[8]) ? node7080 : 8'b10010000;
												assign node7080 = (inp[10]) ? 8'b10010100 : 8'b10010000;
											assign node7083 = (inp[9]) ? node7085 : 8'b10010000;
												assign node7085 = (inp[8]) ? node7087 : 8'b10110000;
													assign node7087 = (inp[10]) ? 8'b10110100 : 8'b10110000;
										assign node7090 = (inp[1]) ? node7106 : node7091;
											assign node7091 = (inp[10]) ? node7097 : node7092;
												assign node7092 = (inp[13]) ? node7094 : 8'b10010000;
													assign node7094 = (inp[9]) ? 8'b10110000 : 8'b10010000;
												assign node7097 = (inp[8]) ? node7101 : node7098;
													assign node7098 = (inp[9]) ? 8'b10110000 : 8'b10010000;
													assign node7101 = (inp[13]) ? node7103 : 8'b10010100;
														assign node7103 = (inp[9]) ? 8'b10110100 : 8'b10010100;
											assign node7106 = (inp[10]) ? node7112 : node7107;
												assign node7107 = (inp[13]) ? node7109 : 8'b10010001;
													assign node7109 = (inp[9]) ? 8'b10110001 : 8'b10010001;
												assign node7112 = (inp[8]) ? node7114 : 8'b10010001;
													assign node7114 = (inp[9]) ? node7116 : 8'b10010101;
														assign node7116 = (inp[13]) ? 8'b11110101 : 8'b10010101;
									assign node7119 = (inp[10]) ? node7131 : node7120;
										assign node7120 = (inp[13]) ? node7126 : node7121;
											assign node7121 = (inp[3]) ? node7123 : 8'b11110101;
												assign node7123 = (inp[8]) ? 8'b11110101 : 8'b10110100;
											assign node7126 = (inp[9]) ? 8'b10010101 : node7127;
												assign node7127 = (inp[1]) ? 8'b10110100 : 8'b11110101;
										assign node7131 = (inp[8]) ? node7139 : node7132;
											assign node7132 = (inp[1]) ? node7134 : 8'b11110101;
												assign node7134 = (inp[9]) ? node7136 : 8'b10110100;
													assign node7136 = (inp[13]) ? 8'b10010100 : 8'b10110100;
											assign node7139 = (inp[1]) ? node7145 : node7140;
												assign node7140 = (inp[13]) ? node7142 : 8'b10110001;
													assign node7142 = (inp[9]) ? 8'b10010001 : 8'b10110001;
												assign node7145 = (inp[3]) ? 8'b10110000 : 8'b10110001;
					assign node7148 = (inp[2]) ? node7250 : node7149;
						assign node7149 = (inp[1]) ? node7183 : node7150;
							assign node7150 = (inp[8]) ? node7158 : node7151;
								assign node7151 = (inp[13]) ? node7153 : 8'b00000010;
									assign node7153 = (inp[5]) ? 8'b10100000 : node7154;
										assign node7154 = (inp[9]) ? 8'b00000010 : 8'b10100000;
								assign node7158 = (inp[5]) ? node7176 : node7159;
									assign node7159 = (inp[10]) ? node7171 : node7160;
										assign node7160 = (inp[11]) ? node7166 : node7161;
											assign node7161 = (inp[13]) ? node7163 : 8'b10000100;
												assign node7163 = (inp[9]) ? 8'b10000100 : 8'b10100100;
											assign node7166 = (inp[13]) ? node7168 : 8'b10100100;
												assign node7168 = (inp[9]) ? 8'b10100100 : 8'b10000100;
										assign node7171 = (inp[13]) ? node7173 : 8'b00000010;
											assign node7173 = (inp[9]) ? 8'b00000010 : 8'b10100000;
									assign node7176 = (inp[13]) ? node7180 : node7177;
										assign node7177 = (inp[11]) ? 8'b10100100 : 8'b10000100;
										assign node7180 = (inp[11]) ? 8'b10000100 : 8'b10100100;
							assign node7183 = (inp[5]) ? node7235 : node7184;
								assign node7184 = (inp[3]) ? node7214 : node7185;
									assign node7185 = (inp[11]) ? node7199 : node7186;
										assign node7186 = (inp[9]) ? node7194 : node7187;
											assign node7187 = (inp[13]) ? node7189 : 8'b10000001;
												assign node7189 = (inp[10]) ? 8'b10100001 : node7190;
													assign node7190 = (inp[8]) ? 8'b10100101 : 8'b10100001;
											assign node7194 = (inp[10]) ? 8'b10000001 : node7195;
												assign node7195 = (inp[8]) ? 8'b10000101 : 8'b10000001;
										assign node7199 = (inp[9]) ? node7209 : node7200;
											assign node7200 = (inp[13]) ? node7204 : node7201;
												assign node7201 = (inp[8]) ? 8'b10100001 : 8'b10100101;
												assign node7204 = (inp[8]) ? node7206 : 8'b10000101;
													assign node7206 = (inp[10]) ? 8'b10000101 : 8'b10000001;
											assign node7209 = (inp[10]) ? 8'b10100101 : node7210;
												assign node7210 = (inp[8]) ? 8'b10100001 : 8'b10100101;
									assign node7214 = (inp[8]) ? node7220 : node7215;
										assign node7215 = (inp[9]) ? 8'b00000010 : node7216;
											assign node7216 = (inp[13]) ? 8'b10100000 : 8'b00000010;
										assign node7220 = (inp[10]) ? node7230 : node7221;
											assign node7221 = (inp[11]) ? node7225 : node7222;
												assign node7222 = (inp[13]) ? 8'b10100100 : 8'b10000100;
												assign node7225 = (inp[9]) ? 8'b10100100 : node7226;
													assign node7226 = (inp[13]) ? 8'b10000100 : 8'b10100100;
											assign node7230 = (inp[9]) ? 8'b00000010 : node7231;
												assign node7231 = (inp[13]) ? 8'b10100000 : 8'b00000010;
								assign node7235 = (inp[11]) ? node7243 : node7236;
									assign node7236 = (inp[8]) ? node7240 : node7237;
										assign node7237 = (inp[13]) ? 8'b10100001 : 8'b10000001;
										assign node7240 = (inp[13]) ? 8'b10100101 : 8'b10000101;
									assign node7243 = (inp[13]) ? node7247 : node7244;
										assign node7244 = (inp[8]) ? 8'b10100001 : 8'b10100101;
										assign node7247 = (inp[8]) ? 8'b10000001 : 8'b10000101;
						assign node7250 = (inp[5]) ? node7394 : node7251;
							assign node7251 = (inp[6]) ? node7323 : node7252;
								assign node7252 = (inp[11]) ? node7286 : node7253;
									assign node7253 = (inp[10]) ? node7273 : node7254;
										assign node7254 = (inp[8]) ? node7264 : node7255;
											assign node7255 = (inp[9]) ? 8'b10010000 : node7256;
												assign node7256 = (inp[13]) ? node7260 : node7257;
													assign node7257 = (inp[1]) ? 8'b10010001 : 8'b10010000;
													assign node7260 = (inp[1]) ? 8'b10110001 : 8'b10110000;
											assign node7264 = (inp[3]) ? node7268 : node7265;
												assign node7265 = (inp[1]) ? 8'b10010101 : 8'b10010100;
												assign node7268 = (inp[13]) ? node7270 : 8'b10010100;
													assign node7270 = (inp[9]) ? 8'b10010100 : 8'b10110100;
										assign node7273 = (inp[1]) ? node7279 : node7274;
											assign node7274 = (inp[13]) ? node7276 : 8'b10010000;
												assign node7276 = (inp[9]) ? 8'b10010000 : 8'b10110000;
											assign node7279 = (inp[3]) ? node7281 : 8'b10010001;
												assign node7281 = (inp[9]) ? 8'b10010000 : node7282;
													assign node7282 = (inp[13]) ? 8'b10110000 : 8'b10010000;
									assign node7286 = (inp[13]) ? node7304 : node7287;
										assign node7287 = (inp[10]) ? node7299 : node7288;
											assign node7288 = (inp[8]) ? node7294 : node7289;
												assign node7289 = (inp[3]) ? 8'b11110101 : node7290;
													assign node7290 = (inp[1]) ? 8'b10110100 : 8'b11110101;
												assign node7294 = (inp[3]) ? 8'b10110001 : node7295;
													assign node7295 = (inp[1]) ? 8'b10110000 : 8'b10110001;
											assign node7299 = (inp[1]) ? node7301 : 8'b11110101;
												assign node7301 = (inp[3]) ? 8'b11110101 : 8'b10110100;
										assign node7304 = (inp[9]) ? node7314 : node7305;
											assign node7305 = (inp[8]) ? node7311 : node7306;
												assign node7306 = (inp[3]) ? 8'b10010101 : node7307;
													assign node7307 = (inp[1]) ? 8'b10010100 : 8'b10010101;
												assign node7311 = (inp[10]) ? 8'b10010101 : 8'b10010001;
											assign node7314 = (inp[3]) ? node7318 : node7315;
												assign node7315 = (inp[1]) ? 8'b10110100 : 8'b11110101;
												assign node7318 = (inp[10]) ? 8'b11110101 : node7319;
													assign node7319 = (inp[8]) ? 8'b10110001 : 8'b11110101;
								assign node7323 = (inp[8]) ? node7347 : node7324;
									assign node7324 = (inp[1]) ? node7330 : node7325;
										assign node7325 = (inp[9]) ? 8'b00000010 : node7326;
											assign node7326 = (inp[13]) ? 8'b10100000 : 8'b00000010;
										assign node7330 = (inp[3]) ? node7342 : node7331;
											assign node7331 = (inp[11]) ? node7337 : node7332;
												assign node7332 = (inp[9]) ? 8'b10000001 : node7333;
													assign node7333 = (inp[13]) ? 8'b10100001 : 8'b10000001;
												assign node7337 = (inp[13]) ? node7339 : 8'b10100101;
													assign node7339 = (inp[10]) ? 8'b10100101 : 8'b10000101;
											assign node7342 = (inp[9]) ? 8'b00000010 : node7343;
												assign node7343 = (inp[13]) ? 8'b10100000 : 8'b00000010;
									assign node7347 = (inp[10]) ? node7375 : node7348;
										assign node7348 = (inp[1]) ? node7360 : node7349;
											assign node7349 = (inp[11]) ? node7355 : node7350;
												assign node7350 = (inp[13]) ? node7352 : 8'b10000100;
													assign node7352 = (inp[9]) ? 8'b10000100 : 8'b10100100;
												assign node7355 = (inp[9]) ? 8'b10100100 : node7356;
													assign node7356 = (inp[3]) ? 8'b10000100 : 8'b10100100;
											assign node7360 = (inp[3]) ? node7370 : node7361;
												assign node7361 = (inp[11]) ? node7367 : node7362;
													assign node7362 = (inp[9]) ? 8'b10000101 : node7363;
														assign node7363 = (inp[13]) ? 8'b10100101 : 8'b10000101;
													assign node7367 = (inp[9]) ? 8'b10100001 : 8'b10000001;
												assign node7370 = (inp[9]) ? 8'b10100100 : node7371;
													assign node7371 = (inp[13]) ? 8'b10000100 : 8'b10100100;
										assign node7375 = (inp[9]) ? node7387 : node7376;
											assign node7376 = (inp[13]) ? node7382 : node7377;
												assign node7377 = (inp[3]) ? 8'b00000010 : node7378;
													assign node7378 = (inp[1]) ? 8'b10100101 : 8'b00000010;
												assign node7382 = (inp[11]) ? node7384 : 8'b10100000;
													assign node7384 = (inp[1]) ? 8'b10000101 : 8'b10100000;
											assign node7387 = (inp[13]) ? node7389 : 8'b00000010;
												assign node7389 = (inp[11]) ? 8'b00000010 : node7390;
													assign node7390 = (inp[3]) ? 8'b00000010 : 8'b10000001;
							assign node7394 = (inp[6]) ? node7426 : node7395;
								assign node7395 = (inp[8]) ? node7411 : node7396;
									assign node7396 = (inp[11]) ? node7404 : node7397;
										assign node7397 = (inp[1]) ? node7401 : node7398;
											assign node7398 = (inp[13]) ? 8'b10110000 : 8'b10010000;
											assign node7401 = (inp[13]) ? 8'b10110001 : 8'b10010001;
										assign node7404 = (inp[1]) ? node7408 : node7405;
											assign node7405 = (inp[13]) ? 8'b10010101 : 8'b11110101;
											assign node7408 = (inp[13]) ? 8'b10010100 : 8'b10110100;
									assign node7411 = (inp[11]) ? node7419 : node7412;
										assign node7412 = (inp[13]) ? node7416 : node7413;
											assign node7413 = (inp[1]) ? 8'b10010101 : 8'b10010100;
											assign node7416 = (inp[1]) ? 8'b11110101 : 8'b10110100;
										assign node7419 = (inp[1]) ? node7423 : node7420;
											assign node7420 = (inp[13]) ? 8'b10010001 : 8'b10110001;
											assign node7423 = (inp[13]) ? 8'b10010000 : 8'b10110000;
								assign node7426 = (inp[10]) ? node7458 : node7427;
									assign node7427 = (inp[13]) ? node7443 : node7428;
										assign node7428 = (inp[11]) ? node7436 : node7429;
											assign node7429 = (inp[8]) ? node7433 : node7430;
												assign node7430 = (inp[1]) ? 8'b10010001 : 8'b10010000;
												assign node7433 = (inp[1]) ? 8'b10010101 : 8'b10010100;
											assign node7436 = (inp[8]) ? node7440 : node7437;
												assign node7437 = (inp[1]) ? 8'b10110100 : 8'b11110101;
												assign node7440 = (inp[1]) ? 8'b10110000 : 8'b10110001;
										assign node7443 = (inp[11]) ? node7451 : node7444;
											assign node7444 = (inp[8]) ? node7448 : node7445;
												assign node7445 = (inp[1]) ? 8'b10110001 : 8'b10110000;
												assign node7448 = (inp[1]) ? 8'b11110101 : 8'b10110100;
											assign node7451 = (inp[8]) ? node7455 : node7452;
												assign node7452 = (inp[1]) ? 8'b10010100 : 8'b10010101;
												assign node7455 = (inp[1]) ? 8'b10010000 : 8'b10010001;
									assign node7458 = (inp[13]) ? node7474 : node7459;
										assign node7459 = (inp[11]) ? node7467 : node7460;
											assign node7460 = (inp[1]) ? node7464 : node7461;
												assign node7461 = (inp[8]) ? 8'b10010100 : 8'b10010000;
												assign node7464 = (inp[8]) ? 8'b10010101 : 8'b10010001;
											assign node7467 = (inp[1]) ? node7471 : node7468;
												assign node7468 = (inp[8]) ? 8'b10110001 : 8'b11110101;
												assign node7471 = (inp[8]) ? 8'b10110000 : 8'b10110100;
										assign node7474 = (inp[11]) ? node7482 : node7475;
											assign node7475 = (inp[1]) ? node7479 : node7476;
												assign node7476 = (inp[8]) ? 8'b10110100 : 8'b10110000;
												assign node7479 = (inp[8]) ? 8'b11110101 : 8'b10110001;
											assign node7482 = (inp[8]) ? node7486 : node7483;
												assign node7483 = (inp[1]) ? 8'b10010100 : 8'b10010101;
												assign node7486 = (inp[1]) ? 8'b10010000 : 8'b10010001;

endmodule